module basic_3000_30000_3500_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2172,In_1004);
xnor U1 (N_1,In_898,In_978);
nand U2 (N_2,In_1325,In_1056);
or U3 (N_3,In_2344,In_1040);
or U4 (N_4,In_1238,In_1990);
and U5 (N_5,In_156,In_2654);
nor U6 (N_6,In_2576,In_1305);
or U7 (N_7,In_2783,In_1998);
or U8 (N_8,In_2176,In_2279);
or U9 (N_9,In_130,In_326);
nand U10 (N_10,In_1596,In_1367);
nand U11 (N_11,In_2968,In_373);
nand U12 (N_12,In_2212,In_313);
xnor U13 (N_13,In_1250,In_2633);
nand U14 (N_14,In_2864,In_1132);
or U15 (N_15,In_2733,In_2425);
xor U16 (N_16,In_983,In_1117);
nor U17 (N_17,In_1219,In_654);
or U18 (N_18,In_2025,In_371);
nand U19 (N_19,In_1949,In_580);
xor U20 (N_20,In_1186,In_2362);
and U21 (N_21,In_778,In_1463);
nor U22 (N_22,In_2415,In_2996);
or U23 (N_23,In_2985,In_1717);
and U24 (N_24,In_1648,In_2655);
or U25 (N_25,In_2014,In_2874);
nor U26 (N_26,In_821,In_819);
and U27 (N_27,In_2159,In_248);
xnor U28 (N_28,In_1271,In_1360);
nor U29 (N_29,In_2787,In_483);
and U30 (N_30,In_2095,In_2630);
xnor U31 (N_31,In_1289,In_2717);
and U32 (N_32,In_28,In_1541);
nand U33 (N_33,In_91,In_1458);
or U34 (N_34,In_452,In_1549);
nor U35 (N_35,In_1881,In_1165);
xor U36 (N_36,In_1939,In_647);
nand U37 (N_37,In_2522,In_1506);
or U38 (N_38,In_1461,In_1175);
nand U39 (N_39,In_784,In_1850);
nand U40 (N_40,In_1296,In_1788);
and U41 (N_41,In_1265,In_1602);
or U42 (N_42,In_2225,In_257);
xnor U43 (N_43,In_1443,In_1932);
nor U44 (N_44,In_1335,In_1194);
or U45 (N_45,In_1198,In_844);
nor U46 (N_46,In_2183,In_2908);
nand U47 (N_47,In_1757,In_2677);
and U48 (N_48,In_22,In_1083);
and U49 (N_49,In_2177,In_935);
or U50 (N_50,In_2674,In_2647);
nor U51 (N_51,In_2338,In_595);
nor U52 (N_52,In_552,In_1827);
and U53 (N_53,In_502,In_2136);
xor U54 (N_54,In_2353,In_2949);
or U55 (N_55,In_1590,In_1502);
nor U56 (N_56,In_2537,In_2430);
nor U57 (N_57,In_2644,In_1306);
nand U58 (N_58,In_510,In_615);
or U59 (N_59,In_9,In_826);
xor U60 (N_60,In_1753,In_1387);
and U61 (N_61,In_1770,In_2170);
xor U62 (N_62,In_1798,In_2565);
nor U63 (N_63,In_669,In_2347);
and U64 (N_64,In_2959,In_2946);
xnor U65 (N_65,In_2967,In_2632);
and U66 (N_66,In_1014,In_2020);
xnor U67 (N_67,In_136,In_1038);
nor U68 (N_68,In_2847,In_2640);
xor U69 (N_69,In_1046,In_512);
and U70 (N_70,In_2107,In_1503);
or U71 (N_71,In_956,In_410);
and U72 (N_72,In_1828,In_2732);
nand U73 (N_73,In_58,In_707);
xor U74 (N_74,In_2913,In_129);
and U75 (N_75,In_1003,In_1294);
xor U76 (N_76,In_2273,In_633);
nand U77 (N_77,In_1136,In_1779);
nand U78 (N_78,In_1584,In_150);
nor U79 (N_79,In_177,In_2018);
nor U80 (N_80,In_2198,In_26);
nand U81 (N_81,In_1483,In_584);
xnor U82 (N_82,In_1350,In_2178);
and U83 (N_83,In_815,In_1893);
and U84 (N_84,In_210,In_1634);
nor U85 (N_85,In_2068,In_2998);
xor U86 (N_86,In_906,In_397);
and U87 (N_87,In_662,In_916);
nor U88 (N_88,In_2307,In_1459);
nor U89 (N_89,In_2157,In_269);
nor U90 (N_90,In_937,In_1910);
and U91 (N_91,In_2373,In_114);
and U92 (N_92,In_2502,In_539);
nor U93 (N_93,In_1169,In_2120);
nand U94 (N_94,In_742,In_2317);
nand U95 (N_95,In_325,In_2324);
nor U96 (N_96,In_2762,In_2560);
or U97 (N_97,In_630,In_1599);
xor U98 (N_98,In_2870,In_557);
and U99 (N_99,In_886,In_69);
nand U100 (N_100,In_1865,In_2991);
xnor U101 (N_101,In_417,In_550);
xor U102 (N_102,In_2849,In_1532);
nand U103 (N_103,In_2272,In_2501);
nand U104 (N_104,In_2906,In_2485);
or U105 (N_105,In_1775,In_2639);
nor U106 (N_106,In_641,In_1287);
or U107 (N_107,In_631,In_1669);
nor U108 (N_108,In_1478,In_266);
nand U109 (N_109,In_2687,In_1254);
nand U110 (N_110,In_2971,In_1191);
nor U111 (N_111,In_207,In_1394);
xor U112 (N_112,In_1516,In_1122);
or U113 (N_113,In_1741,In_2545);
nor U114 (N_114,In_2993,In_2734);
xnor U115 (N_115,In_2758,In_1232);
nand U116 (N_116,In_1301,In_2327);
xor U117 (N_117,In_816,In_594);
xnor U118 (N_118,In_2500,In_693);
or U119 (N_119,In_1748,In_2541);
nand U120 (N_120,In_2599,In_51);
nor U121 (N_121,In_2749,In_532);
nand U122 (N_122,In_2603,In_831);
nor U123 (N_123,In_974,In_708);
or U124 (N_124,In_888,In_49);
xnor U125 (N_125,In_426,In_1552);
or U126 (N_126,In_2166,In_1563);
nand U127 (N_127,In_219,In_2323);
or U128 (N_128,In_208,In_2466);
xor U129 (N_129,In_2770,In_475);
nand U130 (N_130,In_2715,In_212);
xor U131 (N_131,In_567,In_88);
and U132 (N_132,In_1667,In_1268);
nand U133 (N_133,In_1654,In_202);
and U134 (N_134,In_1534,In_2461);
nand U135 (N_135,In_2050,In_802);
or U136 (N_136,In_501,In_1149);
xnor U137 (N_137,In_220,In_2316);
or U138 (N_138,In_193,In_1120);
nand U139 (N_139,In_1135,In_1057);
xor U140 (N_140,In_195,In_702);
xnor U141 (N_141,In_1639,In_1189);
xnor U142 (N_142,In_1069,In_1575);
nand U143 (N_143,In_2479,In_2840);
nor U144 (N_144,In_1744,In_1288);
xnor U145 (N_145,In_2671,In_2151);
and U146 (N_146,In_198,In_1550);
xor U147 (N_147,In_2547,In_2072);
and U148 (N_148,In_736,In_1846);
nor U149 (N_149,In_2422,In_950);
xor U150 (N_150,In_21,In_574);
or U151 (N_151,In_1433,In_2217);
xnor U152 (N_152,In_454,In_64);
nor U153 (N_153,In_1233,In_1486);
nor U154 (N_154,In_1172,In_1222);
or U155 (N_155,In_2828,In_2478);
or U156 (N_156,In_1774,In_1213);
xnor U157 (N_157,In_321,In_598);
xnor U158 (N_158,In_2100,In_1687);
nor U159 (N_159,In_1002,In_2322);
nand U160 (N_160,In_482,In_1264);
xor U161 (N_161,In_1344,In_60);
or U162 (N_162,In_790,In_846);
nand U163 (N_163,In_1855,In_2363);
and U164 (N_164,In_2296,In_2423);
and U165 (N_165,In_1454,In_2061);
nor U166 (N_166,In_139,In_2085);
and U167 (N_167,In_309,In_30);
or U168 (N_168,In_1036,In_1784);
and U169 (N_169,In_2337,In_2613);
nand U170 (N_170,In_2402,In_2044);
and U171 (N_171,In_667,In_1908);
xor U172 (N_172,In_2258,In_806);
nor U173 (N_173,In_1961,In_2480);
or U174 (N_174,In_1338,In_1638);
nand U175 (N_175,In_2079,In_853);
and U176 (N_176,In_2440,In_2702);
xnor U177 (N_177,In_1522,In_2574);
nand U178 (N_178,In_880,In_770);
nand U179 (N_179,In_1256,In_666);
nand U180 (N_180,In_132,In_2761);
or U181 (N_181,In_684,In_1391);
or U182 (N_182,In_2333,In_356);
and U183 (N_183,In_663,In_2407);
nand U184 (N_184,In_2167,In_1916);
and U185 (N_185,In_834,In_432);
nor U186 (N_186,In_20,In_2054);
and U187 (N_187,In_2988,In_2452);
xnor U188 (N_188,In_2231,In_1032);
nand U189 (N_189,In_1592,In_1684);
nand U190 (N_190,In_133,In_490);
and U191 (N_191,In_968,In_931);
nor U192 (N_192,In_2990,In_2298);
nor U193 (N_193,In_2028,In_610);
xor U194 (N_194,In_2016,In_1464);
xor U195 (N_195,In_710,In_2306);
or U196 (N_196,In_2340,In_1446);
nand U197 (N_197,In_1363,In_2150);
nand U198 (N_198,In_32,In_1691);
xnor U199 (N_199,In_342,In_1204);
nand U200 (N_200,In_351,In_1432);
nor U201 (N_201,In_2449,In_1772);
or U202 (N_202,In_2303,In_290);
xor U203 (N_203,In_1714,In_786);
xor U204 (N_204,In_749,In_733);
and U205 (N_205,In_79,In_244);
nand U206 (N_206,In_920,In_186);
xnor U207 (N_207,In_913,In_750);
xor U208 (N_208,In_1523,In_160);
xnor U209 (N_209,In_1969,In_153);
and U210 (N_210,In_2330,In_521);
nand U211 (N_211,In_1632,In_2263);
and U212 (N_212,In_2725,In_1630);
and U213 (N_213,In_1600,In_830);
and U214 (N_214,In_1157,In_360);
or U215 (N_215,In_2741,In_1514);
or U216 (N_216,In_1399,In_1096);
or U217 (N_217,In_1314,In_839);
and U218 (N_218,In_2123,In_973);
nand U219 (N_219,In_71,In_1824);
xor U220 (N_220,In_2372,In_1508);
nor U221 (N_221,In_2934,In_2726);
nor U222 (N_222,In_1412,In_2437);
nand U223 (N_223,In_1031,In_2714);
or U224 (N_224,In_2370,In_315);
and U225 (N_225,In_458,In_2048);
nand U226 (N_226,In_436,In_2692);
nor U227 (N_227,In_1723,In_120);
xor U228 (N_228,In_1938,In_355);
xnor U229 (N_229,In_2135,In_1809);
nor U230 (N_230,In_2591,In_1569);
nand U231 (N_231,In_2209,In_2510);
and U232 (N_232,In_2800,In_2257);
and U233 (N_233,In_1831,In_1776);
and U234 (N_234,In_2341,In_180);
xor U235 (N_235,In_370,In_489);
and U236 (N_236,In_1535,In_1322);
nor U237 (N_237,In_239,In_1043);
nand U238 (N_238,In_465,In_1517);
nor U239 (N_239,In_1139,In_624);
nand U240 (N_240,In_369,In_542);
or U241 (N_241,In_1123,In_1303);
or U242 (N_242,In_767,In_2262);
and U243 (N_243,In_1261,In_1479);
and U244 (N_244,In_72,In_1022);
or U245 (N_245,In_2109,In_1718);
and U246 (N_246,In_2181,In_1329);
and U247 (N_247,In_1641,In_1848);
and U248 (N_248,In_506,In_2852);
nand U249 (N_249,In_2582,In_1429);
and U250 (N_250,In_2983,In_2361);
nor U251 (N_251,In_1722,In_1284);
and U252 (N_252,In_1366,In_1073);
nand U253 (N_253,In_2794,In_1988);
and U254 (N_254,In_1635,In_723);
nor U255 (N_255,In_627,In_855);
nor U256 (N_256,In_587,In_1889);
and U257 (N_257,In_704,In_35);
nor U258 (N_258,In_1763,In_466);
xor U259 (N_259,In_2237,In_1469);
xor U260 (N_260,In_528,In_1524);
nand U261 (N_261,In_1343,In_398);
nand U262 (N_262,In_1390,In_2943);
xnor U263 (N_263,In_15,In_927);
and U264 (N_264,In_2266,In_1904);
nand U265 (N_265,In_1981,In_2684);
or U266 (N_266,In_1959,In_2679);
xnor U267 (N_267,In_444,In_2807);
nand U268 (N_268,In_1739,In_1864);
xor U269 (N_269,In_2234,In_2464);
or U270 (N_270,In_1234,In_586);
nand U271 (N_271,In_963,In_2477);
nand U272 (N_272,In_2657,In_656);
nand U273 (N_273,In_2778,In_1414);
nor U274 (N_274,In_2888,In_86);
or U275 (N_275,In_304,In_1001);
xnor U276 (N_276,In_1487,In_1808);
nor U277 (N_277,In_1312,In_457);
nand U278 (N_278,In_2859,In_1688);
nor U279 (N_279,In_1041,In_2976);
nor U280 (N_280,In_2301,In_1504);
nand U281 (N_281,In_803,In_412);
and U282 (N_282,In_664,In_1629);
nor U283 (N_283,In_2954,In_1033);
or U284 (N_284,In_2763,In_1019);
nor U285 (N_285,In_866,In_1088);
nor U286 (N_286,In_2948,In_1193);
nand U287 (N_287,In_2282,In_213);
nand U288 (N_288,In_876,In_1823);
or U289 (N_289,In_459,In_2809);
and U290 (N_290,In_1407,In_2346);
nand U291 (N_291,In_2666,In_1293);
nand U292 (N_292,In_2359,In_1890);
or U293 (N_293,In_225,In_2682);
nand U294 (N_294,In_516,In_845);
and U295 (N_295,In_828,In_2270);
xor U296 (N_296,In_2543,In_1931);
xnor U297 (N_297,In_1365,In_1993);
or U298 (N_298,In_1045,In_553);
nor U299 (N_299,In_2869,In_2618);
nand U300 (N_300,In_544,In_2454);
nor U301 (N_301,In_1114,In_520);
and U302 (N_302,In_697,In_1530);
or U303 (N_303,In_1372,In_1614);
nand U304 (N_304,In_1983,In_78);
and U305 (N_305,In_358,In_2345);
or U306 (N_306,In_2116,In_1126);
and U307 (N_307,In_1460,In_2131);
nor U308 (N_308,In_525,In_1124);
or U309 (N_309,In_2535,In_622);
nand U310 (N_310,In_840,In_1593);
xnor U311 (N_311,In_2804,In_2445);
nand U312 (N_312,In_409,In_348);
or U313 (N_313,In_1564,In_1374);
nor U314 (N_314,In_798,In_289);
xnor U315 (N_315,In_1173,In_965);
and U316 (N_316,In_2163,In_2049);
nand U317 (N_317,In_1184,In_124);
and U318 (N_318,In_1199,In_1903);
and U319 (N_319,In_1520,In_1274);
or U320 (N_320,In_1963,In_1105);
nor U321 (N_321,In_2751,In_299);
or U322 (N_322,In_546,In_1397);
nand U323 (N_323,In_1279,In_993);
and U324 (N_324,In_897,In_1146);
or U325 (N_325,In_2469,In_2436);
nand U326 (N_326,In_157,In_2488);
or U327 (N_327,In_357,In_1162);
xnor U328 (N_328,In_2861,In_854);
xor U329 (N_329,In_576,In_365);
nand U330 (N_330,In_445,In_343);
xor U331 (N_331,In_229,In_1385);
xor U332 (N_332,In_2053,In_2635);
xor U333 (N_333,In_825,In_2788);
and U334 (N_334,In_1767,In_1352);
or U335 (N_335,In_2841,In_1392);
nand U336 (N_336,In_665,In_2928);
xor U337 (N_337,In_2705,In_1104);
and U338 (N_338,In_675,In_1950);
or U339 (N_339,In_1286,In_901);
nor U340 (N_340,In_2592,In_275);
and U341 (N_341,In_1396,In_566);
or U342 (N_342,In_141,In_2070);
or U343 (N_343,In_2111,In_147);
nor U344 (N_344,In_2190,In_1710);
or U345 (N_345,In_2977,In_2314);
and U346 (N_346,In_1769,In_564);
nand U347 (N_347,In_2706,In_969);
and U348 (N_348,In_638,In_2408);
and U349 (N_349,In_2838,In_1121);
nand U350 (N_350,In_2332,In_1176);
and U351 (N_351,In_1016,In_431);
nor U352 (N_352,In_1877,In_2607);
xor U353 (N_353,In_2696,In_81);
nand U354 (N_354,In_685,In_1768);
nand U355 (N_355,In_440,In_914);
and U356 (N_356,In_366,In_2058);
nor U357 (N_357,In_2649,In_590);
nor U358 (N_358,In_1834,In_1462);
xnor U359 (N_359,In_2130,In_218);
nand U360 (N_360,In_2989,In_2811);
nor U361 (N_361,In_2304,In_2069);
and U362 (N_362,In_2785,In_2094);
and U363 (N_363,In_1456,In_893);
and U364 (N_364,In_2052,In_1512);
nor U365 (N_365,In_628,In_1738);
or U366 (N_366,In_1851,In_1644);
xor U367 (N_367,In_2339,In_2113);
and U368 (N_368,In_719,In_2772);
nor U369 (N_369,In_1061,In_2115);
nand U370 (N_370,In_1854,In_860);
nand U371 (N_371,In_1997,In_1160);
or U372 (N_372,In_2595,In_1485);
and U373 (N_373,In_1900,In_560);
or U374 (N_374,In_581,In_895);
and U375 (N_375,In_2970,In_2222);
xnor U376 (N_376,In_1490,In_1295);
xor U377 (N_377,In_1106,In_1473);
and U378 (N_378,In_2561,In_1507);
nor U379 (N_379,In_77,In_2816);
xnor U380 (N_380,In_2686,In_2268);
and U381 (N_381,In_894,In_1451);
nor U382 (N_382,In_1536,In_2134);
nor U383 (N_383,In_1472,In_649);
and U384 (N_384,In_1861,In_464);
nor U385 (N_385,In_1039,In_256);
or U386 (N_386,In_1928,In_1488);
and U387 (N_387,In_1230,In_818);
nor U388 (N_388,In_555,In_43);
and U389 (N_389,In_2830,In_1426);
nand U390 (N_390,In_1337,In_2597);
and U391 (N_391,In_2004,In_462);
nand U392 (N_392,In_2865,In_480);
or U393 (N_393,In_722,In_1844);
nor U394 (N_394,In_728,In_2931);
and U395 (N_395,In_2244,In_961);
and U396 (N_396,In_2042,In_1428);
and U397 (N_397,In_1578,In_2155);
nor U398 (N_398,In_849,In_1170);
xor U399 (N_399,In_776,In_1996);
and U400 (N_400,In_2146,In_1421);
xnor U401 (N_401,In_1181,In_2627);
nand U402 (N_402,In_703,In_804);
and U403 (N_403,In_944,In_2264);
xor U404 (N_404,In_972,In_2662);
xnor U405 (N_405,In_478,In_2559);
xor U406 (N_406,In_907,In_2017);
nand U407 (N_407,In_2277,In_1849);
and U408 (N_408,In_2707,In_2295);
nand U409 (N_409,In_1558,In_1869);
nand U410 (N_410,In_903,In_2680);
and U411 (N_411,In_1821,In_1099);
nand U412 (N_412,In_899,In_2133);
xnor U413 (N_413,In_2676,In_1804);
xor U414 (N_414,In_883,In_2200);
nand U415 (N_415,In_2238,In_497);
xor U416 (N_416,In_161,In_2621);
and U417 (N_417,In_2216,In_190);
nand U418 (N_418,In_1663,In_541);
nor U419 (N_419,In_2005,In_1955);
nand U420 (N_420,In_1567,In_1166);
nand U421 (N_421,In_2256,In_1);
or U422 (N_422,In_1946,In_2428);
or U423 (N_423,In_1612,In_2585);
xnor U424 (N_424,In_2494,In_154);
nand U425 (N_425,In_2392,In_1690);
and U426 (N_426,In_1237,In_1859);
nand U427 (N_427,In_1304,In_2568);
xnor U428 (N_428,In_1972,In_2174);
nand U429 (N_429,In_2031,In_771);
nor U430 (N_430,In_286,In_2067);
xnor U431 (N_431,In_508,In_453);
nand U432 (N_432,In_183,In_1084);
nor U433 (N_433,In_294,In_984);
or U434 (N_434,In_2360,In_2775);
xnor U435 (N_435,In_1212,In_942);
xnor U436 (N_436,In_1449,In_2584);
nor U437 (N_437,In_1979,In_2802);
nor U438 (N_438,In_354,In_1049);
xor U439 (N_439,In_2416,In_469);
xnor U440 (N_440,In_987,In_1027);
and U441 (N_441,In_1090,In_1430);
xor U442 (N_442,In_1918,In_339);
or U443 (N_443,In_1349,In_347);
or U444 (N_444,In_499,In_1205);
nor U445 (N_445,In_2528,In_2207);
or U446 (N_446,In_970,In_2080);
nand U447 (N_447,In_1499,In_1403);
and U448 (N_448,In_394,In_588);
and U449 (N_449,In_1163,In_0);
nor U450 (N_450,In_632,In_6);
and U451 (N_451,In_1994,In_2299);
xnor U452 (N_452,In_2420,In_1856);
or U453 (N_453,In_1661,In_1554);
or U454 (N_454,In_1275,In_245);
and U455 (N_455,In_1902,In_115);
nor U456 (N_456,In_250,In_2564);
xnor U457 (N_457,In_2719,In_2197);
or U458 (N_458,In_1659,In_376);
nor U459 (N_459,In_1214,In_2187);
and U460 (N_460,In_1929,In_1225);
xnor U461 (N_461,In_1773,In_882);
xnor U462 (N_462,In_389,In_2140);
xnor U463 (N_463,In_332,In_1899);
xnor U464 (N_464,In_2090,In_2383);
nand U465 (N_465,In_2318,In_1072);
or U466 (N_466,In_735,In_117);
nor U467 (N_467,In_1130,In_2458);
or U468 (N_468,In_2944,In_781);
nor U469 (N_469,In_1476,In_2819);
nor U470 (N_470,In_892,In_2619);
xnor U471 (N_471,In_2076,In_1450);
xnor U472 (N_472,In_1044,In_90);
xnor U473 (N_473,In_303,In_2409);
and U474 (N_474,In_2995,In_138);
and U475 (N_475,In_939,In_1964);
nor U476 (N_476,In_1777,In_89);
xor U477 (N_477,In_434,In_600);
nor U478 (N_478,In_2942,In_441);
nand U479 (N_479,In_2395,In_2589);
nand U480 (N_480,In_1319,In_2448);
and U481 (N_481,In_2315,In_850);
xor U482 (N_482,In_2259,In_1885);
or U483 (N_483,In_2697,In_137);
nor U484 (N_484,In_199,In_2508);
nor U485 (N_485,In_695,In_813);
nand U486 (N_486,In_1064,In_2043);
xnor U487 (N_487,In_1062,In_1542);
and U488 (N_488,In_1974,In_1074);
and U489 (N_489,In_748,In_1252);
nor U490 (N_490,In_926,In_1574);
nor U491 (N_491,In_585,In_2355);
and U492 (N_492,In_990,In_2118);
and U493 (N_493,In_423,In_573);
nor U494 (N_494,In_548,In_1431);
or U495 (N_495,In_173,In_1050);
or U496 (N_496,In_395,In_650);
nor U497 (N_497,In_1422,In_2594);
or U498 (N_498,In_1771,In_2401);
nor U499 (N_499,In_236,In_1551);
nand U500 (N_500,In_668,In_755);
or U501 (N_501,In_1799,In_2010);
nand U502 (N_502,In_2860,In_655);
and U503 (N_503,In_2201,In_887);
nor U504 (N_504,In_2128,In_769);
nor U505 (N_505,In_2210,In_2737);
xor U506 (N_506,In_1028,In_381);
or U507 (N_507,In_865,In_2419);
or U508 (N_508,In_2986,In_2798);
nor U509 (N_509,In_2795,In_337);
xor U510 (N_510,In_267,In_2443);
or U511 (N_511,In_1381,In_252);
nor U512 (N_512,In_2064,In_915);
nand U513 (N_513,In_2290,In_1424);
or U514 (N_514,In_329,In_2921);
or U515 (N_515,In_2211,In_1406);
nand U516 (N_516,In_1326,In_82);
or U517 (N_517,In_639,In_636);
and U518 (N_518,In_2175,In_1342);
nand U519 (N_519,In_258,In_2941);
or U520 (N_520,In_2412,In_2185);
nand U521 (N_521,In_2624,In_2570);
xnor U522 (N_522,In_2586,In_285);
nand U523 (N_523,In_1196,In_1317);
nor U524 (N_524,In_1379,In_2144);
xnor U525 (N_525,In_446,In_2291);
nor U526 (N_526,In_611,In_2081);
nand U527 (N_527,In_113,In_2801);
nand U528 (N_528,In_1448,In_2935);
xnor U529 (N_529,In_2121,In_33);
or U530 (N_530,In_1701,In_959);
nand U531 (N_531,In_2202,In_2265);
and U532 (N_532,In_529,In_1680);
nand U533 (N_533,In_163,In_450);
and U534 (N_534,In_1615,In_323);
and U535 (N_535,In_2831,In_1709);
and U536 (N_536,In_2953,In_2156);
nand U537 (N_537,In_2404,In_2558);
xnor U538 (N_538,In_1605,In_1220);
or U539 (N_539,In_2927,In_2767);
nor U540 (N_540,In_1420,In_1207);
or U541 (N_541,In_380,In_146);
nand U542 (N_542,In_2368,In_2792);
and U543 (N_543,In_2255,In_715);
nand U544 (N_544,In_2057,In_1333);
or U545 (N_545,In_1948,In_1236);
nor U546 (N_546,In_2651,In_2451);
nand U547 (N_547,In_2148,In_2837);
nand U548 (N_548,In_1470,In_2406);
xor U549 (N_549,In_2235,In_1501);
nor U550 (N_550,In_689,In_148);
xor U551 (N_551,In_925,In_1670);
nor U552 (N_552,In_1556,In_2722);
xor U553 (N_553,In_794,In_718);
xor U554 (N_554,In_55,In_683);
nand U555 (N_555,In_928,In_2472);
xnor U556 (N_556,In_374,In_2773);
or U557 (N_557,In_2875,In_1082);
or U558 (N_558,In_1618,In_463);
nand U559 (N_559,In_2089,In_1671);
or U560 (N_560,In_27,In_877);
or U561 (N_561,In_2759,In_701);
nand U562 (N_562,In_172,In_2509);
or U563 (N_563,In_2367,In_2895);
xnor U564 (N_564,In_178,In_2139);
xnor U565 (N_565,In_4,In_1110);
nor U566 (N_566,In_1947,In_1907);
nor U567 (N_567,In_2497,In_396);
or U568 (N_568,In_1962,In_1692);
and U569 (N_569,In_1307,In_2387);
nand U570 (N_570,In_859,In_492);
nor U571 (N_571,In_407,In_1498);
nor U572 (N_572,In_411,In_948);
xnor U573 (N_573,In_421,In_2384);
and U574 (N_574,In_673,In_85);
or U575 (N_575,In_1382,In_1359);
nand U576 (N_576,In_982,In_2192);
nor U577 (N_577,In_583,In_1762);
nand U578 (N_578,In_2499,In_455);
nand U579 (N_579,In_2938,In_1395);
xnor U580 (N_580,In_1624,In_2742);
and U581 (N_581,In_1491,In_1030);
or U582 (N_582,In_1971,In_1562);
and U583 (N_583,In_2835,In_793);
nand U584 (N_584,In_2455,In_2284);
nor U585 (N_585,In_1797,In_2041);
nand U586 (N_586,In_1790,In_2780);
nor U587 (N_587,In_1633,In_1310);
or U588 (N_588,In_558,In_1883);
xor U589 (N_589,In_2336,In_2769);
xor U590 (N_590,In_2484,In_1133);
xor U591 (N_591,In_659,In_2723);
or U592 (N_592,In_292,In_2029);
or U593 (N_593,In_39,In_795);
xnor U594 (N_594,In_863,In_1140);
or U595 (N_595,In_2369,In_827);
and U596 (N_596,In_318,In_958);
nor U597 (N_597,In_1521,In_308);
nand U598 (N_598,In_383,In_2305);
or U599 (N_599,In_1566,In_1007);
and U600 (N_600,In_1277,In_1698);
and U601 (N_601,In_791,In_929);
or U602 (N_602,In_2879,In_2721);
or U603 (N_603,In_1837,In_1868);
nor U604 (N_604,In_2180,In_1005);
nand U605 (N_605,In_111,In_2429);
nor U606 (N_606,In_596,In_368);
and U607 (N_607,In_559,In_569);
xor U608 (N_608,In_44,In_851);
and U609 (N_609,In_2129,In_1200);
or U610 (N_610,In_765,In_2781);
xnor U611 (N_611,In_1740,In_2260);
nand U612 (N_612,In_1571,In_255);
nand U613 (N_613,In_1111,In_1628);
or U614 (N_614,In_1715,In_941);
or U615 (N_615,In_1724,In_2786);
or U616 (N_616,In_2239,In_2376);
and U617 (N_617,In_428,In_2973);
xnor U618 (N_618,In_2527,In_1818);
nor U619 (N_619,In_1138,In_367);
nand U620 (N_620,In_829,In_23);
nand U621 (N_621,In_2313,In_232);
or U622 (N_622,In_919,In_1743);
or U623 (N_623,In_524,In_2963);
nand U624 (N_624,In_2810,In_716);
or U625 (N_625,In_2598,In_1968);
nor U626 (N_626,In_2542,In_536);
nand U627 (N_627,In_1258,In_1666);
nor U628 (N_628,In_328,In_1273);
nor U629 (N_629,In_1276,In_1154);
and U630 (N_630,In_1065,In_2907);
and U631 (N_631,In_2374,In_1283);
or U632 (N_632,In_2743,In_2951);
xnor U633 (N_633,In_2024,In_674);
nand U634 (N_634,In_125,In_1477);
xor U635 (N_635,In_1023,In_1785);
nor U636 (N_636,In_2171,In_796);
nor U637 (N_637,In_832,In_2065);
xor U638 (N_638,In_1298,In_601);
xor U639 (N_639,In_2824,In_1453);
nor U640 (N_640,In_1547,In_1197);
xor U641 (N_641,In_938,In_2033);
or U642 (N_642,In_391,In_743);
nand U643 (N_643,In_1711,In_260);
and U644 (N_644,In_2731,In_182);
or U645 (N_645,In_2579,In_2311);
and U646 (N_646,In_1812,In_1142);
nand U647 (N_647,In_2482,In_1015);
xnor U648 (N_648,In_1010,In_1086);
and U649 (N_649,In_327,In_485);
nand U650 (N_650,In_1909,In_1914);
xor U651 (N_651,In_1822,In_676);
or U652 (N_652,In_2735,In_2650);
and U653 (N_653,In_2213,In_1249);
or U654 (N_654,In_2283,In_991);
or U655 (N_655,In_1920,In_2514);
nand U656 (N_656,In_1009,In_2612);
and U657 (N_657,In_1857,In_2799);
nor U658 (N_658,In_319,In_1291);
nand U659 (N_659,In_364,In_2059);
nand U660 (N_660,In_1936,In_543);
xor U661 (N_661,In_1223,In_295);
nand U662 (N_662,In_1465,In_1548);
nor U663 (N_663,In_2668,In_2453);
or U664 (N_664,In_2890,In_2342);
and U665 (N_665,In_1021,In_2920);
nand U666 (N_666,In_2750,In_1789);
xor U667 (N_667,In_1467,In_1841);
nand U668 (N_668,In_1353,In_134);
xor U669 (N_669,In_1315,In_2538);
or U670 (N_670,In_1604,In_320);
nand U671 (N_671,In_1802,In_997);
nand U672 (N_672,In_112,In_2771);
and U673 (N_673,In_951,In_2739);
nor U674 (N_674,In_498,In_2932);
nand U675 (N_675,In_672,In_1655);
nand U676 (N_676,In_1853,In_2903);
xnor U677 (N_677,In_317,In_175);
xor U678 (N_678,In_2507,In_783);
nor U679 (N_679,In_1585,In_954);
or U680 (N_680,In_1697,In_2587);
xnor U681 (N_681,In_814,In_2611);
nand U682 (N_682,In_1966,In_2729);
xor U683 (N_683,In_1606,In_609);
or U684 (N_684,In_87,In_2540);
nand U685 (N_685,In_2470,In_1647);
xor U686 (N_686,In_989,In_884);
nor U687 (N_687,In_1119,In_1330);
xnor U688 (N_688,In_2459,In_1080);
nor U689 (N_689,In_556,In_1076);
or U690 (N_690,In_1839,In_108);
xor U691 (N_691,In_1079,In_1863);
xnor U692 (N_692,In_1063,In_413);
xor U693 (N_693,In_2912,In_1405);
or U694 (N_694,In_2073,In_1887);
xor U695 (N_695,In_1267,In_981);
nor U696 (N_696,In_95,In_1713);
or U697 (N_697,In_451,In_1206);
or U698 (N_698,In_1047,In_896);
nor U699 (N_699,In_616,In_1787);
nand U700 (N_700,In_921,In_2766);
or U701 (N_701,In_1526,In_1417);
nand U702 (N_702,In_999,In_2006);
or U703 (N_703,In_37,In_1597);
and U704 (N_704,In_1737,In_336);
or U705 (N_705,In_2021,In_2164);
nor U706 (N_706,In_2797,In_2997);
and U707 (N_707,In_234,In_2269);
xnor U708 (N_708,In_1336,In_2987);
and U709 (N_709,In_2834,In_1115);
xor U710 (N_710,In_1656,In_384);
and U711 (N_711,In_2881,In_2827);
xnor U712 (N_712,In_74,In_1765);
nand U713 (N_713,In_2926,In_670);
and U714 (N_714,In_1894,In_2275);
nor U715 (N_715,In_1364,In_1402);
xnor U716 (N_716,In_1702,In_378);
xor U717 (N_717,In_1978,In_1935);
nor U718 (N_718,In_2556,In_1726);
or U719 (N_719,In_460,In_1209);
nor U720 (N_720,In_1208,In_123);
xor U721 (N_721,In_31,In_1805);
nand U722 (N_722,In_25,In_2498);
nand U723 (N_723,In_960,In_2974);
or U724 (N_724,In_2125,In_1813);
or U725 (N_725,In_1678,In_1623);
nand U726 (N_726,In_251,In_1611);
nor U727 (N_727,In_2410,In_551);
nor U728 (N_728,In_1539,In_1708);
and U729 (N_729,In_2698,In_2911);
xor U730 (N_730,In_1401,In_747);
xnor U731 (N_731,In_1649,In_2348);
or U732 (N_732,In_1591,In_2473);
nor U733 (N_733,In_1174,In_2851);
and U734 (N_734,In_1339,In_477);
nand U735 (N_735,In_2665,In_2536);
or U736 (N_736,In_900,In_41);
xor U737 (N_737,In_404,In_1361);
xnor U738 (N_738,In_842,In_579);
nand U739 (N_739,In_2475,In_2378);
nand U740 (N_740,In_362,In_1842);
or U741 (N_741,In_1573,In_660);
and U742 (N_742,In_545,In_2030);
or U743 (N_743,In_2593,In_1484);
or U744 (N_744,In_1653,In_936);
nand U745 (N_745,In_2220,In_1494);
nand U746 (N_746,In_678,In_758);
nor U747 (N_747,In_2380,In_2960);
and U748 (N_748,In_745,In_562);
nor U749 (N_749,In_2385,In_2727);
and U750 (N_750,In_762,In_2441);
nor U751 (N_751,In_511,In_2352);
or U752 (N_752,In_142,In_1355);
xor U753 (N_753,In_18,In_311);
xnor U754 (N_754,In_879,In_437);
or U755 (N_755,In_262,In_1589);
nor U756 (N_756,In_2718,In_1282);
nor U757 (N_757,In_377,In_1876);
nor U758 (N_758,In_1247,In_1505);
nand U759 (N_759,In_2087,In_2823);
nor U760 (N_760,In_439,In_1995);
or U761 (N_761,In_1674,In_589);
and U762 (N_762,In_2228,In_1263);
xor U763 (N_763,In_637,In_1243);
nor U764 (N_764,In_73,In_2703);
or U765 (N_765,In_2247,In_241);
nand U766 (N_766,In_2439,In_2646);
xnor U767 (N_767,In_2814,In_679);
or U768 (N_768,In_29,In_2300);
xor U769 (N_769,In_1327,In_179);
nand U770 (N_770,In_1754,In_1107);
and U771 (N_771,In_2999,In_2078);
or U772 (N_772,In_158,In_1742);
nand U773 (N_773,In_1217,In_2724);
or U774 (N_774,In_2637,In_2168);
or U775 (N_775,In_2994,In_2980);
and U776 (N_776,In_768,In_1527);
nand U777 (N_777,In_1034,In_65);
and U778 (N_778,In_2900,In_330);
xnor U779 (N_779,In_1308,In_1384);
nand U780 (N_780,In_2562,In_789);
xor U781 (N_781,In_1091,In_2701);
nor U782 (N_782,In_2261,In_1643);
or U783 (N_783,In_943,In_305);
or U784 (N_784,In_861,In_504);
nor U785 (N_785,In_291,In_2002);
nand U786 (N_786,In_152,In_1255);
or U787 (N_787,In_261,In_2424);
or U788 (N_788,In_1210,In_1435);
and U789 (N_789,In_1786,In_2467);
xor U790 (N_790,In_2546,In_1884);
or U791 (N_791,In_692,In_96);
or U792 (N_792,In_2250,In_1098);
xnor U793 (N_793,In_2754,In_2503);
nand U794 (N_794,In_908,In_1934);
nand U795 (N_795,In_2992,In_2015);
nor U796 (N_796,In_2752,In_1755);
nor U797 (N_797,In_1346,In_1187);
or U798 (N_798,In_1257,In_2450);
nor U799 (N_799,In_363,In_918);
xnor U800 (N_800,In_912,In_1324);
nand U801 (N_801,In_1081,In_824);
nor U802 (N_802,In_1179,In_836);
or U803 (N_803,In_1756,In_1758);
nor U804 (N_804,In_2520,In_2622);
xnor U805 (N_805,In_1537,In_2631);
xnor U806 (N_806,In_811,In_2492);
or U807 (N_807,In_403,In_400);
xor U808 (N_808,In_858,In_634);
nand U809 (N_809,In_2035,In_1719);
or U810 (N_810,In_296,In_744);
xor U811 (N_811,In_976,In_1682);
nor U812 (N_812,In_2978,In_246);
nor U813 (N_813,In_513,In_191);
nor U814 (N_814,In_2098,In_118);
or U815 (N_815,In_2008,In_2511);
or U816 (N_816,In_97,In_1393);
xnor U817 (N_817,In_2525,In_169);
nor U818 (N_818,In_419,In_1489);
and U819 (N_819,In_2740,In_240);
nor U820 (N_820,In_2636,In_2460);
or U821 (N_821,In_777,In_1511);
nand U822 (N_822,In_1278,In_2939);
nor U823 (N_823,In_2418,In_2101);
xor U824 (N_824,In_2523,In_2685);
and U825 (N_825,In_2884,In_923);
nand U826 (N_826,In_1101,In_2531);
or U827 (N_827,In_1244,In_1311);
and U828 (N_828,In_418,In_449);
and U829 (N_829,In_1796,In_306);
or U830 (N_830,In_1118,In_424);
and U831 (N_831,In_955,In_467);
and U832 (N_832,In_852,In_2887);
nor U833 (N_833,In_334,In_2689);
nor U834 (N_834,In_1398,In_316);
xor U835 (N_835,In_2614,In_2389);
or U836 (N_836,In_233,In_773);
xor U837 (N_837,In_1075,In_657);
nor U838 (N_838,In_1806,In_1982);
and U839 (N_839,In_2575,In_514);
nor U840 (N_840,In_1269,In_2516);
or U841 (N_841,In_2003,In_194);
or U842 (N_842,In_1313,In_756);
nor U843 (N_843,In_287,In_216);
nor U844 (N_844,In_2400,In_799);
or U845 (N_845,In_905,In_1577);
xnor U846 (N_846,In_2141,In_1270);
nand U847 (N_847,In_375,In_881);
and U848 (N_848,In_625,In_231);
and U849 (N_849,In_414,In_1297);
xor U850 (N_850,In_2456,In_338);
or U851 (N_851,In_530,In_1144);
or U852 (N_852,In_2218,In_549);
and U853 (N_853,In_166,In_998);
and U854 (N_854,In_2405,In_1555);
nand U855 (N_855,In_1218,In_2634);
nand U856 (N_856,In_760,In_1515);
and U857 (N_857,In_751,In_438);
and U858 (N_858,In_197,In_340);
xor U859 (N_859,In_995,In_472);
and U860 (N_860,In_1976,In_869);
nand U861 (N_861,In_1747,In_2950);
xor U862 (N_862,In_1582,In_1557);
nor U863 (N_863,In_2060,In_151);
or U864 (N_864,In_1188,In_1053);
nor U865 (N_865,In_2179,In_924);
or U866 (N_866,In_2032,In_2661);
or U867 (N_867,In_2249,In_729);
or U868 (N_868,In_753,In_2364);
and U869 (N_869,In_346,In_1727);
or U870 (N_870,In_2557,In_1705);
and U871 (N_871,In_1735,In_211);
or U872 (N_872,In_2391,In_2670);
or U873 (N_873,In_282,In_242);
nand U874 (N_874,In_2426,In_1127);
nand U875 (N_875,In_2746,In_75);
xnor U876 (N_876,In_68,In_277);
nor U877 (N_877,In_2084,In_2169);
nand U878 (N_878,In_1921,In_1419);
nand U879 (N_879,In_992,In_204);
nor U880 (N_880,In_2486,In_2544);
and U881 (N_881,In_2208,In_385);
xnor U882 (N_882,In_1272,In_1474);
or U883 (N_883,In_227,In_2699);
and U884 (N_884,In_2667,In_2716);
nand U885 (N_885,In_677,In_2242);
or U886 (N_886,In_274,In_724);
xnor U887 (N_887,In_2901,In_1897);
nand U888 (N_888,In_2227,In_1035);
or U889 (N_889,In_63,In_415);
nand U890 (N_890,In_2403,In_617);
nand U891 (N_891,In_1227,In_1561);
and U892 (N_892,In_500,In_1538);
and U893 (N_893,In_2349,In_92);
or U894 (N_894,In_2957,In_2356);
nor U895 (N_895,In_1168,In_2096);
xor U896 (N_896,In_1646,In_2142);
nor U897 (N_897,In_721,In_738);
nor U898 (N_898,In_1356,In_1681);
or U899 (N_899,In_1370,In_109);
xnor U900 (N_900,In_1369,In_2581);
or U901 (N_901,In_1960,In_2104);
nand U902 (N_902,In_2165,In_2675);
and U903 (N_903,In_1509,In_1299);
nand U904 (N_904,In_2124,In_2496);
and U905 (N_905,In_288,In_1059);
nor U906 (N_906,In_2329,In_2793);
and U907 (N_907,In_1341,In_1782);
nand U908 (N_908,In_1260,In_1803);
nor U909 (N_909,In_2471,In_2534);
xor U910 (N_910,In_2082,In_2825);
or U911 (N_911,In_1595,In_2755);
and U912 (N_912,In_2013,In_1546);
or U913 (N_913,In_402,In_2294);
nor U914 (N_914,In_606,In_1087);
xor U915 (N_915,In_300,In_2411);
xnor U916 (N_916,In_875,In_135);
nor U917 (N_917,In_1977,In_1999);
nand U918 (N_918,In_1492,In_484);
nor U919 (N_919,In_1570,In_1637);
nor U920 (N_920,In_144,In_1815);
nor U921 (N_921,In_2267,In_2394);
nor U922 (N_922,In_1875,In_2219);
or U923 (N_923,In_1664,In_519);
xnor U924 (N_924,In_67,In_2483);
nand U925 (N_925,In_1383,In_1533);
nor U926 (N_926,In_1471,In_379);
xor U927 (N_927,In_1572,In_691);
and U928 (N_928,In_2252,In_2023);
nand U929 (N_929,In_2489,In_2427);
nand U930 (N_930,In_870,In_1095);
or U931 (N_931,In_591,In_468);
or U932 (N_932,In_1447,In_1588);
or U933 (N_933,In_249,In_717);
or U934 (N_934,In_2803,In_1576);
nor U935 (N_935,In_2199,In_2083);
xor U936 (N_936,In_1696,In_1650);
nand U937 (N_937,In_1347,In_165);
nor U938 (N_938,In_1444,In_779);
nand U939 (N_939,In_408,In_1871);
xor U940 (N_940,In_1707,In_2276);
and U941 (N_941,In_430,In_2382);
nand U942 (N_942,In_1328,In_1583);
xnor U943 (N_943,In_680,In_1617);
or U944 (N_944,In_714,In_1052);
and U945 (N_945,In_1240,In_810);
xnor U946 (N_946,In_1316,In_966);
xnor U947 (N_947,In_2815,In_2728);
and U948 (N_948,In_2393,In_1544);
or U949 (N_949,In_874,In_2386);
nor U950 (N_950,In_372,In_1943);
xnor U951 (N_951,In_761,In_1673);
nor U952 (N_952,In_2620,In_1024);
xnor U953 (N_953,In_2694,In_2952);
xor U954 (N_954,In_1178,In_2195);
xnor U955 (N_955,In_344,In_578);
or U956 (N_956,In_971,In_1825);
or U957 (N_957,In_102,In_1620);
or U958 (N_958,In_322,In_221);
nor U959 (N_959,In_1989,In_2414);
xnor U960 (N_960,In_699,In_1924);
nor U961 (N_961,In_1266,In_2929);
nand U962 (N_962,In_575,In_189);
or U963 (N_963,In_2051,In_2577);
and U964 (N_964,In_2855,In_280);
nand U965 (N_965,In_687,In_2038);
and U966 (N_966,In_1332,In_1006);
xnor U967 (N_967,In_2910,In_1838);
and U968 (N_968,In_2652,In_253);
or U969 (N_969,In_1445,In_1814);
nor U970 (N_970,In_661,In_1409);
or U971 (N_971,In_2736,In_131);
nor U972 (N_972,In_696,In_2945);
or U973 (N_973,In_2956,In_1965);
nand U974 (N_974,In_2776,In_780);
and U975 (N_975,In_281,In_1975);
or U976 (N_976,In_2610,In_2351);
xor U977 (N_977,In_775,In_2091);
xnor U978 (N_978,In_538,In_1528);
and U979 (N_979,In_493,In_1054);
xnor U980 (N_980,In_2629,In_56);
nand U981 (N_981,In_2898,In_1832);
nand U982 (N_982,In_2077,In_2664);
or U983 (N_983,In_957,In_1880);
xor U984 (N_984,In_1731,In_2334);
nor U985 (N_985,In_1913,In_2966);
or U986 (N_986,In_2805,In_145);
nand U987 (N_987,In_2883,In_737);
xor U988 (N_988,In_1598,In_2604);
nor U989 (N_989,In_1203,In_1211);
nand U990 (N_990,In_2186,In_1733);
nand U991 (N_991,In_1495,In_2066);
xor U992 (N_992,In_254,In_808);
nand U993 (N_993,In_2132,In_2309);
or U994 (N_994,In_947,In_1685);
nor U995 (N_995,In_42,In_1418);
nor U996 (N_996,In_1152,In_1873);
nand U997 (N_997,In_1231,In_2609);
xor U998 (N_998,In_2476,In_1568);
xor U999 (N_999,In_1791,In_2638);
or U1000 (N_1000,In_2036,In_1956);
xor U1001 (N_1001,In_170,In_1020);
nand U1002 (N_1002,In_386,In_2444);
nand U1003 (N_1003,In_1951,In_1794);
nand U1004 (N_1004,In_2325,In_570);
or U1005 (N_1005,In_1862,In_2000);
or U1006 (N_1006,In_1376,In_2434);
nand U1007 (N_1007,In_433,In_476);
or U1008 (N_1008,In_2,In_2286);
and U1009 (N_1009,In_1442,In_1952);
and U1010 (N_1010,In_1565,In_2975);
xor U1011 (N_1011,In_2037,In_868);
nand U1012 (N_1012,In_2969,In_1866);
or U1013 (N_1013,In_1919,In_237);
or U1014 (N_1014,In_1729,In_2243);
and U1015 (N_1015,In_2103,In_2278);
or U1016 (N_1016,In_1242,In_2026);
or U1017 (N_1017,In_273,In_264);
nand U1018 (N_1018,In_2154,In_856);
or U1019 (N_1019,In_48,In_159);
and U1020 (N_1020,In_730,In_215);
nor U1021 (N_1021,In_1886,In_1241);
xor U1022 (N_1022,In_2105,In_1703);
nor U1023 (N_1023,In_1411,In_764);
or U1024 (N_1024,In_1180,In_822);
or U1025 (N_1025,In_2690,In_2871);
xor U1026 (N_1026,In_2137,In_1281);
and U1027 (N_1027,In_1874,In_2979);
xnor U1028 (N_1028,In_1386,In_2173);
nor U1029 (N_1029,In_2700,In_1129);
nand U1030 (N_1030,In_534,In_1750);
or U1031 (N_1031,In_1497,In_801);
nand U1032 (N_1032,In_2768,In_2328);
or U1033 (N_1033,In_2280,In_1321);
nand U1034 (N_1034,In_1795,In_2712);
or U1035 (N_1035,In_1609,In_2616);
nand U1036 (N_1036,In_2947,In_1292);
nand U1037 (N_1037,In_740,In_1531);
or U1038 (N_1038,In_1008,In_8);
nand U1039 (N_1039,In_481,In_620);
and U1040 (N_1040,In_1134,In_2397);
nand U1041 (N_1041,In_1987,In_2233);
or U1042 (N_1042,In_238,In_2075);
and U1043 (N_1043,In_1108,In_2490);
nand U1044 (N_1044,In_1158,In_1318);
nand U1045 (N_1045,In_1425,In_792);
and U1046 (N_1046,In_1870,In_1778);
xnor U1047 (N_1047,In_2319,In_2608);
and U1048 (N_1048,In_1377,In_2071);
nand U1049 (N_1049,In_47,In_2442);
nor U1050 (N_1050,In_2074,In_2839);
nor U1051 (N_1051,In_2893,In_470);
nand U1052 (N_1052,In_1066,In_24);
and U1053 (N_1053,In_301,In_2765);
or U1054 (N_1054,In_1730,In_2566);
and U1055 (N_1055,In_1622,In_910);
nor U1056 (N_1056,In_1940,In_2571);
nand U1057 (N_1057,In_2388,In_1847);
xor U1058 (N_1058,In_531,In_547);
and U1059 (N_1059,In_1323,In_2965);
nor U1060 (N_1060,In_2421,In_127);
nand U1061 (N_1061,In_2379,In_350);
or U1062 (N_1062,In_2463,In_2292);
nor U1063 (N_1063,In_2745,In_107);
nand U1064 (N_1064,In_187,In_720);
or U1065 (N_1065,In_5,In_1362);
nand U1066 (N_1066,In_1927,In_2905);
nand U1067 (N_1067,In_1783,In_324);
or U1068 (N_1068,In_517,In_2431);
xnor U1069 (N_1069,In_1519,In_224);
xor U1070 (N_1070,In_643,In_2465);
or U1071 (N_1071,In_359,In_121);
and U1072 (N_1072,In_1221,In_1957);
nor U1073 (N_1073,In_1378,In_1636);
and U1074 (N_1074,In_509,In_2915);
or U1075 (N_1075,In_2872,In_1819);
nor U1076 (N_1076,In_1967,In_1416);
nand U1077 (N_1077,In_1970,In_1801);
nand U1078 (N_1078,In_2784,In_1389);
nor U1079 (N_1079,In_456,In_1672);
nor U1080 (N_1080,In_2491,In_393);
or U1081 (N_1081,In_1400,In_1898);
and U1082 (N_1082,In_805,In_725);
or U1083 (N_1083,In_946,In_1482);
xor U1084 (N_1084,In_2553,In_2713);
or U1085 (N_1085,In_2972,In_425);
xnor U1086 (N_1086,In_2600,In_1025);
nand U1087 (N_1087,In_2730,In_706);
nand U1088 (N_1088,In_2789,In_1619);
and U1089 (N_1089,In_2326,In_105);
or U1090 (N_1090,In_800,In_1781);
or U1091 (N_1091,In_2796,In_2626);
and U1092 (N_1092,In_732,In_772);
xnor U1093 (N_1093,In_2964,In_1686);
or U1094 (N_1094,In_537,In_2506);
xor U1095 (N_1095,In_949,In_1290);
or U1096 (N_1096,In_2106,In_1060);
nand U1097 (N_1097,In_1177,In_1676);
nor U1098 (N_1098,In_1586,In_1300);
xnor U1099 (N_1099,In_2817,In_1371);
or U1100 (N_1100,In_1594,In_184);
and U1101 (N_1101,In_1017,In_885);
or U1102 (N_1102,In_1695,In_1858);
nand U1103 (N_1103,In_608,In_392);
or U1104 (N_1104,In_734,In_2022);
nor U1105 (N_1105,In_2438,In_2808);
or U1106 (N_1106,In_1380,In_1601);
and U1107 (N_1107,In_93,In_2088);
nor U1108 (N_1108,In_1616,In_2653);
xnor U1109 (N_1109,In_1745,In_1510);
nand U1110 (N_1110,In_1845,In_731);
or U1111 (N_1111,In_645,In_571);
or U1112 (N_1112,In_2708,In_1368);
or U1113 (N_1113,In_1112,In_474);
nor U1114 (N_1114,In_763,In_235);
and U1115 (N_1115,In_265,In_1466);
and U1116 (N_1116,In_2889,In_471);
nor U1117 (N_1117,In_1645,In_1481);
nor U1118 (N_1118,In_1603,In_2396);
xor U1119 (N_1119,In_1156,In_2143);
xnor U1120 (N_1120,In_2709,In_461);
nand U1121 (N_1121,In_2518,In_2310);
nor U1122 (N_1122,In_1734,In_612);
or U1123 (N_1123,In_1164,In_1245);
xnor U1124 (N_1124,In_1145,In_515);
nor U1125 (N_1125,In_99,In_682);
xnor U1126 (N_1126,In_2846,In_1331);
xor U1127 (N_1127,In_2863,In_953);
or U1128 (N_1128,In_1766,In_17);
nand U1129 (N_1129,In_1693,In_1941);
nand U1130 (N_1130,In_2007,In_2093);
and U1131 (N_1131,In_223,In_2184);
nor U1132 (N_1132,In_1480,In_2645);
nor U1133 (N_1133,In_2241,In_2122);
nand U1134 (N_1134,In_2853,In_1000);
xor U1135 (N_1135,In_1092,In_2366);
nor U1136 (N_1136,In_1475,In_788);
and U1137 (N_1137,In_399,In_2205);
or U1138 (N_1138,In_401,In_1026);
or U1139 (N_1139,In_1800,In_642);
nand U1140 (N_1140,In_2274,In_1878);
nand U1141 (N_1141,In_726,In_2009);
nand U1142 (N_1142,In_554,In_1954);
xnor U1143 (N_1143,In_119,In_2481);
xor U1144 (N_1144,In_1354,In_1958);
xnor U1145 (N_1145,In_1089,In_171);
nand U1146 (N_1146,In_2513,In_2462);
xnor U1147 (N_1147,In_2487,In_2764);
nand U1148 (N_1148,In_2602,In_986);
and U1149 (N_1149,In_711,In_1749);
nor U1150 (N_1150,In_709,In_2526);
and U1151 (N_1151,In_561,In_40);
or U1152 (N_1152,In_2854,In_126);
nand U1153 (N_1153,In_1280,In_2027);
and U1154 (N_1154,In_2691,In_1259);
xnor U1155 (N_1155,In_1529,In_1440);
nand U1156 (N_1156,In_1613,In_2821);
and U1157 (N_1157,In_932,In_2399);
xor U1158 (N_1158,In_2517,In_1309);
xor U1159 (N_1159,In_2617,In_162);
and U1160 (N_1160,In_2659,In_618);
nor U1161 (N_1161,In_2162,In_214);
or U1162 (N_1162,In_1579,In_1438);
or U1163 (N_1163,In_2693,In_2214);
or U1164 (N_1164,In_565,In_1917);
nor U1165 (N_1165,In_964,In_2413);
xnor U1166 (N_1166,In_1759,In_2933);
or U1167 (N_1167,In_1608,In_1150);
xor U1168 (N_1168,In_2882,In_2390);
xor U1169 (N_1169,In_1358,In_2474);
nor U1170 (N_1170,In_101,In_390);
nor U1171 (N_1171,In_205,In_2108);
xnor U1172 (N_1172,In_52,In_1642);
xor U1173 (N_1173,In_2161,In_1699);
nor U1174 (N_1174,In_243,In_226);
nand U1175 (N_1175,In_1468,In_2447);
or U1176 (N_1176,In_2433,In_1985);
and U1177 (N_1177,In_1493,In_2930);
xnor U1178 (N_1178,In_1161,In_1137);
nand U1179 (N_1179,In_2850,In_2548);
or U1180 (N_1180,In_83,In_2215);
or U1181 (N_1181,In_345,In_2493);
and U1182 (N_1182,In_2289,In_149);
and U1183 (N_1183,In_688,In_1833);
nor U1184 (N_1184,In_843,In_2435);
xnor U1185 (N_1185,In_1251,In_1843);
nor U1186 (N_1186,In_2826,In_1109);
nand U1187 (N_1187,In_1202,In_1852);
nor U1188 (N_1188,In_1543,In_2695);
nor U1189 (N_1189,In_2744,In_2623);
xnor U1190 (N_1190,In_2138,In_727);
xor U1191 (N_1191,In_766,In_2381);
and U1192 (N_1192,In_871,In_2550);
and U1193 (N_1193,In_1668,In_1992);
nor U1194 (N_1194,In_2529,In_2046);
and U1195 (N_1195,In_230,In_174);
xor U1196 (N_1196,In_712,In_488);
and U1197 (N_1197,In_1116,In_1700);
nand U1198 (N_1198,In_1262,In_934);
xnor U1199 (N_1199,In_222,In_2925);
nand U1200 (N_1200,In_1410,In_122);
nor U1201 (N_1201,In_592,In_1627);
nand U1202 (N_1202,In_185,In_2936);
xnor U1203 (N_1203,In_2271,In_577);
xnor U1204 (N_1204,In_1373,In_1013);
and U1205 (N_1205,In_1102,In_917);
nor U1206 (N_1206,In_104,In_1285);
nand U1207 (N_1207,In_496,In_2293);
xnor U1208 (N_1208,In_1068,In_2062);
nor U1209 (N_1209,In_2012,In_2567);
and U1210 (N_1210,In_2357,In_1817);
nand U1211 (N_1211,In_2232,In_1141);
nand U1212 (N_1212,In_1746,In_1302);
and U1213 (N_1213,In_2224,In_2398);
or U1214 (N_1214,In_2720,In_164);
nor U1215 (N_1215,In_479,In_809);
and U1216 (N_1216,In_353,In_2779);
and U1217 (N_1217,In_2530,In_1860);
nor U1218 (N_1218,In_16,In_2832);
or U1219 (N_1219,In_671,In_2204);
nand U1220 (N_1220,In_817,In_2782);
nor U1221 (N_1221,In_2011,In_1560);
or U1222 (N_1222,In_626,In_217);
or U1223 (N_1223,In_98,In_2056);
xor U1224 (N_1224,In_2524,In_1679);
nor U1225 (N_1225,In_1437,In_1048);
nand U1226 (N_1226,In_700,In_1439);
and U1227 (N_1227,In_1388,In_2191);
nand U1228 (N_1228,In_629,In_302);
and U1229 (N_1229,In_2539,In_2588);
and U1230 (N_1230,In_2981,In_19);
or U1231 (N_1231,In_2230,In_2757);
nand U1232 (N_1232,In_526,In_1725);
xnor U1233 (N_1233,In_2747,In_298);
or U1234 (N_1234,In_443,In_2877);
or U1235 (N_1235,In_904,In_975);
and U1236 (N_1236,In_1704,In_1228);
xor U1237 (N_1237,In_34,In_838);
or U1238 (N_1238,In_201,In_2656);
or U1239 (N_1239,In_2320,In_646);
nand U1240 (N_1240,In_2158,In_1100);
nand U1241 (N_1241,In_106,In_1525);
nor U1242 (N_1242,In_1085,In_1915);
nand U1243 (N_1243,In_1235,In_2055);
or U1244 (N_1244,In_658,In_2554);
nor U1245 (N_1245,In_382,In_2606);
or U1246 (N_1246,In_694,In_2918);
nand U1247 (N_1247,In_422,In_80);
nor U1248 (N_1248,In_1159,In_2288);
xor U1249 (N_1249,In_1070,In_1216);
or U1250 (N_1250,In_268,In_1732);
nand U1251 (N_1251,In_2446,In_1621);
nor U1252 (N_1252,In_2774,In_1067);
xor U1253 (N_1253,In_1518,In_635);
nor U1254 (N_1254,In_746,In_1192);
nand U1255 (N_1255,In_70,In_2573);
nor U1256 (N_1256,In_1042,In_2897);
xnor U1257 (N_1257,In_774,In_614);
and U1258 (N_1258,In_518,In_945);
xnor U1259 (N_1259,In_2615,In_1942);
and U1260 (N_1260,In_527,In_279);
nand U1261 (N_1261,In_2880,In_607);
and U1262 (N_1262,In_505,In_2601);
nand U1263 (N_1263,In_2240,In_889);
or U1264 (N_1264,In_2791,In_335);
xor U1265 (N_1265,In_2563,In_1752);
xor U1266 (N_1266,In_1689,In_1182);
and U1267 (N_1267,In_2688,In_1901);
nand U1268 (N_1268,In_1375,In_2833);
xnor U1269 (N_1269,In_2285,In_593);
nand U1270 (N_1270,In_2092,In_820);
nand U1271 (N_1271,In_2916,In_1826);
and U1272 (N_1272,In_2958,In_2063);
nor U1273 (N_1273,In_1018,In_2182);
xnor U1274 (N_1274,In_1226,In_1652);
and U1275 (N_1275,In_867,In_1215);
nand U1276 (N_1276,In_1925,In_2873);
and U1277 (N_1277,In_1657,In_619);
nor U1278 (N_1278,In_2862,In_1706);
and U1279 (N_1279,In_1513,In_1888);
nand U1280 (N_1280,In_752,In_1148);
xnor U1281 (N_1281,In_980,In_782);
xor U1282 (N_1282,In_181,In_2160);
nand U1283 (N_1283,In_2813,In_2822);
nand U1284 (N_1284,In_785,In_2253);
and U1285 (N_1285,In_605,In_2287);
nor U1286 (N_1286,In_823,In_2521);
nand U1287 (N_1287,In_940,In_11);
xnor U1288 (N_1288,In_2365,In_2312);
xor U1289 (N_1289,In_681,In_705);
nor U1290 (N_1290,In_2642,In_361);
nand U1291 (N_1291,In_2350,In_1545);
xnor U1292 (N_1292,In_1944,In_1665);
nor U1293 (N_1293,In_2923,In_54);
and U1294 (N_1294,In_2354,In_57);
and U1295 (N_1295,In_2097,In_420);
xnor U1296 (N_1296,In_1071,In_1077);
or U1297 (N_1297,In_2229,In_1113);
and U1298 (N_1298,In_2110,In_62);
xnor U1299 (N_1299,In_807,In_1348);
xor U1300 (N_1300,In_2909,In_930);
and U1301 (N_1301,In_1728,In_2532);
or U1302 (N_1302,In_66,In_2955);
nor U1303 (N_1303,In_2226,In_2515);
or U1304 (N_1304,In_1423,In_1345);
nor U1305 (N_1305,In_2672,In_2867);
xnor U1306 (N_1306,In_864,In_582);
nor U1307 (N_1307,In_698,In_787);
nand U1308 (N_1308,In_2628,In_2878);
nand U1309 (N_1309,In_2982,In_2885);
or U1310 (N_1310,In_1201,In_1351);
nor U1311 (N_1311,In_1093,In_2504);
xnor U1312 (N_1312,In_1128,In_2886);
xnor U1313 (N_1313,In_1640,In_196);
nor U1314 (N_1314,In_494,In_2648);
or U1315 (N_1315,In_2663,In_1830);
or U1316 (N_1316,In_962,In_271);
nand U1317 (N_1317,In_1651,In_405);
or U1318 (N_1318,In_103,In_427);
nor U1319 (N_1319,In_2836,In_996);
or U1320 (N_1320,In_1625,In_952);
or U1321 (N_1321,In_140,In_2845);
xor U1322 (N_1322,In_1895,In_2034);
nor U1323 (N_1323,In_1581,In_522);
and U1324 (N_1324,In_206,In_2738);
or U1325 (N_1325,In_1736,In_602);
nand U1326 (N_1326,In_1540,In_1973);
and U1327 (N_1327,In_1811,In_2753);
nor U1328 (N_1328,In_128,In_523);
nor U1329 (N_1329,In_686,In_985);
xor U1330 (N_1330,In_1810,In_7);
or U1331 (N_1331,In_603,In_2102);
or U1332 (N_1332,In_1559,In_994);
xnor U1333 (N_1333,In_1183,In_2126);
xor U1334 (N_1334,In_2711,In_2019);
or U1335 (N_1335,In_1694,In_1829);
nand U1336 (N_1336,In_10,In_487);
nand U1337 (N_1337,In_1631,In_2678);
nand U1338 (N_1338,In_1427,In_1103);
and U1339 (N_1339,In_2643,In_1151);
nor U1340 (N_1340,In_2914,In_1721);
or U1341 (N_1341,In_272,In_209);
nand U1342 (N_1342,In_2505,In_653);
or U1343 (N_1343,In_1155,In_1125);
and U1344 (N_1344,In_1760,In_2331);
xor U1345 (N_1345,In_1793,In_1675);
or U1346 (N_1346,In_2039,In_2555);
or U1347 (N_1347,In_14,In_1896);
nand U1348 (N_1348,In_623,In_1012);
nand U1349 (N_1349,In_2193,In_563);
nor U1350 (N_1350,In_797,In_1923);
xnor U1351 (N_1351,In_2924,In_1764);
xnor U1352 (N_1352,In_94,In_1930);
nand U1353 (N_1353,In_2673,In_2114);
or U1354 (N_1354,In_406,In_967);
and U1355 (N_1355,In_535,In_284);
nand U1356 (N_1356,In_495,In_192);
and U1357 (N_1357,In_2302,In_1751);
nor U1358 (N_1358,In_533,In_2669);
or U1359 (N_1359,In_100,In_228);
nand U1360 (N_1360,In_1436,In_1922);
xor U1361 (N_1361,In_283,In_2876);
xnor U1362 (N_1362,In_1761,In_739);
nand U1363 (N_1363,In_835,In_857);
xnor U1364 (N_1364,In_2590,In_2457);
and U1365 (N_1365,In_333,In_2152);
xnor U1366 (N_1366,In_2904,In_276);
and U1367 (N_1367,In_644,In_507);
nor U1368 (N_1368,In_2045,In_2856);
nor U1369 (N_1369,In_1253,In_38);
nor U1370 (N_1370,In_651,In_597);
nor U1371 (N_1371,In_435,In_713);
or U1372 (N_1372,In_2919,In_2818);
and U1373 (N_1373,In_1320,In_2281);
nor U1374 (N_1374,In_2681,In_1078);
or U1375 (N_1375,In_12,In_2321);
nand U1376 (N_1376,In_2641,In_2417);
xnor U1377 (N_1377,In_759,In_2189);
xor U1378 (N_1378,In_2099,In_2512);
xor U1379 (N_1379,In_2086,In_1792);
xor U1380 (N_1380,In_1097,In_2892);
nor U1381 (N_1381,In_2777,In_599);
xor U1382 (N_1382,In_2552,In_293);
nor U1383 (N_1383,In_2127,In_247);
or U1384 (N_1384,In_640,In_2549);
and U1385 (N_1385,In_988,In_2145);
nor U1386 (N_1386,In_1683,In_2899);
and U1387 (N_1387,In_307,In_872);
or U1388 (N_1388,In_2683,In_2248);
or U1389 (N_1389,In_2844,In_1051);
xor U1390 (N_1390,In_1662,In_1867);
nand U1391 (N_1391,In_2820,In_13);
nor U1392 (N_1392,In_45,In_572);
xnor U1393 (N_1393,In_621,In_568);
nor U1394 (N_1394,In_1334,In_2857);
nor U1395 (N_1395,In_155,In_1716);
nand U1396 (N_1396,In_341,In_1340);
or U1397 (N_1397,In_1239,In_2940);
or U1398 (N_1398,In_2917,In_1906);
nand U1399 (N_1399,In_110,In_1587);
and U1400 (N_1400,In_837,In_2047);
and U1401 (N_1401,In_2829,In_1246);
and U1402 (N_1402,In_841,In_61);
nand U1403 (N_1403,In_50,In_1658);
xnor U1404 (N_1404,In_862,In_848);
nor U1405 (N_1405,In_278,In_84);
or U1406 (N_1406,In_1820,In_1872);
and U1407 (N_1407,In_2221,In_416);
or U1408 (N_1408,In_1905,In_387);
nand U1409 (N_1409,In_1720,In_2153);
and U1410 (N_1410,In_1413,In_188);
and U1411 (N_1411,In_1434,In_1911);
or U1412 (N_1412,In_2961,In_754);
nand U1413 (N_1413,In_2468,In_46);
xnor U1414 (N_1414,In_833,In_652);
or U1415 (N_1415,In_1610,In_741);
or U1416 (N_1416,In_2194,In_2660);
or U1417 (N_1417,In_2848,In_604);
xnor U1418 (N_1418,In_922,In_1912);
nand U1419 (N_1419,In_1408,In_1248);
and U1420 (N_1420,In_3,In_2519);
and U1421 (N_1421,In_312,In_2371);
or U1422 (N_1422,In_143,In_2896);
nor U1423 (N_1423,In_690,In_2806);
and U1424 (N_1424,In_263,In_167);
xnor U1425 (N_1425,In_977,In_447);
or U1426 (N_1426,In_2377,In_203);
and U1427 (N_1427,In_757,In_2495);
xnor U1428 (N_1428,In_486,In_2605);
and U1429 (N_1429,In_1937,In_648);
xnor U1430 (N_1430,In_2868,In_812);
nand U1431 (N_1431,In_847,In_2297);
nor U1432 (N_1432,In_429,In_613);
nand U1433 (N_1433,In_176,In_2858);
xor U1434 (N_1434,In_1147,In_1780);
nand U1435 (N_1435,In_1224,In_902);
nand U1436 (N_1436,In_2246,In_1415);
xnor U1437 (N_1437,In_2625,In_448);
and U1438 (N_1438,In_2760,In_53);
nand U1439 (N_1439,In_2984,In_2308);
nor U1440 (N_1440,In_2572,In_1953);
and U1441 (N_1441,In_873,In_1835);
and U1442 (N_1442,In_979,In_1229);
or U1443 (N_1443,In_59,In_1153);
nand U1444 (N_1444,In_2432,In_1807);
and U1445 (N_1445,In_2245,In_349);
nor U1446 (N_1446,In_1980,In_1167);
nor U1447 (N_1447,In_2251,In_2001);
or U1448 (N_1448,In_1457,In_388);
or U1449 (N_1449,In_1029,In_1496);
xor U1450 (N_1450,In_2112,In_1037);
nand U1451 (N_1451,In_1926,In_2580);
xnor U1452 (N_1452,In_2254,In_1580);
or U1453 (N_1453,In_116,In_1055);
nor U1454 (N_1454,In_2937,In_1892);
xnor U1455 (N_1455,In_1840,In_1357);
nor U1456 (N_1456,In_1660,In_1991);
and U1457 (N_1457,In_2223,In_1011);
nor U1458 (N_1458,In_1404,In_2843);
or U1459 (N_1459,In_1441,In_1945);
nor U1460 (N_1460,In_2583,In_1933);
and U1461 (N_1461,In_2335,In_2149);
and U1462 (N_1462,In_2790,In_2206);
nor U1463 (N_1463,In_168,In_1094);
xnor U1464 (N_1464,In_310,In_2842);
and U1465 (N_1465,In_2866,In_2147);
or U1466 (N_1466,In_1171,In_491);
nor U1467 (N_1467,In_1452,In_2533);
nand U1468 (N_1468,In_331,In_352);
and U1469 (N_1469,In_933,In_2902);
and U1470 (N_1470,In_1816,In_1185);
and U1471 (N_1471,In_890,In_1986);
nor U1472 (N_1472,In_1195,In_1882);
or U1473 (N_1473,In_259,In_1836);
or U1474 (N_1474,In_2203,In_878);
or U1475 (N_1475,In_2551,In_891);
nor U1476 (N_1476,In_2196,In_1607);
and U1477 (N_1477,In_1879,In_1058);
xnor U1478 (N_1478,In_2569,In_1712);
or U1479 (N_1479,In_2578,In_1455);
xor U1480 (N_1480,In_1891,In_1984);
nand U1481 (N_1481,In_911,In_473);
and U1482 (N_1482,In_2658,In_1143);
nand U1483 (N_1483,In_2812,In_2748);
or U1484 (N_1484,In_2358,In_2117);
nand U1485 (N_1485,In_2704,In_36);
xnor U1486 (N_1486,In_297,In_2375);
or U1487 (N_1487,In_503,In_2710);
nand U1488 (N_1488,In_2119,In_2188);
and U1489 (N_1489,In_540,In_1131);
or U1490 (N_1490,In_1190,In_2596);
nand U1491 (N_1491,In_200,In_2756);
xor U1492 (N_1492,In_2922,In_76);
and U1493 (N_1493,In_1553,In_2040);
xor U1494 (N_1494,In_270,In_2343);
nand U1495 (N_1495,In_2236,In_1626);
xnor U1496 (N_1496,In_1677,In_2894);
xnor U1497 (N_1497,In_2962,In_1500);
nor U1498 (N_1498,In_442,In_314);
xnor U1499 (N_1499,In_2891,In_909);
nand U1500 (N_1500,In_1688,In_895);
and U1501 (N_1501,In_2986,In_1585);
xnor U1502 (N_1502,In_2126,In_1254);
xnor U1503 (N_1503,In_995,In_157);
nand U1504 (N_1504,In_2050,In_1488);
nand U1505 (N_1505,In_330,In_2984);
nand U1506 (N_1506,In_2461,In_2230);
nand U1507 (N_1507,In_1073,In_1618);
nand U1508 (N_1508,In_1534,In_2000);
xnor U1509 (N_1509,In_1293,In_419);
and U1510 (N_1510,In_993,In_1333);
and U1511 (N_1511,In_2808,In_1550);
or U1512 (N_1512,In_411,In_354);
or U1513 (N_1513,In_2596,In_1979);
nand U1514 (N_1514,In_1165,In_932);
and U1515 (N_1515,In_608,In_1686);
and U1516 (N_1516,In_1832,In_519);
xor U1517 (N_1517,In_568,In_691);
nor U1518 (N_1518,In_715,In_2475);
xnor U1519 (N_1519,In_2903,In_84);
xnor U1520 (N_1520,In_1767,In_2103);
nor U1521 (N_1521,In_1483,In_1614);
nor U1522 (N_1522,In_1014,In_562);
xor U1523 (N_1523,In_1413,In_2740);
or U1524 (N_1524,In_506,In_502);
and U1525 (N_1525,In_968,In_2283);
nor U1526 (N_1526,In_2586,In_1662);
xor U1527 (N_1527,In_2356,In_446);
or U1528 (N_1528,In_1370,In_126);
xnor U1529 (N_1529,In_2265,In_1757);
xnor U1530 (N_1530,In_1436,In_218);
nor U1531 (N_1531,In_2417,In_2978);
nor U1532 (N_1532,In_339,In_336);
and U1533 (N_1533,In_1717,In_2846);
and U1534 (N_1534,In_2812,In_784);
nor U1535 (N_1535,In_1781,In_428);
nand U1536 (N_1536,In_462,In_1837);
xor U1537 (N_1537,In_2417,In_531);
and U1538 (N_1538,In_2742,In_471);
nand U1539 (N_1539,In_1921,In_1711);
nor U1540 (N_1540,In_614,In_848);
or U1541 (N_1541,In_1318,In_1984);
nand U1542 (N_1542,In_2000,In_1252);
and U1543 (N_1543,In_2133,In_1502);
nand U1544 (N_1544,In_398,In_1545);
or U1545 (N_1545,In_476,In_2426);
xor U1546 (N_1546,In_2574,In_2016);
nor U1547 (N_1547,In_1135,In_1195);
or U1548 (N_1548,In_173,In_2896);
nor U1549 (N_1549,In_1265,In_1918);
or U1550 (N_1550,In_2167,In_1000);
xor U1551 (N_1551,In_855,In_1100);
and U1552 (N_1552,In_2891,In_2703);
nor U1553 (N_1553,In_509,In_293);
xor U1554 (N_1554,In_1271,In_15);
nor U1555 (N_1555,In_2690,In_299);
and U1556 (N_1556,In_2995,In_2485);
and U1557 (N_1557,In_2474,In_536);
or U1558 (N_1558,In_768,In_1387);
or U1559 (N_1559,In_1081,In_1391);
nor U1560 (N_1560,In_738,In_2267);
nand U1561 (N_1561,In_2780,In_935);
nand U1562 (N_1562,In_2399,In_445);
nand U1563 (N_1563,In_1047,In_427);
xor U1564 (N_1564,In_1057,In_1663);
nor U1565 (N_1565,In_1940,In_317);
nor U1566 (N_1566,In_2201,In_2755);
xnor U1567 (N_1567,In_1290,In_1678);
xnor U1568 (N_1568,In_2348,In_721);
and U1569 (N_1569,In_2029,In_529);
nand U1570 (N_1570,In_383,In_729);
or U1571 (N_1571,In_2581,In_2841);
xor U1572 (N_1572,In_2416,In_2804);
xor U1573 (N_1573,In_20,In_1748);
nor U1574 (N_1574,In_911,In_1173);
and U1575 (N_1575,In_2152,In_2015);
or U1576 (N_1576,In_2695,In_1512);
nand U1577 (N_1577,In_1581,In_1918);
xor U1578 (N_1578,In_1966,In_2820);
nand U1579 (N_1579,In_2641,In_1891);
nor U1580 (N_1580,In_352,In_2065);
or U1581 (N_1581,In_2120,In_2341);
nor U1582 (N_1582,In_2514,In_2211);
xor U1583 (N_1583,In_1519,In_1727);
nor U1584 (N_1584,In_752,In_2127);
xor U1585 (N_1585,In_1578,In_2958);
xnor U1586 (N_1586,In_1276,In_1928);
nand U1587 (N_1587,In_1304,In_2564);
nand U1588 (N_1588,In_2432,In_1344);
and U1589 (N_1589,In_2482,In_918);
nand U1590 (N_1590,In_254,In_10);
xor U1591 (N_1591,In_859,In_531);
and U1592 (N_1592,In_2806,In_2687);
or U1593 (N_1593,In_1682,In_521);
nor U1594 (N_1594,In_501,In_1021);
or U1595 (N_1595,In_1067,In_2050);
nand U1596 (N_1596,In_2072,In_534);
or U1597 (N_1597,In_2105,In_748);
nand U1598 (N_1598,In_396,In_1075);
and U1599 (N_1599,In_2117,In_185);
or U1600 (N_1600,In_2463,In_2889);
xor U1601 (N_1601,In_1479,In_2441);
nand U1602 (N_1602,In_1025,In_2877);
nand U1603 (N_1603,In_2096,In_2451);
nor U1604 (N_1604,In_1764,In_2868);
or U1605 (N_1605,In_2725,In_1736);
nand U1606 (N_1606,In_1850,In_2996);
and U1607 (N_1607,In_1208,In_31);
nor U1608 (N_1608,In_2001,In_775);
nand U1609 (N_1609,In_1207,In_880);
nor U1610 (N_1610,In_1338,In_2688);
or U1611 (N_1611,In_1756,In_1556);
xnor U1612 (N_1612,In_1793,In_1052);
nor U1613 (N_1613,In_336,In_1907);
and U1614 (N_1614,In_2634,In_2277);
or U1615 (N_1615,In_428,In_946);
xor U1616 (N_1616,In_2935,In_1204);
xnor U1617 (N_1617,In_890,In_2167);
xor U1618 (N_1618,In_2826,In_2621);
nand U1619 (N_1619,In_1058,In_2913);
nor U1620 (N_1620,In_2673,In_1857);
nand U1621 (N_1621,In_2372,In_242);
xor U1622 (N_1622,In_2873,In_2670);
xor U1623 (N_1623,In_1530,In_1302);
nand U1624 (N_1624,In_1567,In_1400);
nor U1625 (N_1625,In_949,In_2716);
or U1626 (N_1626,In_2118,In_2760);
or U1627 (N_1627,In_1220,In_1096);
nor U1628 (N_1628,In_909,In_379);
and U1629 (N_1629,In_2260,In_2451);
nor U1630 (N_1630,In_2329,In_501);
or U1631 (N_1631,In_929,In_2565);
nor U1632 (N_1632,In_317,In_2727);
and U1633 (N_1633,In_2428,In_849);
or U1634 (N_1634,In_232,In_39);
and U1635 (N_1635,In_2301,In_1519);
and U1636 (N_1636,In_840,In_910);
nor U1637 (N_1637,In_231,In_1585);
or U1638 (N_1638,In_1442,In_2593);
and U1639 (N_1639,In_519,In_148);
or U1640 (N_1640,In_702,In_1911);
nand U1641 (N_1641,In_537,In_1094);
nor U1642 (N_1642,In_2101,In_2572);
nand U1643 (N_1643,In_1765,In_2381);
nor U1644 (N_1644,In_2784,In_1418);
xor U1645 (N_1645,In_1349,In_1217);
and U1646 (N_1646,In_2946,In_634);
nand U1647 (N_1647,In_1845,In_2071);
xnor U1648 (N_1648,In_2629,In_177);
or U1649 (N_1649,In_2217,In_102);
or U1650 (N_1650,In_472,In_2839);
nor U1651 (N_1651,In_2276,In_2773);
nand U1652 (N_1652,In_1686,In_536);
nor U1653 (N_1653,In_2740,In_2651);
or U1654 (N_1654,In_1117,In_1136);
xor U1655 (N_1655,In_1715,In_551);
and U1656 (N_1656,In_1221,In_2550);
nor U1657 (N_1657,In_1511,In_2929);
and U1658 (N_1658,In_2043,In_1187);
nand U1659 (N_1659,In_877,In_1398);
nand U1660 (N_1660,In_741,In_1489);
or U1661 (N_1661,In_1494,In_811);
xnor U1662 (N_1662,In_1166,In_1667);
or U1663 (N_1663,In_1447,In_1718);
xnor U1664 (N_1664,In_2385,In_686);
nand U1665 (N_1665,In_2893,In_199);
nand U1666 (N_1666,In_2031,In_2674);
or U1667 (N_1667,In_186,In_251);
nand U1668 (N_1668,In_871,In_2041);
nand U1669 (N_1669,In_879,In_1823);
or U1670 (N_1670,In_2473,In_2430);
xor U1671 (N_1671,In_554,In_890);
nor U1672 (N_1672,In_1347,In_1503);
or U1673 (N_1673,In_627,In_2054);
or U1674 (N_1674,In_175,In_1498);
or U1675 (N_1675,In_2819,In_2121);
or U1676 (N_1676,In_594,In_1313);
nor U1677 (N_1677,In_2253,In_1670);
nand U1678 (N_1678,In_2428,In_2298);
xor U1679 (N_1679,In_751,In_373);
nand U1680 (N_1680,In_1556,In_376);
nand U1681 (N_1681,In_1514,In_1576);
nand U1682 (N_1682,In_2795,In_1239);
and U1683 (N_1683,In_2337,In_526);
nor U1684 (N_1684,In_1352,In_777);
nand U1685 (N_1685,In_347,In_2168);
nand U1686 (N_1686,In_378,In_1153);
nand U1687 (N_1687,In_1042,In_2466);
and U1688 (N_1688,In_617,In_2620);
or U1689 (N_1689,In_1077,In_1691);
and U1690 (N_1690,In_2387,In_2742);
nand U1691 (N_1691,In_2590,In_874);
xor U1692 (N_1692,In_869,In_2271);
nand U1693 (N_1693,In_1946,In_332);
nor U1694 (N_1694,In_2745,In_2406);
or U1695 (N_1695,In_2295,In_1390);
nand U1696 (N_1696,In_1838,In_2034);
nor U1697 (N_1697,In_1505,In_912);
nand U1698 (N_1698,In_2991,In_2409);
nand U1699 (N_1699,In_596,In_598);
xor U1700 (N_1700,In_1154,In_2352);
or U1701 (N_1701,In_61,In_1420);
xor U1702 (N_1702,In_2642,In_2120);
or U1703 (N_1703,In_2617,In_2767);
nor U1704 (N_1704,In_1595,In_2563);
or U1705 (N_1705,In_2568,In_2683);
xor U1706 (N_1706,In_2596,In_2030);
xor U1707 (N_1707,In_487,In_1939);
nand U1708 (N_1708,In_2247,In_141);
and U1709 (N_1709,In_1959,In_2178);
nand U1710 (N_1710,In_876,In_903);
nand U1711 (N_1711,In_236,In_1721);
nand U1712 (N_1712,In_500,In_1197);
nor U1713 (N_1713,In_524,In_1575);
nand U1714 (N_1714,In_497,In_772);
nor U1715 (N_1715,In_608,In_2397);
and U1716 (N_1716,In_2556,In_1375);
xor U1717 (N_1717,In_865,In_2463);
nand U1718 (N_1718,In_1687,In_956);
xor U1719 (N_1719,In_501,In_2791);
nand U1720 (N_1720,In_23,In_604);
xnor U1721 (N_1721,In_485,In_1260);
nand U1722 (N_1722,In_2701,In_1258);
xnor U1723 (N_1723,In_889,In_225);
nor U1724 (N_1724,In_1433,In_2700);
and U1725 (N_1725,In_280,In_1619);
xor U1726 (N_1726,In_2893,In_805);
nor U1727 (N_1727,In_1248,In_1171);
xnor U1728 (N_1728,In_1794,In_1540);
nand U1729 (N_1729,In_2203,In_1418);
or U1730 (N_1730,In_1826,In_426);
nand U1731 (N_1731,In_560,In_629);
nand U1732 (N_1732,In_1103,In_1167);
nand U1733 (N_1733,In_214,In_2381);
nand U1734 (N_1734,In_1337,In_1843);
nand U1735 (N_1735,In_1417,In_797);
nand U1736 (N_1736,In_2042,In_1853);
nand U1737 (N_1737,In_623,In_380);
or U1738 (N_1738,In_1286,In_2218);
nand U1739 (N_1739,In_1264,In_1853);
and U1740 (N_1740,In_2344,In_820);
xor U1741 (N_1741,In_1871,In_2313);
or U1742 (N_1742,In_2685,In_1404);
xor U1743 (N_1743,In_288,In_2563);
nand U1744 (N_1744,In_2012,In_1965);
and U1745 (N_1745,In_1218,In_619);
xor U1746 (N_1746,In_963,In_1018);
and U1747 (N_1747,In_1718,In_1782);
nor U1748 (N_1748,In_2854,In_829);
and U1749 (N_1749,In_2103,In_1936);
nand U1750 (N_1750,In_615,In_1623);
or U1751 (N_1751,In_314,In_42);
nand U1752 (N_1752,In_1654,In_2986);
nor U1753 (N_1753,In_2274,In_1497);
and U1754 (N_1754,In_2033,In_2184);
xor U1755 (N_1755,In_73,In_1249);
nor U1756 (N_1756,In_1898,In_2737);
nand U1757 (N_1757,In_2493,In_2225);
and U1758 (N_1758,In_749,In_1069);
or U1759 (N_1759,In_1845,In_2824);
or U1760 (N_1760,In_1225,In_2319);
or U1761 (N_1761,In_2266,In_2755);
and U1762 (N_1762,In_458,In_1930);
nand U1763 (N_1763,In_643,In_1928);
xor U1764 (N_1764,In_1129,In_2941);
or U1765 (N_1765,In_1591,In_612);
or U1766 (N_1766,In_2271,In_74);
xnor U1767 (N_1767,In_1960,In_2574);
or U1768 (N_1768,In_1880,In_1247);
xor U1769 (N_1769,In_247,In_2274);
or U1770 (N_1770,In_2313,In_1196);
nand U1771 (N_1771,In_1733,In_1323);
nand U1772 (N_1772,In_1208,In_330);
nor U1773 (N_1773,In_2189,In_2144);
nand U1774 (N_1774,In_641,In_2631);
nor U1775 (N_1775,In_1929,In_100);
xnor U1776 (N_1776,In_1985,In_1915);
nor U1777 (N_1777,In_1885,In_2698);
xnor U1778 (N_1778,In_801,In_889);
nand U1779 (N_1779,In_777,In_1242);
or U1780 (N_1780,In_361,In_1215);
and U1781 (N_1781,In_690,In_1198);
nand U1782 (N_1782,In_2860,In_1639);
and U1783 (N_1783,In_709,In_1327);
nand U1784 (N_1784,In_456,In_1560);
xor U1785 (N_1785,In_2407,In_1478);
and U1786 (N_1786,In_2691,In_2484);
nand U1787 (N_1787,In_2300,In_1345);
nand U1788 (N_1788,In_1005,In_2146);
or U1789 (N_1789,In_773,In_698);
nand U1790 (N_1790,In_1677,In_375);
nand U1791 (N_1791,In_1353,In_190);
nor U1792 (N_1792,In_2466,In_950);
xnor U1793 (N_1793,In_536,In_2173);
or U1794 (N_1794,In_91,In_1997);
xnor U1795 (N_1795,In_1159,In_380);
nand U1796 (N_1796,In_969,In_2460);
or U1797 (N_1797,In_568,In_1873);
and U1798 (N_1798,In_2311,In_2457);
or U1799 (N_1799,In_1171,In_2697);
xor U1800 (N_1800,In_214,In_2094);
or U1801 (N_1801,In_502,In_2536);
and U1802 (N_1802,In_2841,In_1311);
xnor U1803 (N_1803,In_2071,In_1818);
nand U1804 (N_1804,In_689,In_1144);
nand U1805 (N_1805,In_1634,In_2470);
xor U1806 (N_1806,In_2146,In_2874);
and U1807 (N_1807,In_2589,In_2428);
xnor U1808 (N_1808,In_113,In_50);
or U1809 (N_1809,In_817,In_2628);
and U1810 (N_1810,In_253,In_1228);
nand U1811 (N_1811,In_729,In_332);
nor U1812 (N_1812,In_2085,In_356);
xnor U1813 (N_1813,In_1750,In_2197);
or U1814 (N_1814,In_185,In_589);
xnor U1815 (N_1815,In_2388,In_1415);
and U1816 (N_1816,In_151,In_97);
nand U1817 (N_1817,In_1764,In_1759);
and U1818 (N_1818,In_1390,In_2072);
or U1819 (N_1819,In_606,In_2352);
or U1820 (N_1820,In_909,In_810);
xor U1821 (N_1821,In_2655,In_304);
nor U1822 (N_1822,In_229,In_1773);
or U1823 (N_1823,In_485,In_2045);
or U1824 (N_1824,In_821,In_300);
nor U1825 (N_1825,In_1373,In_331);
xor U1826 (N_1826,In_451,In_1202);
nor U1827 (N_1827,In_1139,In_254);
nand U1828 (N_1828,In_2107,In_325);
xnor U1829 (N_1829,In_2001,In_1096);
or U1830 (N_1830,In_2786,In_1566);
nand U1831 (N_1831,In_1580,In_1132);
and U1832 (N_1832,In_1558,In_2501);
or U1833 (N_1833,In_1269,In_401);
or U1834 (N_1834,In_2606,In_2065);
nor U1835 (N_1835,In_825,In_2537);
and U1836 (N_1836,In_295,In_1653);
or U1837 (N_1837,In_2286,In_262);
xor U1838 (N_1838,In_1391,In_807);
xnor U1839 (N_1839,In_2327,In_961);
xnor U1840 (N_1840,In_2820,In_2290);
and U1841 (N_1841,In_1840,In_1090);
and U1842 (N_1842,In_590,In_2796);
nor U1843 (N_1843,In_1039,In_1568);
xor U1844 (N_1844,In_1793,In_914);
nor U1845 (N_1845,In_1471,In_1600);
or U1846 (N_1846,In_341,In_1069);
xor U1847 (N_1847,In_2356,In_1666);
xnor U1848 (N_1848,In_64,In_811);
nor U1849 (N_1849,In_1428,In_1204);
or U1850 (N_1850,In_606,In_1821);
nor U1851 (N_1851,In_133,In_1484);
nor U1852 (N_1852,In_1415,In_2070);
nand U1853 (N_1853,In_2762,In_2971);
nor U1854 (N_1854,In_776,In_2903);
nand U1855 (N_1855,In_1414,In_488);
or U1856 (N_1856,In_834,In_1847);
nand U1857 (N_1857,In_2348,In_2346);
nand U1858 (N_1858,In_2298,In_2394);
nor U1859 (N_1859,In_445,In_1762);
and U1860 (N_1860,In_761,In_1012);
nand U1861 (N_1861,In_210,In_206);
or U1862 (N_1862,In_2789,In_2713);
xnor U1863 (N_1863,In_2123,In_818);
xnor U1864 (N_1864,In_916,In_1178);
xor U1865 (N_1865,In_501,In_812);
or U1866 (N_1866,In_1270,In_2735);
nor U1867 (N_1867,In_2129,In_2580);
and U1868 (N_1868,In_98,In_481);
or U1869 (N_1869,In_2181,In_1377);
or U1870 (N_1870,In_2625,In_663);
or U1871 (N_1871,In_2541,In_2436);
nor U1872 (N_1872,In_2355,In_1682);
xnor U1873 (N_1873,In_689,In_1356);
nand U1874 (N_1874,In_2593,In_227);
xor U1875 (N_1875,In_1308,In_2828);
xnor U1876 (N_1876,In_177,In_2181);
or U1877 (N_1877,In_2897,In_1160);
and U1878 (N_1878,In_1337,In_2901);
or U1879 (N_1879,In_355,In_1252);
xnor U1880 (N_1880,In_1307,In_2283);
nor U1881 (N_1881,In_2902,In_742);
xnor U1882 (N_1882,In_1766,In_434);
xor U1883 (N_1883,In_778,In_2301);
nor U1884 (N_1884,In_19,In_2899);
or U1885 (N_1885,In_2981,In_1033);
nor U1886 (N_1886,In_2686,In_2611);
xnor U1887 (N_1887,In_2932,In_1148);
and U1888 (N_1888,In_733,In_1653);
nand U1889 (N_1889,In_2610,In_274);
nand U1890 (N_1890,In_1714,In_808);
nor U1891 (N_1891,In_1744,In_973);
nand U1892 (N_1892,In_2077,In_2837);
and U1893 (N_1893,In_2719,In_1163);
nand U1894 (N_1894,In_2974,In_2369);
or U1895 (N_1895,In_509,In_1611);
nor U1896 (N_1896,In_429,In_434);
and U1897 (N_1897,In_2348,In_692);
and U1898 (N_1898,In_2414,In_1109);
and U1899 (N_1899,In_811,In_1122);
nand U1900 (N_1900,In_1105,In_2498);
or U1901 (N_1901,In_2627,In_383);
and U1902 (N_1902,In_1942,In_638);
xor U1903 (N_1903,In_2383,In_1638);
xor U1904 (N_1904,In_2330,In_2239);
nand U1905 (N_1905,In_2922,In_857);
nor U1906 (N_1906,In_1638,In_2622);
or U1907 (N_1907,In_520,In_209);
xnor U1908 (N_1908,In_2819,In_1978);
or U1909 (N_1909,In_497,In_1153);
nor U1910 (N_1910,In_1187,In_13);
and U1911 (N_1911,In_1662,In_2252);
xnor U1912 (N_1912,In_2132,In_1787);
xor U1913 (N_1913,In_370,In_514);
and U1914 (N_1914,In_1759,In_1431);
nor U1915 (N_1915,In_658,In_199);
or U1916 (N_1916,In_2013,In_2730);
nor U1917 (N_1917,In_1699,In_270);
xnor U1918 (N_1918,In_30,In_2378);
and U1919 (N_1919,In_264,In_1212);
nor U1920 (N_1920,In_1369,In_422);
or U1921 (N_1921,In_2591,In_1927);
xnor U1922 (N_1922,In_2313,In_1801);
nor U1923 (N_1923,In_1616,In_2206);
xnor U1924 (N_1924,In_2777,In_2378);
nand U1925 (N_1925,In_766,In_189);
or U1926 (N_1926,In_1933,In_2741);
and U1927 (N_1927,In_177,In_658);
nor U1928 (N_1928,In_1626,In_2832);
nand U1929 (N_1929,In_2545,In_2463);
and U1930 (N_1930,In_754,In_534);
nor U1931 (N_1931,In_2951,In_2100);
or U1932 (N_1932,In_235,In_2882);
and U1933 (N_1933,In_2190,In_2222);
or U1934 (N_1934,In_264,In_2021);
and U1935 (N_1935,In_1382,In_2975);
nor U1936 (N_1936,In_940,In_2530);
or U1937 (N_1937,In_2937,In_1560);
and U1938 (N_1938,In_2298,In_160);
or U1939 (N_1939,In_1887,In_863);
and U1940 (N_1940,In_2044,In_738);
and U1941 (N_1941,In_1607,In_414);
and U1942 (N_1942,In_16,In_584);
xnor U1943 (N_1943,In_1247,In_1259);
or U1944 (N_1944,In_2589,In_1040);
xor U1945 (N_1945,In_1836,In_1220);
nor U1946 (N_1946,In_2789,In_558);
nor U1947 (N_1947,In_2117,In_739);
xor U1948 (N_1948,In_2705,In_2843);
nand U1949 (N_1949,In_2293,In_2741);
nand U1950 (N_1950,In_2926,In_913);
or U1951 (N_1951,In_1118,In_187);
and U1952 (N_1952,In_1356,In_2291);
or U1953 (N_1953,In_2046,In_2282);
nor U1954 (N_1954,In_2466,In_1819);
xnor U1955 (N_1955,In_2816,In_431);
and U1956 (N_1956,In_1819,In_2718);
xor U1957 (N_1957,In_1964,In_1131);
nand U1958 (N_1958,In_1255,In_2550);
nor U1959 (N_1959,In_2057,In_1341);
and U1960 (N_1960,In_118,In_1520);
xnor U1961 (N_1961,In_2742,In_2501);
nand U1962 (N_1962,In_2640,In_2600);
nor U1963 (N_1963,In_1082,In_2650);
nor U1964 (N_1964,In_1460,In_1744);
nor U1965 (N_1965,In_2619,In_1456);
xnor U1966 (N_1966,In_1723,In_1856);
or U1967 (N_1967,In_443,In_1725);
nand U1968 (N_1968,In_1804,In_2250);
and U1969 (N_1969,In_1932,In_1605);
xnor U1970 (N_1970,In_1154,In_2495);
nand U1971 (N_1971,In_555,In_2262);
nor U1972 (N_1972,In_146,In_671);
nor U1973 (N_1973,In_655,In_1718);
or U1974 (N_1974,In_2874,In_2260);
nor U1975 (N_1975,In_2583,In_1306);
or U1976 (N_1976,In_2548,In_2515);
or U1977 (N_1977,In_1677,In_802);
nor U1978 (N_1978,In_973,In_110);
xnor U1979 (N_1979,In_2819,In_1258);
xor U1980 (N_1980,In_2614,In_1025);
nor U1981 (N_1981,In_945,In_270);
nand U1982 (N_1982,In_451,In_2053);
nand U1983 (N_1983,In_2501,In_1004);
or U1984 (N_1984,In_782,In_1309);
nor U1985 (N_1985,In_876,In_650);
or U1986 (N_1986,In_1555,In_590);
or U1987 (N_1987,In_362,In_1083);
xor U1988 (N_1988,In_585,In_1879);
nor U1989 (N_1989,In_1275,In_2206);
xor U1990 (N_1990,In_2085,In_564);
nor U1991 (N_1991,In_1591,In_1652);
nor U1992 (N_1992,In_2658,In_545);
and U1993 (N_1993,In_1583,In_2165);
nand U1994 (N_1994,In_409,In_495);
xnor U1995 (N_1995,In_1827,In_2193);
nand U1996 (N_1996,In_1789,In_2528);
and U1997 (N_1997,In_753,In_44);
and U1998 (N_1998,In_2855,In_1950);
or U1999 (N_1999,In_1578,In_474);
nand U2000 (N_2000,In_1725,In_2274);
and U2001 (N_2001,In_2514,In_886);
xor U2002 (N_2002,In_2680,In_2139);
or U2003 (N_2003,In_2707,In_922);
nor U2004 (N_2004,In_2988,In_1072);
nor U2005 (N_2005,In_1159,In_2575);
nand U2006 (N_2006,In_442,In_27);
xnor U2007 (N_2007,In_1408,In_1423);
xnor U2008 (N_2008,In_2335,In_1656);
xor U2009 (N_2009,In_2342,In_489);
nand U2010 (N_2010,In_950,In_2518);
nand U2011 (N_2011,In_1385,In_1340);
and U2012 (N_2012,In_2433,In_967);
and U2013 (N_2013,In_228,In_367);
nand U2014 (N_2014,In_1006,In_894);
or U2015 (N_2015,In_1345,In_2807);
xor U2016 (N_2016,In_1914,In_2933);
xnor U2017 (N_2017,In_1116,In_2109);
nor U2018 (N_2018,In_338,In_333);
nor U2019 (N_2019,In_2537,In_1549);
xnor U2020 (N_2020,In_1644,In_1141);
xor U2021 (N_2021,In_2903,In_2309);
or U2022 (N_2022,In_13,In_2192);
and U2023 (N_2023,In_2470,In_491);
nand U2024 (N_2024,In_2414,In_2848);
or U2025 (N_2025,In_1737,In_1297);
and U2026 (N_2026,In_2280,In_727);
xor U2027 (N_2027,In_2383,In_308);
nand U2028 (N_2028,In_1224,In_1271);
xor U2029 (N_2029,In_2135,In_1475);
nand U2030 (N_2030,In_530,In_1909);
or U2031 (N_2031,In_702,In_1175);
nor U2032 (N_2032,In_2890,In_2);
xnor U2033 (N_2033,In_2974,In_53);
or U2034 (N_2034,In_1355,In_56);
nor U2035 (N_2035,In_1486,In_409);
nor U2036 (N_2036,In_302,In_2519);
xor U2037 (N_2037,In_1267,In_2168);
nor U2038 (N_2038,In_1379,In_2461);
and U2039 (N_2039,In_1962,In_2668);
nor U2040 (N_2040,In_1702,In_1108);
and U2041 (N_2041,In_724,In_1856);
and U2042 (N_2042,In_1777,In_1710);
nor U2043 (N_2043,In_683,In_2863);
nand U2044 (N_2044,In_1475,In_1876);
or U2045 (N_2045,In_912,In_140);
or U2046 (N_2046,In_1267,In_2216);
xnor U2047 (N_2047,In_2984,In_717);
nand U2048 (N_2048,In_27,In_2266);
nand U2049 (N_2049,In_744,In_1565);
and U2050 (N_2050,In_166,In_1744);
nand U2051 (N_2051,In_2673,In_1309);
nor U2052 (N_2052,In_1738,In_2138);
xnor U2053 (N_2053,In_1095,In_2180);
or U2054 (N_2054,In_1938,In_554);
and U2055 (N_2055,In_908,In_1378);
nor U2056 (N_2056,In_44,In_624);
nand U2057 (N_2057,In_1926,In_2170);
nand U2058 (N_2058,In_2856,In_1989);
and U2059 (N_2059,In_2266,In_632);
or U2060 (N_2060,In_1312,In_164);
nand U2061 (N_2061,In_415,In_2937);
nor U2062 (N_2062,In_1507,In_1988);
nor U2063 (N_2063,In_1799,In_1265);
and U2064 (N_2064,In_924,In_1462);
and U2065 (N_2065,In_1395,In_1192);
or U2066 (N_2066,In_1950,In_648);
xor U2067 (N_2067,In_242,In_2388);
nor U2068 (N_2068,In_321,In_1142);
nand U2069 (N_2069,In_979,In_530);
xor U2070 (N_2070,In_1577,In_1449);
nand U2071 (N_2071,In_1808,In_1092);
xor U2072 (N_2072,In_1544,In_555);
xor U2073 (N_2073,In_2666,In_2753);
or U2074 (N_2074,In_2330,In_384);
and U2075 (N_2075,In_1110,In_212);
nand U2076 (N_2076,In_1259,In_2873);
xnor U2077 (N_2077,In_508,In_2154);
nor U2078 (N_2078,In_1671,In_2836);
and U2079 (N_2079,In_1004,In_2830);
nand U2080 (N_2080,In_2432,In_2119);
or U2081 (N_2081,In_2043,In_1117);
xnor U2082 (N_2082,In_1852,In_1820);
xnor U2083 (N_2083,In_2011,In_851);
or U2084 (N_2084,In_623,In_535);
nor U2085 (N_2085,In_2365,In_384);
or U2086 (N_2086,In_2279,In_2923);
and U2087 (N_2087,In_895,In_2054);
and U2088 (N_2088,In_866,In_2493);
nor U2089 (N_2089,In_923,In_797);
and U2090 (N_2090,In_2253,In_1933);
or U2091 (N_2091,In_1544,In_1725);
or U2092 (N_2092,In_2825,In_184);
nand U2093 (N_2093,In_1398,In_812);
xnor U2094 (N_2094,In_2372,In_1232);
and U2095 (N_2095,In_1018,In_43);
nand U2096 (N_2096,In_1606,In_271);
nand U2097 (N_2097,In_1003,In_2483);
and U2098 (N_2098,In_862,In_2062);
and U2099 (N_2099,In_2335,In_2847);
nor U2100 (N_2100,In_1837,In_1164);
nand U2101 (N_2101,In_1448,In_507);
nand U2102 (N_2102,In_1898,In_2976);
nor U2103 (N_2103,In_787,In_1936);
nand U2104 (N_2104,In_716,In_1466);
or U2105 (N_2105,In_501,In_1988);
nor U2106 (N_2106,In_194,In_2779);
xnor U2107 (N_2107,In_466,In_435);
xnor U2108 (N_2108,In_1755,In_545);
and U2109 (N_2109,In_1312,In_1565);
nor U2110 (N_2110,In_2931,In_2563);
xnor U2111 (N_2111,In_1701,In_2784);
nor U2112 (N_2112,In_787,In_164);
nand U2113 (N_2113,In_2578,In_515);
xor U2114 (N_2114,In_2799,In_739);
xor U2115 (N_2115,In_2533,In_307);
nor U2116 (N_2116,In_1933,In_1080);
nor U2117 (N_2117,In_1572,In_221);
and U2118 (N_2118,In_2549,In_8);
or U2119 (N_2119,In_1880,In_903);
nor U2120 (N_2120,In_2259,In_2970);
nor U2121 (N_2121,In_2261,In_364);
nand U2122 (N_2122,In_622,In_1780);
nor U2123 (N_2123,In_2854,In_2783);
nand U2124 (N_2124,In_1438,In_119);
and U2125 (N_2125,In_1708,In_1061);
and U2126 (N_2126,In_1266,In_1738);
and U2127 (N_2127,In_1646,In_2913);
or U2128 (N_2128,In_984,In_2443);
nand U2129 (N_2129,In_1993,In_408);
and U2130 (N_2130,In_2324,In_753);
or U2131 (N_2131,In_220,In_1106);
or U2132 (N_2132,In_854,In_138);
nor U2133 (N_2133,In_1224,In_1508);
nor U2134 (N_2134,In_1736,In_2253);
xor U2135 (N_2135,In_2074,In_318);
xnor U2136 (N_2136,In_2538,In_406);
nor U2137 (N_2137,In_1383,In_1947);
nand U2138 (N_2138,In_1227,In_871);
nand U2139 (N_2139,In_1741,In_1822);
nor U2140 (N_2140,In_720,In_1799);
nor U2141 (N_2141,In_1625,In_2234);
or U2142 (N_2142,In_1868,In_851);
nand U2143 (N_2143,In_690,In_413);
and U2144 (N_2144,In_1706,In_2);
nor U2145 (N_2145,In_602,In_1057);
or U2146 (N_2146,In_2548,In_746);
or U2147 (N_2147,In_40,In_1822);
nor U2148 (N_2148,In_1626,In_2632);
xor U2149 (N_2149,In_707,In_289);
or U2150 (N_2150,In_623,In_1229);
and U2151 (N_2151,In_2331,In_1943);
or U2152 (N_2152,In_2021,In_193);
and U2153 (N_2153,In_2737,In_2948);
and U2154 (N_2154,In_274,In_1799);
nand U2155 (N_2155,In_424,In_854);
nor U2156 (N_2156,In_376,In_994);
nor U2157 (N_2157,In_1747,In_2582);
and U2158 (N_2158,In_1959,In_2935);
nor U2159 (N_2159,In_50,In_1595);
or U2160 (N_2160,In_40,In_1467);
or U2161 (N_2161,In_323,In_444);
or U2162 (N_2162,In_702,In_1673);
xnor U2163 (N_2163,In_1284,In_602);
or U2164 (N_2164,In_393,In_408);
or U2165 (N_2165,In_254,In_756);
nor U2166 (N_2166,In_2220,In_873);
and U2167 (N_2167,In_204,In_2045);
and U2168 (N_2168,In_355,In_2906);
nand U2169 (N_2169,In_2341,In_798);
nor U2170 (N_2170,In_2786,In_2117);
xor U2171 (N_2171,In_1179,In_352);
and U2172 (N_2172,In_285,In_1666);
and U2173 (N_2173,In_1028,In_1276);
nand U2174 (N_2174,In_1807,In_2153);
and U2175 (N_2175,In_1076,In_2985);
and U2176 (N_2176,In_2310,In_2983);
xor U2177 (N_2177,In_1170,In_1843);
nand U2178 (N_2178,In_1241,In_2337);
xnor U2179 (N_2179,In_1650,In_1979);
or U2180 (N_2180,In_1333,In_2643);
and U2181 (N_2181,In_771,In_1873);
and U2182 (N_2182,In_1996,In_1339);
or U2183 (N_2183,In_932,In_2682);
nor U2184 (N_2184,In_1753,In_433);
or U2185 (N_2185,In_1182,In_2346);
nor U2186 (N_2186,In_2440,In_171);
nor U2187 (N_2187,In_1630,In_416);
or U2188 (N_2188,In_1295,In_1720);
nand U2189 (N_2189,In_52,In_799);
or U2190 (N_2190,In_476,In_2637);
or U2191 (N_2191,In_2335,In_303);
nand U2192 (N_2192,In_241,In_829);
and U2193 (N_2193,In_1317,In_120);
xnor U2194 (N_2194,In_2674,In_81);
or U2195 (N_2195,In_2727,In_1412);
xnor U2196 (N_2196,In_486,In_1974);
nor U2197 (N_2197,In_1608,In_2575);
nand U2198 (N_2198,In_2789,In_2485);
xor U2199 (N_2199,In_2947,In_731);
and U2200 (N_2200,In_986,In_2250);
nand U2201 (N_2201,In_2368,In_747);
or U2202 (N_2202,In_2705,In_1651);
nand U2203 (N_2203,In_26,In_480);
nor U2204 (N_2204,In_1021,In_2479);
xor U2205 (N_2205,In_2873,In_2321);
nand U2206 (N_2206,In_1813,In_2617);
or U2207 (N_2207,In_1403,In_2);
nor U2208 (N_2208,In_2090,In_2958);
or U2209 (N_2209,In_1977,In_1771);
or U2210 (N_2210,In_1117,In_2929);
nand U2211 (N_2211,In_2862,In_1775);
or U2212 (N_2212,In_1851,In_2652);
or U2213 (N_2213,In_497,In_2948);
nand U2214 (N_2214,In_1102,In_2063);
and U2215 (N_2215,In_1003,In_2771);
and U2216 (N_2216,In_2408,In_1078);
or U2217 (N_2217,In_423,In_1008);
or U2218 (N_2218,In_442,In_2764);
nor U2219 (N_2219,In_1672,In_2375);
nor U2220 (N_2220,In_447,In_2962);
nand U2221 (N_2221,In_856,In_2616);
nor U2222 (N_2222,In_2990,In_2107);
or U2223 (N_2223,In_159,In_1586);
nand U2224 (N_2224,In_1597,In_1212);
or U2225 (N_2225,In_1507,In_2464);
and U2226 (N_2226,In_1516,In_1954);
nand U2227 (N_2227,In_951,In_2306);
or U2228 (N_2228,In_162,In_2869);
nand U2229 (N_2229,In_228,In_2316);
xor U2230 (N_2230,In_1827,In_2846);
xnor U2231 (N_2231,In_431,In_307);
nor U2232 (N_2232,In_466,In_913);
nand U2233 (N_2233,In_2171,In_363);
nor U2234 (N_2234,In_1732,In_690);
nor U2235 (N_2235,In_1990,In_577);
or U2236 (N_2236,In_2741,In_744);
nand U2237 (N_2237,In_1797,In_2130);
xor U2238 (N_2238,In_1693,In_1946);
nor U2239 (N_2239,In_1865,In_1336);
nand U2240 (N_2240,In_153,In_2010);
or U2241 (N_2241,In_2815,In_345);
nand U2242 (N_2242,In_1262,In_1768);
nor U2243 (N_2243,In_998,In_735);
xor U2244 (N_2244,In_288,In_1888);
or U2245 (N_2245,In_716,In_2288);
xor U2246 (N_2246,In_672,In_1295);
or U2247 (N_2247,In_653,In_1042);
xnor U2248 (N_2248,In_802,In_954);
or U2249 (N_2249,In_797,In_2621);
and U2250 (N_2250,In_2636,In_533);
nor U2251 (N_2251,In_888,In_128);
nand U2252 (N_2252,In_887,In_871);
and U2253 (N_2253,In_1759,In_2981);
nand U2254 (N_2254,In_998,In_1107);
or U2255 (N_2255,In_2897,In_171);
nand U2256 (N_2256,In_656,In_1242);
and U2257 (N_2257,In_2933,In_415);
and U2258 (N_2258,In_383,In_1645);
nand U2259 (N_2259,In_2900,In_211);
nand U2260 (N_2260,In_210,In_2036);
nor U2261 (N_2261,In_2131,In_2772);
xnor U2262 (N_2262,In_1879,In_2185);
or U2263 (N_2263,In_2585,In_2422);
nor U2264 (N_2264,In_114,In_1151);
or U2265 (N_2265,In_2601,In_498);
xnor U2266 (N_2266,In_2494,In_1011);
nor U2267 (N_2267,In_2194,In_1658);
nand U2268 (N_2268,In_208,In_1501);
nand U2269 (N_2269,In_1862,In_35);
and U2270 (N_2270,In_2703,In_827);
and U2271 (N_2271,In_2656,In_501);
xnor U2272 (N_2272,In_2743,In_1263);
nor U2273 (N_2273,In_359,In_1876);
nor U2274 (N_2274,In_1742,In_911);
and U2275 (N_2275,In_1706,In_2636);
nor U2276 (N_2276,In_1134,In_1746);
xor U2277 (N_2277,In_2961,In_479);
nand U2278 (N_2278,In_2080,In_307);
or U2279 (N_2279,In_211,In_2845);
xnor U2280 (N_2280,In_1546,In_1210);
or U2281 (N_2281,In_425,In_1524);
or U2282 (N_2282,In_2255,In_2023);
and U2283 (N_2283,In_2157,In_1415);
xnor U2284 (N_2284,In_1393,In_1237);
xnor U2285 (N_2285,In_700,In_935);
nor U2286 (N_2286,In_287,In_566);
nand U2287 (N_2287,In_1688,In_2268);
and U2288 (N_2288,In_2487,In_2236);
nor U2289 (N_2289,In_70,In_157);
and U2290 (N_2290,In_220,In_2885);
nor U2291 (N_2291,In_1168,In_1928);
or U2292 (N_2292,In_1894,In_1956);
xnor U2293 (N_2293,In_843,In_1116);
nand U2294 (N_2294,In_1817,In_1752);
or U2295 (N_2295,In_2097,In_2868);
xnor U2296 (N_2296,In_2365,In_143);
xnor U2297 (N_2297,In_2179,In_1814);
or U2298 (N_2298,In_1889,In_746);
or U2299 (N_2299,In_1463,In_1473);
xor U2300 (N_2300,In_1700,In_1110);
and U2301 (N_2301,In_2519,In_274);
xnor U2302 (N_2302,In_2970,In_2033);
xor U2303 (N_2303,In_457,In_930);
nor U2304 (N_2304,In_1437,In_2522);
or U2305 (N_2305,In_1533,In_1109);
xor U2306 (N_2306,In_1075,In_2175);
nor U2307 (N_2307,In_2118,In_2267);
nand U2308 (N_2308,In_1652,In_412);
xor U2309 (N_2309,In_116,In_1292);
nor U2310 (N_2310,In_157,In_185);
xnor U2311 (N_2311,In_350,In_2996);
and U2312 (N_2312,In_1,In_1494);
xnor U2313 (N_2313,In_1228,In_2876);
and U2314 (N_2314,In_588,In_1199);
xnor U2315 (N_2315,In_2560,In_1360);
and U2316 (N_2316,In_2451,In_859);
and U2317 (N_2317,In_2816,In_2752);
or U2318 (N_2318,In_2984,In_292);
and U2319 (N_2319,In_695,In_2272);
nand U2320 (N_2320,In_2150,In_814);
xnor U2321 (N_2321,In_2671,In_1652);
nand U2322 (N_2322,In_1951,In_939);
and U2323 (N_2323,In_2318,In_1124);
nor U2324 (N_2324,In_932,In_700);
nor U2325 (N_2325,In_2887,In_1377);
xnor U2326 (N_2326,In_2581,In_829);
xnor U2327 (N_2327,In_887,In_1569);
or U2328 (N_2328,In_2189,In_1471);
xnor U2329 (N_2329,In_2079,In_784);
nor U2330 (N_2330,In_292,In_907);
nand U2331 (N_2331,In_2520,In_2466);
nor U2332 (N_2332,In_2481,In_2408);
nor U2333 (N_2333,In_2484,In_255);
and U2334 (N_2334,In_296,In_834);
nor U2335 (N_2335,In_2694,In_1678);
and U2336 (N_2336,In_71,In_2157);
nor U2337 (N_2337,In_1070,In_1390);
or U2338 (N_2338,In_360,In_1551);
nor U2339 (N_2339,In_516,In_950);
and U2340 (N_2340,In_93,In_1209);
xor U2341 (N_2341,In_2445,In_961);
xnor U2342 (N_2342,In_1371,In_1200);
xor U2343 (N_2343,In_700,In_2418);
or U2344 (N_2344,In_672,In_2605);
xnor U2345 (N_2345,In_957,In_1227);
and U2346 (N_2346,In_441,In_1098);
xor U2347 (N_2347,In_2958,In_2084);
xor U2348 (N_2348,In_561,In_614);
nand U2349 (N_2349,In_229,In_609);
nand U2350 (N_2350,In_516,In_2744);
and U2351 (N_2351,In_2864,In_2728);
and U2352 (N_2352,In_581,In_1779);
or U2353 (N_2353,In_2870,In_2217);
xor U2354 (N_2354,In_2468,In_2274);
nand U2355 (N_2355,In_737,In_2690);
nor U2356 (N_2356,In_2763,In_1416);
and U2357 (N_2357,In_2105,In_125);
and U2358 (N_2358,In_1016,In_122);
and U2359 (N_2359,In_2690,In_887);
nand U2360 (N_2360,In_897,In_2203);
xnor U2361 (N_2361,In_10,In_1428);
or U2362 (N_2362,In_1268,In_1462);
nor U2363 (N_2363,In_360,In_619);
xnor U2364 (N_2364,In_2926,In_95);
nand U2365 (N_2365,In_1682,In_896);
nor U2366 (N_2366,In_869,In_2468);
or U2367 (N_2367,In_2951,In_728);
or U2368 (N_2368,In_2421,In_520);
xor U2369 (N_2369,In_2602,In_816);
nand U2370 (N_2370,In_1849,In_2527);
and U2371 (N_2371,In_1235,In_1211);
nand U2372 (N_2372,In_2959,In_2487);
nand U2373 (N_2373,In_2537,In_1720);
xnor U2374 (N_2374,In_2403,In_1677);
and U2375 (N_2375,In_534,In_910);
or U2376 (N_2376,In_2599,In_2045);
nor U2377 (N_2377,In_672,In_147);
nor U2378 (N_2378,In_155,In_2680);
xnor U2379 (N_2379,In_424,In_1693);
xor U2380 (N_2380,In_1929,In_2222);
nor U2381 (N_2381,In_2978,In_2233);
xor U2382 (N_2382,In_2584,In_1292);
and U2383 (N_2383,In_2744,In_2584);
nor U2384 (N_2384,In_2704,In_243);
xnor U2385 (N_2385,In_933,In_2871);
xnor U2386 (N_2386,In_1268,In_2138);
and U2387 (N_2387,In_1861,In_1812);
or U2388 (N_2388,In_1975,In_2105);
nor U2389 (N_2389,In_2365,In_404);
or U2390 (N_2390,In_1777,In_2217);
and U2391 (N_2391,In_288,In_398);
or U2392 (N_2392,In_2088,In_508);
xor U2393 (N_2393,In_2666,In_2246);
or U2394 (N_2394,In_2794,In_2236);
nand U2395 (N_2395,In_2537,In_169);
xnor U2396 (N_2396,In_1566,In_1548);
xnor U2397 (N_2397,In_2966,In_838);
nor U2398 (N_2398,In_1348,In_1413);
nor U2399 (N_2399,In_2681,In_2926);
nor U2400 (N_2400,In_1254,In_925);
nand U2401 (N_2401,In_2786,In_2751);
nand U2402 (N_2402,In_755,In_406);
nor U2403 (N_2403,In_515,In_2985);
xor U2404 (N_2404,In_56,In_1120);
xor U2405 (N_2405,In_925,In_1851);
nand U2406 (N_2406,In_1619,In_2552);
nand U2407 (N_2407,In_86,In_1973);
or U2408 (N_2408,In_1333,In_778);
xnor U2409 (N_2409,In_663,In_1541);
or U2410 (N_2410,In_1767,In_427);
nand U2411 (N_2411,In_264,In_1413);
and U2412 (N_2412,In_1061,In_313);
xnor U2413 (N_2413,In_2168,In_1236);
nand U2414 (N_2414,In_398,In_2504);
and U2415 (N_2415,In_1298,In_635);
and U2416 (N_2416,In_1175,In_1356);
nor U2417 (N_2417,In_2583,In_2402);
and U2418 (N_2418,In_691,In_2538);
xnor U2419 (N_2419,In_1187,In_514);
nor U2420 (N_2420,In_450,In_1314);
xnor U2421 (N_2421,In_714,In_1314);
nand U2422 (N_2422,In_1895,In_2773);
nor U2423 (N_2423,In_98,In_338);
or U2424 (N_2424,In_1042,In_2818);
nor U2425 (N_2425,In_155,In_426);
nand U2426 (N_2426,In_246,In_1302);
xnor U2427 (N_2427,In_1423,In_530);
nor U2428 (N_2428,In_294,In_2327);
and U2429 (N_2429,In_1128,In_363);
or U2430 (N_2430,In_2390,In_848);
nor U2431 (N_2431,In_2377,In_716);
or U2432 (N_2432,In_1961,In_1462);
nor U2433 (N_2433,In_2647,In_575);
nand U2434 (N_2434,In_1027,In_2795);
or U2435 (N_2435,In_2153,In_975);
or U2436 (N_2436,In_1208,In_699);
and U2437 (N_2437,In_2155,In_248);
and U2438 (N_2438,In_2474,In_1167);
or U2439 (N_2439,In_496,In_2644);
xnor U2440 (N_2440,In_1159,In_343);
nor U2441 (N_2441,In_875,In_775);
and U2442 (N_2442,In_684,In_2509);
nor U2443 (N_2443,In_422,In_609);
or U2444 (N_2444,In_924,In_1858);
xor U2445 (N_2445,In_1299,In_750);
xor U2446 (N_2446,In_462,In_441);
nor U2447 (N_2447,In_2255,In_2995);
nor U2448 (N_2448,In_1616,In_2316);
nor U2449 (N_2449,In_190,In_1308);
xor U2450 (N_2450,In_221,In_1150);
or U2451 (N_2451,In_1346,In_2223);
xnor U2452 (N_2452,In_2644,In_1589);
nor U2453 (N_2453,In_1303,In_2035);
nor U2454 (N_2454,In_1227,In_2426);
nand U2455 (N_2455,In_1811,In_2525);
or U2456 (N_2456,In_819,In_992);
nor U2457 (N_2457,In_183,In_932);
nand U2458 (N_2458,In_2630,In_2395);
or U2459 (N_2459,In_2337,In_2228);
nand U2460 (N_2460,In_2476,In_2778);
nor U2461 (N_2461,In_1447,In_529);
nor U2462 (N_2462,In_387,In_2596);
nor U2463 (N_2463,In_2473,In_1912);
or U2464 (N_2464,In_1545,In_1255);
or U2465 (N_2465,In_818,In_1332);
nor U2466 (N_2466,In_635,In_1093);
and U2467 (N_2467,In_2317,In_340);
and U2468 (N_2468,In_772,In_1264);
nand U2469 (N_2469,In_2709,In_433);
xnor U2470 (N_2470,In_981,In_407);
and U2471 (N_2471,In_2145,In_2060);
nand U2472 (N_2472,In_1238,In_1174);
nand U2473 (N_2473,In_590,In_617);
xor U2474 (N_2474,In_2460,In_2486);
and U2475 (N_2475,In_742,In_2675);
and U2476 (N_2476,In_2799,In_2912);
or U2477 (N_2477,In_42,In_2633);
xor U2478 (N_2478,In_2263,In_1123);
nand U2479 (N_2479,In_986,In_2529);
xor U2480 (N_2480,In_90,In_871);
xor U2481 (N_2481,In_2219,In_451);
xor U2482 (N_2482,In_1135,In_1153);
nor U2483 (N_2483,In_2563,In_1447);
and U2484 (N_2484,In_1501,In_885);
xor U2485 (N_2485,In_2863,In_2073);
or U2486 (N_2486,In_846,In_2947);
nand U2487 (N_2487,In_1588,In_130);
xnor U2488 (N_2488,In_1291,In_2061);
nor U2489 (N_2489,In_2758,In_833);
nor U2490 (N_2490,In_1847,In_2987);
or U2491 (N_2491,In_119,In_1032);
or U2492 (N_2492,In_950,In_1705);
nand U2493 (N_2493,In_1606,In_2475);
nand U2494 (N_2494,In_535,In_506);
xnor U2495 (N_2495,In_345,In_2789);
or U2496 (N_2496,In_2092,In_1056);
or U2497 (N_2497,In_1511,In_1555);
and U2498 (N_2498,In_1975,In_1763);
nor U2499 (N_2499,In_578,In_2587);
xor U2500 (N_2500,In_988,In_1897);
xnor U2501 (N_2501,In_2256,In_1673);
nor U2502 (N_2502,In_610,In_2997);
or U2503 (N_2503,In_295,In_552);
xor U2504 (N_2504,In_2060,In_206);
or U2505 (N_2505,In_2284,In_2506);
and U2506 (N_2506,In_401,In_2424);
nor U2507 (N_2507,In_2260,In_1327);
and U2508 (N_2508,In_2765,In_1462);
nor U2509 (N_2509,In_1393,In_2141);
xnor U2510 (N_2510,In_2102,In_1295);
xnor U2511 (N_2511,In_2498,In_2152);
nand U2512 (N_2512,In_937,In_175);
xnor U2513 (N_2513,In_81,In_559);
and U2514 (N_2514,In_736,In_1716);
nor U2515 (N_2515,In_2513,In_2422);
nor U2516 (N_2516,In_1091,In_2784);
nor U2517 (N_2517,In_1437,In_626);
nand U2518 (N_2518,In_2223,In_2199);
and U2519 (N_2519,In_1198,In_246);
nor U2520 (N_2520,In_2734,In_2140);
nand U2521 (N_2521,In_1770,In_1181);
nor U2522 (N_2522,In_2002,In_1476);
or U2523 (N_2523,In_1722,In_502);
nand U2524 (N_2524,In_1331,In_155);
and U2525 (N_2525,In_1300,In_2311);
nor U2526 (N_2526,In_1269,In_1735);
xor U2527 (N_2527,In_2290,In_1599);
nand U2528 (N_2528,In_1182,In_1570);
nand U2529 (N_2529,In_775,In_154);
nor U2530 (N_2530,In_1528,In_2048);
or U2531 (N_2531,In_2920,In_170);
nand U2532 (N_2532,In_2275,In_2734);
nand U2533 (N_2533,In_815,In_2520);
nor U2534 (N_2534,In_970,In_1421);
xnor U2535 (N_2535,In_263,In_1330);
nor U2536 (N_2536,In_1622,In_1697);
or U2537 (N_2537,In_2142,In_2736);
and U2538 (N_2538,In_1690,In_279);
and U2539 (N_2539,In_829,In_491);
xor U2540 (N_2540,In_1721,In_1160);
or U2541 (N_2541,In_742,In_1256);
and U2542 (N_2542,In_2304,In_357);
xnor U2543 (N_2543,In_503,In_177);
xor U2544 (N_2544,In_1370,In_2161);
xnor U2545 (N_2545,In_1604,In_1504);
xor U2546 (N_2546,In_719,In_2258);
nor U2547 (N_2547,In_1144,In_2483);
nand U2548 (N_2548,In_1024,In_1091);
and U2549 (N_2549,In_952,In_2634);
nand U2550 (N_2550,In_2022,In_2543);
nor U2551 (N_2551,In_2330,In_1165);
nor U2552 (N_2552,In_833,In_1892);
or U2553 (N_2553,In_2196,In_2878);
or U2554 (N_2554,In_768,In_2565);
and U2555 (N_2555,In_2404,In_1385);
nor U2556 (N_2556,In_1553,In_1631);
or U2557 (N_2557,In_1115,In_965);
and U2558 (N_2558,In_334,In_2071);
nor U2559 (N_2559,In_1811,In_1614);
nand U2560 (N_2560,In_376,In_2013);
xor U2561 (N_2561,In_677,In_1773);
nor U2562 (N_2562,In_1147,In_1754);
xor U2563 (N_2563,In_977,In_1340);
nand U2564 (N_2564,In_1915,In_850);
nor U2565 (N_2565,In_571,In_1189);
and U2566 (N_2566,In_1293,In_2320);
xor U2567 (N_2567,In_661,In_1356);
or U2568 (N_2568,In_2494,In_2250);
xor U2569 (N_2569,In_229,In_2179);
xnor U2570 (N_2570,In_1654,In_2100);
and U2571 (N_2571,In_1606,In_2942);
and U2572 (N_2572,In_587,In_2976);
nand U2573 (N_2573,In_1724,In_603);
or U2574 (N_2574,In_1361,In_2802);
or U2575 (N_2575,In_205,In_2239);
nor U2576 (N_2576,In_2654,In_2019);
nand U2577 (N_2577,In_2801,In_1332);
nor U2578 (N_2578,In_366,In_1994);
and U2579 (N_2579,In_1027,In_1767);
and U2580 (N_2580,In_2216,In_1618);
or U2581 (N_2581,In_1853,In_301);
and U2582 (N_2582,In_2268,In_2508);
and U2583 (N_2583,In_284,In_1136);
nand U2584 (N_2584,In_1184,In_518);
and U2585 (N_2585,In_1849,In_2716);
nor U2586 (N_2586,In_197,In_2462);
or U2587 (N_2587,In_1239,In_242);
and U2588 (N_2588,In_1694,In_665);
or U2589 (N_2589,In_2395,In_722);
or U2590 (N_2590,In_641,In_2151);
nor U2591 (N_2591,In_2625,In_2682);
or U2592 (N_2592,In_2314,In_1470);
or U2593 (N_2593,In_2926,In_1235);
xnor U2594 (N_2594,In_950,In_1798);
nand U2595 (N_2595,In_805,In_2007);
xor U2596 (N_2596,In_1880,In_1895);
or U2597 (N_2597,In_493,In_613);
nor U2598 (N_2598,In_620,In_2451);
or U2599 (N_2599,In_1208,In_1041);
nand U2600 (N_2600,In_1640,In_1563);
nor U2601 (N_2601,In_2493,In_2631);
xor U2602 (N_2602,In_648,In_1236);
nor U2603 (N_2603,In_993,In_2753);
and U2604 (N_2604,In_1597,In_1908);
and U2605 (N_2605,In_2186,In_457);
xor U2606 (N_2606,In_2159,In_2427);
or U2607 (N_2607,In_400,In_2849);
and U2608 (N_2608,In_147,In_343);
or U2609 (N_2609,In_1476,In_752);
nand U2610 (N_2610,In_1243,In_2659);
nand U2611 (N_2611,In_1376,In_855);
or U2612 (N_2612,In_34,In_1607);
nor U2613 (N_2613,In_605,In_160);
and U2614 (N_2614,In_1492,In_500);
or U2615 (N_2615,In_2354,In_1401);
and U2616 (N_2616,In_74,In_1407);
or U2617 (N_2617,In_2745,In_1964);
and U2618 (N_2618,In_2714,In_1950);
or U2619 (N_2619,In_2260,In_1968);
xor U2620 (N_2620,In_2497,In_379);
or U2621 (N_2621,In_1854,In_157);
nand U2622 (N_2622,In_1189,In_1704);
or U2623 (N_2623,In_602,In_1463);
nand U2624 (N_2624,In_2424,In_1235);
and U2625 (N_2625,In_618,In_1819);
and U2626 (N_2626,In_1683,In_2701);
xnor U2627 (N_2627,In_879,In_1950);
or U2628 (N_2628,In_1810,In_2083);
xnor U2629 (N_2629,In_888,In_880);
nor U2630 (N_2630,In_671,In_820);
nand U2631 (N_2631,In_2312,In_186);
nand U2632 (N_2632,In_2502,In_2193);
and U2633 (N_2633,In_1807,In_2161);
nor U2634 (N_2634,In_1660,In_2405);
or U2635 (N_2635,In_336,In_2429);
xnor U2636 (N_2636,In_230,In_1088);
nor U2637 (N_2637,In_2654,In_906);
or U2638 (N_2638,In_2496,In_114);
and U2639 (N_2639,In_2510,In_959);
and U2640 (N_2640,In_1733,In_209);
and U2641 (N_2641,In_2417,In_2753);
nor U2642 (N_2642,In_1571,In_2076);
or U2643 (N_2643,In_133,In_315);
or U2644 (N_2644,In_541,In_2304);
xor U2645 (N_2645,In_1122,In_1141);
nor U2646 (N_2646,In_1369,In_2378);
nor U2647 (N_2647,In_1142,In_2912);
and U2648 (N_2648,In_1304,In_1115);
xor U2649 (N_2649,In_1001,In_2817);
xnor U2650 (N_2650,In_987,In_1034);
nor U2651 (N_2651,In_2891,In_674);
and U2652 (N_2652,In_1585,In_2310);
and U2653 (N_2653,In_95,In_1318);
nand U2654 (N_2654,In_1210,In_549);
nand U2655 (N_2655,In_569,In_2899);
nor U2656 (N_2656,In_288,In_2652);
and U2657 (N_2657,In_351,In_588);
and U2658 (N_2658,In_1002,In_1507);
and U2659 (N_2659,In_1807,In_2449);
nand U2660 (N_2660,In_1758,In_2451);
nand U2661 (N_2661,In_1376,In_2049);
nand U2662 (N_2662,In_55,In_2529);
nor U2663 (N_2663,In_2933,In_1549);
nor U2664 (N_2664,In_2757,In_1313);
nor U2665 (N_2665,In_1887,In_672);
or U2666 (N_2666,In_241,In_550);
or U2667 (N_2667,In_2776,In_2285);
or U2668 (N_2668,In_1930,In_1247);
nand U2669 (N_2669,In_1249,In_1454);
and U2670 (N_2670,In_426,In_328);
nand U2671 (N_2671,In_2727,In_1809);
nor U2672 (N_2672,In_1720,In_451);
and U2673 (N_2673,In_2170,In_134);
xnor U2674 (N_2674,In_1061,In_1449);
xor U2675 (N_2675,In_779,In_1856);
xnor U2676 (N_2676,In_1782,In_671);
or U2677 (N_2677,In_2921,In_2618);
and U2678 (N_2678,In_858,In_1538);
xnor U2679 (N_2679,In_183,In_2923);
xnor U2680 (N_2680,In_2975,In_1205);
nand U2681 (N_2681,In_1076,In_409);
nand U2682 (N_2682,In_2038,In_329);
nor U2683 (N_2683,In_1133,In_1869);
nor U2684 (N_2684,In_1856,In_1835);
and U2685 (N_2685,In_2981,In_1742);
or U2686 (N_2686,In_2403,In_840);
and U2687 (N_2687,In_1446,In_634);
and U2688 (N_2688,In_1554,In_2351);
nor U2689 (N_2689,In_1732,In_1468);
nand U2690 (N_2690,In_1664,In_791);
nand U2691 (N_2691,In_515,In_115);
nor U2692 (N_2692,In_576,In_792);
xor U2693 (N_2693,In_1973,In_679);
and U2694 (N_2694,In_2731,In_161);
or U2695 (N_2695,In_1663,In_987);
and U2696 (N_2696,In_4,In_916);
and U2697 (N_2697,In_2278,In_1362);
or U2698 (N_2698,In_1542,In_1515);
xor U2699 (N_2699,In_2676,In_340);
nor U2700 (N_2700,In_767,In_2831);
or U2701 (N_2701,In_1567,In_2052);
xnor U2702 (N_2702,In_118,In_2280);
nor U2703 (N_2703,In_1104,In_1165);
and U2704 (N_2704,In_2344,In_2764);
nand U2705 (N_2705,In_2346,In_2806);
or U2706 (N_2706,In_1881,In_1639);
nand U2707 (N_2707,In_2372,In_813);
nand U2708 (N_2708,In_2326,In_2078);
or U2709 (N_2709,In_2448,In_1779);
or U2710 (N_2710,In_235,In_804);
xnor U2711 (N_2711,In_1650,In_633);
nor U2712 (N_2712,In_858,In_1463);
xor U2713 (N_2713,In_402,In_450);
nand U2714 (N_2714,In_40,In_953);
and U2715 (N_2715,In_756,In_569);
and U2716 (N_2716,In_2008,In_1062);
nand U2717 (N_2717,In_2766,In_2884);
and U2718 (N_2718,In_289,In_577);
or U2719 (N_2719,In_1505,In_2430);
nor U2720 (N_2720,In_2570,In_2191);
or U2721 (N_2721,In_1525,In_1977);
nor U2722 (N_2722,In_2573,In_2834);
nor U2723 (N_2723,In_2092,In_1838);
or U2724 (N_2724,In_1075,In_1932);
or U2725 (N_2725,In_2245,In_2172);
or U2726 (N_2726,In_638,In_786);
nor U2727 (N_2727,In_172,In_738);
or U2728 (N_2728,In_1812,In_1109);
nand U2729 (N_2729,In_547,In_1094);
and U2730 (N_2730,In_2347,In_1126);
nand U2731 (N_2731,In_60,In_913);
or U2732 (N_2732,In_46,In_465);
or U2733 (N_2733,In_2630,In_1896);
or U2734 (N_2734,In_1697,In_2733);
nor U2735 (N_2735,In_2182,In_867);
and U2736 (N_2736,In_817,In_2361);
and U2737 (N_2737,In_28,In_865);
or U2738 (N_2738,In_995,In_1738);
nand U2739 (N_2739,In_1027,In_1246);
nor U2740 (N_2740,In_78,In_650);
nor U2741 (N_2741,In_441,In_2177);
and U2742 (N_2742,In_1518,In_643);
nor U2743 (N_2743,In_1051,In_339);
nor U2744 (N_2744,In_1264,In_2440);
nand U2745 (N_2745,In_355,In_169);
nand U2746 (N_2746,In_13,In_2854);
xor U2747 (N_2747,In_211,In_1822);
or U2748 (N_2748,In_481,In_1318);
nor U2749 (N_2749,In_824,In_716);
xnor U2750 (N_2750,In_1996,In_2888);
nand U2751 (N_2751,In_1068,In_421);
or U2752 (N_2752,In_1429,In_1522);
and U2753 (N_2753,In_1740,In_1059);
nor U2754 (N_2754,In_1626,In_1149);
or U2755 (N_2755,In_2060,In_2339);
nor U2756 (N_2756,In_1414,In_352);
nor U2757 (N_2757,In_2829,In_504);
nor U2758 (N_2758,In_2210,In_561);
or U2759 (N_2759,In_2800,In_1448);
nand U2760 (N_2760,In_2887,In_672);
xnor U2761 (N_2761,In_1209,In_291);
and U2762 (N_2762,In_2135,In_1992);
xor U2763 (N_2763,In_220,In_2513);
or U2764 (N_2764,In_566,In_353);
and U2765 (N_2765,In_2680,In_967);
nor U2766 (N_2766,In_140,In_881);
or U2767 (N_2767,In_472,In_268);
xor U2768 (N_2768,In_1162,In_777);
xnor U2769 (N_2769,In_1021,In_705);
nor U2770 (N_2770,In_1635,In_813);
or U2771 (N_2771,In_2654,In_2342);
nand U2772 (N_2772,In_795,In_2997);
xor U2773 (N_2773,In_920,In_2934);
or U2774 (N_2774,In_1986,In_409);
or U2775 (N_2775,In_823,In_147);
nor U2776 (N_2776,In_985,In_243);
and U2777 (N_2777,In_68,In_845);
nand U2778 (N_2778,In_1004,In_37);
and U2779 (N_2779,In_735,In_1685);
nand U2780 (N_2780,In_790,In_1838);
xnor U2781 (N_2781,In_1218,In_2247);
or U2782 (N_2782,In_2847,In_112);
and U2783 (N_2783,In_382,In_2465);
or U2784 (N_2784,In_2947,In_1436);
xnor U2785 (N_2785,In_121,In_1485);
xnor U2786 (N_2786,In_2295,In_812);
nand U2787 (N_2787,In_1890,In_2898);
and U2788 (N_2788,In_543,In_2422);
nor U2789 (N_2789,In_1255,In_108);
or U2790 (N_2790,In_881,In_1095);
and U2791 (N_2791,In_226,In_503);
and U2792 (N_2792,In_2595,In_934);
nor U2793 (N_2793,In_1017,In_2108);
xor U2794 (N_2794,In_1441,In_764);
nand U2795 (N_2795,In_323,In_2521);
and U2796 (N_2796,In_1214,In_2936);
and U2797 (N_2797,In_2256,In_1932);
nor U2798 (N_2798,In_628,In_2671);
xor U2799 (N_2799,In_627,In_2824);
or U2800 (N_2800,In_897,In_2372);
xnor U2801 (N_2801,In_2717,In_2037);
or U2802 (N_2802,In_1457,In_869);
nor U2803 (N_2803,In_733,In_948);
or U2804 (N_2804,In_2504,In_836);
nor U2805 (N_2805,In_150,In_1519);
or U2806 (N_2806,In_1508,In_2006);
xor U2807 (N_2807,In_163,In_2385);
nor U2808 (N_2808,In_1259,In_2967);
nand U2809 (N_2809,In_2787,In_1783);
nor U2810 (N_2810,In_2356,In_409);
and U2811 (N_2811,In_811,In_102);
or U2812 (N_2812,In_1891,In_601);
and U2813 (N_2813,In_2924,In_2956);
and U2814 (N_2814,In_2817,In_715);
nand U2815 (N_2815,In_1612,In_1071);
and U2816 (N_2816,In_545,In_169);
nand U2817 (N_2817,In_595,In_1730);
nand U2818 (N_2818,In_716,In_830);
or U2819 (N_2819,In_780,In_932);
or U2820 (N_2820,In_2273,In_631);
xnor U2821 (N_2821,In_219,In_953);
nand U2822 (N_2822,In_2806,In_81);
or U2823 (N_2823,In_971,In_232);
nor U2824 (N_2824,In_1665,In_2807);
or U2825 (N_2825,In_307,In_2806);
and U2826 (N_2826,In_258,In_1073);
and U2827 (N_2827,In_835,In_344);
nand U2828 (N_2828,In_776,In_2208);
or U2829 (N_2829,In_2207,In_416);
nor U2830 (N_2830,In_2064,In_1688);
nor U2831 (N_2831,In_173,In_2544);
xnor U2832 (N_2832,In_2401,In_1117);
or U2833 (N_2833,In_556,In_2552);
and U2834 (N_2834,In_1822,In_147);
nor U2835 (N_2835,In_2652,In_1055);
nor U2836 (N_2836,In_2773,In_2704);
or U2837 (N_2837,In_2618,In_2383);
and U2838 (N_2838,In_277,In_912);
nand U2839 (N_2839,In_498,In_1903);
or U2840 (N_2840,In_2090,In_2469);
xor U2841 (N_2841,In_2420,In_1404);
or U2842 (N_2842,In_1434,In_2905);
and U2843 (N_2843,In_1936,In_1701);
nand U2844 (N_2844,In_173,In_1757);
or U2845 (N_2845,In_1459,In_1606);
nor U2846 (N_2846,In_2031,In_693);
nand U2847 (N_2847,In_1754,In_2026);
and U2848 (N_2848,In_2692,In_1014);
xor U2849 (N_2849,In_2428,In_312);
xnor U2850 (N_2850,In_517,In_999);
nor U2851 (N_2851,In_571,In_2758);
and U2852 (N_2852,In_2560,In_2802);
and U2853 (N_2853,In_1113,In_448);
xor U2854 (N_2854,In_2032,In_1505);
nand U2855 (N_2855,In_1480,In_876);
and U2856 (N_2856,In_905,In_2010);
xor U2857 (N_2857,In_2606,In_454);
nor U2858 (N_2858,In_2524,In_2969);
nor U2859 (N_2859,In_1881,In_466);
xor U2860 (N_2860,In_2431,In_2965);
xor U2861 (N_2861,In_1321,In_2882);
nor U2862 (N_2862,In_905,In_764);
and U2863 (N_2863,In_2940,In_2147);
nor U2864 (N_2864,In_2802,In_402);
or U2865 (N_2865,In_660,In_1798);
nand U2866 (N_2866,In_2458,In_1598);
nor U2867 (N_2867,In_2844,In_2634);
nand U2868 (N_2868,In_300,In_883);
xnor U2869 (N_2869,In_2206,In_2771);
nand U2870 (N_2870,In_1216,In_2088);
nor U2871 (N_2871,In_962,In_1051);
or U2872 (N_2872,In_1389,In_288);
xnor U2873 (N_2873,In_2955,In_1883);
and U2874 (N_2874,In_933,In_2383);
nor U2875 (N_2875,In_1905,In_2282);
xnor U2876 (N_2876,In_1232,In_1802);
nor U2877 (N_2877,In_129,In_1844);
nand U2878 (N_2878,In_999,In_1041);
nand U2879 (N_2879,In_1070,In_2487);
and U2880 (N_2880,In_1292,In_1376);
nor U2881 (N_2881,In_1734,In_2229);
or U2882 (N_2882,In_1622,In_1537);
nand U2883 (N_2883,In_2361,In_2140);
nor U2884 (N_2884,In_1462,In_443);
xnor U2885 (N_2885,In_772,In_2099);
xnor U2886 (N_2886,In_855,In_1616);
xor U2887 (N_2887,In_2236,In_2585);
or U2888 (N_2888,In_63,In_216);
and U2889 (N_2889,In_800,In_1219);
and U2890 (N_2890,In_1776,In_76);
xnor U2891 (N_2891,In_1174,In_2384);
and U2892 (N_2892,In_1383,In_1208);
nor U2893 (N_2893,In_2236,In_2728);
xnor U2894 (N_2894,In_274,In_2354);
and U2895 (N_2895,In_88,In_885);
or U2896 (N_2896,In_93,In_1976);
nand U2897 (N_2897,In_101,In_2535);
or U2898 (N_2898,In_1922,In_98);
xor U2899 (N_2899,In_1147,In_1862);
xnor U2900 (N_2900,In_1983,In_419);
nor U2901 (N_2901,In_1247,In_2640);
xor U2902 (N_2902,In_1835,In_684);
or U2903 (N_2903,In_1355,In_2336);
or U2904 (N_2904,In_2027,In_2231);
and U2905 (N_2905,In_2844,In_1823);
and U2906 (N_2906,In_1284,In_233);
xor U2907 (N_2907,In_808,In_414);
nand U2908 (N_2908,In_2856,In_717);
xor U2909 (N_2909,In_783,In_738);
nor U2910 (N_2910,In_1291,In_677);
or U2911 (N_2911,In_199,In_685);
nor U2912 (N_2912,In_540,In_1574);
nand U2913 (N_2913,In_627,In_899);
or U2914 (N_2914,In_1638,In_34);
nand U2915 (N_2915,In_2202,In_397);
nor U2916 (N_2916,In_2673,In_487);
nor U2917 (N_2917,In_324,In_260);
or U2918 (N_2918,In_1274,In_1617);
xnor U2919 (N_2919,In_405,In_731);
and U2920 (N_2920,In_1755,In_749);
or U2921 (N_2921,In_919,In_2452);
and U2922 (N_2922,In_1180,In_1748);
xor U2923 (N_2923,In_1702,In_435);
and U2924 (N_2924,In_2576,In_1571);
and U2925 (N_2925,In_796,In_1802);
and U2926 (N_2926,In_589,In_1033);
nand U2927 (N_2927,In_1886,In_466);
nor U2928 (N_2928,In_897,In_344);
nand U2929 (N_2929,In_2295,In_163);
or U2930 (N_2930,In_752,In_2646);
xor U2931 (N_2931,In_2297,In_704);
nor U2932 (N_2932,In_2643,In_2225);
nand U2933 (N_2933,In_24,In_130);
nand U2934 (N_2934,In_2065,In_1655);
nand U2935 (N_2935,In_1952,In_2322);
or U2936 (N_2936,In_2081,In_2823);
nor U2937 (N_2937,In_1180,In_2433);
nor U2938 (N_2938,In_1915,In_2402);
and U2939 (N_2939,In_2676,In_360);
nand U2940 (N_2940,In_270,In_132);
nor U2941 (N_2941,In_1150,In_1816);
nor U2942 (N_2942,In_2045,In_1729);
nor U2943 (N_2943,In_348,In_2661);
xor U2944 (N_2944,In_2641,In_824);
nand U2945 (N_2945,In_1259,In_1018);
and U2946 (N_2946,In_848,In_2037);
nor U2947 (N_2947,In_1141,In_1174);
nor U2948 (N_2948,In_2935,In_2477);
or U2949 (N_2949,In_382,In_1867);
and U2950 (N_2950,In_2383,In_339);
or U2951 (N_2951,In_1447,In_2092);
and U2952 (N_2952,In_242,In_254);
nand U2953 (N_2953,In_2959,In_152);
nor U2954 (N_2954,In_1233,In_557);
nor U2955 (N_2955,In_452,In_951);
nor U2956 (N_2956,In_1511,In_1512);
and U2957 (N_2957,In_706,In_624);
nor U2958 (N_2958,In_535,In_1101);
nor U2959 (N_2959,In_144,In_979);
nor U2960 (N_2960,In_118,In_484);
nor U2961 (N_2961,In_1064,In_2976);
nor U2962 (N_2962,In_2826,In_2331);
xor U2963 (N_2963,In_1407,In_1675);
and U2964 (N_2964,In_2229,In_1003);
and U2965 (N_2965,In_1371,In_1330);
xor U2966 (N_2966,In_1907,In_603);
or U2967 (N_2967,In_367,In_2286);
xnor U2968 (N_2968,In_957,In_1092);
xor U2969 (N_2969,In_1982,In_63);
xor U2970 (N_2970,In_1827,In_2830);
and U2971 (N_2971,In_35,In_314);
nor U2972 (N_2972,In_1286,In_747);
xnor U2973 (N_2973,In_81,In_1890);
nor U2974 (N_2974,In_459,In_1537);
nor U2975 (N_2975,In_2089,In_1023);
xnor U2976 (N_2976,In_2635,In_2857);
and U2977 (N_2977,In_2308,In_930);
and U2978 (N_2978,In_2583,In_806);
xnor U2979 (N_2979,In_308,In_2316);
xnor U2980 (N_2980,In_1322,In_1680);
nor U2981 (N_2981,In_172,In_2958);
nand U2982 (N_2982,In_1271,In_328);
and U2983 (N_2983,In_133,In_1972);
xor U2984 (N_2984,In_2090,In_978);
and U2985 (N_2985,In_1003,In_1041);
nand U2986 (N_2986,In_1812,In_354);
nor U2987 (N_2987,In_2620,In_1402);
nor U2988 (N_2988,In_862,In_29);
xor U2989 (N_2989,In_1083,In_1015);
nand U2990 (N_2990,In_1262,In_431);
nor U2991 (N_2991,In_2644,In_1849);
and U2992 (N_2992,In_50,In_526);
and U2993 (N_2993,In_1744,In_2789);
or U2994 (N_2994,In_1239,In_2703);
nor U2995 (N_2995,In_1964,In_2347);
xor U2996 (N_2996,In_536,In_2803);
nand U2997 (N_2997,In_134,In_2783);
and U2998 (N_2998,In_759,In_2336);
nor U2999 (N_2999,In_306,In_926);
nand U3000 (N_3000,N_1712,N_1861);
or U3001 (N_3001,N_2222,N_933);
or U3002 (N_3002,N_2166,N_2826);
and U3003 (N_3003,N_2308,N_1073);
nor U3004 (N_3004,N_1442,N_1935);
xnor U3005 (N_3005,N_2515,N_1584);
and U3006 (N_3006,N_1688,N_2824);
or U3007 (N_3007,N_132,N_1803);
nor U3008 (N_3008,N_974,N_387);
or U3009 (N_3009,N_1109,N_1618);
or U3010 (N_3010,N_2958,N_2794);
and U3011 (N_3011,N_2013,N_1387);
and U3012 (N_3012,N_1320,N_1280);
or U3013 (N_3013,N_2056,N_1605);
xor U3014 (N_3014,N_2366,N_2118);
and U3015 (N_3015,N_491,N_1385);
or U3016 (N_3016,N_547,N_2832);
and U3017 (N_3017,N_2537,N_1922);
xnor U3018 (N_3018,N_1526,N_347);
or U3019 (N_3019,N_668,N_2005);
xor U3020 (N_3020,N_2564,N_1423);
or U3021 (N_3021,N_736,N_1431);
or U3022 (N_3022,N_1613,N_1382);
nand U3023 (N_3023,N_879,N_1196);
and U3024 (N_3024,N_1041,N_499);
or U3025 (N_3025,N_613,N_232);
nor U3026 (N_3026,N_1979,N_774);
xor U3027 (N_3027,N_792,N_2018);
and U3028 (N_3028,N_2187,N_1198);
or U3029 (N_3029,N_689,N_2896);
xnor U3030 (N_3030,N_766,N_1507);
nand U3031 (N_3031,N_409,N_2230);
xnor U3032 (N_3032,N_1728,N_2511);
xnor U3033 (N_3033,N_1469,N_399);
or U3034 (N_3034,N_2711,N_2943);
and U3035 (N_3035,N_2531,N_684);
nand U3036 (N_3036,N_1181,N_2120);
nand U3037 (N_3037,N_2545,N_847);
nand U3038 (N_3038,N_2093,N_1800);
and U3039 (N_3039,N_1975,N_1719);
nand U3040 (N_3040,N_1790,N_1833);
or U3041 (N_3041,N_1404,N_1807);
xnor U3042 (N_3042,N_75,N_1380);
nor U3043 (N_3043,N_1889,N_1984);
or U3044 (N_3044,N_382,N_1753);
or U3045 (N_3045,N_640,N_2264);
nor U3046 (N_3046,N_2393,N_2940);
nand U3047 (N_3047,N_997,N_1437);
and U3048 (N_3048,N_2936,N_1053);
nand U3049 (N_3049,N_1286,N_2052);
xor U3050 (N_3050,N_200,N_964);
and U3051 (N_3051,N_1251,N_1815);
nor U3052 (N_3052,N_2612,N_26);
nand U3053 (N_3053,N_2575,N_1106);
nor U3054 (N_3054,N_1457,N_1313);
and U3055 (N_3055,N_1042,N_2599);
or U3056 (N_3056,N_864,N_2695);
or U3057 (N_3057,N_2977,N_809);
and U3058 (N_3058,N_2781,N_811);
and U3059 (N_3059,N_2964,N_1865);
nor U3060 (N_3060,N_2050,N_1103);
nand U3061 (N_3061,N_561,N_2126);
nor U3062 (N_3062,N_1598,N_685);
and U3063 (N_3063,N_1119,N_2810);
or U3064 (N_3064,N_1545,N_2925);
nor U3065 (N_3065,N_1446,N_616);
or U3066 (N_3066,N_2967,N_1377);
nand U3067 (N_3067,N_23,N_2779);
and U3068 (N_3068,N_1642,N_2662);
xor U3069 (N_3069,N_1232,N_1187);
xor U3070 (N_3070,N_1152,N_1144);
and U3071 (N_3071,N_840,N_621);
nor U3072 (N_3072,N_487,N_2757);
and U3073 (N_3073,N_1600,N_1652);
nor U3074 (N_3074,N_832,N_2196);
xnor U3075 (N_3075,N_374,N_1905);
nor U3076 (N_3076,N_998,N_906);
or U3077 (N_3077,N_165,N_749);
and U3078 (N_3078,N_1947,N_1319);
nand U3079 (N_3079,N_496,N_1189);
xnor U3080 (N_3080,N_240,N_1099);
and U3081 (N_3081,N_89,N_167);
nand U3082 (N_3082,N_2540,N_1236);
nand U3083 (N_3083,N_1562,N_464);
or U3084 (N_3084,N_1468,N_2233);
nor U3085 (N_3085,N_1915,N_492);
xnor U3086 (N_3086,N_1448,N_2414);
xnor U3087 (N_3087,N_1764,N_1250);
or U3088 (N_3088,N_451,N_803);
xor U3089 (N_3089,N_1765,N_897);
and U3090 (N_3090,N_1130,N_1341);
nor U3091 (N_3091,N_1031,N_204);
xor U3092 (N_3092,N_2706,N_2415);
xor U3093 (N_3093,N_597,N_397);
and U3094 (N_3094,N_131,N_618);
nor U3095 (N_3095,N_1517,N_2494);
xor U3096 (N_3096,N_2541,N_406);
and U3097 (N_3097,N_2316,N_1116);
nand U3098 (N_3098,N_2817,N_2270);
nor U3099 (N_3099,N_1410,N_1497);
or U3100 (N_3100,N_914,N_2804);
or U3101 (N_3101,N_2713,N_793);
xor U3102 (N_3102,N_1824,N_77);
and U3103 (N_3103,N_2960,N_256);
xnor U3104 (N_3104,N_2950,N_1994);
and U3105 (N_3105,N_1773,N_57);
or U3106 (N_3106,N_291,N_1972);
nor U3107 (N_3107,N_1316,N_748);
xnor U3108 (N_3108,N_1756,N_432);
and U3109 (N_3109,N_485,N_1893);
xor U3110 (N_3110,N_2199,N_1619);
and U3111 (N_3111,N_2178,N_2948);
and U3112 (N_3112,N_1094,N_1669);
nand U3113 (N_3113,N_817,N_1456);
nand U3114 (N_3114,N_140,N_2659);
nor U3115 (N_3115,N_2693,N_2190);
nand U3116 (N_3116,N_959,N_656);
nor U3117 (N_3117,N_2933,N_151);
nor U3118 (N_3118,N_13,N_110);
or U3119 (N_3119,N_2859,N_2402);
xnor U3120 (N_3120,N_296,N_206);
or U3121 (N_3121,N_1681,N_1911);
xor U3122 (N_3122,N_1447,N_521);
or U3123 (N_3123,N_437,N_2150);
or U3124 (N_3124,N_545,N_2866);
and U3125 (N_3125,N_1230,N_2040);
nand U3126 (N_3126,N_144,N_2800);
and U3127 (N_3127,N_377,N_290);
nor U3128 (N_3128,N_1853,N_2517);
nor U3129 (N_3129,N_677,N_2953);
nor U3130 (N_3130,N_1025,N_2888);
xor U3131 (N_3131,N_2766,N_2407);
nor U3132 (N_3132,N_642,N_960);
nand U3133 (N_3133,N_1943,N_842);
xor U3134 (N_3134,N_288,N_2247);
or U3135 (N_3135,N_1503,N_2821);
nand U3136 (N_3136,N_884,N_1542);
nor U3137 (N_3137,N_731,N_2136);
and U3138 (N_3138,N_2796,N_1019);
xor U3139 (N_3139,N_1967,N_2700);
or U3140 (N_3140,N_2828,N_2176);
nand U3141 (N_3141,N_1521,N_1259);
nor U3142 (N_3142,N_693,N_1100);
or U3143 (N_3143,N_2211,N_572);
xnor U3144 (N_3144,N_976,N_135);
nor U3145 (N_3145,N_41,N_130);
or U3146 (N_3146,N_761,N_1817);
nand U3147 (N_3147,N_2142,N_1916);
or U3148 (N_3148,N_2401,N_367);
nand U3149 (N_3149,N_1030,N_1634);
and U3150 (N_3150,N_2219,N_1869);
nand U3151 (N_3151,N_1878,N_1485);
nor U3152 (N_3152,N_791,N_2942);
nor U3153 (N_3153,N_1034,N_1586);
xor U3154 (N_3154,N_2974,N_8);
xnor U3155 (N_3155,N_2084,N_2356);
and U3156 (N_3156,N_423,N_2555);
nor U3157 (N_3157,N_1304,N_2727);
nand U3158 (N_3158,N_2076,N_546);
or U3159 (N_3159,N_2019,N_1093);
nor U3160 (N_3160,N_2482,N_401);
xor U3161 (N_3161,N_2111,N_703);
nor U3162 (N_3162,N_862,N_2636);
nor U3163 (N_3163,N_2945,N_695);
or U3164 (N_3164,N_2582,N_2554);
nand U3165 (N_3165,N_2444,N_2914);
nand U3166 (N_3166,N_1327,N_1964);
or U3167 (N_3167,N_2365,N_2512);
or U3168 (N_3168,N_501,N_1996);
nor U3169 (N_3169,N_2472,N_2637);
nor U3170 (N_3170,N_2294,N_1338);
xnor U3171 (N_3171,N_829,N_1062);
nand U3172 (N_3172,N_1257,N_1283);
nand U3173 (N_3173,N_539,N_512);
and U3174 (N_3174,N_1705,N_1139);
nand U3175 (N_3175,N_2218,N_529);
or U3176 (N_3176,N_2091,N_2073);
nand U3177 (N_3177,N_2742,N_2969);
or U3178 (N_3178,N_2855,N_602);
xor U3179 (N_3179,N_405,N_541);
or U3180 (N_3180,N_2321,N_1054);
nand U3181 (N_3181,N_567,N_2317);
nor U3182 (N_3182,N_2788,N_152);
and U3183 (N_3183,N_1581,N_1427);
or U3184 (N_3184,N_1298,N_161);
xnor U3185 (N_3185,N_1604,N_1300);
and U3186 (N_3186,N_2231,N_1394);
or U3187 (N_3187,N_2115,N_2453);
nor U3188 (N_3188,N_2207,N_73);
nand U3189 (N_3189,N_885,N_1510);
and U3190 (N_3190,N_1822,N_944);
xor U3191 (N_3191,N_2849,N_883);
and U3192 (N_3192,N_2476,N_1081);
nor U3193 (N_3193,N_1247,N_648);
nor U3194 (N_3194,N_538,N_2372);
nand U3195 (N_3195,N_2499,N_1347);
nor U3196 (N_3196,N_2023,N_1021);
nand U3197 (N_3197,N_1265,N_500);
or U3198 (N_3198,N_2216,N_138);
xnor U3199 (N_3199,N_1525,N_1527);
nand U3200 (N_3200,N_1821,N_2623);
or U3201 (N_3201,N_1571,N_908);
or U3202 (N_3202,N_1848,N_2833);
xor U3203 (N_3203,N_1621,N_1176);
nor U3204 (N_3204,N_634,N_1675);
nand U3205 (N_3205,N_1594,N_2615);
xnor U3206 (N_3206,N_143,N_1593);
or U3207 (N_3207,N_969,N_860);
nand U3208 (N_3208,N_2851,N_1723);
nand U3209 (N_3209,N_2744,N_2431);
nor U3210 (N_3210,N_315,N_2962);
nand U3211 (N_3211,N_2139,N_35);
or U3212 (N_3212,N_1488,N_2085);
and U3213 (N_3213,N_1095,N_1227);
or U3214 (N_3214,N_318,N_261);
nand U3215 (N_3215,N_556,N_1234);
or U3216 (N_3216,N_2813,N_2333);
nor U3217 (N_3217,N_156,N_72);
nand U3218 (N_3218,N_1684,N_579);
nor U3219 (N_3219,N_1412,N_2310);
xnor U3220 (N_3220,N_1355,N_1885);
nor U3221 (N_3221,N_2376,N_1046);
nand U3222 (N_3222,N_2437,N_394);
nand U3223 (N_3223,N_2456,N_54);
and U3224 (N_3224,N_963,N_566);
nand U3225 (N_3225,N_623,N_452);
nand U3226 (N_3226,N_2236,N_1160);
and U3227 (N_3227,N_1153,N_365);
nand U3228 (N_3228,N_2524,N_818);
nor U3229 (N_3229,N_497,N_1059);
nor U3230 (N_3230,N_2463,N_2282);
or U3231 (N_3231,N_2957,N_2811);
nor U3232 (N_3232,N_2138,N_2075);
nor U3233 (N_3233,N_2159,N_558);
xnor U3234 (N_3234,N_51,N_229);
xnor U3235 (N_3235,N_84,N_1577);
xor U3236 (N_3236,N_1354,N_1069);
nand U3237 (N_3237,N_2055,N_1532);
xnor U3238 (N_3238,N_543,N_475);
nand U3239 (N_3239,N_308,N_2065);
nor U3240 (N_3240,N_1426,N_2635);
nand U3241 (N_3241,N_1462,N_1262);
and U3242 (N_3242,N_2587,N_671);
nand U3243 (N_3243,N_734,N_2217);
nor U3244 (N_3244,N_2568,N_804);
and U3245 (N_3245,N_2507,N_1284);
nor U3246 (N_3246,N_276,N_2751);
nor U3247 (N_3247,N_1435,N_1246);
xnor U3248 (N_3248,N_2227,N_776);
and U3249 (N_3249,N_2323,N_858);
and U3250 (N_3250,N_2956,N_1311);
or U3251 (N_3251,N_834,N_2736);
xnor U3252 (N_3252,N_21,N_1209);
and U3253 (N_3253,N_2273,N_590);
nand U3254 (N_3254,N_2763,N_1074);
nor U3255 (N_3255,N_246,N_1886);
nor U3256 (N_3256,N_1292,N_18);
nand U3257 (N_3257,N_641,N_2307);
nor U3258 (N_3258,N_248,N_1750);
or U3259 (N_3259,N_2123,N_346);
nand U3260 (N_3260,N_2949,N_662);
nor U3261 (N_3261,N_2860,N_2006);
nand U3262 (N_3262,N_1294,N_19);
or U3263 (N_3263,N_444,N_852);
and U3264 (N_3264,N_923,N_304);
and U3265 (N_3265,N_2331,N_1709);
nor U3266 (N_3266,N_714,N_2926);
or U3267 (N_3267,N_1482,N_2262);
nand U3268 (N_3268,N_2593,N_869);
or U3269 (N_3269,N_50,N_2899);
nand U3270 (N_3270,N_1249,N_905);
nor U3271 (N_3271,N_956,N_1459);
xnor U3272 (N_3272,N_1882,N_1067);
nor U3273 (N_3273,N_1986,N_1992);
nand U3274 (N_3274,N_2080,N_2816);
xor U3275 (N_3275,N_2108,N_2296);
xor U3276 (N_3276,N_2732,N_920);
nand U3277 (N_3277,N_2750,N_509);
nand U3278 (N_3278,N_939,N_989);
and U3279 (N_3279,N_2382,N_163);
nor U3280 (N_3280,N_1540,N_183);
and U3281 (N_3281,N_2028,N_238);
and U3282 (N_3282,N_767,N_2666);
xor U3283 (N_3283,N_510,N_478);
or U3284 (N_3284,N_1453,N_392);
nand U3285 (N_3285,N_2480,N_1832);
or U3286 (N_3286,N_1364,N_1504);
nand U3287 (N_3287,N_2092,N_2867);
xnor U3288 (N_3288,N_2137,N_1474);
and U3289 (N_3289,N_220,N_626);
nor U3290 (N_3290,N_148,N_1239);
xnor U3291 (N_3291,N_342,N_1818);
xor U3292 (N_3292,N_1836,N_239);
or U3293 (N_3293,N_2398,N_2586);
nor U3294 (N_3294,N_2761,N_1721);
or U3295 (N_3295,N_861,N_2206);
and U3296 (N_3296,N_1786,N_1625);
or U3297 (N_3297,N_2620,N_350);
and U3298 (N_3298,N_195,N_81);
nand U3299 (N_3299,N_2889,N_1299);
nor U3300 (N_3300,N_1923,N_1666);
or U3301 (N_3301,N_559,N_2753);
nand U3302 (N_3302,N_1976,N_585);
nand U3303 (N_3303,N_787,N_1151);
xor U3304 (N_3304,N_2493,N_1509);
and U3305 (N_3305,N_1702,N_1658);
xor U3306 (N_3306,N_2959,N_2058);
nor U3307 (N_3307,N_713,N_210);
nand U3308 (N_3308,N_1508,N_985);
nand U3309 (N_3309,N_786,N_2876);
nand U3310 (N_3310,N_754,N_2525);
nor U3311 (N_3311,N_2772,N_2773);
nor U3312 (N_3312,N_1700,N_2184);
nor U3313 (N_3313,N_463,N_2634);
and U3314 (N_3314,N_2213,N_2681);
xor U3315 (N_3315,N_42,N_1543);
and U3316 (N_3316,N_65,N_1252);
nand U3317 (N_3317,N_2991,N_790);
and U3318 (N_3318,N_527,N_80);
nor U3319 (N_3319,N_2968,N_1632);
nor U3320 (N_3320,N_768,N_63);
and U3321 (N_3321,N_1438,N_2172);
nor U3322 (N_3322,N_2117,N_2355);
nand U3323 (N_3323,N_1724,N_1443);
nor U3324 (N_3324,N_2007,N_353);
nor U3325 (N_3325,N_214,N_1798);
and U3326 (N_3326,N_1293,N_2924);
nand U3327 (N_3327,N_1592,N_2601);
or U3328 (N_3328,N_1463,N_1432);
nand U3329 (N_3329,N_106,N_1961);
and U3330 (N_3330,N_1999,N_1129);
nor U3331 (N_3331,N_87,N_1607);
and U3332 (N_3332,N_1133,N_1221);
xor U3333 (N_3333,N_2938,N_1258);
xor U3334 (N_3334,N_800,N_1413);
or U3335 (N_3335,N_596,N_2526);
or U3336 (N_3336,N_870,N_863);
and U3337 (N_3337,N_2687,N_1809);
and U3338 (N_3338,N_2265,N_2992);
and U3339 (N_3339,N_2379,N_2716);
or U3340 (N_3340,N_719,N_854);
nor U3341 (N_3341,N_2034,N_332);
xor U3342 (N_3342,N_617,N_986);
nand U3343 (N_3343,N_343,N_789);
and U3344 (N_3344,N_1868,N_357);
or U3345 (N_3345,N_2774,N_2975);
xnor U3346 (N_3346,N_917,N_941);
nand U3347 (N_3347,N_1222,N_1194);
nand U3348 (N_3348,N_1157,N_1348);
and U3349 (N_3349,N_1216,N_2677);
xor U3350 (N_3350,N_609,N_218);
or U3351 (N_3351,N_1963,N_1203);
and U3352 (N_3352,N_2679,N_1623);
nand U3353 (N_3353,N_1883,N_1726);
or U3354 (N_3354,N_1585,N_2543);
nor U3355 (N_3355,N_2424,N_1396);
nand U3356 (N_3356,N_2802,N_2605);
and U3357 (N_3357,N_781,N_1378);
or U3358 (N_3358,N_1927,N_2647);
xor U3359 (N_3359,N_2078,N_2303);
nand U3360 (N_3360,N_796,N_1450);
nor U3361 (N_3361,N_937,N_1012);
and U3362 (N_3362,N_711,N_1941);
xor U3363 (N_3363,N_275,N_2200);
nand U3364 (N_3364,N_2897,N_1148);
xnor U3365 (N_3365,N_1601,N_1372);
and U3366 (N_3366,N_524,N_1890);
nand U3367 (N_3367,N_1091,N_1624);
nor U3368 (N_3368,N_2249,N_2253);
nor U3369 (N_3369,N_1391,N_2237);
and U3370 (N_3370,N_1329,N_1622);
nand U3371 (N_3371,N_2739,N_1971);
and U3372 (N_3372,N_2468,N_2251);
and U3373 (N_3373,N_2286,N_2894);
nand U3374 (N_3374,N_563,N_1210);
nor U3375 (N_3375,N_1027,N_1774);
and U3376 (N_3376,N_1529,N_1533);
nand U3377 (N_3377,N_273,N_2892);
nand U3378 (N_3378,N_515,N_856);
xnor U3379 (N_3379,N_1872,N_1495);
and U3380 (N_3380,N_822,N_2557);
xnor U3381 (N_3381,N_2399,N_2426);
xnor U3382 (N_3382,N_1352,N_2151);
or U3383 (N_3383,N_853,N_755);
nand U3384 (N_3384,N_310,N_7);
xor U3385 (N_3385,N_2429,N_1627);
nand U3386 (N_3386,N_2241,N_2010);
and U3387 (N_3387,N_2754,N_1989);
or U3388 (N_3388,N_2565,N_2322);
and U3389 (N_3389,N_2054,N_333);
or U3390 (N_3390,N_1796,N_1309);
or U3391 (N_3391,N_1858,N_1661);
or U3392 (N_3392,N_2063,N_2539);
or U3393 (N_3393,N_359,N_2931);
xnor U3394 (N_3394,N_1939,N_1717);
nor U3395 (N_3395,N_1820,N_1184);
xnor U3396 (N_3396,N_368,N_369);
nor U3397 (N_3397,N_2168,N_1128);
nand U3398 (N_3398,N_2442,N_201);
and U3399 (N_3399,N_1070,N_867);
and U3400 (N_3400,N_2629,N_661);
or U3401 (N_3401,N_1180,N_1155);
xnor U3402 (N_3402,N_2884,N_1193);
xor U3403 (N_3403,N_1557,N_1659);
nor U3404 (N_3404,N_2342,N_1914);
nor U3405 (N_3405,N_2795,N_1754);
or U3406 (N_3406,N_1743,N_2371);
nand U3407 (N_3407,N_2096,N_1114);
and U3408 (N_3408,N_2287,N_830);
and U3409 (N_3409,N_1548,N_2721);
and U3410 (N_3410,N_2246,N_1272);
nor U3411 (N_3411,N_922,N_2595);
and U3412 (N_3412,N_20,N_2302);
nor U3413 (N_3413,N_1780,N_2728);
nor U3414 (N_3414,N_1146,N_2209);
nand U3415 (N_3415,N_1425,N_2986);
xnor U3416 (N_3416,N_2809,N_2069);
or U3417 (N_3417,N_1932,N_101);
and U3418 (N_3418,N_172,N_812);
xnor U3419 (N_3419,N_2141,N_2718);
and U3420 (N_3420,N_1860,N_2979);
nor U3421 (N_3421,N_253,N_2818);
nor U3422 (N_3422,N_2250,N_2907);
nor U3423 (N_3423,N_1710,N_2027);
and U3424 (N_3424,N_2223,N_913);
or U3425 (N_3425,N_2970,N_1925);
nand U3426 (N_3426,N_433,N_2893);
or U3427 (N_3427,N_270,N_1268);
and U3428 (N_3428,N_580,N_780);
nor U3429 (N_3429,N_1863,N_1064);
xnor U3430 (N_3430,N_2192,N_2664);
and U3431 (N_3431,N_1711,N_2153);
nor U3432 (N_3432,N_2838,N_1206);
nor U3433 (N_3433,N_2737,N_2983);
or U3434 (N_3434,N_436,N_486);
nand U3435 (N_3435,N_2961,N_875);
and U3436 (N_3436,N_1223,N_1930);
and U3437 (N_3437,N_2835,N_1703);
and U3438 (N_3438,N_1839,N_660);
nand U3439 (N_3439,N_2697,N_64);
nor U3440 (N_3440,N_2394,N_1770);
nor U3441 (N_3441,N_2709,N_871);
and U3442 (N_3442,N_1403,N_213);
nand U3443 (N_3443,N_2690,N_1016);
nand U3444 (N_3444,N_1841,N_1475);
xor U3445 (N_3445,N_2090,N_657);
and U3446 (N_3446,N_1440,N_980);
xor U3447 (N_3447,N_2848,N_2457);
and U3448 (N_3448,N_2361,N_2665);
xor U3449 (N_3449,N_476,N_1536);
nand U3450 (N_3450,N_1047,N_12);
nand U3451 (N_3451,N_1955,N_141);
and U3452 (N_3452,N_1814,N_1043);
nor U3453 (N_3453,N_1940,N_1813);
or U3454 (N_3454,N_2688,N_2416);
nor U3455 (N_3455,N_469,N_2145);
nor U3456 (N_3456,N_355,N_2783);
nand U3457 (N_3457,N_231,N_1125);
or U3458 (N_3458,N_1639,N_2806);
or U3459 (N_3459,N_2592,N_2127);
xor U3460 (N_3460,N_1359,N_385);
xnor U3461 (N_3461,N_1416,N_2060);
or U3462 (N_3462,N_1386,N_297);
and U3463 (N_3463,N_1892,N_1720);
nor U3464 (N_3464,N_209,N_582);
nor U3465 (N_3465,N_203,N_2167);
nor U3466 (N_3466,N_2022,N_225);
and U3467 (N_3467,N_2715,N_2895);
nand U3468 (N_3468,N_2067,N_345);
or U3469 (N_3469,N_1910,N_358);
and U3470 (N_3470,N_1350,N_1217);
nor U3471 (N_3471,N_1240,N_1178);
xor U3472 (N_3472,N_877,N_542);
or U3473 (N_3473,N_197,N_705);
and U3474 (N_3474,N_32,N_1334);
or U3475 (N_3475,N_1086,N_2608);
xnor U3476 (N_3476,N_321,N_2485);
or U3477 (N_3477,N_1270,N_1875);
nand U3478 (N_3478,N_785,N_2692);
or U3479 (N_3479,N_1077,N_1797);
nor U3480 (N_3480,N_2584,N_395);
nand U3481 (N_3481,N_1235,N_993);
nand U3482 (N_3482,N_772,N_2663);
or U3483 (N_3483,N_943,N_709);
nor U3484 (N_3484,N_2822,N_1375);
and U3485 (N_3485,N_1037,N_1212);
or U3486 (N_3486,N_2850,N_2104);
xor U3487 (N_3487,N_2489,N_2102);
nor U3488 (N_3488,N_707,N_1127);
and U3489 (N_3489,N_931,N_743);
nor U3490 (N_3490,N_2182,N_1161);
nor U3491 (N_3491,N_1722,N_483);
nand U3492 (N_3492,N_1757,N_1225);
xnor U3493 (N_3493,N_2505,N_2455);
nand U3494 (N_3494,N_1366,N_2865);
nor U3495 (N_3495,N_302,N_2406);
xor U3496 (N_3496,N_571,N_2973);
and U3497 (N_3497,N_2724,N_1897);
nand U3498 (N_3498,N_2735,N_1260);
and U3499 (N_3499,N_1101,N_1145);
nand U3500 (N_3500,N_1969,N_2491);
nor U3501 (N_3501,N_1397,N_1523);
and U3502 (N_3502,N_1573,N_2955);
xnor U3503 (N_3503,N_2873,N_727);
and U3504 (N_3504,N_187,N_336);
nor U3505 (N_3505,N_1117,N_2459);
and U3506 (N_3506,N_2320,N_2644);
xnor U3507 (N_3507,N_925,N_857);
and U3508 (N_3508,N_1835,N_2281);
nand U3509 (N_3509,N_2173,N_921);
nand U3510 (N_3510,N_2645,N_1572);
xnor U3511 (N_3511,N_126,N_1881);
or U3512 (N_3512,N_2870,N_1501);
nand U3513 (N_3513,N_349,N_1358);
or U3514 (N_3514,N_978,N_2965);
xnor U3515 (N_3515,N_1179,N_1421);
nor U3516 (N_3516,N_2513,N_1670);
or U3517 (N_3517,N_2465,N_425);
xor U3518 (N_3518,N_362,N_2087);
or U3519 (N_3519,N_453,N_1379);
nor U3520 (N_3520,N_1657,N_1524);
and U3521 (N_3521,N_2238,N_179);
xnor U3522 (N_3522,N_967,N_2508);
nand U3523 (N_3523,N_667,N_1195);
or U3524 (N_3524,N_2392,N_2466);
and U3525 (N_3525,N_1906,N_954);
nor U3526 (N_3526,N_1531,N_1645);
and U3527 (N_3527,N_2312,N_718);
and U3528 (N_3528,N_257,N_1381);
nor U3529 (N_3529,N_2257,N_2439);
or U3530 (N_3530,N_522,N_2920);
nand U3531 (N_3531,N_977,N_1891);
and U3532 (N_3532,N_2003,N_2155);
nand U3533 (N_3533,N_2550,N_473);
and U3534 (N_3534,N_2882,N_2911);
xor U3535 (N_3535,N_2110,N_1748);
or U3536 (N_3536,N_1326,N_252);
xnor U3537 (N_3537,N_1401,N_265);
or U3538 (N_3538,N_1991,N_2883);
nor U3539 (N_3539,N_2755,N_2261);
or U3540 (N_3540,N_2352,N_1981);
xor U3541 (N_3541,N_1873,N_1331);
xnor U3542 (N_3542,N_2068,N_2083);
or U3543 (N_3543,N_1977,N_2169);
xnor U3544 (N_3544,N_27,N_1777);
and U3545 (N_3545,N_2617,N_2328);
nand U3546 (N_3546,N_278,N_250);
or U3547 (N_3547,N_174,N_182);
or U3548 (N_3548,N_1197,N_2288);
or U3549 (N_3549,N_957,N_2741);
nand U3550 (N_3550,N_987,N_716);
and U3551 (N_3551,N_2578,N_2135);
nand U3552 (N_3552,N_282,N_2497);
nand U3553 (N_3553,N_947,N_1570);
nor U3554 (N_3554,N_622,N_251);
xnor U3555 (N_3555,N_2191,N_983);
nand U3556 (N_3556,N_564,N_150);
xor U3557 (N_3557,N_1982,N_2639);
xnor U3558 (N_3558,N_1244,N_2864);
xor U3559 (N_3559,N_324,N_1630);
nor U3560 (N_3560,N_940,N_1749);
or U3561 (N_3561,N_553,N_673);
or U3562 (N_3562,N_1328,N_109);
and U3563 (N_3563,N_1182,N_2396);
or U3564 (N_3564,N_619,N_262);
and U3565 (N_3565,N_1318,N_1392);
nor U3566 (N_3566,N_25,N_2919);
nand U3567 (N_3567,N_2079,N_1233);
nor U3568 (N_3568,N_891,N_850);
and U3569 (N_3569,N_872,N_1170);
xor U3570 (N_3570,N_2738,N_1097);
and U3571 (N_3571,N_1055,N_2613);
or U3572 (N_3572,N_2332,N_2904);
nor U3573 (N_3573,N_445,N_388);
and U3574 (N_3574,N_2343,N_1399);
or U3575 (N_3575,N_813,N_31);
xnor U3576 (N_3576,N_1778,N_2435);
nand U3577 (N_3577,N_10,N_2768);
nor U3578 (N_3578,N_2758,N_127);
nor U3579 (N_3579,N_1032,N_784);
xor U3580 (N_3580,N_71,N_119);
or U3581 (N_3581,N_1455,N_1199);
or U3582 (N_3582,N_1165,N_1422);
nor U3583 (N_3583,N_2450,N_2520);
nand U3584 (N_3584,N_2205,N_2988);
or U3585 (N_3585,N_2654,N_1900);
nor U3586 (N_3586,N_1200,N_2045);
nor U3587 (N_3587,N_91,N_975);
nor U3588 (N_3588,N_2387,N_1654);
nand U3589 (N_3589,N_2694,N_1599);
and U3590 (N_3590,N_142,N_2682);
nand U3591 (N_3591,N_2267,N_173);
nor U3592 (N_3592,N_2107,N_2720);
nand U3593 (N_3593,N_1691,N_752);
xor U3594 (N_3594,N_1275,N_1918);
xnor U3595 (N_3595,N_28,N_259);
and U3596 (N_3596,N_85,N_701);
nand U3597 (N_3597,N_2255,N_412);
or U3598 (N_3598,N_2419,N_2551);
xor U3599 (N_3599,N_2842,N_2852);
and U3600 (N_3600,N_2702,N_653);
nand U3601 (N_3601,N_2775,N_422);
and U3602 (N_3602,N_402,N_2917);
and U3603 (N_3603,N_2872,N_1776);
or U3604 (N_3604,N_86,N_1650);
xor U3605 (N_3605,N_2295,N_2131);
xnor U3606 (N_3606,N_2290,N_1384);
and U3607 (N_3607,N_1433,N_694);
xor U3608 (N_3608,N_1603,N_893);
nand U3609 (N_3609,N_525,N_1678);
xor U3610 (N_3610,N_2618,N_886);
nand U3611 (N_3611,N_981,N_1123);
and U3612 (N_3612,N_699,N_2843);
nor U3613 (N_3613,N_598,N_1278);
nand U3614 (N_3614,N_1802,N_2330);
and U3615 (N_3615,N_664,N_1306);
or U3616 (N_3616,N_788,N_2874);
or U3617 (N_3617,N_2935,N_228);
nand U3618 (N_3618,N_372,N_102);
nor U3619 (N_3619,N_2053,N_237);
and U3620 (N_3620,N_1132,N_2194);
or U3621 (N_3621,N_1357,N_1213);
or U3622 (N_3622,N_2861,N_1242);
nand U3623 (N_3623,N_2357,N_1395);
nand U3624 (N_3624,N_489,N_189);
and U3625 (N_3625,N_540,N_1002);
or U3626 (N_3626,N_593,N_1009);
and U3627 (N_3627,N_247,N_1732);
or U3628 (N_3628,N_2999,N_2051);
nor U3629 (N_3629,N_351,N_2641);
xor U3630 (N_3630,N_2204,N_1924);
and U3631 (N_3631,N_2015,N_1692);
nand U3632 (N_3632,N_769,N_1301);
or U3633 (N_3633,N_294,N_900);
and U3634 (N_3634,N_1725,N_697);
xor U3635 (N_3635,N_477,N_1502);
nand U3636 (N_3636,N_927,N_326);
or U3637 (N_3637,N_2600,N_2676);
or U3638 (N_3638,N_526,N_926);
nand U3639 (N_3639,N_95,N_2031);
or U3640 (N_3640,N_2650,N_2385);
nand U3641 (N_3641,N_777,N_407);
xnor U3642 (N_3642,N_1373,N_942);
and U3643 (N_3643,N_2912,N_894);
nor U3644 (N_3644,N_2916,N_435);
and U3645 (N_3645,N_2119,N_1274);
nand U3646 (N_3646,N_2981,N_160);
xnor U3647 (N_3647,N_122,N_1816);
nor U3648 (N_3648,N_2701,N_1111);
nor U3649 (N_3649,N_466,N_810);
or U3650 (N_3650,N_1574,N_2891);
xor U3651 (N_3651,N_2179,N_1698);
or U3652 (N_3652,N_111,N_205);
or U3653 (N_3653,N_1966,N_1282);
and U3654 (N_3654,N_1931,N_1325);
and U3655 (N_3655,N_390,N_583);
nor U3656 (N_3656,N_1794,N_1799);
or U3657 (N_3657,N_159,N_298);
xor U3658 (N_3658,N_2890,N_1285);
xnor U3659 (N_3659,N_1844,N_1556);
and U3660 (N_3660,N_1828,N_651);
xor U3661 (N_3661,N_2594,N_1740);
or U3662 (N_3662,N_1115,N_2232);
xor U3663 (N_3663,N_1324,N_2789);
nor U3664 (N_3664,N_948,N_1050);
xor U3665 (N_3665,N_2823,N_2391);
nor U3666 (N_3666,N_726,N_737);
nor U3667 (N_3667,N_314,N_2336);
and U3668 (N_3668,N_514,N_649);
and U3669 (N_3669,N_2181,N_708);
nand U3670 (N_3670,N_2460,N_2180);
xnor U3671 (N_3671,N_1978,N_120);
nor U3672 (N_3672,N_2799,N_1192);
nor U3673 (N_3673,N_1168,N_379);
nor U3674 (N_3674,N_404,N_625);
nor U3675 (N_3675,N_2898,N_575);
xnor U3676 (N_3676,N_2354,N_1689);
xor U3677 (N_3677,N_1563,N_1631);
or U3678 (N_3678,N_1188,N_2625);
nand U3679 (N_3679,N_2527,N_313);
nor U3680 (N_3680,N_224,N_1988);
or U3681 (N_3681,N_2017,N_254);
nand U3682 (N_3682,N_2004,N_226);
nor U3683 (N_3683,N_2797,N_319);
and U3684 (N_3684,N_607,N_272);
nor U3685 (N_3685,N_1370,N_1149);
or U3686 (N_3686,N_1314,N_2881);
xnor U3687 (N_3687,N_1159,N_456);
and U3688 (N_3688,N_2059,N_1228);
or U3689 (N_3689,N_1400,N_1884);
and U3690 (N_3690,N_2252,N_137);
or U3691 (N_3691,N_1205,N_307);
xnor U3692 (N_3692,N_639,N_1360);
nor U3693 (N_3693,N_2989,N_2671);
nand U3694 (N_3694,N_1460,N_2163);
and U3695 (N_3695,N_2900,N_1124);
or U3696 (N_3696,N_1676,N_439);
nand U3697 (N_3697,N_1183,N_1664);
and U3698 (N_3698,N_1795,N_208);
nand U3699 (N_3699,N_1107,N_2616);
nand U3700 (N_3700,N_2954,N_446);
and U3701 (N_3701,N_1201,N_814);
nor U3702 (N_3702,N_507,N_2140);
nor U3703 (N_3703,N_2837,N_1483);
and U3704 (N_3704,N_170,N_1218);
xnor U3705 (N_3705,N_2927,N_2869);
nand U3706 (N_3706,N_1850,N_1950);
xnor U3707 (N_3707,N_1954,N_281);
or U3708 (N_3708,N_2,N_169);
and U3709 (N_3709,N_698,N_2740);
or U3710 (N_3710,N_973,N_1345);
or U3711 (N_3711,N_1004,N_1045);
or U3712 (N_3712,N_2160,N_408);
and U3713 (N_3713,N_650,N_1056);
nor U3714 (N_3714,N_2628,N_1353);
or U3715 (N_3715,N_299,N_2814);
nand U3716 (N_3716,N_675,N_2012);
nor U3717 (N_3717,N_1060,N_672);
and U3718 (N_3718,N_2825,N_1024);
nor U3719 (N_3719,N_1473,N_2001);
xnor U3720 (N_3720,N_2438,N_1864);
or U3721 (N_3721,N_1958,N_2349);
or U3722 (N_3722,N_1470,N_1003);
nor U3723 (N_3723,N_1983,N_441);
nand U3724 (N_3724,N_2915,N_1596);
xnor U3725 (N_3725,N_2162,N_1638);
and U3726 (N_3726,N_2674,N_2124);
or U3727 (N_3727,N_899,N_2934);
xor U3728 (N_3728,N_264,N_756);
xor U3729 (N_3729,N_1229,N_2846);
nor U3730 (N_3730,N_2631,N_370);
nand U3731 (N_3731,N_775,N_523);
nor U3732 (N_3732,N_532,N_1957);
and U3733 (N_3733,N_1340,N_1785);
or U3734 (N_3734,N_2239,N_2780);
or U3735 (N_3735,N_1303,N_1597);
or U3736 (N_3736,N_1811,N_1738);
xnor U3737 (N_3737,N_2212,N_2787);
and U3738 (N_3738,N_2684,N_717);
or U3739 (N_3739,N_2360,N_2305);
xor U3740 (N_3740,N_1083,N_1617);
nand U3741 (N_3741,N_2475,N_325);
nor U3742 (N_3742,N_9,N_1933);
or U3743 (N_3743,N_470,N_1512);
nor U3744 (N_3744,N_462,N_1953);
or U3745 (N_3745,N_484,N_1855);
or U3746 (N_3746,N_46,N_696);
and U3747 (N_3747,N_1026,N_1685);
and U3748 (N_3748,N_1766,N_1346);
xnor U3749 (N_3749,N_1143,N_995);
nand U3750 (N_3750,N_1829,N_1461);
or U3751 (N_3751,N_460,N_1428);
xnor U3752 (N_3752,N_1444,N_568);
xnor U3753 (N_3753,N_824,N_2458);
and U3754 (N_3754,N_1789,N_1699);
xnor U3755 (N_3755,N_2521,N_191);
nor U3756 (N_3756,N_1744,N_2128);
nand U3757 (N_3757,N_1248,N_577);
or U3758 (N_3758,N_2770,N_1902);
or U3759 (N_3759,N_2602,N_2388);
and U3760 (N_3760,N_982,N_1874);
xor U3761 (N_3761,N_386,N_1823);
xor U3762 (N_3762,N_794,N_2909);
or U3763 (N_3763,N_1945,N_2885);
xnor U3764 (N_3764,N_1843,N_418);
nand U3765 (N_3765,N_1122,N_1960);
nand U3766 (N_3766,N_1831,N_1819);
and U3767 (N_3767,N_2443,N_1376);
and U3768 (N_3768,N_2445,N_1806);
and U3769 (N_3769,N_2669,N_1471);
or U3770 (N_3770,N_233,N_1142);
and U3771 (N_3771,N_2375,N_1405);
xnor U3772 (N_3772,N_584,N_837);
and U3773 (N_3773,N_2614,N_958);
xnor U3774 (N_3774,N_826,N_2523);
or U3775 (N_3775,N_2363,N_129);
nand U3776 (N_3776,N_624,N_2235);
xnor U3777 (N_3777,N_1907,N_2289);
nand U3778 (N_3778,N_471,N_560);
and U3779 (N_3779,N_1477,N_341);
xor U3780 (N_3780,N_1655,N_1134);
and U3781 (N_3781,N_2980,N_1842);
or U3782 (N_3782,N_287,N_2283);
nand U3783 (N_3783,N_1520,N_928);
or U3784 (N_3784,N_178,N_2077);
nor U3785 (N_3785,N_1321,N_1704);
nand U3786 (N_3786,N_2234,N_2767);
nor U3787 (N_3787,N_2717,N_601);
and U3788 (N_3788,N_24,N_1852);
or U3789 (N_3789,N_2484,N_815);
or U3790 (N_3790,N_544,N_38);
xor U3791 (N_3791,N_202,N_274);
or U3792 (N_3792,N_548,N_1342);
xor U3793 (N_3793,N_44,N_627);
xor U3794 (N_3794,N_2082,N_773);
nor U3795 (N_3795,N_1085,N_2106);
nand U3796 (N_3796,N_2805,N_728);
nand U3797 (N_3797,N_1174,N_1315);
nand U3798 (N_3798,N_1788,N_2114);
and U3799 (N_3799,N_2952,N_2462);
or U3800 (N_3800,N_2097,N_2488);
nand U3801 (N_3801,N_1772,N_5);
nand U3802 (N_3802,N_448,N_2020);
or U3803 (N_3803,N_1602,N_902);
xnor U3804 (N_3804,N_2390,N_1516);
nor U3805 (N_3805,N_1667,N_295);
nand U3806 (N_3806,N_916,N_2268);
or U3807 (N_3807,N_936,N_2221);
xnor U3808 (N_3808,N_1333,N_770);
xnor U3809 (N_3809,N_2492,N_2686);
nor U3810 (N_3810,N_2224,N_633);
or U3811 (N_3811,N_1787,N_2269);
and U3812 (N_3812,N_79,N_45);
nor U3813 (N_3813,N_1231,N_1879);
nor U3814 (N_3814,N_2566,N_2725);
nand U3815 (N_3815,N_1793,N_2712);
nand U3816 (N_3816,N_2756,N_962);
or U3817 (N_3817,N_2129,N_292);
or U3818 (N_3818,N_62,N_2315);
xor U3819 (N_3819,N_2042,N_1108);
and U3820 (N_3820,N_746,N_2177);
nor U3821 (N_3821,N_171,N_890);
and U3822 (N_3822,N_1838,N_2946);
or U3823 (N_3823,N_1565,N_279);
nor U3824 (N_3824,N_2368,N_2430);
or U3825 (N_3825,N_271,N_2877);
nor U3826 (N_3826,N_1888,N_442);
or U3827 (N_3827,N_1576,N_2793);
xor U3828 (N_3828,N_2622,N_1974);
or U3829 (N_3829,N_2143,N_2146);
xnor U3830 (N_3830,N_1965,N_2518);
nand U3831 (N_3831,N_2562,N_434);
or U3832 (N_3832,N_37,N_1066);
nor U3833 (N_3833,N_2171,N_53);
nand U3834 (N_3834,N_646,N_1014);
or U3835 (N_3835,N_186,N_1131);
or U3836 (N_3836,N_2803,N_43);
nor U3837 (N_3837,N_2378,N_1048);
or U3838 (N_3838,N_2026,N_1589);
nor U3839 (N_3839,N_1349,N_2530);
nor U3840 (N_3840,N_2573,N_1166);
nor U3841 (N_3841,N_909,N_2188);
xnor U3842 (N_3842,N_380,N_2008);
nand U3843 (N_3843,N_2529,N_738);
and U3844 (N_3844,N_94,N_2404);
nand U3845 (N_3845,N_991,N_1612);
xor U3846 (N_3846,N_1289,N_1936);
xor U3847 (N_3847,N_2689,N_74);
nor U3848 (N_3848,N_1804,N_33);
or U3849 (N_3849,N_1288,N_2556);
nor U3850 (N_3850,N_2847,N_2504);
nand U3851 (N_3851,N_2879,N_910);
nand U3852 (N_3852,N_1614,N_2242);
and U3853 (N_3853,N_2798,N_1690);
or U3854 (N_3854,N_494,N_1013);
nand U3855 (N_3855,N_682,N_2638);
nor U3856 (N_3856,N_1253,N_474);
nor U3857 (N_3857,N_1080,N_396);
xnor U3858 (N_3858,N_1267,N_831);
or U3859 (N_3859,N_1901,N_1310);
xnor U3860 (N_3860,N_1998,N_1277);
nand U3861 (N_3861,N_1569,N_1715);
nand U3862 (N_3862,N_517,N_427);
and U3863 (N_3863,N_1011,N_878);
xor U3864 (N_3864,N_2384,N_1126);
nor U3865 (N_3865,N_2563,N_168);
or U3866 (N_3866,N_2134,N_1997);
nor U3867 (N_3867,N_1948,N_1039);
or U3868 (N_3868,N_2158,N_39);
nor U3869 (N_3869,N_1162,N_403);
xor U3870 (N_3870,N_970,N_2362);
and U3871 (N_3871,N_599,N_757);
nor U3872 (N_3872,N_429,N_2364);
or U3873 (N_3873,N_2778,N_2340);
and U3874 (N_3874,N_588,N_378);
and U3875 (N_3875,N_2432,N_562);
or U3876 (N_3876,N_2533,N_739);
nor U3877 (N_3877,N_1419,N_1862);
nand U3878 (N_3878,N_22,N_2157);
xor U3879 (N_3879,N_2284,N_552);
or U3880 (N_3880,N_1028,N_1337);
nand U3881 (N_3881,N_680,N_2144);
or U3882 (N_3882,N_683,N_2478);
and U3883 (N_3883,N_2880,N_589);
nor U3884 (N_3884,N_1567,N_1827);
or U3885 (N_3885,N_2071,N_2292);
xor U3886 (N_3886,N_2335,N_592);
or U3887 (N_3887,N_966,N_1980);
nor U3888 (N_3888,N_2519,N_600);
and U3889 (N_3889,N_825,N_929);
or U3890 (N_3890,N_1949,N_628);
nand U3891 (N_3891,N_2642,N_1629);
xor U3892 (N_3892,N_990,N_591);
and U3893 (N_3893,N_1135,N_1088);
nand U3894 (N_3894,N_2189,N_889);
and U3895 (N_3895,N_1220,N_992);
xor U3896 (N_3896,N_1706,N_2947);
xor U3897 (N_3897,N_216,N_2776);
or U3898 (N_3898,N_1051,N_1480);
xnor U3899 (N_3899,N_1591,N_2112);
and U3900 (N_3900,N_2777,N_915);
xor U3901 (N_3901,N_17,N_1487);
and U3902 (N_3902,N_2571,N_1092);
nand U3903 (N_3903,N_2486,N_821);
nand U3904 (N_3904,N_1643,N_2229);
nand U3905 (N_3905,N_2923,N_329);
and U3906 (N_3906,N_2658,N_1547);
or U3907 (N_3907,N_364,N_366);
nor U3908 (N_3908,N_1465,N_2417);
nor U3909 (N_3909,N_534,N_2619);
and U3910 (N_3910,N_1609,N_1044);
and U3911 (N_3911,N_1010,N_93);
or U3912 (N_3912,N_504,N_1751);
nand U3913 (N_3913,N_659,N_2350);
and U3914 (N_3914,N_1904,N_828);
xnor U3915 (N_3915,N_1564,N_912);
nor U3916 (N_3916,N_1186,N_1215);
and U3917 (N_3917,N_2760,N_1001);
and U3918 (N_3918,N_2678,N_1015);
nor U3919 (N_3919,N_2280,N_1937);
and U3920 (N_3920,N_1241,N_2812);
and U3921 (N_3921,N_2500,N_635);
or U3922 (N_3922,N_83,N_2831);
xnor U3923 (N_3923,N_1322,N_2344);
xor U3924 (N_3924,N_2538,N_1017);
nand U3925 (N_3925,N_2061,N_2918);
or U3926 (N_3926,N_260,N_493);
xnor U3927 (N_3927,N_98,N_2723);
xor U3928 (N_3928,N_2820,N_2910);
and U3929 (N_3929,N_177,N_2348);
nor U3930 (N_3930,N_2655,N_1367);
and U3931 (N_3931,N_1637,N_153);
and U3932 (N_3932,N_637,N_2696);
nand U3933 (N_3933,N_1481,N_300);
nand U3934 (N_3934,N_2995,N_2649);
or U3935 (N_3935,N_1237,N_245);
nand U3936 (N_3936,N_2609,N_2759);
or U3937 (N_3937,N_2990,N_503);
nand U3938 (N_3938,N_1336,N_2708);
nand U3939 (N_3939,N_1388,N_762);
and U3940 (N_3940,N_1245,N_2560);
or U3941 (N_3941,N_1078,N_1578);
and U3942 (N_3942,N_1492,N_1136);
and U3943 (N_3943,N_166,N_612);
xnor U3944 (N_3944,N_334,N_243);
or U3945 (N_3945,N_1708,N_2749);
nand U3946 (N_3946,N_1332,N_865);
nor U3947 (N_3947,N_1454,N_1295);
nand U3948 (N_3948,N_323,N_158);
nor U3949 (N_3949,N_1568,N_1987);
nor U3950 (N_3950,N_1452,N_2161);
nor U3951 (N_3951,N_2839,N_819);
or U3952 (N_3952,N_361,N_311);
or U3953 (N_3953,N_480,N_2422);
and U3954 (N_3954,N_2829,N_459);
xnor U3955 (N_3955,N_1281,N_1745);
or U3956 (N_3956,N_479,N_2558);
or U3957 (N_3957,N_1775,N_1393);
or U3958 (N_3958,N_481,N_1163);
and U3959 (N_3959,N_222,N_2130);
and U3960 (N_3960,N_636,N_841);
nand U3961 (N_3961,N_2621,N_972);
nor U3962 (N_3962,N_2220,N_574);
or U3963 (N_3963,N_2747,N_2997);
and U3964 (N_3964,N_1291,N_2256);
nor U3965 (N_3965,N_1022,N_176);
xor U3966 (N_3966,N_2278,N_196);
or U3967 (N_3967,N_482,N_113);
nor U3968 (N_3968,N_283,N_2703);
nand U3969 (N_3969,N_1686,N_1305);
or U3970 (N_3970,N_2427,N_1737);
or U3971 (N_3971,N_1912,N_2039);
nor U3972 (N_3972,N_2887,N_2844);
xnor U3973 (N_3973,N_1990,N_2306);
nor U3974 (N_3974,N_55,N_833);
xor U3975 (N_3975,N_90,N_2868);
or U3976 (N_3976,N_988,N_2395);
xor U3977 (N_3977,N_2370,N_1434);
xnor U3978 (N_3978,N_104,N_1323);
and U3979 (N_3979,N_1651,N_348);
nor U3980 (N_3980,N_2791,N_66);
nand U3981 (N_3981,N_2845,N_2921);
or U3982 (N_3982,N_1020,N_851);
nand U3983 (N_3983,N_2966,N_1845);
nor U3984 (N_3984,N_1491,N_2830);
xnor U3985 (N_3985,N_2996,N_1254);
nand U3986 (N_3986,N_1513,N_932);
and U3987 (N_3987,N_1727,N_1071);
nand U3988 (N_3988,N_155,N_945);
nand U3989 (N_3989,N_1138,N_2611);
and U3990 (N_3990,N_565,N_1418);
nand U3991 (N_3991,N_1537,N_2035);
and U3992 (N_3992,N_193,N_528);
nand U3993 (N_3993,N_1494,N_645);
or U3994 (N_3994,N_1919,N_2185);
and U3995 (N_3995,N_2707,N_604);
nand U3996 (N_3996,N_2581,N_2436);
and U3997 (N_3997,N_2583,N_631);
nor U3998 (N_3998,N_461,N_513);
xor U3999 (N_3999,N_2987,N_2447);
nor U4000 (N_4000,N_555,N_2580);
or U4001 (N_4001,N_1734,N_417);
and U4002 (N_4002,N_2553,N_1110);
nor U4003 (N_4003,N_2433,N_454);
xor U4004 (N_4004,N_330,N_1279);
and U4005 (N_4005,N_1587,N_1680);
and U4006 (N_4006,N_2038,N_2745);
or U4007 (N_4007,N_1867,N_2099);
or U4008 (N_4008,N_1826,N_1036);
or U4009 (N_4009,N_1758,N_704);
xor U4010 (N_4010,N_128,N_2412);
xnor U4011 (N_4011,N_949,N_1409);
nor U4012 (N_4012,N_215,N_2369);
or U4013 (N_4013,N_384,N_1484);
nand U4014 (N_4014,N_805,N_157);
and U4015 (N_4015,N_1583,N_2057);
nand U4016 (N_4016,N_2863,N_449);
nor U4017 (N_4017,N_2125,N_1713);
nor U4018 (N_4018,N_918,N_1479);
or U4019 (N_4019,N_2345,N_2673);
xnor U4020 (N_4020,N_1506,N_2577);
nand U4021 (N_4021,N_2116,N_2905);
and U4022 (N_4022,N_1716,N_2474);
xnor U4023 (N_4023,N_1608,N_1538);
or U4024 (N_4024,N_2807,N_430);
and U4025 (N_4025,N_1805,N_2490);
or U4026 (N_4026,N_2483,N_2858);
or U4027 (N_4027,N_1307,N_1118);
nor U4028 (N_4028,N_1561,N_2132);
xor U4029 (N_4029,N_700,N_1424);
or U4030 (N_4030,N_745,N_164);
or U4031 (N_4031,N_424,N_2498);
nand U4032 (N_4032,N_2072,N_859);
nand U4033 (N_4033,N_2680,N_1171);
and U4034 (N_4034,N_1243,N_1441);
nand U4035 (N_4035,N_352,N_644);
and U4036 (N_4036,N_1866,N_2792);
xor U4037 (N_4037,N_2726,N_1812);
and U4038 (N_4038,N_1356,N_70);
nor U4039 (N_4039,N_946,N_1089);
xnor U4040 (N_4040,N_2471,N_1402);
and U4041 (N_4041,N_1052,N_2451);
xor U4042 (N_4042,N_550,N_255);
and U4043 (N_4043,N_2886,N_2413);
and U4044 (N_4044,N_676,N_1934);
nand U4045 (N_4045,N_398,N_393);
xor U4046 (N_4046,N_1825,N_1847);
xor U4047 (N_4047,N_2226,N_2495);
or U4048 (N_4048,N_2397,N_1928);
or U4049 (N_4049,N_895,N_2309);
xnor U4050 (N_4050,N_2786,N_147);
nor U4051 (N_4051,N_2047,N_907);
and U4052 (N_4052,N_1660,N_1120);
xor U4053 (N_4053,N_1951,N_67);
xnor U4054 (N_4054,N_994,N_1760);
nor U4055 (N_4055,N_930,N_40);
and U4056 (N_4056,N_6,N_277);
and U4057 (N_4057,N_2748,N_1344);
and U4058 (N_4058,N_438,N_2467);
nor U4059 (N_4059,N_2285,N_901);
or U4060 (N_4060,N_192,N_455);
and U4061 (N_4061,N_2510,N_2719);
nor U4062 (N_4062,N_244,N_1856);
and U4063 (N_4063,N_1635,N_1451);
xor U4064 (N_4064,N_381,N_679);
nor U4065 (N_4065,N_1741,N_654);
or U4066 (N_4066,N_1755,N_549);
nand U4067 (N_4067,N_1414,N_78);
xor U4068 (N_4068,N_188,N_2266);
and U4069 (N_4069,N_2002,N_2148);
nand U4070 (N_4070,N_2448,N_1970);
xor U4071 (N_4071,N_2646,N_312);
nand U4072 (N_4072,N_802,N_2293);
nand U4073 (N_4073,N_2552,N_2913);
or U4074 (N_4074,N_533,N_1335);
and U4075 (N_4075,N_1579,N_554);
nor U4076 (N_4076,N_416,N_2291);
nor U4077 (N_4077,N_1164,N_36);
or U4078 (N_4078,N_375,N_795);
nor U4079 (N_4079,N_2532,N_904);
xor U4080 (N_4080,N_2016,N_59);
and U4081 (N_4081,N_2441,N_2259);
or U4082 (N_4082,N_2941,N_207);
and U4083 (N_4083,N_2274,N_306);
or U4084 (N_4084,N_2359,N_2066);
nand U4085 (N_4085,N_535,N_420);
xnor U4086 (N_4086,N_1390,N_1061);
or U4087 (N_4087,N_836,N_1389);
nand U4088 (N_4088,N_1747,N_1466);
or U4089 (N_4089,N_2790,N_344);
nand U4090 (N_4090,N_638,N_320);
xnor U4091 (N_4091,N_1544,N_2100);
and U4092 (N_4092,N_1000,N_608);
nor U4093 (N_4093,N_280,N_0);
xor U4094 (N_4094,N_2542,N_1580);
xor U4095 (N_4095,N_4,N_2652);
and U4096 (N_4096,N_706,N_2771);
or U4097 (N_4097,N_1880,N_2311);
and U4098 (N_4098,N_2930,N_2656);
nand U4099 (N_4099,N_1752,N_955);
nor U4100 (N_4100,N_2329,N_1895);
nand U4101 (N_4101,N_117,N_751);
and U4102 (N_4102,N_1665,N_2875);
or U4103 (N_4103,N_880,N_1784);
and U4104 (N_4104,N_1411,N_2346);
or U4105 (N_4105,N_603,N_663);
nand U4106 (N_4106,N_2929,N_58);
xor U4107 (N_4107,N_2561,N_2386);
xor U4108 (N_4108,N_1068,N_2501);
and U4109 (N_4109,N_2972,N_286);
nand U4110 (N_4110,N_2901,N_2840);
xnor U4111 (N_4111,N_2514,N_1830);
and U4112 (N_4112,N_2277,N_1662);
nor U4113 (N_4113,N_1742,N_1896);
xor U4114 (N_4114,N_670,N_868);
or U4115 (N_4115,N_1926,N_658);
xor U4116 (N_4116,N_2699,N_1007);
and U4117 (N_4117,N_702,N_519);
or U4118 (N_4118,N_1290,N_2627);
nor U4119 (N_4119,N_154,N_518);
nor U4120 (N_4120,N_2011,N_371);
xor U4121 (N_4121,N_2165,N_2547);
or U4122 (N_4122,N_1445,N_1112);
xnor U4123 (N_4123,N_1739,N_2103);
nand U4124 (N_4124,N_2088,N_2374);
nor U4125 (N_4125,N_2062,N_1172);
nand U4126 (N_4126,N_971,N_2408);
or U4127 (N_4127,N_1312,N_1296);
or U4128 (N_4128,N_816,N_2670);
nor U4129 (N_4129,N_1942,N_1371);
xor U4130 (N_4130,N_953,N_595);
nor U4131 (N_4131,N_88,N_2420);
xnor U4132 (N_4132,N_1496,N_666);
nand U4133 (N_4133,N_2095,N_938);
and U4134 (N_4134,N_866,N_2871);
xnor U4135 (N_4135,N_1464,N_1909);
nor U4136 (N_4136,N_2313,N_1683);
nor U4137 (N_4137,N_2170,N_2590);
and U4138 (N_4138,N_2318,N_1610);
and U4139 (N_4139,N_2548,N_2089);
and U4140 (N_4140,N_2341,N_49);
and U4141 (N_4141,N_1287,N_2245);
xnor U4142 (N_4142,N_303,N_356);
xnor U4143 (N_4143,N_2668,N_2383);
and U4144 (N_4144,N_984,N_2326);
nand U4145 (N_4145,N_531,N_1505);
and U4146 (N_4146,N_2481,N_2854);
or U4147 (N_4147,N_145,N_2714);
nor U4148 (N_4148,N_2036,N_1595);
xor U4149 (N_4149,N_722,N_1150);
or U4150 (N_4150,N_1736,N_1141);
and U4151 (N_4151,N_414,N_799);
nor U4152 (N_4152,N_903,N_1696);
xnor U4153 (N_4153,N_1640,N_68);
nor U4154 (N_4154,N_581,N_2380);
and U4155 (N_4155,N_181,N_2908);
nor U4156 (N_4156,N_1735,N_996);
nand U4157 (N_4157,N_56,N_1177);
and U4158 (N_4158,N_2228,N_1266);
nor U4159 (N_4159,N_219,N_335);
nor U4160 (N_4160,N_1649,N_2186);
nand U4161 (N_4161,N_2377,N_1175);
nor U4162 (N_4162,N_2698,N_652);
and U4163 (N_4163,N_655,N_1633);
or U4164 (N_4164,N_2651,N_2819);
and U4165 (N_4165,N_230,N_594);
nand U4166 (N_4166,N_2324,N_750);
nand U4167 (N_4167,N_2784,N_741);
and U4168 (N_4168,N_316,N_2574);
or U4169 (N_4169,N_783,N_691);
nor U4170 (N_4170,N_1190,N_415);
and U4171 (N_4171,N_1472,N_2630);
or U4172 (N_4172,N_1467,N_2856);
and U4173 (N_4173,N_2009,N_2014);
nor U4174 (N_4174,N_1096,N_753);
nor U4175 (N_4175,N_2536,N_1993);
nand U4176 (N_4176,N_2522,N_92);
and U4177 (N_4177,N_1499,N_1489);
xnor U4178 (N_4178,N_537,N_1672);
nor U4179 (N_4179,N_105,N_710);
xnor U4180 (N_4180,N_1674,N_2133);
or U4181 (N_4181,N_61,N_2452);
xnor U4182 (N_4182,N_1191,N_1208);
nand U4183 (N_4183,N_1476,N_1552);
nor U4184 (N_4184,N_1641,N_2752);
nand U4185 (N_4185,N_1718,N_1302);
nor U4186 (N_4186,N_1308,N_1255);
nand U4187 (N_4187,N_1606,N_968);
and U4188 (N_4188,N_919,N_2046);
nand U4189 (N_4189,N_1944,N_1204);
xnor U4190 (N_4190,N_103,N_965);
and U4191 (N_4191,N_2113,N_1558);
nor U4192 (N_4192,N_29,N_1458);
nor U4193 (N_4193,N_2477,N_759);
or U4194 (N_4194,N_820,N_1801);
nor U4195 (N_4195,N_123,N_1620);
nand U4196 (N_4196,N_2509,N_1490);
nor U4197 (N_4197,N_1782,N_1729);
nand U4198 (N_4198,N_723,N_426);
nor U4199 (N_4199,N_1018,N_1771);
and U4200 (N_4200,N_1261,N_2993);
or U4201 (N_4201,N_2024,N_1768);
and U4202 (N_4202,N_669,N_2576);
xnor U4203 (N_4203,N_887,N_69);
xor U4204 (N_4204,N_450,N_2597);
nor U4205 (N_4205,N_2319,N_82);
nand U4206 (N_4206,N_502,N_198);
nand U4207 (N_4207,N_2338,N_185);
nor U4208 (N_4208,N_2603,N_2951);
xnor U4209 (N_4209,N_2225,N_2403);
xnor U4210 (N_4210,N_1057,N_2624);
or U4211 (N_4211,N_1877,N_1962);
nor U4212 (N_4212,N_2203,N_1899);
or U4213 (N_4213,N_2215,N_1156);
or U4214 (N_4214,N_2411,N_2661);
and U4215 (N_4215,N_1113,N_1876);
nand U4216 (N_4216,N_1362,N_258);
xnor U4217 (N_4217,N_845,N_1554);
xor U4218 (N_4218,N_2762,N_1167);
and U4219 (N_4219,N_1498,N_2279);
and U4220 (N_4220,N_447,N_1528);
nor U4221 (N_4221,N_1663,N_431);
nor U4222 (N_4222,N_1522,N_136);
nor U4223 (N_4223,N_896,N_2633);
or U4224 (N_4224,N_2464,N_2971);
nor U4225 (N_4225,N_846,N_1121);
nand U4226 (N_4226,N_843,N_520);
nor U4227 (N_4227,N_2195,N_413);
xor U4228 (N_4228,N_2801,N_892);
nand U4229 (N_4229,N_1500,N_2301);
xnor U4230 (N_4230,N_732,N_194);
and U4231 (N_4231,N_2549,N_2339);
or U4232 (N_4232,N_2409,N_1330);
or U4233 (N_4233,N_1214,N_2963);
nor U4234 (N_4234,N_2300,N_935);
nor U4235 (N_4235,N_2086,N_1854);
or U4236 (N_4236,N_1644,N_268);
or U4237 (N_4237,N_2049,N_1264);
nor U4238 (N_4238,N_242,N_1072);
nor U4239 (N_4239,N_363,N_1226);
or U4240 (N_4240,N_118,N_2598);
or U4241 (N_4241,N_688,N_2528);
xnor U4242 (N_4242,N_2782,N_2982);
nand U4243 (N_4243,N_2648,N_1647);
nand U4244 (N_4244,N_1514,N_1084);
and U4245 (N_4245,N_1559,N_2604);
and U4246 (N_4246,N_530,N_2903);
or U4247 (N_4247,N_1140,N_797);
nor U4248 (N_4248,N_2258,N_108);
nand U4249 (N_4249,N_457,N_2567);
nor U4250 (N_4250,N_1730,N_227);
and U4251 (N_4251,N_1276,N_844);
and U4252 (N_4252,N_2976,N_2579);
and U4253 (N_4253,N_411,N_712);
xor U4254 (N_4254,N_807,N_1551);
nand U4255 (N_4255,N_60,N_839);
or U4256 (N_4256,N_331,N_443);
nor U4257 (N_4257,N_134,N_1887);
xor U4258 (N_4258,N_2730,N_2208);
and U4259 (N_4259,N_2535,N_1908);
xnor U4260 (N_4260,N_2109,N_999);
nor U4261 (N_4261,N_876,N_1493);
and U4262 (N_4262,N_1929,N_2240);
xnor U4263 (N_4263,N_801,N_2685);
and U4264 (N_4264,N_1256,N_715);
or U4265 (N_4265,N_1098,N_1546);
nand U4266 (N_4266,N_2094,N_2098);
or U4267 (N_4267,N_2610,N_1636);
and U4268 (N_4268,N_2197,N_1065);
xnor U4269 (N_4269,N_2469,N_2731);
nor U4270 (N_4270,N_2428,N_1952);
xnor U4271 (N_4271,N_2502,N_234);
and U4272 (N_4272,N_1076,N_2487);
and U4273 (N_4273,N_1648,N_2588);
nand U4274 (N_4274,N_180,N_2410);
nor U4275 (N_4275,N_665,N_1857);
nor U4276 (N_4276,N_578,N_97);
and U4277 (N_4277,N_495,N_2446);
nor U4278 (N_4278,N_1408,N_2434);
xor U4279 (N_4279,N_2902,N_1588);
xnor U4280 (N_4280,N_410,N_573);
and U4281 (N_4281,N_1439,N_125);
nand U4282 (N_4282,N_2149,N_1530);
or U4283 (N_4283,N_373,N_175);
nor U4284 (N_4284,N_2198,N_1781);
or U4285 (N_4285,N_2733,N_1687);
and U4286 (N_4286,N_2994,N_211);
xnor U4287 (N_4287,N_615,N_1946);
nor U4288 (N_4288,N_2202,N_1343);
nor U4289 (N_4289,N_1779,N_729);
and U4290 (N_4290,N_2496,N_328);
nand U4291 (N_4291,N_162,N_2834);
nand U4292 (N_4292,N_305,N_1398);
xor U4293 (N_4293,N_632,N_2922);
nor U4294 (N_4294,N_1519,N_2351);
and U4295 (N_4295,N_389,N_1238);
and U4296 (N_4296,N_516,N_2862);
nor U4297 (N_4297,N_2808,N_2461);
nand U4298 (N_4298,N_1102,N_2653);
xor U4299 (N_4299,N_1363,N_267);
xor U4300 (N_4300,N_1846,N_2373);
and U4301 (N_4301,N_1763,N_611);
xnor U4302 (N_4302,N_1697,N_2785);
or U4303 (N_4303,N_1539,N_301);
xor U4304 (N_4304,N_2516,N_1515);
xor U4305 (N_4305,N_674,N_99);
nor U4306 (N_4306,N_1008,N_2029);
nand U4307 (N_4307,N_285,N_3);
or U4308 (N_4308,N_1714,N_629);
nand U4309 (N_4309,N_2254,N_2334);
and U4310 (N_4310,N_838,N_2939);
and U4311 (N_4311,N_2033,N_888);
nand U4312 (N_4312,N_2878,N_2297);
and U4313 (N_4313,N_606,N_1429);
nor U4314 (N_4314,N_376,N_2299);
nor U4315 (N_4315,N_1035,N_1769);
nand U4316 (N_4316,N_1921,N_1870);
and U4317 (N_4317,N_1029,N_2421);
nand U4318 (N_4318,N_2164,N_2201);
nor U4319 (N_4319,N_2734,N_421);
nor U4320 (N_4320,N_760,N_2156);
and U4321 (N_4321,N_1365,N_11);
and U4322 (N_4322,N_979,N_2070);
and U4323 (N_4323,N_2032,N_2479);
nand U4324 (N_4324,N_322,N_107);
nor U4325 (N_4325,N_2353,N_1271);
or U4326 (N_4326,N_1079,N_2025);
nand U4327 (N_4327,N_2906,N_2667);
and U4328 (N_4328,N_1534,N_647);
nor U4329 (N_4329,N_76,N_881);
nand U4330 (N_4330,N_1023,N_1810);
nand U4331 (N_4331,N_765,N_2746);
or U4332 (N_4332,N_2691,N_2672);
or U4333 (N_4333,N_586,N_551);
xor U4334 (N_4334,N_2243,N_2041);
and U4335 (N_4335,N_1808,N_2440);
xor U4336 (N_4336,N_1616,N_961);
nor U4337 (N_4337,N_2607,N_1090);
xor U4338 (N_4338,N_614,N_2260);
nand U4339 (N_4339,N_2152,N_52);
nand U4340 (N_4340,N_1406,N_1693);
xor U4341 (N_4341,N_720,N_1903);
xnor U4342 (N_4342,N_1677,N_505);
and U4343 (N_4343,N_1436,N_1154);
or U4344 (N_4344,N_1834,N_472);
and U4345 (N_4345,N_2546,N_2248);
nor U4346 (N_4346,N_1415,N_1369);
xor U4347 (N_4347,N_2841,N_1);
or U4348 (N_4348,N_1733,N_339);
and U4349 (N_4349,N_730,N_124);
nor U4350 (N_4350,N_1985,N_569);
nand U4351 (N_4351,N_630,N_882);
and U4352 (N_4352,N_835,N_2932);
nand U4353 (N_4353,N_468,N_1535);
nand U4354 (N_4354,N_2325,N_400);
or U4355 (N_4355,N_690,N_848);
nand U4356 (N_4356,N_1849,N_338);
nor U4357 (N_4357,N_1792,N_2705);
nor U4358 (N_4358,N_236,N_1449);
nand U4359 (N_4359,N_2928,N_1695);
and U4360 (N_4360,N_490,N_747);
and U4361 (N_4361,N_2122,N_1518);
or U4362 (N_4362,N_2836,N_2021);
nor U4363 (N_4363,N_1759,N_2154);
and U4364 (N_4364,N_2298,N_293);
nor U4365 (N_4365,N_678,N_114);
nand U4366 (N_4366,N_1701,N_1511);
or U4367 (N_4367,N_2626,N_2381);
nor U4368 (N_4368,N_2314,N_2815);
xnor U4369 (N_4369,N_1656,N_2174);
nand U4370 (N_4370,N_849,N_2675);
or U4371 (N_4371,N_1707,N_2037);
nand U4372 (N_4372,N_874,N_1575);
or U4373 (N_4373,N_1555,N_309);
xnor U4374 (N_4374,N_2722,N_2304);
nand U4375 (N_4375,N_2632,N_2183);
nor U4376 (N_4376,N_146,N_337);
and U4377 (N_4377,N_2534,N_2210);
nand U4378 (N_4378,N_1063,N_1104);
and U4379 (N_4379,N_620,N_2389);
and U4380 (N_4380,N_2978,N_2657);
nand U4381 (N_4381,N_1005,N_1673);
nand U4382 (N_4382,N_1938,N_763);
nor U4383 (N_4383,N_133,N_1430);
or U4384 (N_4384,N_1202,N_263);
xnor U4385 (N_4385,N_1269,N_2064);
nor U4386 (N_4386,N_1968,N_2043);
nand U4387 (N_4387,N_681,N_1339);
and U4388 (N_4388,N_217,N_235);
and U4389 (N_4389,N_488,N_1087);
and U4390 (N_4390,N_2853,N_2589);
or U4391 (N_4391,N_511,N_692);
and U4392 (N_4392,N_2743,N_2764);
and U4393 (N_4393,N_1549,N_1297);
or U4394 (N_4394,N_1973,N_1767);
nand U4395 (N_4395,N_1898,N_2425);
or U4396 (N_4396,N_1137,N_2473);
xnor U4397 (N_4397,N_1541,N_419);
or U4398 (N_4398,N_911,N_1219);
nand U4399 (N_4399,N_100,N_806);
and U4400 (N_4400,N_1913,N_1560);
or U4401 (N_4401,N_855,N_1006);
nand U4402 (N_4402,N_771,N_778);
or U4403 (N_4403,N_498,N_2643);
nor U4404 (N_4404,N_1871,N_1956);
and U4405 (N_4405,N_2769,N_354);
nand U4406 (N_4406,N_740,N_1368);
or U4407 (N_4407,N_1590,N_2470);
xor U4408 (N_4408,N_2423,N_2765);
nor U4409 (N_4409,N_576,N_1224);
xnor U4410 (N_4410,N_2984,N_1791);
xnor U4411 (N_4411,N_440,N_2585);
and U4412 (N_4412,N_1553,N_223);
nor U4413 (N_4413,N_1783,N_289);
nor U4414 (N_4414,N_725,N_1185);
nor U4415 (N_4415,N_686,N_2275);
and U4416 (N_4416,N_2044,N_1351);
xor U4417 (N_4417,N_115,N_1263);
nor U4418 (N_4418,N_465,N_2937);
and U4419 (N_4419,N_2358,N_1158);
nor U4420 (N_4420,N_96,N_2827);
xor U4421 (N_4421,N_1550,N_2729);
or U4422 (N_4422,N_149,N_2544);
and U4423 (N_4423,N_2105,N_508);
and U4424 (N_4424,N_808,N_1679);
and U4425 (N_4425,N_735,N_2367);
nand U4426 (N_4426,N_1917,N_2074);
nor U4427 (N_4427,N_764,N_2704);
nor U4428 (N_4428,N_1851,N_16);
xor U4429 (N_4429,N_1040,N_2998);
and U4430 (N_4430,N_827,N_1615);
nand U4431 (N_4431,N_2506,N_317);
nor U4432 (N_4432,N_2569,N_2559);
nor U4433 (N_4433,N_2710,N_1762);
nor U4434 (N_4434,N_1169,N_467);
nand U4435 (N_4435,N_1840,N_610);
and U4436 (N_4436,N_587,N_1173);
xor U4437 (N_4437,N_2640,N_2147);
xor U4438 (N_4438,N_2606,N_1920);
nor U4439 (N_4439,N_1582,N_2570);
or U4440 (N_4440,N_241,N_1626);
nor U4441 (N_4441,N_1959,N_924);
nor U4442 (N_4442,N_1486,N_1478);
or U4443 (N_4443,N_2683,N_249);
nand U4444 (N_4444,N_557,N_744);
xor U4445 (N_4445,N_952,N_1082);
and U4446 (N_4446,N_212,N_2347);
nor U4447 (N_4447,N_121,N_1207);
nor U4448 (N_4448,N_14,N_758);
nor U4449 (N_4449,N_2193,N_1420);
xor U4450 (N_4450,N_2081,N_1671);
nor U4451 (N_4451,N_383,N_605);
and U4452 (N_4452,N_48,N_742);
xnor U4453 (N_4453,N_391,N_2000);
nand U4454 (N_4454,N_2263,N_1147);
xnor U4455 (N_4455,N_15,N_1075);
nand U4456 (N_4456,N_1033,N_1731);
nor U4457 (N_4457,N_1746,N_30);
or U4458 (N_4458,N_184,N_898);
nand U4459 (N_4459,N_733,N_458);
xnor U4460 (N_4460,N_2030,N_139);
xor U4461 (N_4461,N_340,N_798);
nand U4462 (N_4462,N_2405,N_2591);
xor U4463 (N_4463,N_1682,N_190);
nor U4464 (N_4464,N_1694,N_2175);
nand U4465 (N_4465,N_2944,N_1995);
xor U4466 (N_4466,N_1211,N_327);
nand U4467 (N_4467,N_2660,N_1837);
nand U4468 (N_4468,N_779,N_221);
xor U4469 (N_4469,N_2327,N_1049);
nand U4470 (N_4470,N_2400,N_1374);
or U4471 (N_4471,N_269,N_1894);
xnor U4472 (N_4472,N_1038,N_2337);
xor U4473 (N_4473,N_950,N_1668);
xnor U4474 (N_4474,N_2985,N_112);
nand U4475 (N_4475,N_2214,N_1646);
and U4476 (N_4476,N_2418,N_506);
nor U4477 (N_4477,N_284,N_1653);
xnor U4478 (N_4478,N_1566,N_360);
nand U4479 (N_4479,N_687,N_266);
nor U4480 (N_4480,N_951,N_2454);
nor U4481 (N_4481,N_1859,N_1628);
or U4482 (N_4482,N_721,N_570);
or U4483 (N_4483,N_2271,N_34);
nor U4484 (N_4484,N_1407,N_536);
nand U4485 (N_4485,N_782,N_724);
or U4486 (N_4486,N_2572,N_2503);
and U4487 (N_4487,N_1611,N_2272);
nand U4488 (N_4488,N_428,N_2048);
xor U4489 (N_4489,N_2449,N_873);
or U4490 (N_4490,N_823,N_1361);
nand U4491 (N_4491,N_1273,N_2101);
xor U4492 (N_4492,N_47,N_2121);
nor U4493 (N_4493,N_1383,N_1058);
nor U4494 (N_4494,N_2596,N_1105);
nor U4495 (N_4495,N_2244,N_199);
or U4496 (N_4496,N_1761,N_934);
xor U4497 (N_4497,N_116,N_643);
nand U4498 (N_4498,N_1317,N_2857);
or U4499 (N_4499,N_1417,N_2276);
or U4500 (N_4500,N_2769,N_477);
xor U4501 (N_4501,N_2246,N_999);
nor U4502 (N_4502,N_971,N_2633);
nand U4503 (N_4503,N_1249,N_18);
xor U4504 (N_4504,N_2294,N_918);
nor U4505 (N_4505,N_2678,N_1780);
nor U4506 (N_4506,N_1827,N_2353);
or U4507 (N_4507,N_2946,N_2598);
xnor U4508 (N_4508,N_1363,N_1256);
nand U4509 (N_4509,N_717,N_1421);
xnor U4510 (N_4510,N_1459,N_1446);
nand U4511 (N_4511,N_2345,N_1382);
and U4512 (N_4512,N_711,N_2085);
and U4513 (N_4513,N_1170,N_2878);
and U4514 (N_4514,N_90,N_635);
xnor U4515 (N_4515,N_2248,N_349);
nor U4516 (N_4516,N_44,N_2846);
xnor U4517 (N_4517,N_550,N_743);
xnor U4518 (N_4518,N_651,N_2201);
nor U4519 (N_4519,N_2201,N_2146);
nor U4520 (N_4520,N_1686,N_2166);
xor U4521 (N_4521,N_805,N_925);
xor U4522 (N_4522,N_1962,N_382);
xnor U4523 (N_4523,N_1226,N_1941);
and U4524 (N_4524,N_2044,N_747);
xor U4525 (N_4525,N_983,N_2004);
nor U4526 (N_4526,N_2026,N_999);
nand U4527 (N_4527,N_2769,N_1685);
nor U4528 (N_4528,N_2299,N_2046);
or U4529 (N_4529,N_662,N_1224);
or U4530 (N_4530,N_2676,N_530);
and U4531 (N_4531,N_2466,N_2717);
nor U4532 (N_4532,N_2821,N_1992);
xor U4533 (N_4533,N_2089,N_1784);
and U4534 (N_4534,N_1443,N_2358);
nor U4535 (N_4535,N_860,N_624);
or U4536 (N_4536,N_2828,N_15);
xor U4537 (N_4537,N_758,N_742);
xnor U4538 (N_4538,N_689,N_1436);
nor U4539 (N_4539,N_1253,N_2968);
xor U4540 (N_4540,N_1360,N_115);
xnor U4541 (N_4541,N_2695,N_2316);
or U4542 (N_4542,N_1509,N_1587);
xor U4543 (N_4543,N_2934,N_706);
xnor U4544 (N_4544,N_2317,N_1605);
or U4545 (N_4545,N_1083,N_812);
or U4546 (N_4546,N_1999,N_2047);
or U4547 (N_4547,N_455,N_2350);
and U4548 (N_4548,N_1129,N_414);
nand U4549 (N_4549,N_1249,N_555);
nor U4550 (N_4550,N_2137,N_2572);
xor U4551 (N_4551,N_418,N_2812);
and U4552 (N_4552,N_826,N_168);
xor U4553 (N_4553,N_899,N_724);
nor U4554 (N_4554,N_23,N_16);
xor U4555 (N_4555,N_2571,N_824);
nor U4556 (N_4556,N_2585,N_1539);
or U4557 (N_4557,N_1833,N_1230);
and U4558 (N_4558,N_2120,N_2826);
nand U4559 (N_4559,N_1487,N_567);
xnor U4560 (N_4560,N_352,N_1364);
xnor U4561 (N_4561,N_1572,N_1217);
and U4562 (N_4562,N_332,N_1531);
or U4563 (N_4563,N_2285,N_0);
xnor U4564 (N_4564,N_2378,N_208);
xor U4565 (N_4565,N_144,N_489);
nor U4566 (N_4566,N_750,N_2752);
nor U4567 (N_4567,N_1161,N_2200);
xor U4568 (N_4568,N_2509,N_816);
or U4569 (N_4569,N_2658,N_1353);
nor U4570 (N_4570,N_2121,N_988);
or U4571 (N_4571,N_743,N_245);
nor U4572 (N_4572,N_2057,N_1915);
nand U4573 (N_4573,N_1422,N_2364);
xor U4574 (N_4574,N_1158,N_2839);
nand U4575 (N_4575,N_541,N_707);
xor U4576 (N_4576,N_2349,N_1020);
and U4577 (N_4577,N_1371,N_896);
nand U4578 (N_4578,N_1913,N_1241);
nor U4579 (N_4579,N_851,N_2832);
and U4580 (N_4580,N_2611,N_1576);
xnor U4581 (N_4581,N_1657,N_2053);
nor U4582 (N_4582,N_2887,N_98);
or U4583 (N_4583,N_168,N_2387);
and U4584 (N_4584,N_1251,N_2858);
nand U4585 (N_4585,N_776,N_2532);
xnor U4586 (N_4586,N_967,N_1459);
or U4587 (N_4587,N_541,N_1723);
or U4588 (N_4588,N_2438,N_681);
nand U4589 (N_4589,N_1345,N_281);
xnor U4590 (N_4590,N_1995,N_2284);
and U4591 (N_4591,N_1838,N_2764);
nor U4592 (N_4592,N_630,N_660);
or U4593 (N_4593,N_2803,N_887);
xor U4594 (N_4594,N_2170,N_2088);
or U4595 (N_4595,N_366,N_93);
nand U4596 (N_4596,N_2838,N_504);
and U4597 (N_4597,N_2641,N_1878);
and U4598 (N_4598,N_2129,N_958);
xor U4599 (N_4599,N_2903,N_449);
or U4600 (N_4600,N_1303,N_2939);
nand U4601 (N_4601,N_2465,N_765);
and U4602 (N_4602,N_636,N_542);
and U4603 (N_4603,N_401,N_730);
nor U4604 (N_4604,N_247,N_1633);
or U4605 (N_4605,N_576,N_1725);
nor U4606 (N_4606,N_1948,N_2212);
and U4607 (N_4607,N_648,N_1239);
and U4608 (N_4608,N_16,N_2338);
or U4609 (N_4609,N_694,N_2220);
xnor U4610 (N_4610,N_1527,N_798);
and U4611 (N_4611,N_903,N_2584);
nand U4612 (N_4612,N_801,N_1571);
nor U4613 (N_4613,N_2621,N_106);
and U4614 (N_4614,N_2605,N_639);
or U4615 (N_4615,N_225,N_2842);
and U4616 (N_4616,N_2418,N_784);
nor U4617 (N_4617,N_1835,N_1914);
nor U4618 (N_4618,N_1518,N_92);
nand U4619 (N_4619,N_2616,N_1127);
xnor U4620 (N_4620,N_2877,N_141);
or U4621 (N_4621,N_1568,N_669);
nor U4622 (N_4622,N_1030,N_1173);
xnor U4623 (N_4623,N_1571,N_985);
or U4624 (N_4624,N_1591,N_1014);
nand U4625 (N_4625,N_403,N_2308);
nand U4626 (N_4626,N_1930,N_1403);
xor U4627 (N_4627,N_1803,N_1468);
and U4628 (N_4628,N_2491,N_2617);
nor U4629 (N_4629,N_51,N_2562);
and U4630 (N_4630,N_703,N_2904);
and U4631 (N_4631,N_2947,N_1881);
xnor U4632 (N_4632,N_1331,N_2540);
nor U4633 (N_4633,N_569,N_2008);
xnor U4634 (N_4634,N_570,N_2044);
nor U4635 (N_4635,N_512,N_2009);
nor U4636 (N_4636,N_1308,N_2225);
xor U4637 (N_4637,N_923,N_2715);
xor U4638 (N_4638,N_1428,N_2551);
nor U4639 (N_4639,N_80,N_1545);
xnor U4640 (N_4640,N_1909,N_959);
xor U4641 (N_4641,N_2436,N_438);
nor U4642 (N_4642,N_2840,N_327);
xnor U4643 (N_4643,N_421,N_1686);
nor U4644 (N_4644,N_2655,N_329);
nand U4645 (N_4645,N_582,N_1336);
nand U4646 (N_4646,N_1948,N_74);
nor U4647 (N_4647,N_1540,N_219);
nand U4648 (N_4648,N_401,N_1723);
nor U4649 (N_4649,N_1776,N_1198);
nor U4650 (N_4650,N_322,N_1954);
and U4651 (N_4651,N_280,N_1531);
nand U4652 (N_4652,N_515,N_1643);
nor U4653 (N_4653,N_2543,N_1221);
or U4654 (N_4654,N_948,N_2698);
nand U4655 (N_4655,N_4,N_1715);
nand U4656 (N_4656,N_1419,N_807);
xnor U4657 (N_4657,N_2462,N_513);
xnor U4658 (N_4658,N_1573,N_2342);
and U4659 (N_4659,N_1070,N_402);
nand U4660 (N_4660,N_527,N_1017);
or U4661 (N_4661,N_2729,N_2119);
or U4662 (N_4662,N_964,N_590);
nor U4663 (N_4663,N_2610,N_2734);
xnor U4664 (N_4664,N_1173,N_83);
nor U4665 (N_4665,N_472,N_453);
nor U4666 (N_4666,N_2505,N_1080);
or U4667 (N_4667,N_2241,N_123);
and U4668 (N_4668,N_947,N_181);
or U4669 (N_4669,N_1878,N_2843);
and U4670 (N_4670,N_1575,N_2588);
nor U4671 (N_4671,N_1662,N_2894);
or U4672 (N_4672,N_1431,N_1560);
nor U4673 (N_4673,N_2721,N_2670);
xnor U4674 (N_4674,N_1603,N_1766);
or U4675 (N_4675,N_1994,N_1897);
and U4676 (N_4676,N_1941,N_2270);
xor U4677 (N_4677,N_2634,N_168);
nor U4678 (N_4678,N_436,N_2152);
nor U4679 (N_4679,N_1720,N_1990);
nand U4680 (N_4680,N_1822,N_1969);
nand U4681 (N_4681,N_1878,N_1819);
and U4682 (N_4682,N_1851,N_1485);
or U4683 (N_4683,N_1053,N_2202);
nor U4684 (N_4684,N_1112,N_806);
nor U4685 (N_4685,N_1003,N_2424);
or U4686 (N_4686,N_2353,N_1546);
or U4687 (N_4687,N_2240,N_458);
and U4688 (N_4688,N_639,N_2468);
and U4689 (N_4689,N_906,N_1318);
nand U4690 (N_4690,N_2185,N_1004);
nand U4691 (N_4691,N_2427,N_1659);
or U4692 (N_4692,N_1798,N_805);
nand U4693 (N_4693,N_164,N_1316);
nor U4694 (N_4694,N_2392,N_2671);
and U4695 (N_4695,N_534,N_1432);
or U4696 (N_4696,N_2480,N_753);
nor U4697 (N_4697,N_2099,N_2860);
and U4698 (N_4698,N_2477,N_181);
nand U4699 (N_4699,N_1780,N_1013);
nand U4700 (N_4700,N_2008,N_1717);
or U4701 (N_4701,N_749,N_43);
nor U4702 (N_4702,N_143,N_2672);
xor U4703 (N_4703,N_870,N_2010);
and U4704 (N_4704,N_814,N_1604);
or U4705 (N_4705,N_1714,N_576);
nor U4706 (N_4706,N_2898,N_486);
nor U4707 (N_4707,N_2533,N_2148);
or U4708 (N_4708,N_2279,N_850);
nand U4709 (N_4709,N_798,N_628);
xnor U4710 (N_4710,N_1879,N_2191);
or U4711 (N_4711,N_439,N_404);
or U4712 (N_4712,N_2454,N_1751);
nand U4713 (N_4713,N_1970,N_2652);
and U4714 (N_4714,N_209,N_1876);
or U4715 (N_4715,N_1051,N_884);
nand U4716 (N_4716,N_1273,N_2461);
and U4717 (N_4717,N_602,N_2033);
and U4718 (N_4718,N_748,N_2813);
nor U4719 (N_4719,N_735,N_1777);
nor U4720 (N_4720,N_2729,N_2507);
and U4721 (N_4721,N_1709,N_576);
and U4722 (N_4722,N_864,N_2437);
or U4723 (N_4723,N_572,N_177);
nor U4724 (N_4724,N_1257,N_863);
nand U4725 (N_4725,N_131,N_1647);
xnor U4726 (N_4726,N_1206,N_929);
nand U4727 (N_4727,N_1981,N_2763);
or U4728 (N_4728,N_1723,N_750);
nor U4729 (N_4729,N_915,N_2747);
nand U4730 (N_4730,N_1345,N_1400);
nor U4731 (N_4731,N_1159,N_139);
nand U4732 (N_4732,N_2572,N_2019);
nor U4733 (N_4733,N_1568,N_594);
xor U4734 (N_4734,N_2218,N_1668);
nand U4735 (N_4735,N_2193,N_2648);
nand U4736 (N_4736,N_1133,N_818);
nand U4737 (N_4737,N_2492,N_192);
nand U4738 (N_4738,N_2111,N_206);
and U4739 (N_4739,N_268,N_1605);
or U4740 (N_4740,N_1650,N_1647);
nand U4741 (N_4741,N_386,N_1151);
and U4742 (N_4742,N_1920,N_2926);
nor U4743 (N_4743,N_2779,N_2765);
xnor U4744 (N_4744,N_258,N_226);
or U4745 (N_4745,N_1276,N_2812);
xor U4746 (N_4746,N_2411,N_1968);
xnor U4747 (N_4747,N_2561,N_11);
or U4748 (N_4748,N_1899,N_729);
nor U4749 (N_4749,N_1459,N_1485);
and U4750 (N_4750,N_1892,N_1307);
xnor U4751 (N_4751,N_813,N_2455);
or U4752 (N_4752,N_1405,N_187);
nor U4753 (N_4753,N_2595,N_578);
xnor U4754 (N_4754,N_2296,N_1833);
and U4755 (N_4755,N_1973,N_919);
or U4756 (N_4756,N_2652,N_1729);
nand U4757 (N_4757,N_507,N_730);
or U4758 (N_4758,N_699,N_505);
or U4759 (N_4759,N_2840,N_2586);
xnor U4760 (N_4760,N_1161,N_453);
xnor U4761 (N_4761,N_394,N_835);
and U4762 (N_4762,N_2024,N_1069);
nand U4763 (N_4763,N_2070,N_562);
nor U4764 (N_4764,N_1821,N_910);
nand U4765 (N_4765,N_626,N_600);
nand U4766 (N_4766,N_700,N_685);
nand U4767 (N_4767,N_1864,N_827);
nand U4768 (N_4768,N_1261,N_1701);
nand U4769 (N_4769,N_1695,N_2626);
and U4770 (N_4770,N_1891,N_1644);
and U4771 (N_4771,N_94,N_220);
or U4772 (N_4772,N_2636,N_1658);
nand U4773 (N_4773,N_633,N_1826);
xor U4774 (N_4774,N_1801,N_2279);
and U4775 (N_4775,N_646,N_1338);
xor U4776 (N_4776,N_1165,N_832);
and U4777 (N_4777,N_2973,N_1163);
and U4778 (N_4778,N_1763,N_48);
xnor U4779 (N_4779,N_2027,N_2260);
xnor U4780 (N_4780,N_2654,N_725);
nand U4781 (N_4781,N_2724,N_1523);
or U4782 (N_4782,N_2759,N_2138);
nor U4783 (N_4783,N_2704,N_561);
nor U4784 (N_4784,N_1721,N_1798);
nand U4785 (N_4785,N_921,N_912);
xor U4786 (N_4786,N_2647,N_242);
nor U4787 (N_4787,N_1994,N_1484);
xnor U4788 (N_4788,N_756,N_912);
nor U4789 (N_4789,N_1870,N_1172);
or U4790 (N_4790,N_2165,N_2329);
and U4791 (N_4791,N_274,N_19);
xor U4792 (N_4792,N_485,N_2901);
nand U4793 (N_4793,N_806,N_2087);
or U4794 (N_4794,N_1212,N_1329);
xor U4795 (N_4795,N_254,N_1522);
nor U4796 (N_4796,N_574,N_669);
nand U4797 (N_4797,N_1140,N_778);
xor U4798 (N_4798,N_2202,N_11);
or U4799 (N_4799,N_300,N_1130);
nor U4800 (N_4800,N_2678,N_2755);
nor U4801 (N_4801,N_24,N_1702);
xnor U4802 (N_4802,N_1122,N_954);
or U4803 (N_4803,N_842,N_78);
and U4804 (N_4804,N_2257,N_959);
nand U4805 (N_4805,N_1792,N_672);
nor U4806 (N_4806,N_1715,N_1043);
xor U4807 (N_4807,N_2947,N_2232);
xor U4808 (N_4808,N_2135,N_809);
and U4809 (N_4809,N_1262,N_2807);
nand U4810 (N_4810,N_2375,N_1665);
xor U4811 (N_4811,N_1893,N_1886);
xor U4812 (N_4812,N_2655,N_864);
nor U4813 (N_4813,N_1268,N_306);
or U4814 (N_4814,N_2454,N_2023);
xor U4815 (N_4815,N_728,N_1483);
nand U4816 (N_4816,N_832,N_1107);
or U4817 (N_4817,N_2334,N_1867);
nor U4818 (N_4818,N_1365,N_63);
nor U4819 (N_4819,N_1067,N_53);
nand U4820 (N_4820,N_556,N_2680);
nor U4821 (N_4821,N_1600,N_456);
and U4822 (N_4822,N_1215,N_309);
nor U4823 (N_4823,N_2437,N_324);
and U4824 (N_4824,N_2682,N_2686);
and U4825 (N_4825,N_1723,N_1397);
nand U4826 (N_4826,N_2300,N_1241);
xor U4827 (N_4827,N_1142,N_274);
or U4828 (N_4828,N_2098,N_573);
or U4829 (N_4829,N_352,N_156);
nor U4830 (N_4830,N_1069,N_1808);
nor U4831 (N_4831,N_702,N_438);
xnor U4832 (N_4832,N_2788,N_2212);
and U4833 (N_4833,N_1599,N_1021);
and U4834 (N_4834,N_495,N_2586);
nand U4835 (N_4835,N_2038,N_593);
xor U4836 (N_4836,N_1619,N_378);
nand U4837 (N_4837,N_2928,N_30);
xnor U4838 (N_4838,N_331,N_539);
nor U4839 (N_4839,N_1746,N_1778);
nand U4840 (N_4840,N_48,N_599);
and U4841 (N_4841,N_2225,N_659);
or U4842 (N_4842,N_2606,N_2692);
nor U4843 (N_4843,N_2764,N_1446);
or U4844 (N_4844,N_2324,N_704);
nor U4845 (N_4845,N_2164,N_2620);
xor U4846 (N_4846,N_1486,N_597);
nand U4847 (N_4847,N_610,N_1870);
and U4848 (N_4848,N_156,N_742);
nand U4849 (N_4849,N_335,N_1452);
or U4850 (N_4850,N_459,N_2132);
xor U4851 (N_4851,N_885,N_1377);
or U4852 (N_4852,N_233,N_2530);
and U4853 (N_4853,N_2991,N_119);
nand U4854 (N_4854,N_227,N_1470);
xnor U4855 (N_4855,N_2155,N_2739);
xor U4856 (N_4856,N_962,N_973);
nand U4857 (N_4857,N_937,N_2439);
nor U4858 (N_4858,N_2143,N_2868);
xor U4859 (N_4859,N_481,N_2538);
xor U4860 (N_4860,N_882,N_2860);
and U4861 (N_4861,N_2223,N_348);
or U4862 (N_4862,N_2821,N_2425);
or U4863 (N_4863,N_2330,N_1188);
and U4864 (N_4864,N_2744,N_572);
or U4865 (N_4865,N_1657,N_2971);
xor U4866 (N_4866,N_1091,N_336);
and U4867 (N_4867,N_814,N_1348);
and U4868 (N_4868,N_1778,N_1213);
nand U4869 (N_4869,N_737,N_580);
nor U4870 (N_4870,N_2012,N_2927);
or U4871 (N_4871,N_2129,N_591);
and U4872 (N_4872,N_2702,N_1505);
nand U4873 (N_4873,N_1532,N_2339);
nor U4874 (N_4874,N_2259,N_972);
nor U4875 (N_4875,N_1248,N_1885);
nand U4876 (N_4876,N_1286,N_576);
nand U4877 (N_4877,N_2307,N_1185);
xnor U4878 (N_4878,N_1915,N_791);
nor U4879 (N_4879,N_1653,N_1183);
nor U4880 (N_4880,N_448,N_1774);
xor U4881 (N_4881,N_966,N_1819);
xnor U4882 (N_4882,N_1800,N_772);
or U4883 (N_4883,N_2557,N_80);
xor U4884 (N_4884,N_2917,N_1022);
and U4885 (N_4885,N_97,N_2555);
xor U4886 (N_4886,N_2717,N_318);
xnor U4887 (N_4887,N_2708,N_2289);
xor U4888 (N_4888,N_305,N_2025);
and U4889 (N_4889,N_2500,N_321);
or U4890 (N_4890,N_1761,N_1274);
or U4891 (N_4891,N_2875,N_1701);
nand U4892 (N_4892,N_2172,N_716);
xnor U4893 (N_4893,N_545,N_2173);
and U4894 (N_4894,N_2968,N_1500);
nand U4895 (N_4895,N_1656,N_1003);
or U4896 (N_4896,N_1244,N_1267);
nor U4897 (N_4897,N_1441,N_1789);
nand U4898 (N_4898,N_1976,N_1685);
or U4899 (N_4899,N_2101,N_2292);
nand U4900 (N_4900,N_1596,N_2513);
nor U4901 (N_4901,N_1605,N_2452);
xor U4902 (N_4902,N_1563,N_2984);
xor U4903 (N_4903,N_1468,N_2849);
or U4904 (N_4904,N_139,N_2916);
nor U4905 (N_4905,N_673,N_1179);
xor U4906 (N_4906,N_2896,N_842);
xor U4907 (N_4907,N_2226,N_2177);
or U4908 (N_4908,N_1877,N_1208);
or U4909 (N_4909,N_2364,N_1970);
nor U4910 (N_4910,N_2062,N_2458);
nor U4911 (N_4911,N_1788,N_2415);
and U4912 (N_4912,N_375,N_1113);
nor U4913 (N_4913,N_1040,N_166);
nor U4914 (N_4914,N_2979,N_543);
xnor U4915 (N_4915,N_2467,N_2340);
nor U4916 (N_4916,N_1642,N_2810);
or U4917 (N_4917,N_1627,N_2806);
xnor U4918 (N_4918,N_720,N_1286);
xnor U4919 (N_4919,N_2958,N_2949);
xnor U4920 (N_4920,N_1060,N_103);
or U4921 (N_4921,N_2155,N_791);
and U4922 (N_4922,N_2355,N_1822);
and U4923 (N_4923,N_2041,N_847);
nor U4924 (N_4924,N_2863,N_1210);
and U4925 (N_4925,N_1193,N_907);
or U4926 (N_4926,N_1009,N_2533);
xnor U4927 (N_4927,N_1075,N_2325);
xnor U4928 (N_4928,N_351,N_2938);
or U4929 (N_4929,N_2722,N_1480);
nand U4930 (N_4930,N_1668,N_2957);
nand U4931 (N_4931,N_1642,N_1360);
and U4932 (N_4932,N_493,N_2277);
xnor U4933 (N_4933,N_1598,N_112);
xor U4934 (N_4934,N_2277,N_1963);
or U4935 (N_4935,N_1807,N_1428);
nor U4936 (N_4936,N_2786,N_1955);
nor U4937 (N_4937,N_1577,N_2213);
nor U4938 (N_4938,N_2604,N_1623);
nand U4939 (N_4939,N_1,N_2603);
and U4940 (N_4940,N_1353,N_2744);
xor U4941 (N_4941,N_1190,N_2369);
nand U4942 (N_4942,N_1439,N_988);
or U4943 (N_4943,N_1190,N_701);
xnor U4944 (N_4944,N_487,N_1649);
or U4945 (N_4945,N_1355,N_2707);
nor U4946 (N_4946,N_1291,N_531);
nor U4947 (N_4947,N_1744,N_1613);
or U4948 (N_4948,N_174,N_1631);
and U4949 (N_4949,N_574,N_2903);
nand U4950 (N_4950,N_2002,N_71);
or U4951 (N_4951,N_2354,N_871);
and U4952 (N_4952,N_2553,N_2757);
or U4953 (N_4953,N_1976,N_1053);
xor U4954 (N_4954,N_1680,N_476);
and U4955 (N_4955,N_1901,N_1371);
and U4956 (N_4956,N_888,N_782);
nand U4957 (N_4957,N_1637,N_2876);
xnor U4958 (N_4958,N_2778,N_1362);
xor U4959 (N_4959,N_2330,N_346);
nand U4960 (N_4960,N_1091,N_2343);
nand U4961 (N_4961,N_1295,N_702);
and U4962 (N_4962,N_1614,N_995);
nor U4963 (N_4963,N_777,N_2121);
and U4964 (N_4964,N_1855,N_161);
and U4965 (N_4965,N_2795,N_2704);
or U4966 (N_4966,N_1441,N_2062);
nand U4967 (N_4967,N_1392,N_1772);
xor U4968 (N_4968,N_931,N_2025);
nor U4969 (N_4969,N_1743,N_487);
or U4970 (N_4970,N_2559,N_2067);
nor U4971 (N_4971,N_1965,N_251);
and U4972 (N_4972,N_2764,N_978);
xnor U4973 (N_4973,N_13,N_2691);
nand U4974 (N_4974,N_581,N_1928);
nor U4975 (N_4975,N_416,N_2954);
xnor U4976 (N_4976,N_907,N_192);
xnor U4977 (N_4977,N_1585,N_2231);
nor U4978 (N_4978,N_1576,N_301);
nand U4979 (N_4979,N_549,N_224);
and U4980 (N_4980,N_1558,N_2222);
xnor U4981 (N_4981,N_2536,N_895);
xor U4982 (N_4982,N_2821,N_1412);
xnor U4983 (N_4983,N_2609,N_2446);
xnor U4984 (N_4984,N_2065,N_451);
nor U4985 (N_4985,N_332,N_2947);
nor U4986 (N_4986,N_633,N_1158);
or U4987 (N_4987,N_181,N_830);
or U4988 (N_4988,N_677,N_465);
or U4989 (N_4989,N_1921,N_918);
xnor U4990 (N_4990,N_261,N_1274);
nand U4991 (N_4991,N_2036,N_883);
or U4992 (N_4992,N_1129,N_2345);
and U4993 (N_4993,N_2221,N_2195);
and U4994 (N_4994,N_1032,N_952);
and U4995 (N_4995,N_1738,N_149);
or U4996 (N_4996,N_2288,N_872);
nand U4997 (N_4997,N_1087,N_1040);
and U4998 (N_4998,N_113,N_2298);
or U4999 (N_4999,N_2770,N_1003);
nor U5000 (N_5000,N_2705,N_2728);
and U5001 (N_5001,N_1180,N_363);
xor U5002 (N_5002,N_375,N_632);
and U5003 (N_5003,N_2269,N_680);
and U5004 (N_5004,N_2097,N_233);
xor U5005 (N_5005,N_640,N_562);
nand U5006 (N_5006,N_1018,N_1550);
and U5007 (N_5007,N_247,N_1847);
or U5008 (N_5008,N_1573,N_1813);
nand U5009 (N_5009,N_53,N_2344);
nor U5010 (N_5010,N_2516,N_87);
xnor U5011 (N_5011,N_1361,N_2740);
nand U5012 (N_5012,N_2052,N_2479);
xnor U5013 (N_5013,N_1204,N_2515);
xnor U5014 (N_5014,N_1237,N_1861);
nand U5015 (N_5015,N_2656,N_2968);
nor U5016 (N_5016,N_701,N_846);
and U5017 (N_5017,N_1451,N_337);
xor U5018 (N_5018,N_189,N_118);
or U5019 (N_5019,N_589,N_987);
or U5020 (N_5020,N_2250,N_2031);
or U5021 (N_5021,N_8,N_1286);
nor U5022 (N_5022,N_1366,N_2933);
or U5023 (N_5023,N_1765,N_1990);
xor U5024 (N_5024,N_1830,N_1711);
nor U5025 (N_5025,N_1446,N_2896);
xor U5026 (N_5026,N_192,N_1235);
or U5027 (N_5027,N_2607,N_2023);
nor U5028 (N_5028,N_418,N_265);
nor U5029 (N_5029,N_670,N_2927);
nand U5030 (N_5030,N_109,N_1610);
xor U5031 (N_5031,N_9,N_2098);
xor U5032 (N_5032,N_1716,N_1900);
or U5033 (N_5033,N_930,N_1482);
nand U5034 (N_5034,N_1358,N_807);
xor U5035 (N_5035,N_2622,N_6);
and U5036 (N_5036,N_771,N_2570);
xnor U5037 (N_5037,N_615,N_1670);
nor U5038 (N_5038,N_443,N_883);
or U5039 (N_5039,N_920,N_1437);
xor U5040 (N_5040,N_2408,N_2497);
nand U5041 (N_5041,N_1534,N_1124);
or U5042 (N_5042,N_403,N_1504);
xor U5043 (N_5043,N_1447,N_984);
xnor U5044 (N_5044,N_1928,N_8);
and U5045 (N_5045,N_2037,N_1994);
nor U5046 (N_5046,N_221,N_1310);
or U5047 (N_5047,N_2678,N_2343);
and U5048 (N_5048,N_39,N_1469);
or U5049 (N_5049,N_1957,N_1300);
and U5050 (N_5050,N_2058,N_1847);
xnor U5051 (N_5051,N_2299,N_1836);
or U5052 (N_5052,N_303,N_830);
nand U5053 (N_5053,N_858,N_761);
or U5054 (N_5054,N_2948,N_2113);
or U5055 (N_5055,N_782,N_221);
xor U5056 (N_5056,N_1151,N_2507);
or U5057 (N_5057,N_702,N_1070);
or U5058 (N_5058,N_581,N_352);
xor U5059 (N_5059,N_735,N_2836);
or U5060 (N_5060,N_1982,N_637);
or U5061 (N_5061,N_1460,N_89);
or U5062 (N_5062,N_2407,N_172);
nor U5063 (N_5063,N_2067,N_669);
xnor U5064 (N_5064,N_2919,N_1691);
nor U5065 (N_5065,N_284,N_1344);
nor U5066 (N_5066,N_593,N_573);
nand U5067 (N_5067,N_1813,N_1853);
and U5068 (N_5068,N_2482,N_2320);
xnor U5069 (N_5069,N_790,N_385);
xor U5070 (N_5070,N_2417,N_1979);
nor U5071 (N_5071,N_1651,N_2864);
nand U5072 (N_5072,N_1479,N_2995);
and U5073 (N_5073,N_2513,N_1478);
and U5074 (N_5074,N_642,N_1129);
xnor U5075 (N_5075,N_375,N_706);
and U5076 (N_5076,N_1011,N_2136);
or U5077 (N_5077,N_1167,N_2265);
nand U5078 (N_5078,N_745,N_283);
nand U5079 (N_5079,N_1253,N_288);
nand U5080 (N_5080,N_1504,N_652);
and U5081 (N_5081,N_1708,N_2623);
or U5082 (N_5082,N_1479,N_1089);
xnor U5083 (N_5083,N_2316,N_1858);
xor U5084 (N_5084,N_2619,N_2657);
or U5085 (N_5085,N_1968,N_2841);
or U5086 (N_5086,N_2149,N_1248);
xnor U5087 (N_5087,N_2966,N_2086);
or U5088 (N_5088,N_2129,N_2063);
and U5089 (N_5089,N_708,N_1743);
or U5090 (N_5090,N_74,N_283);
or U5091 (N_5091,N_2327,N_1907);
or U5092 (N_5092,N_2538,N_1974);
and U5093 (N_5093,N_1864,N_1859);
nor U5094 (N_5094,N_1169,N_177);
xor U5095 (N_5095,N_962,N_803);
and U5096 (N_5096,N_2425,N_2513);
and U5097 (N_5097,N_913,N_658);
and U5098 (N_5098,N_2197,N_1848);
xor U5099 (N_5099,N_563,N_805);
or U5100 (N_5100,N_1263,N_1975);
and U5101 (N_5101,N_1442,N_472);
nand U5102 (N_5102,N_257,N_100);
and U5103 (N_5103,N_1266,N_183);
nand U5104 (N_5104,N_252,N_2004);
xor U5105 (N_5105,N_2274,N_2943);
nor U5106 (N_5106,N_1755,N_1836);
xor U5107 (N_5107,N_1271,N_780);
or U5108 (N_5108,N_1327,N_2706);
or U5109 (N_5109,N_519,N_411);
or U5110 (N_5110,N_381,N_1410);
nand U5111 (N_5111,N_744,N_2399);
or U5112 (N_5112,N_2370,N_2699);
xor U5113 (N_5113,N_2415,N_1917);
nand U5114 (N_5114,N_344,N_1840);
xnor U5115 (N_5115,N_590,N_343);
nor U5116 (N_5116,N_618,N_1124);
xor U5117 (N_5117,N_670,N_1511);
nand U5118 (N_5118,N_2130,N_517);
nor U5119 (N_5119,N_8,N_2780);
or U5120 (N_5120,N_6,N_2114);
and U5121 (N_5121,N_1089,N_2336);
and U5122 (N_5122,N_1743,N_1724);
nor U5123 (N_5123,N_363,N_265);
nor U5124 (N_5124,N_1332,N_857);
nor U5125 (N_5125,N_1824,N_689);
and U5126 (N_5126,N_2981,N_2425);
xor U5127 (N_5127,N_1508,N_1417);
and U5128 (N_5128,N_1404,N_522);
xnor U5129 (N_5129,N_2802,N_2864);
and U5130 (N_5130,N_2655,N_713);
or U5131 (N_5131,N_1597,N_1409);
and U5132 (N_5132,N_1550,N_952);
nand U5133 (N_5133,N_679,N_2948);
xor U5134 (N_5134,N_46,N_2915);
nand U5135 (N_5135,N_1684,N_339);
nor U5136 (N_5136,N_2011,N_2221);
and U5137 (N_5137,N_861,N_2451);
or U5138 (N_5138,N_2173,N_1958);
nand U5139 (N_5139,N_2252,N_873);
nand U5140 (N_5140,N_2979,N_2067);
nor U5141 (N_5141,N_2818,N_2057);
nand U5142 (N_5142,N_2867,N_1738);
xnor U5143 (N_5143,N_874,N_260);
or U5144 (N_5144,N_1211,N_2702);
or U5145 (N_5145,N_721,N_2112);
nand U5146 (N_5146,N_2457,N_2725);
nor U5147 (N_5147,N_2981,N_342);
or U5148 (N_5148,N_2354,N_1923);
xor U5149 (N_5149,N_2137,N_1879);
xnor U5150 (N_5150,N_1935,N_2722);
or U5151 (N_5151,N_924,N_2478);
or U5152 (N_5152,N_2489,N_2431);
nor U5153 (N_5153,N_2548,N_2082);
or U5154 (N_5154,N_1835,N_1818);
xor U5155 (N_5155,N_2461,N_1344);
nor U5156 (N_5156,N_1565,N_1177);
nand U5157 (N_5157,N_2164,N_124);
or U5158 (N_5158,N_215,N_1129);
and U5159 (N_5159,N_302,N_1626);
or U5160 (N_5160,N_1537,N_1096);
and U5161 (N_5161,N_503,N_282);
nor U5162 (N_5162,N_1624,N_2513);
nor U5163 (N_5163,N_608,N_2008);
and U5164 (N_5164,N_437,N_886);
nor U5165 (N_5165,N_2586,N_369);
and U5166 (N_5166,N_917,N_1144);
nor U5167 (N_5167,N_1178,N_654);
xnor U5168 (N_5168,N_2075,N_1095);
nand U5169 (N_5169,N_1175,N_547);
and U5170 (N_5170,N_1330,N_2642);
and U5171 (N_5171,N_2620,N_2371);
or U5172 (N_5172,N_82,N_2322);
nor U5173 (N_5173,N_1322,N_156);
and U5174 (N_5174,N_1337,N_708);
and U5175 (N_5175,N_1113,N_1325);
and U5176 (N_5176,N_2070,N_1152);
nand U5177 (N_5177,N_1459,N_2517);
or U5178 (N_5178,N_2081,N_2501);
or U5179 (N_5179,N_1117,N_2099);
xnor U5180 (N_5180,N_1247,N_454);
nand U5181 (N_5181,N_59,N_2279);
or U5182 (N_5182,N_2475,N_513);
nor U5183 (N_5183,N_2702,N_440);
nand U5184 (N_5184,N_2137,N_272);
or U5185 (N_5185,N_1080,N_589);
nand U5186 (N_5186,N_1047,N_1460);
nand U5187 (N_5187,N_1781,N_155);
and U5188 (N_5188,N_1041,N_2562);
and U5189 (N_5189,N_1197,N_157);
nand U5190 (N_5190,N_1055,N_2766);
nor U5191 (N_5191,N_2885,N_1341);
or U5192 (N_5192,N_2725,N_2299);
nand U5193 (N_5193,N_1761,N_250);
xnor U5194 (N_5194,N_897,N_1347);
xor U5195 (N_5195,N_1220,N_2579);
or U5196 (N_5196,N_2003,N_429);
xor U5197 (N_5197,N_2299,N_1886);
or U5198 (N_5198,N_1483,N_2463);
or U5199 (N_5199,N_1640,N_441);
xor U5200 (N_5200,N_1036,N_2060);
nor U5201 (N_5201,N_1937,N_1026);
or U5202 (N_5202,N_1273,N_746);
or U5203 (N_5203,N_1318,N_1080);
or U5204 (N_5204,N_879,N_2039);
or U5205 (N_5205,N_1155,N_151);
or U5206 (N_5206,N_549,N_897);
nor U5207 (N_5207,N_1191,N_1958);
xnor U5208 (N_5208,N_1932,N_1510);
nor U5209 (N_5209,N_549,N_2181);
and U5210 (N_5210,N_1465,N_1255);
nand U5211 (N_5211,N_2762,N_1425);
xor U5212 (N_5212,N_2197,N_2141);
xor U5213 (N_5213,N_342,N_798);
nor U5214 (N_5214,N_470,N_311);
and U5215 (N_5215,N_2414,N_266);
nand U5216 (N_5216,N_1576,N_2598);
and U5217 (N_5217,N_2159,N_893);
or U5218 (N_5218,N_2559,N_1347);
and U5219 (N_5219,N_1094,N_1684);
nand U5220 (N_5220,N_167,N_2407);
nand U5221 (N_5221,N_546,N_1588);
nand U5222 (N_5222,N_2223,N_2961);
nand U5223 (N_5223,N_112,N_1264);
and U5224 (N_5224,N_2434,N_1244);
or U5225 (N_5225,N_100,N_2753);
nor U5226 (N_5226,N_727,N_2626);
nor U5227 (N_5227,N_1752,N_194);
and U5228 (N_5228,N_1847,N_2834);
or U5229 (N_5229,N_2984,N_285);
nor U5230 (N_5230,N_1491,N_2101);
xnor U5231 (N_5231,N_118,N_459);
and U5232 (N_5232,N_2073,N_40);
xor U5233 (N_5233,N_1017,N_2647);
nor U5234 (N_5234,N_2609,N_468);
xor U5235 (N_5235,N_628,N_836);
nor U5236 (N_5236,N_2649,N_1445);
nor U5237 (N_5237,N_2857,N_1382);
xor U5238 (N_5238,N_2369,N_471);
or U5239 (N_5239,N_2475,N_178);
xnor U5240 (N_5240,N_902,N_1738);
and U5241 (N_5241,N_64,N_1257);
nand U5242 (N_5242,N_2408,N_1423);
xnor U5243 (N_5243,N_600,N_1775);
or U5244 (N_5244,N_200,N_1150);
nor U5245 (N_5245,N_1583,N_1918);
xor U5246 (N_5246,N_1925,N_93);
xor U5247 (N_5247,N_1356,N_2625);
nand U5248 (N_5248,N_393,N_366);
or U5249 (N_5249,N_1861,N_2132);
and U5250 (N_5250,N_2251,N_339);
nor U5251 (N_5251,N_816,N_157);
nand U5252 (N_5252,N_2182,N_1163);
or U5253 (N_5253,N_152,N_456);
nor U5254 (N_5254,N_2814,N_1611);
or U5255 (N_5255,N_1935,N_2597);
nor U5256 (N_5256,N_667,N_34);
and U5257 (N_5257,N_302,N_2028);
nand U5258 (N_5258,N_2387,N_2457);
nand U5259 (N_5259,N_1304,N_2404);
xnor U5260 (N_5260,N_2492,N_1716);
xor U5261 (N_5261,N_2736,N_77);
and U5262 (N_5262,N_2769,N_599);
nand U5263 (N_5263,N_1155,N_555);
and U5264 (N_5264,N_2754,N_1858);
nor U5265 (N_5265,N_2713,N_2254);
nand U5266 (N_5266,N_209,N_2054);
xor U5267 (N_5267,N_459,N_292);
or U5268 (N_5268,N_2626,N_216);
or U5269 (N_5269,N_389,N_1792);
and U5270 (N_5270,N_1932,N_1750);
xor U5271 (N_5271,N_1205,N_1624);
or U5272 (N_5272,N_2472,N_486);
and U5273 (N_5273,N_2996,N_1561);
or U5274 (N_5274,N_230,N_629);
nand U5275 (N_5275,N_2809,N_607);
and U5276 (N_5276,N_614,N_139);
xor U5277 (N_5277,N_1111,N_579);
or U5278 (N_5278,N_860,N_2283);
and U5279 (N_5279,N_215,N_662);
or U5280 (N_5280,N_889,N_2824);
or U5281 (N_5281,N_1398,N_1630);
nor U5282 (N_5282,N_386,N_933);
xnor U5283 (N_5283,N_1634,N_1739);
or U5284 (N_5284,N_1174,N_2227);
nand U5285 (N_5285,N_2202,N_2510);
nand U5286 (N_5286,N_2914,N_1183);
nand U5287 (N_5287,N_489,N_181);
nand U5288 (N_5288,N_1444,N_2624);
or U5289 (N_5289,N_459,N_361);
nor U5290 (N_5290,N_2103,N_1969);
nor U5291 (N_5291,N_18,N_2324);
nand U5292 (N_5292,N_1467,N_1470);
nand U5293 (N_5293,N_1994,N_1151);
or U5294 (N_5294,N_9,N_2773);
or U5295 (N_5295,N_2839,N_779);
xnor U5296 (N_5296,N_1304,N_2680);
or U5297 (N_5297,N_2746,N_2208);
nand U5298 (N_5298,N_870,N_2640);
and U5299 (N_5299,N_844,N_2493);
or U5300 (N_5300,N_1737,N_2375);
xor U5301 (N_5301,N_2831,N_1483);
nand U5302 (N_5302,N_1110,N_2797);
and U5303 (N_5303,N_368,N_2698);
or U5304 (N_5304,N_126,N_2870);
xnor U5305 (N_5305,N_631,N_1265);
nand U5306 (N_5306,N_1864,N_2833);
and U5307 (N_5307,N_2502,N_2841);
nor U5308 (N_5308,N_836,N_2462);
or U5309 (N_5309,N_2075,N_141);
xor U5310 (N_5310,N_213,N_1181);
nor U5311 (N_5311,N_1207,N_2627);
xor U5312 (N_5312,N_1212,N_2169);
xnor U5313 (N_5313,N_793,N_1917);
xnor U5314 (N_5314,N_2254,N_1884);
nor U5315 (N_5315,N_1573,N_359);
nor U5316 (N_5316,N_1734,N_339);
or U5317 (N_5317,N_1745,N_1792);
nand U5318 (N_5318,N_487,N_1173);
xnor U5319 (N_5319,N_369,N_1129);
nand U5320 (N_5320,N_259,N_63);
nand U5321 (N_5321,N_527,N_2483);
xor U5322 (N_5322,N_31,N_32);
xnor U5323 (N_5323,N_383,N_12);
nor U5324 (N_5324,N_741,N_2485);
xor U5325 (N_5325,N_820,N_2377);
and U5326 (N_5326,N_1394,N_1493);
or U5327 (N_5327,N_329,N_1340);
nand U5328 (N_5328,N_936,N_1797);
nand U5329 (N_5329,N_2429,N_904);
and U5330 (N_5330,N_1158,N_2887);
xnor U5331 (N_5331,N_125,N_888);
xor U5332 (N_5332,N_114,N_1602);
nor U5333 (N_5333,N_841,N_2958);
and U5334 (N_5334,N_914,N_1265);
xor U5335 (N_5335,N_2591,N_2406);
or U5336 (N_5336,N_2993,N_2497);
or U5337 (N_5337,N_2722,N_57);
and U5338 (N_5338,N_211,N_794);
or U5339 (N_5339,N_2678,N_1108);
or U5340 (N_5340,N_332,N_758);
and U5341 (N_5341,N_1281,N_419);
xor U5342 (N_5342,N_285,N_1367);
or U5343 (N_5343,N_445,N_572);
and U5344 (N_5344,N_695,N_2397);
or U5345 (N_5345,N_2946,N_2386);
nor U5346 (N_5346,N_1467,N_418);
or U5347 (N_5347,N_2002,N_627);
nand U5348 (N_5348,N_1546,N_1110);
and U5349 (N_5349,N_945,N_2595);
xnor U5350 (N_5350,N_82,N_2195);
nor U5351 (N_5351,N_2970,N_2495);
nor U5352 (N_5352,N_2140,N_1383);
nor U5353 (N_5353,N_2224,N_2519);
and U5354 (N_5354,N_2756,N_1606);
xnor U5355 (N_5355,N_964,N_1337);
or U5356 (N_5356,N_2272,N_1434);
nand U5357 (N_5357,N_2799,N_404);
xor U5358 (N_5358,N_2745,N_129);
nor U5359 (N_5359,N_1183,N_564);
or U5360 (N_5360,N_593,N_2511);
nand U5361 (N_5361,N_1658,N_626);
nand U5362 (N_5362,N_2699,N_709);
or U5363 (N_5363,N_1026,N_2867);
nand U5364 (N_5364,N_863,N_906);
nor U5365 (N_5365,N_2279,N_2180);
nor U5366 (N_5366,N_432,N_1917);
and U5367 (N_5367,N_427,N_24);
nor U5368 (N_5368,N_2235,N_1807);
and U5369 (N_5369,N_1714,N_1243);
nor U5370 (N_5370,N_2554,N_2136);
xnor U5371 (N_5371,N_1342,N_1512);
or U5372 (N_5372,N_2482,N_20);
nand U5373 (N_5373,N_488,N_876);
nor U5374 (N_5374,N_1354,N_233);
and U5375 (N_5375,N_1653,N_2033);
and U5376 (N_5376,N_1452,N_2327);
or U5377 (N_5377,N_1391,N_2227);
and U5378 (N_5378,N_943,N_2178);
or U5379 (N_5379,N_2709,N_2300);
nand U5380 (N_5380,N_2835,N_2202);
and U5381 (N_5381,N_1625,N_575);
nand U5382 (N_5382,N_1435,N_2026);
and U5383 (N_5383,N_1617,N_2275);
xnor U5384 (N_5384,N_118,N_254);
nand U5385 (N_5385,N_1958,N_1422);
nor U5386 (N_5386,N_1838,N_2297);
xnor U5387 (N_5387,N_2483,N_1192);
nand U5388 (N_5388,N_800,N_546);
and U5389 (N_5389,N_2967,N_1628);
and U5390 (N_5390,N_2375,N_2780);
and U5391 (N_5391,N_138,N_1580);
and U5392 (N_5392,N_1842,N_1357);
or U5393 (N_5393,N_2126,N_1019);
xnor U5394 (N_5394,N_952,N_1405);
or U5395 (N_5395,N_2133,N_1438);
nor U5396 (N_5396,N_1630,N_1408);
and U5397 (N_5397,N_572,N_123);
xnor U5398 (N_5398,N_2796,N_2393);
or U5399 (N_5399,N_1685,N_639);
or U5400 (N_5400,N_312,N_2665);
xnor U5401 (N_5401,N_2480,N_149);
xor U5402 (N_5402,N_1107,N_565);
nor U5403 (N_5403,N_2116,N_2256);
nand U5404 (N_5404,N_609,N_1592);
nand U5405 (N_5405,N_2144,N_886);
nor U5406 (N_5406,N_2651,N_2429);
nand U5407 (N_5407,N_2981,N_13);
nand U5408 (N_5408,N_259,N_1516);
and U5409 (N_5409,N_163,N_2645);
nor U5410 (N_5410,N_2206,N_2653);
nand U5411 (N_5411,N_722,N_1158);
nor U5412 (N_5412,N_484,N_2502);
nor U5413 (N_5413,N_2089,N_546);
nand U5414 (N_5414,N_2957,N_725);
or U5415 (N_5415,N_124,N_2989);
and U5416 (N_5416,N_131,N_478);
nand U5417 (N_5417,N_2500,N_908);
xnor U5418 (N_5418,N_775,N_96);
or U5419 (N_5419,N_2492,N_2364);
or U5420 (N_5420,N_204,N_2354);
xor U5421 (N_5421,N_2043,N_249);
or U5422 (N_5422,N_500,N_2557);
and U5423 (N_5423,N_964,N_1610);
or U5424 (N_5424,N_1923,N_2336);
nor U5425 (N_5425,N_1528,N_457);
nor U5426 (N_5426,N_335,N_2073);
nand U5427 (N_5427,N_1259,N_1481);
nor U5428 (N_5428,N_1134,N_969);
nor U5429 (N_5429,N_338,N_1125);
nor U5430 (N_5430,N_2753,N_1060);
and U5431 (N_5431,N_1694,N_1842);
xnor U5432 (N_5432,N_2276,N_1597);
and U5433 (N_5433,N_2148,N_1944);
or U5434 (N_5434,N_1972,N_2213);
or U5435 (N_5435,N_794,N_1456);
or U5436 (N_5436,N_1705,N_1453);
xnor U5437 (N_5437,N_1735,N_2416);
xor U5438 (N_5438,N_2610,N_2812);
xor U5439 (N_5439,N_565,N_1295);
and U5440 (N_5440,N_229,N_2591);
and U5441 (N_5441,N_328,N_1159);
nor U5442 (N_5442,N_176,N_2006);
xor U5443 (N_5443,N_2927,N_1369);
xnor U5444 (N_5444,N_990,N_2057);
and U5445 (N_5445,N_2173,N_554);
nor U5446 (N_5446,N_748,N_698);
nor U5447 (N_5447,N_2711,N_2246);
nor U5448 (N_5448,N_438,N_1282);
or U5449 (N_5449,N_1231,N_1314);
nor U5450 (N_5450,N_122,N_1412);
nor U5451 (N_5451,N_2745,N_1374);
xor U5452 (N_5452,N_1195,N_1205);
nor U5453 (N_5453,N_143,N_2472);
xnor U5454 (N_5454,N_536,N_1205);
nand U5455 (N_5455,N_1416,N_2358);
xor U5456 (N_5456,N_1833,N_1089);
xor U5457 (N_5457,N_202,N_1627);
nor U5458 (N_5458,N_2553,N_1065);
nand U5459 (N_5459,N_1767,N_2026);
and U5460 (N_5460,N_1980,N_941);
nor U5461 (N_5461,N_1099,N_317);
nand U5462 (N_5462,N_2507,N_992);
nor U5463 (N_5463,N_2827,N_1092);
nand U5464 (N_5464,N_221,N_1340);
nor U5465 (N_5465,N_2173,N_1500);
or U5466 (N_5466,N_893,N_224);
or U5467 (N_5467,N_1552,N_2565);
nand U5468 (N_5468,N_2032,N_608);
and U5469 (N_5469,N_71,N_1205);
or U5470 (N_5470,N_1090,N_1493);
and U5471 (N_5471,N_1772,N_818);
or U5472 (N_5472,N_1713,N_2520);
or U5473 (N_5473,N_1181,N_1489);
xnor U5474 (N_5474,N_1531,N_2869);
nand U5475 (N_5475,N_1985,N_2187);
and U5476 (N_5476,N_2977,N_66);
nand U5477 (N_5477,N_626,N_2688);
and U5478 (N_5478,N_1082,N_2518);
nand U5479 (N_5479,N_432,N_1713);
nand U5480 (N_5480,N_2650,N_2678);
xor U5481 (N_5481,N_495,N_1753);
xor U5482 (N_5482,N_112,N_818);
nor U5483 (N_5483,N_2021,N_2030);
nand U5484 (N_5484,N_405,N_2551);
xnor U5485 (N_5485,N_96,N_821);
and U5486 (N_5486,N_482,N_1894);
and U5487 (N_5487,N_2734,N_1819);
xnor U5488 (N_5488,N_1374,N_2012);
xnor U5489 (N_5489,N_528,N_132);
and U5490 (N_5490,N_2758,N_2429);
and U5491 (N_5491,N_1838,N_1385);
nand U5492 (N_5492,N_1495,N_2212);
or U5493 (N_5493,N_2531,N_2147);
nor U5494 (N_5494,N_413,N_902);
nor U5495 (N_5495,N_298,N_436);
xnor U5496 (N_5496,N_2081,N_177);
xor U5497 (N_5497,N_1748,N_425);
nand U5498 (N_5498,N_2983,N_2837);
and U5499 (N_5499,N_1323,N_1494);
and U5500 (N_5500,N_934,N_982);
nand U5501 (N_5501,N_224,N_790);
nor U5502 (N_5502,N_96,N_1970);
or U5503 (N_5503,N_1323,N_2091);
nor U5504 (N_5504,N_1311,N_2198);
xor U5505 (N_5505,N_2953,N_1807);
nor U5506 (N_5506,N_2843,N_2233);
nand U5507 (N_5507,N_1173,N_34);
and U5508 (N_5508,N_2392,N_1423);
xor U5509 (N_5509,N_602,N_2197);
or U5510 (N_5510,N_2597,N_1807);
or U5511 (N_5511,N_869,N_1707);
and U5512 (N_5512,N_726,N_2901);
xor U5513 (N_5513,N_2645,N_2049);
nand U5514 (N_5514,N_975,N_2683);
nor U5515 (N_5515,N_2041,N_2004);
xnor U5516 (N_5516,N_733,N_1881);
and U5517 (N_5517,N_940,N_2818);
nand U5518 (N_5518,N_335,N_2864);
and U5519 (N_5519,N_1855,N_1066);
or U5520 (N_5520,N_2198,N_1701);
or U5521 (N_5521,N_1777,N_80);
nor U5522 (N_5522,N_950,N_147);
and U5523 (N_5523,N_1184,N_1359);
xnor U5524 (N_5524,N_2444,N_1183);
xor U5525 (N_5525,N_84,N_2006);
nand U5526 (N_5526,N_2120,N_2055);
or U5527 (N_5527,N_1650,N_335);
or U5528 (N_5528,N_1085,N_2359);
nand U5529 (N_5529,N_1445,N_980);
xnor U5530 (N_5530,N_2730,N_2471);
nand U5531 (N_5531,N_108,N_487);
and U5532 (N_5532,N_1222,N_2193);
or U5533 (N_5533,N_2898,N_510);
and U5534 (N_5534,N_1229,N_133);
nor U5535 (N_5535,N_2040,N_521);
nand U5536 (N_5536,N_1153,N_571);
xor U5537 (N_5537,N_2380,N_539);
and U5538 (N_5538,N_1302,N_2922);
and U5539 (N_5539,N_148,N_2834);
xor U5540 (N_5540,N_2502,N_2057);
nand U5541 (N_5541,N_2729,N_2169);
xor U5542 (N_5542,N_896,N_1895);
or U5543 (N_5543,N_110,N_1652);
and U5544 (N_5544,N_16,N_2852);
nand U5545 (N_5545,N_1797,N_947);
and U5546 (N_5546,N_2503,N_365);
and U5547 (N_5547,N_1805,N_719);
nand U5548 (N_5548,N_1985,N_709);
and U5549 (N_5549,N_2369,N_484);
and U5550 (N_5550,N_1872,N_1236);
and U5551 (N_5551,N_1025,N_2148);
nor U5552 (N_5552,N_2580,N_648);
or U5553 (N_5553,N_2686,N_2216);
or U5554 (N_5554,N_118,N_1619);
and U5555 (N_5555,N_1293,N_1837);
xnor U5556 (N_5556,N_2615,N_851);
nand U5557 (N_5557,N_2044,N_962);
or U5558 (N_5558,N_841,N_972);
or U5559 (N_5559,N_489,N_2611);
or U5560 (N_5560,N_666,N_209);
or U5561 (N_5561,N_139,N_2610);
and U5562 (N_5562,N_194,N_2804);
nand U5563 (N_5563,N_1046,N_665);
xor U5564 (N_5564,N_1325,N_873);
and U5565 (N_5565,N_2982,N_1923);
xor U5566 (N_5566,N_1152,N_341);
or U5567 (N_5567,N_2825,N_2357);
and U5568 (N_5568,N_2231,N_719);
or U5569 (N_5569,N_1732,N_310);
or U5570 (N_5570,N_437,N_1982);
nand U5571 (N_5571,N_789,N_1859);
and U5572 (N_5572,N_2594,N_1954);
nor U5573 (N_5573,N_2435,N_203);
nor U5574 (N_5574,N_1135,N_1652);
nand U5575 (N_5575,N_521,N_828);
xor U5576 (N_5576,N_729,N_1127);
nand U5577 (N_5577,N_2676,N_1957);
nor U5578 (N_5578,N_1252,N_2029);
xor U5579 (N_5579,N_2879,N_1937);
nand U5580 (N_5580,N_2412,N_920);
nor U5581 (N_5581,N_1891,N_2529);
nor U5582 (N_5582,N_1225,N_490);
nor U5583 (N_5583,N_2824,N_2468);
or U5584 (N_5584,N_425,N_2735);
nand U5585 (N_5585,N_651,N_973);
or U5586 (N_5586,N_1884,N_1441);
nand U5587 (N_5587,N_97,N_1750);
xnor U5588 (N_5588,N_2637,N_278);
xor U5589 (N_5589,N_1763,N_2550);
nand U5590 (N_5590,N_1044,N_125);
or U5591 (N_5591,N_634,N_341);
xor U5592 (N_5592,N_204,N_705);
or U5593 (N_5593,N_776,N_1860);
and U5594 (N_5594,N_1160,N_405);
xor U5595 (N_5595,N_2126,N_2536);
or U5596 (N_5596,N_1123,N_2489);
nor U5597 (N_5597,N_2432,N_2773);
and U5598 (N_5598,N_984,N_2338);
or U5599 (N_5599,N_819,N_905);
nor U5600 (N_5600,N_1823,N_365);
nor U5601 (N_5601,N_1540,N_2220);
or U5602 (N_5602,N_2641,N_366);
and U5603 (N_5603,N_771,N_1871);
xor U5604 (N_5604,N_1014,N_264);
or U5605 (N_5605,N_1005,N_2681);
nor U5606 (N_5606,N_2944,N_838);
and U5607 (N_5607,N_1651,N_1890);
nor U5608 (N_5608,N_1817,N_1497);
nand U5609 (N_5609,N_2602,N_654);
xnor U5610 (N_5610,N_990,N_2688);
nor U5611 (N_5611,N_2102,N_1089);
and U5612 (N_5612,N_538,N_1481);
nand U5613 (N_5613,N_17,N_965);
nor U5614 (N_5614,N_817,N_1147);
and U5615 (N_5615,N_2790,N_677);
xnor U5616 (N_5616,N_2273,N_593);
nor U5617 (N_5617,N_1273,N_2810);
and U5618 (N_5618,N_1882,N_1178);
or U5619 (N_5619,N_157,N_2443);
nand U5620 (N_5620,N_1718,N_791);
nor U5621 (N_5621,N_2606,N_1120);
nand U5622 (N_5622,N_1240,N_2360);
and U5623 (N_5623,N_1254,N_1386);
nor U5624 (N_5624,N_1089,N_1336);
or U5625 (N_5625,N_1884,N_427);
or U5626 (N_5626,N_1067,N_1847);
nor U5627 (N_5627,N_1920,N_297);
or U5628 (N_5628,N_1850,N_1134);
nand U5629 (N_5629,N_2446,N_1947);
and U5630 (N_5630,N_862,N_525);
nor U5631 (N_5631,N_2961,N_2937);
or U5632 (N_5632,N_1283,N_46);
and U5633 (N_5633,N_2402,N_801);
nor U5634 (N_5634,N_556,N_2873);
nand U5635 (N_5635,N_1120,N_929);
nor U5636 (N_5636,N_968,N_1951);
nor U5637 (N_5637,N_1977,N_184);
and U5638 (N_5638,N_2832,N_1370);
xor U5639 (N_5639,N_2240,N_852);
nand U5640 (N_5640,N_825,N_2402);
nor U5641 (N_5641,N_2704,N_1860);
and U5642 (N_5642,N_18,N_720);
or U5643 (N_5643,N_1257,N_1385);
or U5644 (N_5644,N_826,N_1005);
and U5645 (N_5645,N_2001,N_1254);
nand U5646 (N_5646,N_1045,N_1538);
nor U5647 (N_5647,N_1326,N_598);
and U5648 (N_5648,N_2460,N_2828);
and U5649 (N_5649,N_1114,N_2621);
and U5650 (N_5650,N_2635,N_2598);
nor U5651 (N_5651,N_1087,N_2601);
or U5652 (N_5652,N_553,N_613);
nor U5653 (N_5653,N_2474,N_1470);
or U5654 (N_5654,N_347,N_1735);
or U5655 (N_5655,N_2209,N_182);
nor U5656 (N_5656,N_1598,N_600);
nor U5657 (N_5657,N_1862,N_2614);
and U5658 (N_5658,N_1087,N_1672);
or U5659 (N_5659,N_1446,N_618);
nor U5660 (N_5660,N_848,N_1156);
nor U5661 (N_5661,N_2284,N_295);
xor U5662 (N_5662,N_747,N_2662);
and U5663 (N_5663,N_1390,N_2619);
xnor U5664 (N_5664,N_1263,N_1581);
nor U5665 (N_5665,N_2023,N_1846);
and U5666 (N_5666,N_296,N_2026);
nand U5667 (N_5667,N_2297,N_2611);
nand U5668 (N_5668,N_630,N_2180);
nor U5669 (N_5669,N_2027,N_1948);
xnor U5670 (N_5670,N_1123,N_1676);
nand U5671 (N_5671,N_1490,N_2532);
and U5672 (N_5672,N_1490,N_699);
and U5673 (N_5673,N_60,N_2831);
or U5674 (N_5674,N_768,N_2471);
or U5675 (N_5675,N_2643,N_2011);
or U5676 (N_5676,N_586,N_2791);
xor U5677 (N_5677,N_2868,N_383);
nor U5678 (N_5678,N_2297,N_1033);
and U5679 (N_5679,N_2616,N_4);
nor U5680 (N_5680,N_1974,N_1657);
or U5681 (N_5681,N_1787,N_2768);
nand U5682 (N_5682,N_2493,N_192);
or U5683 (N_5683,N_2505,N_2085);
or U5684 (N_5684,N_557,N_546);
xnor U5685 (N_5685,N_542,N_918);
and U5686 (N_5686,N_1346,N_2045);
and U5687 (N_5687,N_1234,N_2859);
and U5688 (N_5688,N_2199,N_1284);
xnor U5689 (N_5689,N_1442,N_2790);
nor U5690 (N_5690,N_1221,N_2934);
or U5691 (N_5691,N_192,N_976);
and U5692 (N_5692,N_2350,N_1037);
or U5693 (N_5693,N_1873,N_2845);
xor U5694 (N_5694,N_232,N_1498);
xnor U5695 (N_5695,N_317,N_450);
xor U5696 (N_5696,N_2379,N_2124);
and U5697 (N_5697,N_557,N_2944);
and U5698 (N_5698,N_2598,N_1059);
nand U5699 (N_5699,N_1930,N_2905);
and U5700 (N_5700,N_1780,N_394);
xor U5701 (N_5701,N_2036,N_1812);
or U5702 (N_5702,N_1523,N_1696);
nand U5703 (N_5703,N_2179,N_2218);
nor U5704 (N_5704,N_2264,N_509);
nor U5705 (N_5705,N_2026,N_654);
nand U5706 (N_5706,N_2740,N_2347);
nand U5707 (N_5707,N_657,N_2200);
and U5708 (N_5708,N_1040,N_1685);
nor U5709 (N_5709,N_44,N_2791);
nand U5710 (N_5710,N_2772,N_610);
nand U5711 (N_5711,N_1598,N_1768);
xor U5712 (N_5712,N_2918,N_373);
nor U5713 (N_5713,N_2463,N_787);
and U5714 (N_5714,N_1387,N_436);
or U5715 (N_5715,N_342,N_412);
nand U5716 (N_5716,N_2319,N_1708);
nor U5717 (N_5717,N_545,N_728);
or U5718 (N_5718,N_2140,N_2938);
or U5719 (N_5719,N_928,N_303);
nand U5720 (N_5720,N_253,N_2200);
nand U5721 (N_5721,N_2124,N_1476);
or U5722 (N_5722,N_378,N_1818);
xor U5723 (N_5723,N_1884,N_1633);
xnor U5724 (N_5724,N_2830,N_746);
nor U5725 (N_5725,N_1144,N_2304);
or U5726 (N_5726,N_240,N_560);
nand U5727 (N_5727,N_2852,N_369);
nand U5728 (N_5728,N_2827,N_1101);
xnor U5729 (N_5729,N_1168,N_733);
and U5730 (N_5730,N_157,N_1392);
nand U5731 (N_5731,N_1650,N_634);
or U5732 (N_5732,N_1885,N_1992);
or U5733 (N_5733,N_362,N_1152);
or U5734 (N_5734,N_2412,N_1653);
and U5735 (N_5735,N_2180,N_1110);
nand U5736 (N_5736,N_2721,N_2682);
xor U5737 (N_5737,N_1097,N_520);
xor U5738 (N_5738,N_973,N_300);
nor U5739 (N_5739,N_602,N_567);
nand U5740 (N_5740,N_1766,N_1824);
and U5741 (N_5741,N_1584,N_2875);
nand U5742 (N_5742,N_96,N_873);
and U5743 (N_5743,N_1736,N_1340);
nand U5744 (N_5744,N_375,N_1735);
nor U5745 (N_5745,N_1134,N_1053);
and U5746 (N_5746,N_1333,N_387);
or U5747 (N_5747,N_2174,N_197);
nand U5748 (N_5748,N_562,N_1058);
xor U5749 (N_5749,N_1366,N_895);
nor U5750 (N_5750,N_2634,N_2780);
and U5751 (N_5751,N_1072,N_641);
nand U5752 (N_5752,N_661,N_2224);
xnor U5753 (N_5753,N_147,N_2657);
and U5754 (N_5754,N_2345,N_872);
and U5755 (N_5755,N_2338,N_132);
and U5756 (N_5756,N_1064,N_334);
xor U5757 (N_5757,N_1329,N_1684);
nor U5758 (N_5758,N_2276,N_835);
nor U5759 (N_5759,N_993,N_181);
nand U5760 (N_5760,N_488,N_883);
nor U5761 (N_5761,N_2300,N_1787);
and U5762 (N_5762,N_2258,N_2002);
nor U5763 (N_5763,N_1333,N_174);
or U5764 (N_5764,N_1579,N_2231);
or U5765 (N_5765,N_662,N_371);
and U5766 (N_5766,N_2664,N_2389);
nor U5767 (N_5767,N_2704,N_2591);
xor U5768 (N_5768,N_1565,N_1727);
xor U5769 (N_5769,N_2229,N_1478);
xnor U5770 (N_5770,N_657,N_593);
or U5771 (N_5771,N_1411,N_1570);
nor U5772 (N_5772,N_1864,N_898);
nand U5773 (N_5773,N_1499,N_1227);
and U5774 (N_5774,N_1603,N_2010);
and U5775 (N_5775,N_1130,N_796);
or U5776 (N_5776,N_1293,N_2015);
and U5777 (N_5777,N_2433,N_168);
and U5778 (N_5778,N_2633,N_2038);
xor U5779 (N_5779,N_1129,N_874);
and U5780 (N_5780,N_2044,N_1782);
and U5781 (N_5781,N_765,N_1735);
nor U5782 (N_5782,N_2098,N_1408);
and U5783 (N_5783,N_700,N_1490);
nand U5784 (N_5784,N_2647,N_2241);
nand U5785 (N_5785,N_392,N_599);
and U5786 (N_5786,N_1878,N_1288);
nand U5787 (N_5787,N_472,N_1224);
and U5788 (N_5788,N_667,N_143);
and U5789 (N_5789,N_2935,N_146);
xor U5790 (N_5790,N_2064,N_2950);
or U5791 (N_5791,N_651,N_1022);
nand U5792 (N_5792,N_2311,N_65);
xnor U5793 (N_5793,N_1202,N_584);
xor U5794 (N_5794,N_2693,N_201);
nand U5795 (N_5795,N_1333,N_1832);
nor U5796 (N_5796,N_186,N_315);
and U5797 (N_5797,N_1795,N_685);
nand U5798 (N_5798,N_106,N_665);
and U5799 (N_5799,N_2323,N_1966);
and U5800 (N_5800,N_2645,N_1754);
or U5801 (N_5801,N_1065,N_255);
xnor U5802 (N_5802,N_1381,N_2596);
or U5803 (N_5803,N_1008,N_1199);
xnor U5804 (N_5804,N_2455,N_1648);
nand U5805 (N_5805,N_1350,N_2961);
nand U5806 (N_5806,N_1514,N_1308);
and U5807 (N_5807,N_749,N_1554);
and U5808 (N_5808,N_1482,N_2233);
and U5809 (N_5809,N_553,N_2714);
xnor U5810 (N_5810,N_655,N_1828);
xor U5811 (N_5811,N_2092,N_1046);
nor U5812 (N_5812,N_1059,N_1698);
and U5813 (N_5813,N_2650,N_2153);
nor U5814 (N_5814,N_478,N_2028);
xnor U5815 (N_5815,N_1300,N_1031);
xnor U5816 (N_5816,N_2120,N_1557);
nand U5817 (N_5817,N_961,N_140);
nor U5818 (N_5818,N_2137,N_2032);
nor U5819 (N_5819,N_224,N_1866);
nor U5820 (N_5820,N_1575,N_2228);
and U5821 (N_5821,N_1742,N_674);
or U5822 (N_5822,N_2705,N_2572);
or U5823 (N_5823,N_2153,N_2064);
and U5824 (N_5824,N_631,N_672);
nor U5825 (N_5825,N_2602,N_370);
nand U5826 (N_5826,N_1148,N_290);
nor U5827 (N_5827,N_2591,N_129);
nand U5828 (N_5828,N_1945,N_255);
nor U5829 (N_5829,N_287,N_2670);
nand U5830 (N_5830,N_2782,N_953);
and U5831 (N_5831,N_2020,N_1827);
nor U5832 (N_5832,N_1835,N_2532);
and U5833 (N_5833,N_1264,N_11);
or U5834 (N_5834,N_634,N_1706);
xnor U5835 (N_5835,N_1215,N_1547);
nand U5836 (N_5836,N_147,N_1780);
xor U5837 (N_5837,N_684,N_1748);
nor U5838 (N_5838,N_2011,N_326);
nand U5839 (N_5839,N_1885,N_158);
nand U5840 (N_5840,N_1061,N_55);
xnor U5841 (N_5841,N_1421,N_2583);
or U5842 (N_5842,N_2366,N_1968);
nand U5843 (N_5843,N_362,N_752);
nand U5844 (N_5844,N_2329,N_1876);
and U5845 (N_5845,N_2357,N_424);
or U5846 (N_5846,N_702,N_2791);
or U5847 (N_5847,N_769,N_783);
nand U5848 (N_5848,N_283,N_2634);
nand U5849 (N_5849,N_347,N_2510);
nor U5850 (N_5850,N_568,N_2129);
xnor U5851 (N_5851,N_2036,N_1311);
xnor U5852 (N_5852,N_1095,N_2593);
nor U5853 (N_5853,N_1859,N_2095);
nor U5854 (N_5854,N_437,N_472);
nand U5855 (N_5855,N_1226,N_1303);
xor U5856 (N_5856,N_660,N_1236);
xor U5857 (N_5857,N_2073,N_788);
xor U5858 (N_5858,N_315,N_449);
nand U5859 (N_5859,N_156,N_1869);
nor U5860 (N_5860,N_1250,N_1747);
nand U5861 (N_5861,N_724,N_1961);
and U5862 (N_5862,N_2,N_2551);
xnor U5863 (N_5863,N_1387,N_429);
nor U5864 (N_5864,N_1213,N_2411);
and U5865 (N_5865,N_2808,N_646);
nand U5866 (N_5866,N_882,N_202);
or U5867 (N_5867,N_1399,N_1579);
xor U5868 (N_5868,N_1605,N_2600);
or U5869 (N_5869,N_1914,N_1122);
and U5870 (N_5870,N_2739,N_1940);
nor U5871 (N_5871,N_2691,N_2678);
xor U5872 (N_5872,N_2255,N_2298);
xnor U5873 (N_5873,N_795,N_2491);
nand U5874 (N_5874,N_2520,N_495);
xnor U5875 (N_5875,N_616,N_2064);
xnor U5876 (N_5876,N_596,N_2734);
and U5877 (N_5877,N_1616,N_2706);
or U5878 (N_5878,N_2987,N_952);
or U5879 (N_5879,N_2147,N_1985);
xnor U5880 (N_5880,N_1614,N_1844);
nor U5881 (N_5881,N_555,N_625);
nor U5882 (N_5882,N_1846,N_651);
or U5883 (N_5883,N_1123,N_1886);
and U5884 (N_5884,N_1054,N_1981);
xnor U5885 (N_5885,N_232,N_157);
nand U5886 (N_5886,N_1532,N_2322);
xor U5887 (N_5887,N_1803,N_2970);
or U5888 (N_5888,N_1986,N_1024);
xnor U5889 (N_5889,N_2201,N_2577);
nor U5890 (N_5890,N_787,N_2550);
or U5891 (N_5891,N_1916,N_720);
nand U5892 (N_5892,N_2900,N_2915);
and U5893 (N_5893,N_1443,N_27);
nor U5894 (N_5894,N_1940,N_1373);
xnor U5895 (N_5895,N_54,N_2893);
xnor U5896 (N_5896,N_692,N_1118);
nor U5897 (N_5897,N_549,N_502);
or U5898 (N_5898,N_1184,N_1280);
xor U5899 (N_5899,N_1465,N_2939);
xnor U5900 (N_5900,N_1284,N_1409);
and U5901 (N_5901,N_646,N_2253);
or U5902 (N_5902,N_2960,N_1291);
nand U5903 (N_5903,N_1191,N_118);
or U5904 (N_5904,N_363,N_2183);
nor U5905 (N_5905,N_1940,N_256);
xnor U5906 (N_5906,N_2424,N_328);
or U5907 (N_5907,N_1059,N_90);
and U5908 (N_5908,N_1903,N_1237);
nor U5909 (N_5909,N_2636,N_2933);
nand U5910 (N_5910,N_1300,N_2672);
nor U5911 (N_5911,N_828,N_1634);
or U5912 (N_5912,N_2031,N_637);
nor U5913 (N_5913,N_863,N_616);
xnor U5914 (N_5914,N_520,N_376);
nand U5915 (N_5915,N_2146,N_2762);
and U5916 (N_5916,N_1224,N_1100);
nor U5917 (N_5917,N_340,N_2311);
nor U5918 (N_5918,N_477,N_1295);
and U5919 (N_5919,N_1033,N_2515);
and U5920 (N_5920,N_2999,N_1531);
or U5921 (N_5921,N_1844,N_166);
nand U5922 (N_5922,N_1703,N_2957);
xor U5923 (N_5923,N_2815,N_1271);
xnor U5924 (N_5924,N_2042,N_1311);
nor U5925 (N_5925,N_1417,N_2695);
xnor U5926 (N_5926,N_1683,N_2465);
and U5927 (N_5927,N_1823,N_2400);
or U5928 (N_5928,N_2836,N_1096);
or U5929 (N_5929,N_1197,N_2129);
xnor U5930 (N_5930,N_1969,N_1319);
and U5931 (N_5931,N_1215,N_1256);
nand U5932 (N_5932,N_1007,N_2475);
or U5933 (N_5933,N_1229,N_1602);
nor U5934 (N_5934,N_2350,N_258);
nor U5935 (N_5935,N_2206,N_2453);
nand U5936 (N_5936,N_2708,N_2140);
nand U5937 (N_5937,N_1194,N_950);
xor U5938 (N_5938,N_2858,N_2291);
or U5939 (N_5939,N_1159,N_1643);
xor U5940 (N_5940,N_402,N_1083);
nand U5941 (N_5941,N_1973,N_2877);
nor U5942 (N_5942,N_728,N_12);
xnor U5943 (N_5943,N_142,N_894);
or U5944 (N_5944,N_465,N_1252);
xor U5945 (N_5945,N_167,N_2994);
xnor U5946 (N_5946,N_2508,N_663);
nor U5947 (N_5947,N_1364,N_1953);
and U5948 (N_5948,N_1981,N_2089);
or U5949 (N_5949,N_1645,N_2084);
nor U5950 (N_5950,N_1085,N_2566);
and U5951 (N_5951,N_2694,N_1651);
nor U5952 (N_5952,N_2750,N_1622);
nor U5953 (N_5953,N_79,N_1277);
or U5954 (N_5954,N_2478,N_1509);
nand U5955 (N_5955,N_1374,N_1231);
xor U5956 (N_5956,N_1641,N_266);
and U5957 (N_5957,N_2855,N_1516);
or U5958 (N_5958,N_1911,N_733);
or U5959 (N_5959,N_1104,N_1397);
and U5960 (N_5960,N_1650,N_1764);
nor U5961 (N_5961,N_2136,N_2271);
or U5962 (N_5962,N_2460,N_128);
xor U5963 (N_5963,N_727,N_1573);
and U5964 (N_5964,N_2074,N_409);
and U5965 (N_5965,N_2396,N_672);
nor U5966 (N_5966,N_471,N_844);
nand U5967 (N_5967,N_831,N_966);
or U5968 (N_5968,N_1015,N_2029);
or U5969 (N_5969,N_295,N_312);
or U5970 (N_5970,N_1545,N_2533);
and U5971 (N_5971,N_41,N_1346);
nor U5972 (N_5972,N_1079,N_2491);
xnor U5973 (N_5973,N_2035,N_2487);
or U5974 (N_5974,N_2572,N_2348);
or U5975 (N_5975,N_1592,N_1379);
nor U5976 (N_5976,N_2791,N_806);
xnor U5977 (N_5977,N_654,N_150);
xnor U5978 (N_5978,N_2090,N_2268);
nand U5979 (N_5979,N_2752,N_2153);
nor U5980 (N_5980,N_1087,N_2867);
nor U5981 (N_5981,N_2911,N_1903);
xnor U5982 (N_5982,N_530,N_1410);
or U5983 (N_5983,N_1651,N_2573);
and U5984 (N_5984,N_410,N_1870);
nand U5985 (N_5985,N_1874,N_29);
xor U5986 (N_5986,N_956,N_23);
and U5987 (N_5987,N_1227,N_2572);
and U5988 (N_5988,N_1544,N_2919);
nor U5989 (N_5989,N_2167,N_2395);
or U5990 (N_5990,N_2509,N_23);
and U5991 (N_5991,N_1300,N_2610);
xnor U5992 (N_5992,N_201,N_38);
xnor U5993 (N_5993,N_1538,N_2492);
nor U5994 (N_5994,N_2321,N_777);
nor U5995 (N_5995,N_167,N_1518);
or U5996 (N_5996,N_2777,N_595);
xnor U5997 (N_5997,N_171,N_183);
nor U5998 (N_5998,N_1513,N_2649);
xnor U5999 (N_5999,N_1940,N_1213);
nor U6000 (N_6000,N_5729,N_5206);
or U6001 (N_6001,N_4078,N_5725);
nor U6002 (N_6002,N_5466,N_4682);
nor U6003 (N_6003,N_4520,N_3062);
or U6004 (N_6004,N_4049,N_3572);
or U6005 (N_6005,N_5645,N_5652);
nor U6006 (N_6006,N_3316,N_3673);
nand U6007 (N_6007,N_4949,N_5872);
nor U6008 (N_6008,N_3751,N_4291);
nor U6009 (N_6009,N_4507,N_3594);
nand U6010 (N_6010,N_3386,N_4036);
xor U6011 (N_6011,N_4428,N_5903);
xnor U6012 (N_6012,N_3637,N_3325);
and U6013 (N_6013,N_4243,N_3873);
nor U6014 (N_6014,N_5785,N_3681);
nor U6015 (N_6015,N_3794,N_5797);
nor U6016 (N_6016,N_3631,N_3924);
xnor U6017 (N_6017,N_4936,N_3306);
xnor U6018 (N_6018,N_5748,N_5942);
and U6019 (N_6019,N_4994,N_5258);
or U6020 (N_6020,N_3584,N_3852);
or U6021 (N_6021,N_4090,N_4536);
nand U6022 (N_6022,N_4136,N_4726);
and U6023 (N_6023,N_3516,N_4177);
xor U6024 (N_6024,N_5231,N_3740);
and U6025 (N_6025,N_5602,N_4293);
nor U6026 (N_6026,N_5139,N_5861);
xor U6027 (N_6027,N_4494,N_4436);
and U6028 (N_6028,N_3095,N_4000);
or U6029 (N_6029,N_5863,N_5694);
and U6030 (N_6030,N_4691,N_3253);
or U6031 (N_6031,N_5036,N_5355);
and U6032 (N_6032,N_5562,N_3053);
nand U6033 (N_6033,N_5707,N_4330);
nor U6034 (N_6034,N_5289,N_3267);
or U6035 (N_6035,N_3546,N_3066);
xor U6036 (N_6036,N_5175,N_3091);
and U6037 (N_6037,N_4931,N_3570);
xnor U6038 (N_6038,N_4512,N_4085);
or U6039 (N_6039,N_3587,N_3919);
nor U6040 (N_6040,N_4781,N_4308);
xnor U6041 (N_6041,N_5757,N_5077);
nor U6042 (N_6042,N_4489,N_3636);
and U6043 (N_6043,N_5560,N_5712);
or U6044 (N_6044,N_3562,N_4877);
or U6045 (N_6045,N_5894,N_4445);
nand U6046 (N_6046,N_4688,N_5104);
xor U6047 (N_6047,N_5693,N_5255);
xor U6048 (N_6048,N_3170,N_3033);
xnor U6049 (N_6049,N_5957,N_4007);
or U6050 (N_6050,N_3159,N_4186);
xnor U6051 (N_6051,N_4527,N_5058);
nand U6052 (N_6052,N_5384,N_5333);
xnor U6053 (N_6053,N_3489,N_4582);
and U6054 (N_6054,N_4733,N_3865);
or U6055 (N_6055,N_5558,N_4805);
nor U6056 (N_6056,N_4895,N_3272);
nand U6057 (N_6057,N_5852,N_4125);
nor U6058 (N_6058,N_4277,N_3703);
and U6059 (N_6059,N_4980,N_3819);
or U6060 (N_6060,N_4411,N_4294);
nand U6061 (N_6061,N_3293,N_3204);
or U6062 (N_6062,N_4148,N_5349);
xnor U6063 (N_6063,N_3365,N_4939);
and U6064 (N_6064,N_5097,N_5897);
and U6065 (N_6065,N_4043,N_4273);
xor U6066 (N_6066,N_5492,N_3916);
and U6067 (N_6067,N_4453,N_3655);
nor U6068 (N_6068,N_3164,N_4075);
and U6069 (N_6069,N_4182,N_5163);
or U6070 (N_6070,N_4801,N_5598);
xnor U6071 (N_6071,N_4875,N_3944);
nor U6072 (N_6072,N_5284,N_5716);
nand U6073 (N_6073,N_4127,N_5904);
nor U6074 (N_6074,N_4959,N_4946);
nor U6075 (N_6075,N_3581,N_5969);
nand U6076 (N_6076,N_5345,N_5145);
nor U6077 (N_6077,N_3321,N_4260);
xnor U6078 (N_6078,N_4482,N_3123);
xnor U6079 (N_6079,N_5361,N_4619);
nand U6080 (N_6080,N_4162,N_3448);
xnor U6081 (N_6081,N_5478,N_5490);
xor U6082 (N_6082,N_3298,N_4855);
nand U6083 (N_6083,N_5322,N_3287);
xor U6084 (N_6084,N_5454,N_3447);
xor U6085 (N_6085,N_3592,N_3550);
and U6086 (N_6086,N_4361,N_5120);
and U6087 (N_6087,N_4033,N_5651);
and U6088 (N_6088,N_4888,N_5238);
nor U6089 (N_6089,N_5089,N_3140);
xor U6090 (N_6090,N_4560,N_4054);
or U6091 (N_6091,N_4181,N_3499);
or U6092 (N_6092,N_4005,N_5851);
nor U6093 (N_6093,N_3810,N_3798);
xor U6094 (N_6094,N_5224,N_5703);
or U6095 (N_6095,N_5477,N_5241);
nor U6096 (N_6096,N_3493,N_5338);
and U6097 (N_6097,N_3492,N_3881);
or U6098 (N_6098,N_4381,N_5252);
nand U6099 (N_6099,N_4350,N_5314);
or U6100 (N_6100,N_3741,N_5704);
nor U6101 (N_6101,N_4755,N_3925);
xnor U6102 (N_6102,N_4396,N_4504);
xnor U6103 (N_6103,N_3395,N_4832);
nand U6104 (N_6104,N_3978,N_3048);
and U6105 (N_6105,N_3989,N_3757);
or U6106 (N_6106,N_3509,N_5290);
xnor U6107 (N_6107,N_3464,N_4508);
and U6108 (N_6108,N_5798,N_3056);
nor U6109 (N_6109,N_5399,N_4544);
nand U6110 (N_6110,N_4571,N_4539);
nand U6111 (N_6111,N_3297,N_4803);
nor U6112 (N_6112,N_3407,N_3840);
xnor U6113 (N_6113,N_3472,N_5899);
xnor U6114 (N_6114,N_4267,N_3052);
xor U6115 (N_6115,N_4736,N_4095);
xor U6116 (N_6116,N_5268,N_5625);
nor U6117 (N_6117,N_4687,N_4395);
nor U6118 (N_6118,N_4584,N_4087);
xnor U6119 (N_6119,N_3735,N_4249);
nor U6120 (N_6120,N_4417,N_3228);
nand U6121 (N_6121,N_4552,N_4662);
or U6122 (N_6122,N_3884,N_3586);
xor U6123 (N_6123,N_5871,N_5391);
or U6124 (N_6124,N_4708,N_4140);
nand U6125 (N_6125,N_4768,N_3393);
or U6126 (N_6126,N_5211,N_3177);
nand U6127 (N_6127,N_4616,N_3427);
xor U6128 (N_6128,N_4187,N_4620);
xnor U6129 (N_6129,N_5012,N_3209);
xnor U6130 (N_6130,N_3027,N_5243);
nand U6131 (N_6131,N_4999,N_5291);
nor U6132 (N_6132,N_4548,N_4813);
nand U6133 (N_6133,N_5028,N_5321);
nor U6134 (N_6134,N_4029,N_5368);
or U6135 (N_6135,N_5074,N_4456);
xnor U6136 (N_6136,N_3108,N_3438);
nand U6137 (N_6137,N_5488,N_3877);
or U6138 (N_6138,N_3497,N_5441);
xor U6139 (N_6139,N_3281,N_3823);
nand U6140 (N_6140,N_3402,N_4339);
and U6141 (N_6141,N_4915,N_5075);
or U6142 (N_6142,N_5017,N_5582);
nand U6143 (N_6143,N_3670,N_5144);
or U6144 (N_6144,N_5730,N_4742);
nand U6145 (N_6145,N_4549,N_5468);
xnor U6146 (N_6146,N_3975,N_3397);
nor U6147 (N_6147,N_4357,N_5737);
and U6148 (N_6148,N_5439,N_3992);
nor U6149 (N_6149,N_4046,N_4851);
nor U6150 (N_6150,N_5022,N_5579);
or U6151 (N_6151,N_5829,N_3382);
nor U6152 (N_6152,N_3484,N_4252);
nand U6153 (N_6153,N_4618,N_5929);
and U6154 (N_6154,N_5496,N_4943);
and U6155 (N_6155,N_4869,N_5962);
or U6156 (N_6156,N_4909,N_5661);
xnor U6157 (N_6157,N_5822,N_3022);
nor U6158 (N_6158,N_5698,N_3433);
or U6159 (N_6159,N_3679,N_3582);
xnor U6160 (N_6160,N_5127,N_5029);
or U6161 (N_6161,N_4985,N_3471);
xnor U6162 (N_6162,N_3277,N_3400);
and U6163 (N_6163,N_3233,N_3363);
nor U6164 (N_6164,N_5953,N_5559);
xor U6165 (N_6165,N_3371,N_3351);
xor U6166 (N_6166,N_4759,N_4292);
xnor U6167 (N_6167,N_4522,N_4922);
nand U6168 (N_6168,N_3211,N_3032);
nor U6169 (N_6169,N_4689,N_4088);
nor U6170 (N_6170,N_5100,N_3947);
nand U6171 (N_6171,N_3901,N_5814);
or U6172 (N_6172,N_4656,N_4655);
nor U6173 (N_6173,N_3566,N_3791);
and U6174 (N_6174,N_4991,N_4463);
nand U6175 (N_6175,N_3050,N_3832);
xnor U6176 (N_6176,N_3892,N_5939);
nor U6177 (N_6177,N_5511,N_4315);
xnor U6178 (N_6178,N_4629,N_5323);
xnor U6179 (N_6179,N_5677,N_3934);
nor U6180 (N_6180,N_4421,N_3709);
or U6181 (N_6181,N_4810,N_3846);
nand U6182 (N_6182,N_5298,N_3428);
or U6183 (N_6183,N_3973,N_5763);
nand U6184 (N_6184,N_3307,N_5945);
or U6185 (N_6185,N_3767,N_4254);
and U6186 (N_6186,N_5997,N_5011);
nand U6187 (N_6187,N_4743,N_3031);
and U6188 (N_6188,N_5425,N_4327);
and U6189 (N_6189,N_5073,N_3906);
nand U6190 (N_6190,N_5801,N_4847);
nand U6191 (N_6191,N_4715,N_5586);
nand U6192 (N_6192,N_3990,N_3068);
xor U6193 (N_6193,N_3987,N_5394);
xnor U6194 (N_6194,N_3678,N_5620);
or U6195 (N_6195,N_3003,N_4573);
nor U6196 (N_6196,N_5691,N_3737);
xnor U6197 (N_6197,N_4150,N_5424);
and U6198 (N_6198,N_5644,N_3291);
nand U6199 (N_6199,N_4562,N_5843);
or U6200 (N_6200,N_4367,N_3800);
or U6201 (N_6201,N_5949,N_5180);
or U6202 (N_6202,N_4776,N_3559);
xnor U6203 (N_6203,N_5048,N_3324);
and U6204 (N_6204,N_3049,N_5001);
and U6205 (N_6205,N_3612,N_4849);
nor U6206 (N_6206,N_5970,N_4434);
or U6207 (N_6207,N_4823,N_3409);
and U6208 (N_6208,N_3792,N_3965);
and U6209 (N_6209,N_5156,N_5951);
nand U6210 (N_6210,N_3257,N_4626);
or U6211 (N_6211,N_5222,N_4022);
xnor U6212 (N_6212,N_3044,N_4201);
nor U6213 (N_6213,N_4156,N_4110);
nor U6214 (N_6214,N_4358,N_3651);
or U6215 (N_6215,N_3419,N_4826);
and U6216 (N_6216,N_5570,N_5989);
or U6217 (N_6217,N_5051,N_5160);
nand U6218 (N_6218,N_5606,N_4673);
nor U6219 (N_6219,N_5534,N_4338);
xnor U6220 (N_6220,N_5194,N_4019);
and U6221 (N_6221,N_3163,N_3743);
and U6222 (N_6222,N_5946,N_4961);
nand U6223 (N_6223,N_3208,N_5044);
xor U6224 (N_6224,N_5189,N_3949);
nand U6225 (N_6225,N_3976,N_5523);
and U6226 (N_6226,N_4280,N_5702);
nor U6227 (N_6227,N_3917,N_5084);
or U6228 (N_6228,N_5937,N_5250);
xnor U6229 (N_6229,N_3215,N_3970);
nand U6230 (N_6230,N_5383,N_3706);
xor U6231 (N_6231,N_5995,N_3701);
nor U6232 (N_6232,N_4163,N_4325);
or U6233 (N_6233,N_5616,N_4449);
and U6234 (N_6234,N_4468,N_3956);
nand U6235 (N_6235,N_3860,N_5738);
or U6236 (N_6236,N_3862,N_3756);
xnor U6237 (N_6237,N_5324,N_3436);
and U6238 (N_6238,N_4667,N_5902);
and U6239 (N_6239,N_4312,N_4380);
and U6240 (N_6240,N_5308,N_4950);
nor U6241 (N_6241,N_5706,N_3843);
or U6242 (N_6242,N_4023,N_5142);
xnor U6243 (N_6243,N_5393,N_5402);
and U6244 (N_6244,N_4918,N_3998);
xnor U6245 (N_6245,N_3654,N_5226);
nand U6246 (N_6246,N_4513,N_5799);
nand U6247 (N_6247,N_4606,N_4518);
and U6248 (N_6248,N_4712,N_3809);
nand U6249 (N_6249,N_3431,N_5283);
and U6250 (N_6250,N_3885,N_3274);
nor U6251 (N_6251,N_4757,N_4400);
xor U6252 (N_6252,N_3895,N_3912);
or U6253 (N_6253,N_4105,N_5524);
xor U6254 (N_6254,N_5448,N_3234);
nand U6255 (N_6255,N_4320,N_5068);
or U6256 (N_6256,N_4842,N_4942);
nand U6257 (N_6257,N_3197,N_3218);
nand U6258 (N_6258,N_4318,N_3959);
or U6259 (N_6259,N_3385,N_4214);
nor U6260 (N_6260,N_4890,N_3317);
xnor U6261 (N_6261,N_5791,N_5812);
and U6262 (N_6262,N_3094,N_4485);
nor U6263 (N_6263,N_3980,N_3092);
or U6264 (N_6264,N_4876,N_4223);
or U6265 (N_6265,N_3192,N_3597);
and U6266 (N_6266,N_5469,N_3165);
xnor U6267 (N_6267,N_3732,N_3129);
nor U6268 (N_6268,N_5143,N_3661);
and U6269 (N_6269,N_4542,N_3610);
xor U6270 (N_6270,N_3311,N_3974);
and U6271 (N_6271,N_3205,N_5171);
nand U6272 (N_6272,N_3888,N_5280);
nand U6273 (N_6273,N_4650,N_5889);
and U6274 (N_6274,N_3966,N_4916);
xor U6275 (N_6275,N_5491,N_5159);
or U6276 (N_6276,N_4501,N_4903);
nor U6277 (N_6277,N_3793,N_3485);
and U6278 (N_6278,N_4026,N_5943);
or U6279 (N_6279,N_3278,N_4506);
or U6280 (N_6280,N_5540,N_4818);
and U6281 (N_6281,N_3506,N_3721);
or U6282 (N_6282,N_4676,N_4885);
and U6283 (N_6283,N_5963,N_4464);
or U6284 (N_6284,N_3318,N_5958);
and U6285 (N_6285,N_3927,N_5952);
or U6286 (N_6286,N_5404,N_5619);
nand U6287 (N_6287,N_3951,N_4756);
or U6288 (N_6288,N_4824,N_4138);
xor U6289 (N_6289,N_3627,N_4372);
nand U6290 (N_6290,N_3065,N_4360);
nand U6291 (N_6291,N_3333,N_5772);
xnor U6292 (N_6292,N_4063,N_5650);
nor U6293 (N_6293,N_4304,N_3104);
nor U6294 (N_6294,N_5296,N_4778);
or U6295 (N_6295,N_5646,N_4575);
nor U6296 (N_6296,N_5535,N_5341);
nor U6297 (N_6297,N_5410,N_3239);
nor U6298 (N_6298,N_5631,N_5476);
xnor U6299 (N_6299,N_4311,N_5302);
or U6300 (N_6300,N_5984,N_3615);
or U6301 (N_6301,N_3780,N_3691);
and U6302 (N_6302,N_3685,N_3848);
nand U6303 (N_6303,N_3137,N_4500);
xor U6304 (N_6304,N_3173,N_5453);
xor U6305 (N_6305,N_4427,N_5792);
and U6306 (N_6306,N_4680,N_5183);
xor U6307 (N_6307,N_5618,N_5484);
xnor U6308 (N_6308,N_5293,N_5744);
xnor U6309 (N_6309,N_5660,N_4219);
and U6310 (N_6310,N_4940,N_5042);
or U6311 (N_6311,N_3229,N_3836);
or U6312 (N_6312,N_5487,N_5914);
nor U6313 (N_6313,N_4387,N_5601);
xor U6314 (N_6314,N_3827,N_4265);
or U6315 (N_6315,N_5769,N_3138);
nand U6316 (N_6316,N_4299,N_4640);
nand U6317 (N_6317,N_3547,N_4988);
or U6318 (N_6318,N_4430,N_3081);
nor U6319 (N_6319,N_5990,N_3977);
or U6320 (N_6320,N_5964,N_4382);
nor U6321 (N_6321,N_5106,N_4274);
xor U6322 (N_6322,N_4593,N_3922);
xor U6323 (N_6323,N_5482,N_3717);
or U6324 (N_6324,N_4198,N_5009);
nand U6325 (N_6325,N_4953,N_3752);
xor U6326 (N_6326,N_5656,N_3694);
and U6327 (N_6327,N_3248,N_5372);
xor U6328 (N_6328,N_3265,N_5935);
nand U6329 (N_6329,N_5397,N_5113);
nand U6330 (N_6330,N_4435,N_4565);
or U6331 (N_6331,N_5697,N_3016);
and U6332 (N_6332,N_5876,N_4960);
and U6333 (N_6333,N_4735,N_3552);
nor U6334 (N_6334,N_3360,N_3540);
xnor U6335 (N_6335,N_5126,N_3329);
nand U6336 (N_6336,N_4384,N_4378);
or U6337 (N_6337,N_4161,N_4424);
xnor U6338 (N_6338,N_5191,N_4098);
nor U6339 (N_6339,N_4989,N_4289);
xnor U6340 (N_6340,N_3804,N_3315);
nand U6341 (N_6341,N_5500,N_3357);
and U6342 (N_6342,N_5629,N_3617);
nor U6343 (N_6343,N_4721,N_3761);
xnor U6344 (N_6344,N_5728,N_4647);
nor U6345 (N_6345,N_5149,N_5455);
and U6346 (N_6346,N_4343,N_3666);
and U6347 (N_6347,N_3041,N_3134);
xor U6348 (N_6348,N_3354,N_3598);
nand U6349 (N_6349,N_4100,N_4622);
and U6350 (N_6350,N_3200,N_3090);
xor U6351 (N_6351,N_3075,N_5556);
nand U6352 (N_6352,N_3640,N_5182);
xnor U6353 (N_6353,N_5327,N_4309);
and U6354 (N_6354,N_3122,N_5128);
nand U6355 (N_6355,N_4514,N_5249);
nor U6356 (N_6356,N_4374,N_3705);
nor U6357 (N_6357,N_5105,N_5960);
nand U6358 (N_6358,N_4285,N_3656);
nand U6359 (N_6359,N_5094,N_3674);
and U6360 (N_6360,N_3185,N_5621);
xnor U6361 (N_6361,N_5049,N_4666);
or U6362 (N_6362,N_5389,N_4080);
and U6363 (N_6363,N_3648,N_5202);
or U6364 (N_6364,N_4786,N_3114);
xnor U6365 (N_6365,N_4342,N_3356);
xnor U6366 (N_6366,N_4341,N_3255);
nand U6367 (N_6367,N_4709,N_4144);
or U6368 (N_6368,N_4170,N_4850);
nand U6369 (N_6369,N_5230,N_5121);
xnor U6370 (N_6370,N_3147,N_5396);
xnor U6371 (N_6371,N_3244,N_5765);
and U6372 (N_6372,N_5266,N_3748);
xor U6373 (N_6373,N_4204,N_4625);
xor U6374 (N_6374,N_5810,N_4770);
and U6375 (N_6375,N_5835,N_5195);
or U6376 (N_6376,N_4957,N_4775);
nand U6377 (N_6377,N_3695,N_5634);
and U6378 (N_6378,N_5115,N_5377);
xor U6379 (N_6379,N_3690,N_3549);
and U6380 (N_6380,N_3513,N_5415);
nand U6381 (N_6381,N_3797,N_5103);
nand U6382 (N_6382,N_4365,N_4183);
xor U6383 (N_6383,N_4459,N_3083);
nand U6384 (N_6384,N_5668,N_4797);
xor U6385 (N_6385,N_4597,N_4840);
or U6386 (N_6386,N_4579,N_5854);
or U6387 (N_6387,N_4583,N_4130);
or U6388 (N_6388,N_3968,N_4478);
nand U6389 (N_6389,N_4651,N_3241);
nand U6390 (N_6390,N_4224,N_5329);
nand U6391 (N_6391,N_3188,N_3786);
nor U6392 (N_6392,N_5418,N_5517);
or U6393 (N_6393,N_4921,N_5685);
or U6394 (N_6394,N_3825,N_4264);
or U6395 (N_6395,N_3242,N_4547);
xor U6396 (N_6396,N_4594,N_3432);
or U6397 (N_6397,N_4745,N_4416);
and U6398 (N_6398,N_5024,N_3111);
or U6399 (N_6399,N_4773,N_3025);
xnor U6400 (N_6400,N_5101,N_5592);
nand U6401 (N_6401,N_3560,N_3284);
and U6402 (N_6402,N_3012,N_3611);
xnor U6403 (N_6403,N_4250,N_3870);
xor U6404 (N_6404,N_3829,N_4725);
or U6405 (N_6405,N_5034,N_5367);
xor U6406 (N_6406,N_5658,N_4045);
or U6407 (N_6407,N_3879,N_4008);
nand U6408 (N_6408,N_4995,N_5526);
or U6409 (N_6409,N_3020,N_4612);
nand U6410 (N_6410,N_3346,N_4331);
nand U6411 (N_6411,N_3534,N_5878);
nor U6412 (N_6412,N_5567,N_4058);
nand U6413 (N_6413,N_3555,N_5304);
nor U6414 (N_6414,N_4670,N_4040);
and U6415 (N_6415,N_3942,N_3672);
or U6416 (N_6416,N_3589,N_3982);
and U6417 (N_6417,N_5486,N_4947);
and U6418 (N_6418,N_5254,N_5818);
xor U6419 (N_6419,N_3641,N_5695);
nor U6420 (N_6420,N_5564,N_4053);
and U6421 (N_6421,N_4429,N_5684);
nor U6422 (N_6422,N_4442,N_5247);
and U6423 (N_6423,N_4256,N_3907);
or U6424 (N_6424,N_4066,N_5025);
nor U6425 (N_6425,N_5248,N_4857);
nor U6426 (N_6426,N_4944,N_4383);
nor U6427 (N_6427,N_4748,N_3868);
nand U6428 (N_6428,N_4324,N_5472);
nand U6429 (N_6429,N_5961,N_3929);
xnor U6430 (N_6430,N_4404,N_3366);
nand U6431 (N_6431,N_3437,N_5561);
nor U6432 (N_6432,N_5178,N_5653);
xor U6433 (N_6433,N_3995,N_4754);
or U6434 (N_6434,N_5063,N_3074);
and U6435 (N_6435,N_4215,N_3772);
nor U6436 (N_6436,N_5007,N_4461);
xnor U6437 (N_6437,N_3468,N_5232);
xor U6438 (N_6438,N_4321,N_4510);
nand U6439 (N_6439,N_5082,N_5886);
nand U6440 (N_6440,N_5362,N_5288);
or U6441 (N_6441,N_4557,N_5907);
nor U6442 (N_6442,N_5597,N_5638);
or U6443 (N_6443,N_4119,N_4690);
xor U6444 (N_6444,N_3342,N_5239);
nor U6445 (N_6445,N_4603,N_3957);
xor U6446 (N_6446,N_4845,N_4795);
nand U6447 (N_6447,N_5199,N_3394);
xnor U6448 (N_6448,N_4599,N_5936);
nor U6449 (N_6449,N_4439,N_3084);
or U6450 (N_6450,N_5336,N_3495);
xnor U6451 (N_6451,N_5485,N_4764);
and U6452 (N_6452,N_4997,N_4983);
nor U6453 (N_6453,N_5696,N_4515);
nor U6454 (N_6454,N_3822,N_5422);
nand U6455 (N_6455,N_5427,N_5760);
or U6456 (N_6456,N_5895,N_4523);
xor U6457 (N_6457,N_3406,N_5880);
nor U6458 (N_6458,N_5917,N_3144);
or U6459 (N_6459,N_3923,N_3399);
nor U6460 (N_6460,N_4607,N_3920);
or U6461 (N_6461,N_4096,N_3101);
nand U6462 (N_6462,N_5842,N_4700);
and U6463 (N_6463,N_5932,N_4509);
and U6464 (N_6464,N_5733,N_4861);
and U6465 (N_6465,N_3577,N_5223);
xor U6466 (N_6466,N_5014,N_5317);
xnor U6467 (N_6467,N_5407,N_5830);
nor U6468 (N_6468,N_3725,N_3423);
xnor U6469 (N_6469,N_4278,N_5102);
or U6470 (N_6470,N_3143,N_3216);
or U6471 (N_6471,N_3189,N_4702);
nor U6472 (N_6472,N_5808,N_5213);
xor U6473 (N_6473,N_3174,N_5824);
nor U6474 (N_6474,N_3001,N_3754);
and U6475 (N_6475,N_3347,N_4234);
nand U6476 (N_6476,N_3300,N_4074);
or U6477 (N_6477,N_3454,N_4300);
nor U6478 (N_6478,N_3458,N_4996);
xnor U6479 (N_6479,N_3946,N_5095);
or U6480 (N_6480,N_3926,N_5680);
xor U6481 (N_6481,N_4684,N_4968);
or U6482 (N_6482,N_4055,N_3969);
or U6483 (N_6483,N_3055,N_4705);
nor U6484 (N_6484,N_4568,N_4815);
xnor U6485 (N_6485,N_4971,N_4402);
xor U6486 (N_6486,N_3314,N_4143);
nor U6487 (N_6487,N_4910,N_3210);
nor U6488 (N_6488,N_3259,N_4492);
nor U6489 (N_6489,N_5541,N_4820);
and U6490 (N_6490,N_3087,N_5245);
and U6491 (N_6491,N_5332,N_4354);
nand U6492 (N_6492,N_5528,N_4067);
nor U6493 (N_6493,N_4635,N_3932);
or U6494 (N_6494,N_4638,N_3145);
or U6495 (N_6495,N_4349,N_3520);
or U6496 (N_6496,N_5581,N_3391);
or U6497 (N_6497,N_3872,N_5035);
nor U6498 (N_6498,N_4719,N_3199);
xnor U6499 (N_6499,N_3414,N_4174);
xor U6500 (N_6500,N_5780,N_5110);
or U6501 (N_6501,N_5432,N_3533);
and U6502 (N_6502,N_4247,N_5335);
and U6503 (N_6503,N_4533,N_3908);
nand U6504 (N_6504,N_3813,N_5475);
xnor U6505 (N_6505,N_3283,N_5709);
nand U6506 (N_6506,N_4099,N_4561);
nor U6507 (N_6507,N_3054,N_3806);
or U6508 (N_6508,N_5406,N_3136);
nor U6509 (N_6509,N_4934,N_5996);
nor U6510 (N_6510,N_3345,N_3026);
nor U6511 (N_6511,N_4111,N_5813);
xnor U6512 (N_6512,N_5617,N_3603);
and U6513 (N_6513,N_5648,N_5351);
and U6514 (N_6514,N_5975,N_3728);
xor U6515 (N_6515,N_4858,N_5563);
xor U6516 (N_6516,N_5079,N_5888);
xnor U6517 (N_6517,N_4852,N_3273);
or U6518 (N_6518,N_3130,N_4235);
nand U6519 (N_6519,N_3962,N_5371);
xnor U6520 (N_6520,N_5219,N_4598);
nand U6521 (N_6521,N_4710,N_5360);
xnor U6522 (N_6522,N_3225,N_4344);
nor U6523 (N_6523,N_3441,N_4297);
nand U6524 (N_6524,N_3789,N_5179);
and U6525 (N_6525,N_4697,N_5270);
or U6526 (N_6526,N_4792,N_3779);
xnor U6527 (N_6527,N_3289,N_3430);
and U6528 (N_6528,N_3404,N_5390);
xor U6529 (N_6529,N_3453,N_4255);
xor U6530 (N_6530,N_4452,N_5297);
xnor U6531 (N_6531,N_5318,N_4732);
nor U6532 (N_6532,N_5364,N_4679);
nand U6533 (N_6533,N_5416,N_4195);
nor U6534 (N_6534,N_4038,N_3460);
nor U6535 (N_6535,N_4761,N_3720);
or U6536 (N_6536,N_4222,N_4559);
nor U6537 (N_6537,N_4703,N_3305);
or U6538 (N_6538,N_4821,N_3118);
or U6539 (N_6539,N_5312,N_4481);
xor U6540 (N_6540,N_5005,N_5761);
or U6541 (N_6541,N_3288,N_4269);
nor U6542 (N_6542,N_3785,N_3093);
or U6543 (N_6543,N_5734,N_3422);
nand U6544 (N_6544,N_4444,N_4614);
and U6545 (N_6545,N_3522,N_3258);
nor U6546 (N_6546,N_3563,N_4176);
or U6547 (N_6547,N_4816,N_4769);
nor U6548 (N_6548,N_5456,N_4642);
xnor U6549 (N_6549,N_3426,N_4370);
nand U6550 (N_6550,N_5430,N_4681);
nand U6551 (N_6551,N_5140,N_5169);
and U6552 (N_6552,N_3302,N_3270);
nor U6553 (N_6553,N_5449,N_3689);
nor U6554 (N_6554,N_3326,N_5274);
xnor U6555 (N_6555,N_4333,N_4799);
or U6556 (N_6556,N_3030,N_5926);
nor U6557 (N_6557,N_4017,N_3609);
nor U6558 (N_6558,N_3983,N_5070);
nand U6559 (N_6559,N_3238,N_3839);
nor U6560 (N_6560,N_3963,N_5912);
nor U6561 (N_6561,N_4190,N_4664);
xor U6562 (N_6562,N_4713,N_5513);
and U6563 (N_6563,N_4158,N_3131);
or U6564 (N_6564,N_5030,N_3911);
and U6565 (N_6565,N_3162,N_3119);
nor U6566 (N_6566,N_5806,N_3886);
nand U6567 (N_6567,N_5777,N_5665);
and U6568 (N_6568,N_5429,N_5622);
or U6569 (N_6569,N_4408,N_4796);
nor U6570 (N_6570,N_5311,N_4734);
or U6571 (N_6571,N_3890,N_3390);
nand U6572 (N_6572,N_5405,N_4543);
and U6573 (N_6573,N_3736,N_3544);
nand U6574 (N_6574,N_5584,N_3352);
nand U6575 (N_6575,N_3169,N_3207);
and U6576 (N_6576,N_4572,N_3038);
nor U6577 (N_6577,N_3061,N_3687);
nor U6578 (N_6578,N_4737,N_4897);
xnor U6579 (N_6579,N_3726,N_5979);
xnor U6580 (N_6580,N_3449,N_5901);
xnor U6581 (N_6581,N_4028,N_3688);
xor U6582 (N_6582,N_5098,N_4037);
or U6583 (N_6583,N_5858,N_3341);
nand U6584 (N_6584,N_4668,N_4902);
xnor U6585 (N_6585,N_4240,N_3816);
and U6586 (N_6586,N_4519,N_5776);
nand U6587 (N_6587,N_5479,N_3525);
nand U6588 (N_6588,N_4532,N_4516);
or U6589 (N_6589,N_3388,N_4928);
xor U6590 (N_6590,N_3850,N_3953);
nor U6591 (N_6591,N_3262,N_5553);
and U6592 (N_6592,N_3718,N_5682);
nand U6593 (N_6593,N_4179,N_4018);
nor U6594 (N_6594,N_5352,N_3632);
and U6595 (N_6595,N_3487,N_4927);
nand U6596 (N_6596,N_5092,N_3880);
or U6597 (N_6597,N_5726,N_4345);
or U6598 (N_6598,N_4233,N_3781);
or U6599 (N_6599,N_5956,N_4109);
nor U6600 (N_6600,N_5687,N_3621);
or U6601 (N_6601,N_5420,N_5868);
and U6602 (N_6602,N_4406,N_5610);
xor U6603 (N_6603,N_3713,N_3712);
nand U6604 (N_6604,N_3236,N_3518);
or U6605 (N_6605,N_5385,N_3719);
or U6606 (N_6606,N_3037,N_5471);
xnor U6607 (N_6607,N_5986,N_3193);
and U6608 (N_6608,N_5138,N_4908);
or U6609 (N_6609,N_3716,N_4746);
nor U6610 (N_6610,N_5578,N_4041);
or U6611 (N_6611,N_4437,N_3282);
and U6612 (N_6612,N_3312,N_3601);
or U6613 (N_6613,N_5568,N_3595);
or U6614 (N_6614,N_5119,N_5091);
nor U6615 (N_6615,N_3380,N_4081);
xnor U6616 (N_6616,N_3626,N_3738);
or U6617 (N_6617,N_3760,N_4206);
or U6618 (N_6618,N_4303,N_4356);
or U6619 (N_6619,N_3510,N_5013);
nand U6620 (N_6620,N_4217,N_4498);
or U6621 (N_6621,N_4397,N_5262);
nor U6622 (N_6622,N_3067,N_3077);
or U6623 (N_6623,N_5826,N_3015);
or U6624 (N_6624,N_5735,N_3671);
or U6625 (N_6625,N_3195,N_4574);
or U6626 (N_6626,N_3214,N_5883);
nor U6627 (N_6627,N_5972,N_3799);
nor U6628 (N_6628,N_4904,N_4359);
or U6629 (N_6629,N_3410,N_4975);
xnor U6630 (N_6630,N_5688,N_5664);
nor U6631 (N_6631,N_3630,N_5759);
xor U6632 (N_6632,N_3724,N_4328);
and U6633 (N_6633,N_3796,N_5640);
nand U6634 (N_6634,N_3576,N_5197);
xnor U6635 (N_6635,N_4777,N_5789);
and U6636 (N_6636,N_5585,N_3931);
nor U6637 (N_6637,N_4178,N_3240);
nand U6638 (N_6638,N_5923,N_4843);
nand U6639 (N_6639,N_4930,N_3434);
xnor U6640 (N_6640,N_4554,N_3788);
nand U6641 (N_6641,N_4894,N_5615);
nand U6642 (N_6642,N_5659,N_4924);
nand U6643 (N_6643,N_3355,N_4644);
and U6644 (N_6644,N_5215,N_4399);
and U6645 (N_6645,N_4964,N_4353);
xnor U6646 (N_6646,N_4160,N_5168);
nand U6647 (N_6647,N_4064,N_5630);
and U6648 (N_6648,N_5334,N_4462);
or U6649 (N_6649,N_3266,N_5207);
nor U6650 (N_6650,N_5263,N_3060);
or U6651 (N_6651,N_4883,N_3335);
or U6652 (N_6652,N_3529,N_5131);
nand U6653 (N_6653,N_5272,N_4648);
and U6654 (N_6654,N_4097,N_3802);
or U6655 (N_6655,N_3443,N_4723);
nor U6656 (N_6656,N_5718,N_5740);
nor U6657 (N_6657,N_3271,N_4772);
and U6658 (N_6658,N_4649,N_4152);
or U6659 (N_6659,N_3875,N_3466);
or U6660 (N_6660,N_3076,N_4807);
or U6661 (N_6661,N_5411,N_4076);
or U6662 (N_6662,N_3331,N_5307);
nand U6663 (N_6663,N_4739,N_4470);
nand U6664 (N_6664,N_5857,N_4926);
xor U6665 (N_6665,N_3820,N_5866);
xor U6666 (N_6666,N_5357,N_5569);
nor U6667 (N_6667,N_4422,N_3878);
nand U6668 (N_6668,N_4047,N_3826);
nor U6669 (N_6669,N_3635,N_5315);
nor U6670 (N_6670,N_5636,N_3508);
and U6671 (N_6671,N_4386,N_4804);
xnor U6672 (N_6672,N_5546,N_4203);
nor U6673 (N_6673,N_3985,N_5885);
nor U6674 (N_6674,N_5378,N_4466);
nand U6675 (N_6675,N_5037,N_5060);
and U6676 (N_6676,N_3643,N_4576);
nand U6677 (N_6677,N_3624,N_4329);
nor U6678 (N_6678,N_4368,N_4192);
nand U6679 (N_6679,N_3010,N_5309);
and U6680 (N_6680,N_5286,N_5294);
nand U6681 (N_6681,N_4798,N_3571);
xor U6682 (N_6682,N_4853,N_3080);
and U6683 (N_6683,N_3684,N_5941);
xnor U6684 (N_6684,N_4962,N_3714);
or U6685 (N_6685,N_3416,N_5915);
nand U6686 (N_6686,N_4630,N_4244);
and U6687 (N_6687,N_4491,N_3882);
and U6688 (N_6688,N_5549,N_5123);
and U6689 (N_6689,N_3085,N_4314);
and U6690 (N_6690,N_4941,N_5742);
xnor U6691 (N_6691,N_3425,N_5340);
xnor U6692 (N_6692,N_4765,N_5846);
nand U6693 (N_6693,N_3303,N_4388);
nor U6694 (N_6694,N_5000,N_4929);
xnor U6695 (N_6695,N_3220,N_4282);
or U6696 (N_6696,N_3148,N_5269);
nand U6697 (N_6697,N_3106,N_5519);
xnor U6698 (N_6698,N_4591,N_3183);
nand U6699 (N_6699,N_4137,N_3680);
xor U6700 (N_6700,N_5971,N_4854);
and U6701 (N_6701,N_4727,N_3614);
nand U6702 (N_6702,N_5779,N_5146);
nand U6703 (N_6703,N_4460,N_4643);
or U6704 (N_6704,N_4782,N_5282);
nand U6705 (N_6705,N_5271,N_4671);
xnor U6706 (N_6706,N_4749,N_4567);
or U6707 (N_6707,N_3634,N_5715);
nand U6708 (N_6708,N_4881,N_3524);
xnor U6709 (N_6709,N_4956,N_4062);
nand U6710 (N_6710,N_4958,N_5869);
or U6711 (N_6711,N_4788,N_5234);
nor U6712 (N_6712,N_3972,N_5331);
nor U6713 (N_6713,N_4937,N_5637);
and U6714 (N_6714,N_3904,N_3279);
or U6715 (N_6715,N_3231,N_5811);
and U6716 (N_6716,N_4371,N_5085);
nor U6717 (N_6717,N_3940,N_3871);
nor U6718 (N_6718,N_4337,N_5819);
and U6719 (N_6719,N_5470,N_4373);
or U6720 (N_6720,N_3098,N_5503);
or U6721 (N_6721,N_4431,N_5489);
nand U6722 (N_6722,N_4425,N_5431);
xor U6723 (N_6723,N_5129,N_5494);
xnor U6724 (N_6724,N_3731,N_4476);
nor U6725 (N_6725,N_3378,N_3515);
nor U6726 (N_6726,N_4917,N_5151);
or U6727 (N_6727,N_4348,N_3146);
nor U6728 (N_6728,N_3997,N_3517);
and U6729 (N_6729,N_3269,N_3046);
nor U6730 (N_6730,N_5515,N_5242);
xnor U6731 (N_6731,N_5771,N_4420);
nand U6732 (N_6732,N_3569,N_4210);
nand U6733 (N_6733,N_3112,N_3361);
or U6734 (N_6734,N_4451,N_3369);
and U6735 (N_6735,N_3960,N_3777);
and U6736 (N_6736,N_3535,N_4683);
xor U6737 (N_6737,N_4751,N_4118);
and U6738 (N_6738,N_5264,N_5580);
nand U6739 (N_6739,N_4390,N_3620);
nor U6740 (N_6740,N_3750,N_5910);
nand U6741 (N_6741,N_5170,N_4774);
xor U6742 (N_6742,N_5887,N_4102);
or U6743 (N_6743,N_3439,N_3874);
xor U6744 (N_6744,N_4933,N_5604);
xnor U6745 (N_6745,N_3043,N_5743);
nor U6746 (N_6746,N_5064,N_5505);
xnor U6747 (N_6747,N_5366,N_3585);
and U6748 (N_6748,N_5176,N_5450);
nor U6749 (N_6749,N_4113,N_5948);
nand U6750 (N_6750,N_4628,N_3411);
and U6751 (N_6751,N_4785,N_4027);
and U6752 (N_6752,N_5983,N_3124);
nand U6753 (N_6753,N_4525,N_5276);
xnor U6754 (N_6754,N_3175,N_5708);
xor U6755 (N_6755,N_3759,N_5347);
or U6756 (N_6756,N_3828,N_5594);
or U6757 (N_6757,N_4789,N_5229);
nor U6758 (N_6758,N_3405,N_3139);
nor U6759 (N_6759,N_5240,N_5041);
or U6760 (N_6760,N_3841,N_4653);
and U6761 (N_6761,N_5452,N_4057);
xnor U6762 (N_6762,N_3771,N_5589);
and U6763 (N_6763,N_4225,N_4503);
and U6764 (N_6764,N_4209,N_5614);
and U6765 (N_6765,N_5031,N_5877);
or U6766 (N_6766,N_4101,N_3196);
xor U6767 (N_6767,N_4661,N_3910);
nor U6768 (N_6768,N_3667,N_3523);
nor U6769 (N_6769,N_5973,N_3017);
nand U6770 (N_6770,N_4124,N_5756);
or U6771 (N_6771,N_4147,N_4637);
nor U6772 (N_6772,N_5583,N_4296);
and U6773 (N_6773,N_4856,N_5267);
xnor U6774 (N_6774,N_3778,N_3514);
xnor U6775 (N_6775,N_4084,N_4693);
nor U6776 (N_6776,N_3782,N_3483);
or U6777 (N_6777,N_4270,N_4281);
nand U6778 (N_6778,N_5803,N_4257);
and U6779 (N_6779,N_5825,N_5423);
nor U6780 (N_6780,N_5442,N_5275);
or U6781 (N_6781,N_5193,N_4490);
or U6782 (N_6782,N_5736,N_5992);
or U6783 (N_6783,N_5988,N_4123);
nor U6784 (N_6784,N_3580,N_3817);
nor U6785 (N_6785,N_4391,N_3097);
or U6786 (N_6786,N_5865,N_3775);
nand U6787 (N_6787,N_4440,N_4272);
nand U6788 (N_6788,N_5711,N_3264);
xnor U6789 (N_6789,N_3364,N_3693);
xor U6790 (N_6790,N_4836,N_4724);
xnor U6791 (N_6791,N_5600,N_4295);
xnor U6792 (N_6792,N_4601,N_4878);
or U6793 (N_6793,N_5125,N_3993);
and U6794 (N_6794,N_3002,N_5774);
xor U6795 (N_6795,N_3308,N_4447);
nand U6796 (N_6796,N_5647,N_3647);
or U6797 (N_6797,N_3292,N_5198);
nor U6798 (N_6798,N_3194,N_4238);
nand U6799 (N_6799,N_5676,N_3633);
nor U6800 (N_6800,N_3488,N_3313);
xor U6801 (N_6801,N_3605,N_5766);
xor U6802 (N_6802,N_3994,N_3103);
or U6803 (N_6803,N_3727,N_4283);
xor U6804 (N_6804,N_4692,N_4091);
nand U6805 (N_6805,N_3883,N_5177);
nand U6806 (N_6806,N_5026,N_3217);
nand U6807 (N_6807,N_5875,N_3127);
xor U6808 (N_6808,N_5464,N_4657);
or U6809 (N_6809,N_4919,N_5279);
and U6810 (N_6810,N_3536,N_3490);
and U6811 (N_6811,N_5721,N_4405);
and U6812 (N_6812,N_3702,N_4802);
xnor U6813 (N_6813,N_4563,N_4202);
xor U6814 (N_6814,N_4602,N_3831);
xor U6815 (N_6815,N_4783,N_5504);
and U6816 (N_6816,N_4864,N_4569);
or U6817 (N_6817,N_3979,N_5497);
or U6818 (N_6818,N_4639,N_3838);
nor U6819 (N_6819,N_4731,N_3668);
nand U6820 (N_6820,N_5212,N_4419);
and U6821 (N_6821,N_5705,N_4586);
and U6822 (N_6822,N_5010,N_3186);
nand U6823 (N_6823,N_5537,N_3795);
and U6824 (N_6824,N_5147,N_4446);
or U6825 (N_6825,N_3096,N_3088);
xor U6826 (N_6826,N_3252,N_3996);
xor U6827 (N_6827,N_4287,N_5980);
nor U6828 (N_6828,N_5654,N_5548);
nor U6829 (N_6829,N_5046,N_4717);
nor U6830 (N_6830,N_5722,N_5310);
or U6831 (N_6831,N_4465,N_3486);
and U6832 (N_6832,N_5994,N_3481);
nor U6833 (N_6833,N_5967,N_3421);
nand U6834 (N_6834,N_3105,N_3150);
or U6835 (N_6835,N_5228,N_3936);
or U6836 (N_6836,N_4838,N_4912);
and U6837 (N_6837,N_4900,N_5527);
xor U6838 (N_6838,N_4166,N_5856);
nand U6839 (N_6839,N_4945,N_3638);
or U6840 (N_6840,N_5641,N_3429);
and U6841 (N_6841,N_3156,N_3154);
nor U6842 (N_6842,N_4379,N_3928);
and U6843 (N_6843,N_5746,N_4992);
nor U6844 (N_6844,N_4154,N_5356);
and U6845 (N_6845,N_4993,N_5358);
xnor U6846 (N_6846,N_5019,N_3120);
or U6847 (N_6847,N_4566,N_5052);
or U6848 (N_6848,N_5978,N_5285);
or U6849 (N_6849,N_3867,N_3981);
nand U6850 (N_6850,N_5141,N_3295);
xnor U6851 (N_6851,N_5855,N_5931);
xnor U6852 (N_6852,N_4611,N_4604);
nand U6853 (N_6853,N_3659,N_5954);
xor U6854 (N_6854,N_5130,N_3398);
and U6855 (N_6855,N_4986,N_3501);
and U6856 (N_6856,N_4423,N_3790);
nor U6857 (N_6857,N_5966,N_3954);
nand U6858 (N_6858,N_3408,N_3023);
or U6859 (N_6859,N_3206,N_5575);
or U6860 (N_6860,N_4741,N_5204);
nand U6861 (N_6861,N_3722,N_4313);
nand U6862 (N_6862,N_5108,N_5398);
xor U6863 (N_6863,N_4239,N_3986);
xor U6864 (N_6864,N_3396,N_5020);
or U6865 (N_6865,N_4538,N_3141);
and U6866 (N_6866,N_3024,N_5934);
nand U6867 (N_6867,N_5218,N_3203);
or U6868 (N_6868,N_4212,N_3697);
or U6869 (N_6869,N_3126,N_3178);
or U6870 (N_6870,N_3463,N_5701);
nand U6871 (N_6871,N_5090,N_3505);
xor U6872 (N_6872,N_3613,N_4600);
nor U6873 (N_6873,N_4831,N_5495);
nor U6874 (N_6874,N_4196,N_4592);
or U6875 (N_6875,N_5690,N_3415);
and U6876 (N_6876,N_3301,N_3887);
nand U6877 (N_6877,N_4319,N_4524);
xnor U6878 (N_6878,N_3961,N_5832);
and U6879 (N_6879,N_4394,N_3444);
nor U6880 (N_6880,N_3168,N_5778);
nand U6881 (N_6881,N_5386,N_4812);
nand U6882 (N_6882,N_3686,N_3561);
nand U6883 (N_6883,N_5067,N_4268);
or U6884 (N_6884,N_5062,N_4479);
nor U6885 (N_6885,N_4497,N_3746);
nand U6886 (N_6886,N_3764,N_3230);
nand U6887 (N_6887,N_3461,N_4266);
xnor U6888 (N_6888,N_3268,N_4013);
xor U6889 (N_6889,N_5459,N_5643);
nand U6890 (N_6890,N_4729,N_4332);
nand U6891 (N_6891,N_3275,N_3675);
nor U6892 (N_6892,N_5906,N_4752);
nand U6893 (N_6893,N_4248,N_4410);
nand U6894 (N_6894,N_5236,N_4450);
and U6895 (N_6895,N_3008,N_5122);
or U6896 (N_6896,N_4973,N_5802);
nor U6897 (N_6897,N_5306,N_5790);
and U6898 (N_6898,N_3894,N_3710);
xnor U6899 (N_6899,N_3553,N_5033);
and U6900 (N_6900,N_4587,N_4172);
nor U6901 (N_6901,N_5608,N_3009);
nand U6902 (N_6902,N_5008,N_4534);
xnor U6903 (N_6903,N_5185,N_5018);
nor U6904 (N_6904,N_3323,N_5166);
xnor U6905 (N_6905,N_5251,N_3221);
and U6906 (N_6906,N_4002,N_5328);
or U6907 (N_6907,N_5460,N_4665);
nand U6908 (N_6908,N_3172,N_5981);
and U6909 (N_6909,N_4595,N_4499);
nand U6910 (N_6910,N_3285,N_5518);
and U6911 (N_6911,N_4441,N_5884);
nand U6912 (N_6912,N_4530,N_3747);
nor U6913 (N_6913,N_4596,N_4707);
nand U6914 (N_6914,N_3467,N_4867);
nand U6915 (N_6915,N_5342,N_3372);
and U6916 (N_6916,N_4932,N_3051);
and U6917 (N_6917,N_5574,N_5137);
nand U6918 (N_6918,N_5800,N_4014);
nor U6919 (N_6919,N_3864,N_4699);
and U6920 (N_6920,N_3491,N_4517);
and U6921 (N_6921,N_5635,N_5462);
nor U6922 (N_6922,N_5278,N_4071);
or U6923 (N_6923,N_4487,N_4474);
xor U6924 (N_6924,N_5655,N_5155);
nor U6925 (N_6925,N_5795,N_5419);
or U6926 (N_6926,N_3812,N_3249);
or U6927 (N_6927,N_3201,N_3176);
or U6928 (N_6928,N_4458,N_3557);
xor U6929 (N_6929,N_4862,N_5874);
or U6930 (N_6930,N_5642,N_4433);
xor U6931 (N_6931,N_3336,N_3116);
and U6932 (N_6932,N_5870,N_4385);
nand U6933 (N_6933,N_5510,N_4232);
nor U6934 (N_6934,N_3805,N_3474);
xnor U6935 (N_6935,N_5257,N_3619);
and U6936 (N_6936,N_4077,N_4298);
nand U6937 (N_6937,N_5982,N_4227);
nand U6938 (N_6938,N_4418,N_4794);
nor U6939 (N_6939,N_3893,N_5038);
nor U6940 (N_6940,N_3132,N_3918);
xnor U6941 (N_6941,N_4972,N_5542);
and U6942 (N_6942,N_5134,N_4979);
or U6943 (N_6943,N_5346,N_4245);
nor U6944 (N_6944,N_3280,N_4535);
nor U6945 (N_6945,N_5434,N_3377);
nor U6946 (N_6946,N_5190,N_5922);
nand U6947 (N_6947,N_4711,N_3403);
nand U6948 (N_6948,N_3319,N_3568);
and U6949 (N_6949,N_3191,N_5401);
nor U6950 (N_6950,N_3583,N_3744);
or U6951 (N_6951,N_3526,N_4652);
and U6952 (N_6952,N_3125,N_5719);
nor U6953 (N_6953,N_5363,N_3676);
or U6954 (N_6954,N_3847,N_4954);
xor U6955 (N_6955,N_5532,N_4355);
or U6956 (N_6956,N_4677,N_5925);
xor U6957 (N_6957,N_5853,N_4893);
and U6958 (N_6958,N_5153,N_3459);
xnor U6959 (N_6959,N_4969,N_4173);
or U6960 (N_6960,N_3937,N_5447);
or U6961 (N_6961,N_5538,N_4079);
nor U6962 (N_6962,N_3723,N_3005);
nor U6963 (N_6963,N_5457,N_5947);
xor U6964 (N_6964,N_4990,N_3657);
nor U6965 (N_6965,N_4488,N_5626);
xor U6966 (N_6966,N_3310,N_5867);
and U6967 (N_6967,N_3219,N_3768);
and U6968 (N_6968,N_3824,N_5040);
xnor U6969 (N_6969,N_3991,N_5354);
nor U6970 (N_6970,N_3707,N_4302);
xnor U6971 (N_6971,N_4809,N_3762);
and U6972 (N_6972,N_3392,N_4556);
xor U6973 (N_6973,N_4457,N_5927);
nor U6974 (N_6974,N_4326,N_4696);
or U6975 (N_6975,N_4564,N_5480);
nor U6976 (N_6976,N_4659,N_5339);
and U6977 (N_6977,N_3135,N_5859);
and U6978 (N_6978,N_4747,N_3538);
xor U6979 (N_6979,N_5783,N_3683);
nand U6980 (N_6980,N_3251,N_4199);
nand U6981 (N_6981,N_3155,N_5380);
xnor U6982 (N_6982,N_5930,N_5132);
nor U6983 (N_6983,N_4529,N_3494);
or U6984 (N_6984,N_3339,N_5112);
nor U6985 (N_6985,N_5879,N_3573);
nand U6986 (N_6986,N_5555,N_5821);
nand U6987 (N_6987,N_3149,N_3379);
or U6988 (N_6988,N_5481,N_5529);
or U6989 (N_6989,N_5714,N_4323);
xor U6990 (N_6990,N_4279,N_5543);
nor U6991 (N_6991,N_5689,N_3905);
xnor U6992 (N_6992,N_4258,N_4621);
nand U6993 (N_6993,N_4722,N_4073);
xnor U6994 (N_6994,N_4585,N_4034);
xor U6995 (N_6995,N_4362,N_5864);
nand U6996 (N_6996,N_4819,N_5373);
or U6997 (N_6997,N_4369,N_4263);
nor U6998 (N_6998,N_4882,N_5072);
nor U6999 (N_6999,N_5909,N_5111);
or U7000 (N_7000,N_3368,N_4032);
and U7001 (N_7001,N_3261,N_4555);
xnor U7002 (N_7002,N_3381,N_5287);
xnor U7003 (N_7003,N_4685,N_4175);
and U7004 (N_7004,N_4230,N_3320);
and U7005 (N_7005,N_3801,N_3470);
xor U7006 (N_7006,N_3945,N_4706);
nand U7007 (N_7007,N_4290,N_3035);
nand U7008 (N_7008,N_5662,N_4310);
nor U7009 (N_7009,N_5739,N_3964);
xnor U7010 (N_7010,N_3299,N_5502);
xnor U7011 (N_7011,N_5753,N_4830);
xor U7012 (N_7012,N_4588,N_3729);
nor U7013 (N_7013,N_4213,N_5833);
and U7014 (N_7014,N_5133,N_5438);
and U7015 (N_7015,N_5443,N_3869);
or U7016 (N_7016,N_4006,N_5955);
or U7017 (N_7017,N_3384,N_5148);
or U7018 (N_7018,N_3913,N_3941);
or U7019 (N_7019,N_4716,N_5056);
or U7020 (N_7020,N_4935,N_3413);
nor U7021 (N_7021,N_5292,N_5209);
nand U7022 (N_7022,N_5596,N_4866);
nor U7023 (N_7023,N_3328,N_4526);
and U7024 (N_7024,N_4120,N_5417);
and U7025 (N_7025,N_5571,N_5632);
and U7026 (N_7026,N_4115,N_3604);
xor U7027 (N_7027,N_3036,N_5834);
or U7028 (N_7028,N_3086,N_3507);
xor U7029 (N_7029,N_5850,N_4834);
and U7030 (N_7030,N_5723,N_3153);
nor U7031 (N_7031,N_3142,N_4454);
nor U7032 (N_7032,N_4307,N_3128);
or U7033 (N_7033,N_5135,N_4590);
xnor U7034 (N_7034,N_4865,N_5545);
nor U7035 (N_7035,N_5162,N_5784);
and U7036 (N_7036,N_5050,N_4704);
and U7037 (N_7037,N_3059,N_5458);
or U7038 (N_7038,N_4660,N_3327);
xnor U7039 (N_7039,N_5369,N_3465);
and U7040 (N_7040,N_3682,N_4578);
or U7041 (N_7041,N_3450,N_3889);
xor U7042 (N_7042,N_5301,N_4346);
and U7043 (N_7043,N_5710,N_5816);
or U7044 (N_7044,N_5093,N_5099);
nand U7045 (N_7045,N_4829,N_3376);
nand U7046 (N_7046,N_4484,N_4698);
nor U7047 (N_7047,N_5032,N_5374);
nor U7048 (N_7048,N_3254,N_5244);
nand U7049 (N_7049,N_4645,N_3250);
nor U7050 (N_7050,N_3334,N_4131);
nand U7051 (N_7051,N_4229,N_4376);
nand U7052 (N_7052,N_4389,N_3902);
nor U7053 (N_7053,N_3628,N_5303);
or U7054 (N_7054,N_3029,N_5860);
and U7055 (N_7055,N_5900,N_4920);
nor U7056 (N_7056,N_3930,N_5253);
nor U7057 (N_7057,N_5672,N_4030);
xnor U7058 (N_7058,N_3646,N_5403);
or U7059 (N_7059,N_3608,N_3653);
nor U7060 (N_7060,N_3089,N_4984);
and U7061 (N_7061,N_3622,N_4104);
nand U7062 (N_7062,N_5717,N_5023);
and U7063 (N_7063,N_4546,N_3072);
or U7064 (N_7064,N_3224,N_5467);
xor U7065 (N_7065,N_4718,N_5675);
nand U7066 (N_7066,N_5977,N_4833);
xnor U7067 (N_7067,N_3160,N_3383);
nand U7068 (N_7068,N_4241,N_4553);
xor U7069 (N_7069,N_3018,N_5225);
nand U7070 (N_7070,N_5395,N_5557);
and U7071 (N_7071,N_3237,N_5920);
and U7072 (N_7072,N_4180,N_3476);
nand U7073 (N_7073,N_4200,N_4760);
and U7074 (N_7074,N_4044,N_5300);
and U7075 (N_7075,N_5210,N_5124);
xor U7076 (N_7076,N_5320,N_5379);
nor U7077 (N_7077,N_5508,N_4336);
or U7078 (N_7078,N_4505,N_5613);
xnor U7079 (N_7079,N_4126,N_3455);
nand U7080 (N_7080,N_5770,N_4663);
and U7081 (N_7081,N_5167,N_5277);
or U7082 (N_7082,N_5387,N_4654);
nor U7083 (N_7083,N_3021,N_3309);
nand U7084 (N_7084,N_3418,N_3900);
xnor U7085 (N_7085,N_4477,N_3914);
nand U7086 (N_7086,N_3482,N_5773);
xnor U7087 (N_7087,N_5572,N_4407);
nor U7088 (N_7088,N_4511,N_5588);
or U7089 (N_7089,N_4157,N_5343);
nor U7090 (N_7090,N_4401,N_4617);
and U7091 (N_7091,N_4151,N_4271);
nor U7092 (N_7092,N_4009,N_4251);
nand U7093 (N_7093,N_5627,N_4167);
and U7094 (N_7094,N_4377,N_5590);
nand U7095 (N_7095,N_5221,N_4848);
and U7096 (N_7096,N_4153,N_4624);
xnor U7097 (N_7097,N_5353,N_4286);
or U7098 (N_7098,N_4835,N_3223);
nand U7099 (N_7099,N_4165,N_4169);
and U7100 (N_7100,N_5181,N_3766);
nor U7101 (N_7101,N_5408,N_4306);
nor U7102 (N_7102,N_4970,N_5326);
nand U7103 (N_7103,N_3948,N_5463);
xnor U7104 (N_7104,N_3071,N_3420);
nor U7105 (N_7105,N_4974,N_5412);
and U7106 (N_7106,N_4977,N_4471);
and U7107 (N_7107,N_3663,N_3047);
xor U7108 (N_7108,N_3247,N_4701);
xnor U7109 (N_7109,N_5805,N_3616);
xor U7110 (N_7110,N_4967,N_4189);
nor U7111 (N_7111,N_4228,N_4896);
xor U7112 (N_7112,N_3190,N_3537);
and U7113 (N_7113,N_4237,N_5088);
or U7114 (N_7114,N_5069,N_3833);
xor U7115 (N_7115,N_5437,N_4720);
nand U7116 (N_7116,N_3359,N_3073);
xor U7117 (N_7117,N_5400,N_4694);
or U7118 (N_7118,N_3115,N_5991);
or U7119 (N_7119,N_4364,N_5788);
nor U7120 (N_7120,N_5444,N_4051);
nand U7121 (N_7121,N_3807,N_4955);
or U7122 (N_7122,N_3565,N_5671);
xor U7123 (N_7123,N_5004,N_3532);
nand U7124 (N_7124,N_3642,N_5605);
nand U7125 (N_7125,N_5172,N_4340);
or U7126 (N_7126,N_5976,N_5838);
xor U7127 (N_7127,N_3625,N_3784);
xor U7128 (N_7128,N_4409,N_5547);
and U7129 (N_7129,N_4004,N_4133);
xnor U7130 (N_7130,N_3855,N_3019);
and U7131 (N_7131,N_4844,N_4911);
nand U7132 (N_7132,N_5150,N_3167);
xor U7133 (N_7133,N_4093,N_3599);
nand U7134 (N_7134,N_4753,N_4155);
or U7135 (N_7135,N_4981,N_4475);
or U7136 (N_7136,N_5281,N_4806);
xnor U7137 (N_7137,N_3590,N_3107);
xnor U7138 (N_7138,N_3629,N_5679);
xnor U7139 (N_7139,N_4779,N_3187);
or U7140 (N_7140,N_5188,N_5928);
nand U7141 (N_7141,N_4631,N_5745);
or U7142 (N_7142,N_4021,N_5053);
and U7143 (N_7143,N_4846,N_5674);
or U7144 (N_7144,N_4082,N_3770);
or U7145 (N_7145,N_3245,N_4221);
and U7146 (N_7146,N_3755,N_5413);
and U7147 (N_7147,N_4714,N_4913);
nor U7148 (N_7148,N_5775,N_4072);
and U7149 (N_7149,N_5514,N_3909);
or U7150 (N_7150,N_3607,N_3842);
xnor U7151 (N_7151,N_4363,N_5844);
xnor U7152 (N_7152,N_5501,N_5809);
or U7153 (N_7153,N_5409,N_5762);
xor U7154 (N_7154,N_3574,N_5381);
or U7155 (N_7155,N_5747,N_3440);
nor U7156 (N_7156,N_5796,N_5461);
or U7157 (N_7157,N_5841,N_4092);
xnor U7158 (N_7158,N_3117,N_4868);
nor U7159 (N_7159,N_5237,N_3528);
or U7160 (N_7160,N_5754,N_3939);
nor U7161 (N_7161,N_5924,N_3063);
xnor U7162 (N_7162,N_4056,N_3113);
and U7163 (N_7163,N_5382,N_5965);
and U7164 (N_7164,N_5039,N_3039);
xnor U7165 (N_7165,N_3473,N_5893);
and U7166 (N_7166,N_4873,N_5080);
xnor U7167 (N_7167,N_3496,N_3662);
or U7168 (N_7168,N_3696,N_5118);
or U7169 (N_7169,N_4129,N_4891);
xnor U7170 (N_7170,N_5916,N_3040);
or U7171 (N_7171,N_5587,N_3435);
or U7172 (N_7172,N_5174,N_3830);
nand U7173 (N_7173,N_4750,N_3511);
xnor U7174 (N_7174,N_3350,N_3504);
or U7175 (N_7175,N_4068,N_3332);
nor U7176 (N_7176,N_3353,N_5649);
nor U7177 (N_7177,N_4103,N_4613);
xor U7178 (N_7178,N_3121,N_4859);
xnor U7179 (N_7179,N_4872,N_3500);
nand U7180 (N_7180,N_4011,N_5787);
or U7181 (N_7181,N_3958,N_5533);
xnor U7182 (N_7182,N_4050,N_3863);
or U7183 (N_7183,N_5435,N_3933);
nor U7184 (N_7184,N_3373,N_5261);
nand U7185 (N_7185,N_4048,N_5782);
nand U7186 (N_7186,N_3861,N_5732);
xor U7187 (N_7187,N_4191,N_4860);
or U7188 (N_7188,N_3479,N_5116);
xor U7189 (N_7189,N_4811,N_4392);
xnor U7190 (N_7190,N_5623,N_5692);
nor U7191 (N_7191,N_4414,N_5836);
nand U7192 (N_7192,N_5203,N_4762);
nand U7193 (N_7193,N_4426,N_5891);
nand U7194 (N_7194,N_5720,N_5057);
and U7195 (N_7195,N_5669,N_5862);
xor U7196 (N_7196,N_3971,N_4771);
xor U7197 (N_7197,N_3602,N_4301);
nor U7198 (N_7198,N_4551,N_3999);
or U7199 (N_7199,N_4216,N_4375);
nand U7200 (N_7200,N_4669,N_4218);
and U7201 (N_7201,N_3109,N_5516);
or U7202 (N_7202,N_5933,N_4901);
nand U7203 (N_7203,N_5998,N_3004);
and U7204 (N_7204,N_4636,N_5260);
or U7205 (N_7205,N_5657,N_4185);
or U7206 (N_7206,N_4347,N_5096);
xnor U7207 (N_7207,N_5208,N_3545);
or U7208 (N_7208,N_5165,N_3567);
nand U7209 (N_7209,N_4184,N_3348);
nor U7210 (N_7210,N_3834,N_5065);
nor U7211 (N_7211,N_3057,N_4413);
nor U7212 (N_7212,N_3753,N_4135);
nor U7213 (N_7213,N_3699,N_4863);
and U7214 (N_7214,N_5959,N_4627);
nor U7215 (N_7215,N_4443,N_3227);
and U7216 (N_7216,N_3296,N_4634);
or U7217 (N_7217,N_5473,N_3181);
nand U7218 (N_7218,N_3896,N_5375);
xnor U7219 (N_7219,N_3304,N_4089);
nand U7220 (N_7220,N_3171,N_3692);
nor U7221 (N_7221,N_3564,N_4521);
nand U7222 (N_7222,N_3375,N_4141);
nand U7223 (N_7223,N_5421,N_5550);
and U7224 (N_7224,N_5576,N_5950);
xor U7225 (N_7225,N_5216,N_5205);
xor U7226 (N_7226,N_3212,N_5016);
and U7227 (N_7227,N_3263,N_4261);
nor U7228 (N_7228,N_3330,N_5305);
or U7229 (N_7229,N_4193,N_3915);
or U7230 (N_7230,N_4825,N_5828);
nor U7231 (N_7231,N_5918,N_4016);
xor U7232 (N_7232,N_3007,N_3551);
and U7233 (N_7233,N_5154,N_3226);
xnor U7234 (N_7234,N_4879,N_5273);
nor U7235 (N_7235,N_3556,N_4914);
xnor U7236 (N_7236,N_5544,N_4966);
or U7237 (N_7237,N_5512,N_3337);
nor U7238 (N_7238,N_5908,N_5433);
xor U7239 (N_7239,N_4982,N_3349);
or U7240 (N_7240,N_5881,N_3711);
and U7241 (N_7241,N_5161,N_4134);
xnor U7242 (N_7242,N_4738,N_3166);
nor U7243 (N_7243,N_3456,N_4674);
nand U7244 (N_7244,N_3276,N_3730);
or U7245 (N_7245,N_4952,N_4003);
and U7246 (N_7246,N_3776,N_4145);
nand U7247 (N_7247,N_5987,N_5325);
or U7248 (N_7248,N_3758,N_3401);
xnor U7249 (N_7249,N_3664,N_3180);
and U7250 (N_7250,N_4633,N_3480);
nand U7251 (N_7251,N_3521,N_4086);
xor U7252 (N_7252,N_3658,N_5392);
nand U7253 (N_7253,N_5817,N_5840);
nand U7254 (N_7254,N_3984,N_3202);
nand U7255 (N_7255,N_3078,N_3387);
nand U7256 (N_7256,N_3811,N_5187);
and U7257 (N_7257,N_5522,N_3955);
nor U7258 (N_7258,N_3478,N_5944);
nor U7259 (N_7259,N_3866,N_5681);
nand U7260 (N_7260,N_5003,N_4541);
or U7261 (N_7261,N_4531,N_5603);
xnor U7262 (N_7262,N_3260,N_4024);
or U7263 (N_7263,N_3650,N_4469);
nand U7264 (N_7264,N_4472,N_3815);
and U7265 (N_7265,N_3734,N_5673);
xnor U7266 (N_7266,N_3243,N_3988);
xor U7267 (N_7267,N_5530,N_4907);
nand U7268 (N_7268,N_4412,N_4766);
nor U7269 (N_7269,N_4496,N_3028);
or U7270 (N_7270,N_4106,N_5593);
nand U7271 (N_7271,N_5731,N_4231);
xor U7272 (N_7272,N_3469,N_3821);
nand U7273 (N_7273,N_3935,N_3899);
or U7274 (N_7274,N_4615,N_4871);
and U7275 (N_7275,N_5344,N_4923);
or U7276 (N_7276,N_3222,N_4276);
nor U7277 (N_7277,N_4577,N_4570);
or U7278 (N_7278,N_3849,N_3596);
or U7279 (N_7279,N_5313,N_5235);
or U7280 (N_7280,N_3457,N_4744);
and U7281 (N_7281,N_4194,N_3579);
nor U7282 (N_7282,N_3876,N_4197);
or U7283 (N_7283,N_3445,N_5043);
or U7284 (N_7284,N_5896,N_3769);
nor U7285 (N_7285,N_3070,N_3921);
xnor U7286 (N_7286,N_3854,N_5465);
nor U7287 (N_7287,N_3294,N_3475);
or U7288 (N_7288,N_5873,N_5047);
xnor U7289 (N_7289,N_4976,N_5173);
and U7290 (N_7290,N_4537,N_4758);
or U7291 (N_7291,N_5348,N_5498);
and U7292 (N_7292,N_5751,N_5599);
nand U7293 (N_7293,N_3575,N_4031);
or U7294 (N_7294,N_3745,N_5428);
nand U7295 (N_7295,N_4730,N_4540);
nor U7296 (N_7296,N_4205,N_4112);
nor U7297 (N_7297,N_3542,N_5217);
xor U7298 (N_7298,N_4502,N_4827);
nand U7299 (N_7299,N_3498,N_5002);
nor U7300 (N_7300,N_5845,N_3099);
nor U7301 (N_7301,N_4122,N_4870);
nor U7302 (N_7302,N_4335,N_3256);
nand U7303 (N_7303,N_4393,N_4817);
nand U7304 (N_7304,N_4139,N_4035);
or U7305 (N_7305,N_3903,N_4094);
and U7306 (N_7306,N_3600,N_3950);
or U7307 (N_7307,N_3198,N_4790);
xor U7308 (N_7308,N_3593,N_4107);
or U7309 (N_7309,N_4808,N_4675);
nand U7310 (N_7310,N_5076,N_5882);
or U7311 (N_7311,N_5186,N_5446);
xor U7312 (N_7312,N_4787,N_3715);
xnor U7313 (N_7313,N_4951,N_3417);
nor U7314 (N_7314,N_4938,N_3543);
xor U7315 (N_7315,N_5786,N_3512);
xnor U7316 (N_7316,N_4580,N_5839);
nor U7317 (N_7317,N_4226,N_3042);
nor U7318 (N_7318,N_5233,N_4545);
xor U7319 (N_7319,N_4020,N_4415);
xor U7320 (N_7320,N_4906,N_4432);
and U7321 (N_7321,N_5539,N_3184);
or U7322 (N_7322,N_5849,N_5451);
or U7323 (N_7323,N_4814,N_4132);
and U7324 (N_7324,N_5919,N_4171);
or U7325 (N_7325,N_4448,N_3246);
and U7326 (N_7326,N_4678,N_3645);
nand U7327 (N_7327,N_4039,N_4605);
or U7328 (N_7328,N_5993,N_5499);
and U7329 (N_7329,N_4042,N_5639);
and U7330 (N_7330,N_4672,N_5330);
xnor U7331 (N_7331,N_3853,N_3358);
nand U7332 (N_7332,N_5890,N_3064);
nor U7333 (N_7333,N_3677,N_4211);
or U7334 (N_7334,N_3739,N_3102);
nor U7335 (N_7335,N_3835,N_5999);
and U7336 (N_7336,N_3157,N_4146);
and U7337 (N_7337,N_3618,N_5246);
nor U7338 (N_7338,N_3343,N_3527);
and U7339 (N_7339,N_3698,N_5713);
and U7340 (N_7340,N_4925,N_5227);
nor U7341 (N_7341,N_4366,N_4728);
and U7342 (N_7342,N_5483,N_4128);
and U7343 (N_7343,N_4305,N_3773);
nand U7344 (N_7344,N_5827,N_3079);
xnor U7345 (N_7345,N_4780,N_5823);
and U7346 (N_7346,N_5905,N_5595);
and U7347 (N_7347,N_4246,N_3235);
nor U7348 (N_7348,N_3502,N_3069);
xnor U7349 (N_7349,N_5536,N_5265);
xor U7350 (N_7350,N_5445,N_4322);
xor U7351 (N_7351,N_5666,N_3530);
and U7352 (N_7352,N_4149,N_4483);
or U7353 (N_7353,N_5551,N_3588);
and U7354 (N_7354,N_3708,N_4284);
nor U7355 (N_7355,N_4965,N_4455);
and U7356 (N_7356,N_3856,N_4589);
nor U7357 (N_7357,N_3837,N_5083);
or U7358 (N_7358,N_3897,N_3058);
and U7359 (N_7359,N_3859,N_5078);
xor U7360 (N_7360,N_3531,N_5898);
xor U7361 (N_7361,N_5609,N_5768);
nand U7362 (N_7362,N_3045,N_4012);
xnor U7363 (N_7363,N_5114,N_5913);
xnor U7364 (N_7364,N_3151,N_3034);
or U7365 (N_7365,N_4117,N_4061);
xor U7366 (N_7366,N_4316,N_4352);
and U7367 (N_7367,N_4398,N_5164);
and U7368 (N_7368,N_3006,N_3182);
nand U7369 (N_7369,N_5807,N_5663);
nand U7370 (N_7370,N_4473,N_5921);
nand U7371 (N_7371,N_5678,N_5319);
nand U7372 (N_7372,N_3232,N_4486);
or U7373 (N_7373,N_5087,N_5628);
nand U7374 (N_7374,N_3845,N_4259);
and U7375 (N_7375,N_5370,N_5724);
nand U7376 (N_7376,N_4083,N_3749);
or U7377 (N_7377,N_3286,N_4791);
and U7378 (N_7378,N_3179,N_5892);
nand U7379 (N_7379,N_5752,N_5436);
xor U7380 (N_7380,N_3665,N_5376);
or U7381 (N_7381,N_5521,N_5577);
and U7382 (N_7382,N_3158,N_3477);
and U7383 (N_7383,N_4998,N_4978);
or U7384 (N_7384,N_5350,N_5426);
xor U7385 (N_7385,N_5686,N_4164);
nor U7386 (N_7386,N_3539,N_4793);
nor U7387 (N_7387,N_5337,N_5633);
nor U7388 (N_7388,N_4963,N_3558);
xnor U7389 (N_7389,N_5388,N_5316);
nor U7390 (N_7390,N_5531,N_5848);
nor U7391 (N_7391,N_3389,N_4108);
xnor U7392 (N_7392,N_3424,N_5938);
or U7393 (N_7393,N_4208,N_5152);
nand U7394 (N_7394,N_3591,N_3814);
or U7395 (N_7395,N_4070,N_3787);
and U7396 (N_7396,N_5359,N_3578);
nor U7397 (N_7397,N_5299,N_4767);
or U7398 (N_7398,N_5767,N_4905);
or U7399 (N_7399,N_3110,N_4528);
xnor U7400 (N_7400,N_3606,N_5831);
xor U7401 (N_7401,N_4262,N_3898);
xnor U7402 (N_7402,N_3082,N_4898);
nand U7403 (N_7403,N_5727,N_4142);
xnor U7404 (N_7404,N_3548,N_4403);
nor U7405 (N_7405,N_3519,N_4069);
xnor U7406 (N_7406,N_5591,N_5220);
xor U7407 (N_7407,N_4841,N_4623);
or U7408 (N_7408,N_3503,N_5837);
or U7409 (N_7409,N_3858,N_3133);
xor U7410 (N_7410,N_5054,N_4467);
or U7411 (N_7411,N_5607,N_5109);
xor U7412 (N_7412,N_4060,N_3952);
xor U7413 (N_7413,N_3370,N_5201);
or U7414 (N_7414,N_5764,N_5781);
nand U7415 (N_7415,N_3649,N_3967);
or U7416 (N_7416,N_4641,N_5086);
nor U7417 (N_7417,N_4608,N_5474);
or U7418 (N_7418,N_3340,N_5667);
nand U7419 (N_7419,N_5021,N_4010);
nand U7420 (N_7420,N_4236,N_3938);
nand U7421 (N_7421,N_3152,N_5554);
and U7422 (N_7422,N_5295,N_5506);
xnor U7423 (N_7423,N_5081,N_3844);
nand U7424 (N_7424,N_3644,N_5612);
and U7425 (N_7425,N_5968,N_4275);
or U7426 (N_7426,N_3669,N_4121);
nor U7427 (N_7427,N_4884,N_5566);
nor U7428 (N_7428,N_4242,N_5525);
xor U7429 (N_7429,N_3374,N_5192);
or U7430 (N_7430,N_5755,N_5015);
or U7431 (N_7431,N_3808,N_3100);
and U7432 (N_7432,N_5055,N_3014);
or U7433 (N_7433,N_3462,N_4188);
and U7434 (N_7434,N_5107,N_3765);
and U7435 (N_7435,N_3442,N_5414);
xnor U7436 (N_7436,N_4065,N_3803);
nand U7437 (N_7437,N_5847,N_3857);
nor U7438 (N_7438,N_3013,N_5624);
nor U7439 (N_7439,N_3639,N_3763);
nand U7440 (N_7440,N_4015,N_5509);
nand U7441 (N_7441,N_5136,N_4889);
nand U7442 (N_7442,N_5741,N_5520);
xor U7443 (N_7443,N_5611,N_3943);
or U7444 (N_7444,N_3446,N_3161);
nor U7445 (N_7445,N_3704,N_4159);
xnor U7446 (N_7446,N_5006,N_3000);
or U7447 (N_7447,N_5974,N_5793);
nand U7448 (N_7448,N_5804,N_3338);
xor U7449 (N_7449,N_4114,N_3451);
and U7450 (N_7450,N_4658,N_4480);
nand U7451 (N_7451,N_4581,N_5027);
and U7452 (N_7452,N_4695,N_4220);
xor U7453 (N_7453,N_4493,N_5493);
and U7454 (N_7454,N_4886,N_4495);
xor U7455 (N_7455,N_5117,N_4828);
or U7456 (N_7456,N_3344,N_5066);
or U7457 (N_7457,N_3362,N_3851);
nand U7458 (N_7458,N_5940,N_3700);
xnor U7459 (N_7459,N_4892,N_3660);
and U7460 (N_7460,N_5820,N_4550);
and U7461 (N_7461,N_4168,N_3213);
nor U7462 (N_7462,N_4887,N_4001);
nor U7463 (N_7463,N_4987,N_4874);
nor U7464 (N_7464,N_5259,N_4948);
and U7465 (N_7465,N_4317,N_5700);
nor U7466 (N_7466,N_4609,N_3818);
or U7467 (N_7467,N_4288,N_4837);
nor U7468 (N_7468,N_4052,N_3322);
or U7469 (N_7469,N_3783,N_4253);
and U7470 (N_7470,N_4632,N_3774);
xor U7471 (N_7471,N_5552,N_5184);
xor U7472 (N_7472,N_5365,N_4800);
nor U7473 (N_7473,N_5683,N_4059);
nand U7474 (N_7474,N_4116,N_5911);
xor U7475 (N_7475,N_4025,N_4740);
xnor U7476 (N_7476,N_3541,N_5158);
nand U7477 (N_7477,N_5750,N_4610);
or U7478 (N_7478,N_4351,N_4880);
xor U7479 (N_7479,N_4839,N_5573);
nand U7480 (N_7480,N_5196,N_4334);
and U7481 (N_7481,N_4438,N_3652);
and U7482 (N_7482,N_5157,N_5794);
xor U7483 (N_7483,N_5061,N_4646);
nand U7484 (N_7484,N_3733,N_3290);
nand U7485 (N_7485,N_5985,N_5758);
nor U7486 (N_7486,N_3742,N_5749);
nand U7487 (N_7487,N_5670,N_4822);
nand U7488 (N_7488,N_5565,N_3367);
or U7489 (N_7489,N_5699,N_3554);
xnor U7490 (N_7490,N_5256,N_4686);
nor U7491 (N_7491,N_5045,N_5059);
nand U7492 (N_7492,N_4763,N_4558);
nand U7493 (N_7493,N_3412,N_4899);
and U7494 (N_7494,N_5200,N_5071);
nand U7495 (N_7495,N_3011,N_5440);
or U7496 (N_7496,N_4784,N_3623);
and U7497 (N_7497,N_4207,N_3891);
nor U7498 (N_7498,N_3452,N_5507);
nand U7499 (N_7499,N_5214,N_5815);
xor U7500 (N_7500,N_3671,N_3479);
nand U7501 (N_7501,N_3850,N_5033);
nor U7502 (N_7502,N_3131,N_4300);
or U7503 (N_7503,N_5360,N_5198);
or U7504 (N_7504,N_5671,N_5920);
nor U7505 (N_7505,N_3321,N_3561);
xnor U7506 (N_7506,N_5380,N_5083);
or U7507 (N_7507,N_5377,N_3272);
nor U7508 (N_7508,N_3295,N_3202);
nand U7509 (N_7509,N_4742,N_4120);
and U7510 (N_7510,N_5868,N_3457);
nor U7511 (N_7511,N_5115,N_4794);
and U7512 (N_7512,N_5486,N_5478);
or U7513 (N_7513,N_4510,N_5037);
nor U7514 (N_7514,N_3186,N_5837);
nand U7515 (N_7515,N_3460,N_4322);
nand U7516 (N_7516,N_4912,N_5143);
or U7517 (N_7517,N_5515,N_3735);
nor U7518 (N_7518,N_4209,N_3721);
or U7519 (N_7519,N_4309,N_4925);
nand U7520 (N_7520,N_3420,N_4582);
nand U7521 (N_7521,N_4082,N_3980);
or U7522 (N_7522,N_3745,N_4823);
nand U7523 (N_7523,N_3617,N_3088);
xor U7524 (N_7524,N_3893,N_4219);
and U7525 (N_7525,N_4337,N_4970);
nor U7526 (N_7526,N_3143,N_3557);
xor U7527 (N_7527,N_5606,N_3511);
xnor U7528 (N_7528,N_3628,N_4475);
xor U7529 (N_7529,N_4780,N_4708);
or U7530 (N_7530,N_5334,N_3979);
nor U7531 (N_7531,N_3267,N_3138);
xnor U7532 (N_7532,N_5971,N_5519);
nor U7533 (N_7533,N_5105,N_3915);
or U7534 (N_7534,N_5850,N_5532);
and U7535 (N_7535,N_5935,N_3631);
nand U7536 (N_7536,N_5219,N_5785);
nor U7537 (N_7537,N_3185,N_4328);
and U7538 (N_7538,N_4321,N_5152);
nor U7539 (N_7539,N_3346,N_4419);
nand U7540 (N_7540,N_5615,N_5861);
xnor U7541 (N_7541,N_3539,N_3697);
and U7542 (N_7542,N_4206,N_4105);
or U7543 (N_7543,N_3601,N_4651);
or U7544 (N_7544,N_3255,N_4496);
nand U7545 (N_7545,N_5743,N_4995);
nand U7546 (N_7546,N_5828,N_4526);
nor U7547 (N_7547,N_4730,N_3102);
nor U7548 (N_7548,N_4551,N_5517);
nor U7549 (N_7549,N_5085,N_5078);
nor U7550 (N_7550,N_4034,N_3764);
or U7551 (N_7551,N_5819,N_3943);
nand U7552 (N_7552,N_5543,N_5188);
or U7553 (N_7553,N_4160,N_5999);
or U7554 (N_7554,N_5205,N_3829);
or U7555 (N_7555,N_5136,N_3239);
nand U7556 (N_7556,N_3949,N_3731);
and U7557 (N_7557,N_4617,N_5326);
xnor U7558 (N_7558,N_4352,N_4970);
nor U7559 (N_7559,N_4584,N_4211);
nand U7560 (N_7560,N_3889,N_4793);
or U7561 (N_7561,N_5477,N_3718);
xnor U7562 (N_7562,N_3819,N_5037);
nand U7563 (N_7563,N_3164,N_3379);
nor U7564 (N_7564,N_4886,N_3565);
or U7565 (N_7565,N_4722,N_5543);
nand U7566 (N_7566,N_4070,N_5518);
nor U7567 (N_7567,N_3360,N_5484);
nand U7568 (N_7568,N_5026,N_5999);
or U7569 (N_7569,N_5096,N_5664);
nand U7570 (N_7570,N_5959,N_4796);
and U7571 (N_7571,N_4298,N_3504);
or U7572 (N_7572,N_3141,N_4981);
or U7573 (N_7573,N_5574,N_3727);
xnor U7574 (N_7574,N_4642,N_3267);
nor U7575 (N_7575,N_5199,N_3301);
and U7576 (N_7576,N_4291,N_3420);
nand U7577 (N_7577,N_4000,N_4912);
nor U7578 (N_7578,N_3279,N_3097);
nor U7579 (N_7579,N_3054,N_5143);
nor U7580 (N_7580,N_4948,N_5726);
or U7581 (N_7581,N_5904,N_5341);
nor U7582 (N_7582,N_3608,N_3378);
and U7583 (N_7583,N_4150,N_5254);
and U7584 (N_7584,N_3854,N_3033);
nor U7585 (N_7585,N_4338,N_3854);
or U7586 (N_7586,N_3104,N_3505);
or U7587 (N_7587,N_3102,N_4243);
and U7588 (N_7588,N_3337,N_3414);
nor U7589 (N_7589,N_5591,N_4115);
nor U7590 (N_7590,N_3680,N_4522);
nand U7591 (N_7591,N_3000,N_4335);
nor U7592 (N_7592,N_5173,N_4147);
xor U7593 (N_7593,N_5383,N_3174);
xor U7594 (N_7594,N_4657,N_3045);
nor U7595 (N_7595,N_3707,N_4246);
xor U7596 (N_7596,N_3039,N_3808);
nor U7597 (N_7597,N_5090,N_4629);
or U7598 (N_7598,N_5919,N_4924);
or U7599 (N_7599,N_5866,N_3108);
and U7600 (N_7600,N_3945,N_4408);
or U7601 (N_7601,N_5962,N_5783);
nand U7602 (N_7602,N_3698,N_4040);
and U7603 (N_7603,N_4604,N_3086);
nor U7604 (N_7604,N_5950,N_5226);
nand U7605 (N_7605,N_3683,N_4750);
xor U7606 (N_7606,N_3204,N_5750);
nand U7607 (N_7607,N_5170,N_3610);
or U7608 (N_7608,N_5345,N_4917);
nor U7609 (N_7609,N_3460,N_4489);
or U7610 (N_7610,N_3767,N_3887);
xor U7611 (N_7611,N_4393,N_3290);
or U7612 (N_7612,N_5267,N_3733);
nor U7613 (N_7613,N_3333,N_3495);
nor U7614 (N_7614,N_4666,N_5771);
or U7615 (N_7615,N_4141,N_5781);
or U7616 (N_7616,N_5561,N_4180);
and U7617 (N_7617,N_5616,N_5614);
and U7618 (N_7618,N_5044,N_4586);
or U7619 (N_7619,N_5317,N_4653);
or U7620 (N_7620,N_4411,N_5817);
nand U7621 (N_7621,N_3663,N_5426);
nor U7622 (N_7622,N_5283,N_4672);
or U7623 (N_7623,N_4241,N_3260);
or U7624 (N_7624,N_3426,N_5844);
nor U7625 (N_7625,N_3725,N_4116);
or U7626 (N_7626,N_4043,N_5599);
and U7627 (N_7627,N_3656,N_5396);
and U7628 (N_7628,N_5759,N_5463);
xor U7629 (N_7629,N_4608,N_4993);
or U7630 (N_7630,N_5499,N_5453);
or U7631 (N_7631,N_4380,N_5033);
nand U7632 (N_7632,N_5898,N_3635);
xnor U7633 (N_7633,N_3363,N_4973);
nand U7634 (N_7634,N_5201,N_4880);
and U7635 (N_7635,N_5990,N_5228);
nand U7636 (N_7636,N_3263,N_5309);
and U7637 (N_7637,N_5270,N_3640);
or U7638 (N_7638,N_4011,N_5619);
nand U7639 (N_7639,N_5352,N_4766);
and U7640 (N_7640,N_5314,N_4640);
nor U7641 (N_7641,N_3308,N_5817);
nor U7642 (N_7642,N_4658,N_5477);
or U7643 (N_7643,N_4706,N_4532);
nand U7644 (N_7644,N_5399,N_5453);
and U7645 (N_7645,N_5153,N_5177);
nand U7646 (N_7646,N_4778,N_3022);
nand U7647 (N_7647,N_3487,N_3752);
or U7648 (N_7648,N_3199,N_4195);
or U7649 (N_7649,N_5768,N_3026);
and U7650 (N_7650,N_4765,N_3037);
or U7651 (N_7651,N_4333,N_4901);
or U7652 (N_7652,N_4564,N_5141);
or U7653 (N_7653,N_4794,N_5140);
or U7654 (N_7654,N_5853,N_3148);
xnor U7655 (N_7655,N_5597,N_5331);
nand U7656 (N_7656,N_3593,N_5945);
and U7657 (N_7657,N_5199,N_4638);
and U7658 (N_7658,N_3053,N_5848);
xor U7659 (N_7659,N_5948,N_5080);
and U7660 (N_7660,N_5468,N_3944);
or U7661 (N_7661,N_3940,N_4874);
or U7662 (N_7662,N_4853,N_4642);
nor U7663 (N_7663,N_3593,N_4342);
nor U7664 (N_7664,N_5244,N_4387);
xor U7665 (N_7665,N_5037,N_5232);
xnor U7666 (N_7666,N_5491,N_4583);
nand U7667 (N_7667,N_4629,N_3083);
nor U7668 (N_7668,N_4201,N_4755);
nor U7669 (N_7669,N_5230,N_5959);
and U7670 (N_7670,N_4029,N_5431);
nor U7671 (N_7671,N_3399,N_3351);
or U7672 (N_7672,N_5696,N_4192);
xor U7673 (N_7673,N_5818,N_4337);
and U7674 (N_7674,N_3675,N_3575);
and U7675 (N_7675,N_5584,N_3640);
xor U7676 (N_7676,N_4363,N_4347);
nor U7677 (N_7677,N_5685,N_4751);
nor U7678 (N_7678,N_4522,N_4875);
xnor U7679 (N_7679,N_5138,N_3054);
or U7680 (N_7680,N_3269,N_4116);
nand U7681 (N_7681,N_5722,N_5179);
nand U7682 (N_7682,N_5345,N_5588);
xnor U7683 (N_7683,N_5243,N_5742);
nand U7684 (N_7684,N_4243,N_4513);
or U7685 (N_7685,N_5326,N_4828);
nor U7686 (N_7686,N_5154,N_5075);
or U7687 (N_7687,N_3944,N_4270);
or U7688 (N_7688,N_5291,N_5528);
nand U7689 (N_7689,N_5967,N_4731);
and U7690 (N_7690,N_3999,N_4977);
and U7691 (N_7691,N_4550,N_3451);
xor U7692 (N_7692,N_3576,N_3377);
nor U7693 (N_7693,N_5328,N_3976);
and U7694 (N_7694,N_4642,N_4857);
nand U7695 (N_7695,N_5261,N_5677);
nor U7696 (N_7696,N_4656,N_3844);
or U7697 (N_7697,N_4255,N_4481);
and U7698 (N_7698,N_3964,N_5016);
nand U7699 (N_7699,N_4531,N_3847);
xnor U7700 (N_7700,N_3950,N_3886);
and U7701 (N_7701,N_3504,N_5739);
xnor U7702 (N_7702,N_3932,N_5011);
nor U7703 (N_7703,N_4338,N_3630);
or U7704 (N_7704,N_4627,N_3723);
xor U7705 (N_7705,N_3935,N_5219);
xnor U7706 (N_7706,N_3979,N_5308);
or U7707 (N_7707,N_5457,N_3765);
or U7708 (N_7708,N_5475,N_3912);
xor U7709 (N_7709,N_4440,N_4377);
and U7710 (N_7710,N_5889,N_3405);
and U7711 (N_7711,N_3041,N_5701);
or U7712 (N_7712,N_4335,N_4755);
nand U7713 (N_7713,N_5648,N_5272);
xnor U7714 (N_7714,N_4406,N_4429);
or U7715 (N_7715,N_5344,N_5832);
nor U7716 (N_7716,N_5061,N_4476);
nand U7717 (N_7717,N_5769,N_4648);
or U7718 (N_7718,N_5559,N_5961);
xnor U7719 (N_7719,N_5466,N_4221);
and U7720 (N_7720,N_3358,N_5362);
and U7721 (N_7721,N_5435,N_5625);
and U7722 (N_7722,N_4243,N_5907);
or U7723 (N_7723,N_5209,N_3027);
nand U7724 (N_7724,N_3237,N_5986);
nand U7725 (N_7725,N_3261,N_4266);
and U7726 (N_7726,N_4188,N_4411);
nand U7727 (N_7727,N_3908,N_5782);
and U7728 (N_7728,N_3791,N_3594);
and U7729 (N_7729,N_5169,N_4164);
xnor U7730 (N_7730,N_3229,N_4321);
xnor U7731 (N_7731,N_3240,N_4582);
or U7732 (N_7732,N_3676,N_5697);
nand U7733 (N_7733,N_5993,N_4440);
and U7734 (N_7734,N_4771,N_3044);
nand U7735 (N_7735,N_5540,N_4458);
xnor U7736 (N_7736,N_5646,N_5375);
and U7737 (N_7737,N_3673,N_4473);
and U7738 (N_7738,N_4732,N_3623);
and U7739 (N_7739,N_4630,N_3508);
xnor U7740 (N_7740,N_3649,N_3281);
and U7741 (N_7741,N_3470,N_5948);
nor U7742 (N_7742,N_3077,N_5186);
nor U7743 (N_7743,N_3632,N_5592);
and U7744 (N_7744,N_4146,N_4608);
xor U7745 (N_7745,N_4551,N_5552);
nand U7746 (N_7746,N_3502,N_5175);
and U7747 (N_7747,N_4748,N_5683);
or U7748 (N_7748,N_3618,N_5558);
and U7749 (N_7749,N_5743,N_3794);
nor U7750 (N_7750,N_3852,N_3623);
nor U7751 (N_7751,N_5526,N_3861);
nand U7752 (N_7752,N_4354,N_5736);
or U7753 (N_7753,N_4278,N_5620);
nand U7754 (N_7754,N_3740,N_4486);
nor U7755 (N_7755,N_5662,N_5918);
nand U7756 (N_7756,N_4060,N_3625);
nor U7757 (N_7757,N_3980,N_4049);
nand U7758 (N_7758,N_5471,N_4541);
nor U7759 (N_7759,N_3536,N_5366);
nor U7760 (N_7760,N_4963,N_5241);
or U7761 (N_7761,N_5172,N_3533);
and U7762 (N_7762,N_5814,N_3260);
and U7763 (N_7763,N_5310,N_4386);
nand U7764 (N_7764,N_4952,N_5047);
or U7765 (N_7765,N_4151,N_4561);
xor U7766 (N_7766,N_3411,N_4074);
xor U7767 (N_7767,N_4312,N_5772);
or U7768 (N_7768,N_4262,N_4704);
xnor U7769 (N_7769,N_3974,N_3253);
or U7770 (N_7770,N_5676,N_3204);
nor U7771 (N_7771,N_3842,N_4453);
and U7772 (N_7772,N_3347,N_3147);
nor U7773 (N_7773,N_3873,N_5420);
nor U7774 (N_7774,N_4865,N_5028);
and U7775 (N_7775,N_5483,N_4807);
xnor U7776 (N_7776,N_5966,N_3551);
and U7777 (N_7777,N_5744,N_5879);
nand U7778 (N_7778,N_5797,N_5336);
or U7779 (N_7779,N_5410,N_5176);
or U7780 (N_7780,N_3606,N_5041);
nand U7781 (N_7781,N_4619,N_4416);
and U7782 (N_7782,N_3494,N_3699);
or U7783 (N_7783,N_4833,N_4834);
or U7784 (N_7784,N_4082,N_3189);
nand U7785 (N_7785,N_3168,N_3661);
nor U7786 (N_7786,N_4866,N_4403);
nand U7787 (N_7787,N_5468,N_5612);
nand U7788 (N_7788,N_5077,N_5556);
or U7789 (N_7789,N_3165,N_5548);
xor U7790 (N_7790,N_5256,N_3786);
nand U7791 (N_7791,N_4677,N_5405);
nor U7792 (N_7792,N_3354,N_5774);
nor U7793 (N_7793,N_4979,N_4726);
xor U7794 (N_7794,N_4673,N_3213);
or U7795 (N_7795,N_3551,N_4750);
xnor U7796 (N_7796,N_3869,N_4259);
and U7797 (N_7797,N_3860,N_3015);
nand U7798 (N_7798,N_3477,N_4976);
or U7799 (N_7799,N_3573,N_3161);
and U7800 (N_7800,N_4864,N_4132);
and U7801 (N_7801,N_3338,N_5912);
xnor U7802 (N_7802,N_3276,N_4098);
nand U7803 (N_7803,N_3664,N_5998);
nor U7804 (N_7804,N_4096,N_5961);
nor U7805 (N_7805,N_5348,N_5968);
nand U7806 (N_7806,N_5385,N_4048);
xnor U7807 (N_7807,N_4584,N_4445);
nand U7808 (N_7808,N_4990,N_4670);
or U7809 (N_7809,N_4704,N_4335);
nor U7810 (N_7810,N_4333,N_5453);
nor U7811 (N_7811,N_3026,N_3139);
nand U7812 (N_7812,N_4636,N_4073);
nand U7813 (N_7813,N_5218,N_4715);
and U7814 (N_7814,N_5620,N_4394);
nand U7815 (N_7815,N_3484,N_4268);
xor U7816 (N_7816,N_5027,N_4870);
nand U7817 (N_7817,N_5692,N_5715);
or U7818 (N_7818,N_3568,N_4518);
or U7819 (N_7819,N_5967,N_3667);
and U7820 (N_7820,N_3561,N_4291);
nor U7821 (N_7821,N_3936,N_5226);
or U7822 (N_7822,N_3015,N_5915);
nor U7823 (N_7823,N_4585,N_3469);
nor U7824 (N_7824,N_5584,N_3225);
and U7825 (N_7825,N_4843,N_5168);
nand U7826 (N_7826,N_3210,N_5828);
nor U7827 (N_7827,N_3898,N_5252);
xnor U7828 (N_7828,N_5261,N_4685);
nand U7829 (N_7829,N_5240,N_4036);
xnor U7830 (N_7830,N_3813,N_3933);
or U7831 (N_7831,N_3155,N_3957);
nor U7832 (N_7832,N_5909,N_4293);
or U7833 (N_7833,N_5764,N_3999);
and U7834 (N_7834,N_4387,N_4392);
or U7835 (N_7835,N_4814,N_5413);
or U7836 (N_7836,N_3469,N_3298);
nand U7837 (N_7837,N_3423,N_4632);
or U7838 (N_7838,N_5868,N_4931);
nand U7839 (N_7839,N_4080,N_4043);
xor U7840 (N_7840,N_5783,N_5698);
xor U7841 (N_7841,N_5427,N_3425);
xor U7842 (N_7842,N_4886,N_5626);
xor U7843 (N_7843,N_5633,N_4156);
or U7844 (N_7844,N_4821,N_5476);
and U7845 (N_7845,N_4182,N_3055);
nand U7846 (N_7846,N_3403,N_5869);
nand U7847 (N_7847,N_3963,N_4239);
nand U7848 (N_7848,N_4348,N_3870);
nand U7849 (N_7849,N_3188,N_3717);
xor U7850 (N_7850,N_4642,N_3484);
xnor U7851 (N_7851,N_3490,N_3018);
xnor U7852 (N_7852,N_4289,N_4321);
and U7853 (N_7853,N_3303,N_3749);
nor U7854 (N_7854,N_3210,N_3328);
nand U7855 (N_7855,N_4305,N_4521);
and U7856 (N_7856,N_5037,N_5389);
nor U7857 (N_7857,N_5741,N_3138);
and U7858 (N_7858,N_5416,N_5076);
xnor U7859 (N_7859,N_5671,N_5990);
nand U7860 (N_7860,N_4174,N_4124);
xor U7861 (N_7861,N_4994,N_4570);
and U7862 (N_7862,N_4234,N_3354);
nand U7863 (N_7863,N_4002,N_3335);
xor U7864 (N_7864,N_3748,N_3221);
or U7865 (N_7865,N_5426,N_3455);
nand U7866 (N_7866,N_3060,N_5080);
or U7867 (N_7867,N_4489,N_5408);
or U7868 (N_7868,N_5203,N_5194);
nor U7869 (N_7869,N_5723,N_5486);
xor U7870 (N_7870,N_4540,N_3896);
or U7871 (N_7871,N_4588,N_3538);
nor U7872 (N_7872,N_4907,N_4266);
nor U7873 (N_7873,N_3815,N_3991);
nor U7874 (N_7874,N_4217,N_5902);
or U7875 (N_7875,N_5122,N_5369);
nor U7876 (N_7876,N_3178,N_3179);
and U7877 (N_7877,N_4163,N_3544);
nand U7878 (N_7878,N_3663,N_4961);
nor U7879 (N_7879,N_3822,N_5245);
nor U7880 (N_7880,N_5249,N_4162);
nand U7881 (N_7881,N_4285,N_5370);
and U7882 (N_7882,N_5998,N_3142);
nor U7883 (N_7883,N_5304,N_5998);
and U7884 (N_7884,N_4146,N_3519);
nor U7885 (N_7885,N_5509,N_5076);
or U7886 (N_7886,N_4818,N_4527);
xor U7887 (N_7887,N_5505,N_5733);
or U7888 (N_7888,N_3703,N_5127);
xnor U7889 (N_7889,N_5271,N_3355);
xor U7890 (N_7890,N_5249,N_3960);
nor U7891 (N_7891,N_4355,N_4538);
xnor U7892 (N_7892,N_5755,N_4576);
nand U7893 (N_7893,N_3483,N_3543);
and U7894 (N_7894,N_5600,N_4888);
or U7895 (N_7895,N_3584,N_3715);
or U7896 (N_7896,N_5630,N_5054);
xor U7897 (N_7897,N_3297,N_3600);
xnor U7898 (N_7898,N_5367,N_5432);
nand U7899 (N_7899,N_4101,N_4629);
nor U7900 (N_7900,N_3005,N_5709);
nor U7901 (N_7901,N_4554,N_4300);
nand U7902 (N_7902,N_3596,N_5526);
and U7903 (N_7903,N_5374,N_3476);
and U7904 (N_7904,N_4889,N_3723);
nor U7905 (N_7905,N_3763,N_4327);
or U7906 (N_7906,N_5444,N_3229);
nor U7907 (N_7907,N_3777,N_5665);
nor U7908 (N_7908,N_5506,N_3112);
and U7909 (N_7909,N_3829,N_3468);
or U7910 (N_7910,N_4551,N_5887);
xnor U7911 (N_7911,N_3822,N_5653);
nor U7912 (N_7912,N_5691,N_3510);
or U7913 (N_7913,N_5356,N_5142);
nand U7914 (N_7914,N_4709,N_5812);
or U7915 (N_7915,N_5487,N_3571);
nor U7916 (N_7916,N_5137,N_4785);
nand U7917 (N_7917,N_4679,N_4644);
xnor U7918 (N_7918,N_4136,N_3980);
or U7919 (N_7919,N_4128,N_3140);
or U7920 (N_7920,N_4421,N_5617);
nor U7921 (N_7921,N_4366,N_5020);
xor U7922 (N_7922,N_4009,N_3536);
nor U7923 (N_7923,N_3687,N_4622);
or U7924 (N_7924,N_3708,N_3983);
xnor U7925 (N_7925,N_5013,N_4819);
or U7926 (N_7926,N_3399,N_5690);
nand U7927 (N_7927,N_3677,N_3951);
and U7928 (N_7928,N_5266,N_3467);
nor U7929 (N_7929,N_3249,N_5243);
nor U7930 (N_7930,N_5146,N_3734);
or U7931 (N_7931,N_5168,N_5187);
nor U7932 (N_7932,N_5918,N_4935);
nand U7933 (N_7933,N_3052,N_4431);
or U7934 (N_7934,N_4905,N_3409);
nand U7935 (N_7935,N_3101,N_3348);
and U7936 (N_7936,N_5707,N_5060);
nor U7937 (N_7937,N_5599,N_3488);
nor U7938 (N_7938,N_5847,N_3052);
and U7939 (N_7939,N_4764,N_5190);
nand U7940 (N_7940,N_4045,N_3572);
nand U7941 (N_7941,N_5783,N_3117);
nand U7942 (N_7942,N_3224,N_5330);
nand U7943 (N_7943,N_4341,N_4623);
and U7944 (N_7944,N_5741,N_5458);
nor U7945 (N_7945,N_4080,N_4848);
and U7946 (N_7946,N_5518,N_5429);
nor U7947 (N_7947,N_3469,N_4495);
nand U7948 (N_7948,N_4698,N_4522);
and U7949 (N_7949,N_3441,N_5560);
nand U7950 (N_7950,N_4381,N_3742);
or U7951 (N_7951,N_4487,N_4019);
and U7952 (N_7952,N_4771,N_3276);
and U7953 (N_7953,N_4693,N_5588);
nand U7954 (N_7954,N_4214,N_5814);
xor U7955 (N_7955,N_5071,N_4812);
xnor U7956 (N_7956,N_4050,N_3611);
or U7957 (N_7957,N_3332,N_4154);
or U7958 (N_7958,N_3827,N_5918);
or U7959 (N_7959,N_3422,N_4636);
or U7960 (N_7960,N_3474,N_4911);
or U7961 (N_7961,N_5272,N_5908);
and U7962 (N_7962,N_3943,N_4231);
and U7963 (N_7963,N_4841,N_3151);
nor U7964 (N_7964,N_5081,N_4721);
nand U7965 (N_7965,N_5131,N_4796);
xnor U7966 (N_7966,N_5360,N_4692);
or U7967 (N_7967,N_5417,N_3082);
or U7968 (N_7968,N_4931,N_4216);
nand U7969 (N_7969,N_3766,N_5937);
or U7970 (N_7970,N_5412,N_3154);
nand U7971 (N_7971,N_4935,N_3247);
and U7972 (N_7972,N_5140,N_4836);
xnor U7973 (N_7973,N_5228,N_5501);
nor U7974 (N_7974,N_5716,N_5161);
xor U7975 (N_7975,N_3772,N_3789);
xnor U7976 (N_7976,N_4775,N_5819);
nor U7977 (N_7977,N_4510,N_3416);
nand U7978 (N_7978,N_3795,N_5200);
and U7979 (N_7979,N_4852,N_5357);
xor U7980 (N_7980,N_3920,N_5791);
nand U7981 (N_7981,N_3443,N_5945);
nand U7982 (N_7982,N_4373,N_4096);
and U7983 (N_7983,N_3081,N_3152);
and U7984 (N_7984,N_5255,N_3792);
xor U7985 (N_7985,N_3417,N_3529);
or U7986 (N_7986,N_4374,N_5467);
nor U7987 (N_7987,N_4207,N_3757);
xnor U7988 (N_7988,N_5841,N_3464);
xor U7989 (N_7989,N_5287,N_5991);
and U7990 (N_7990,N_5784,N_3687);
nand U7991 (N_7991,N_4371,N_5559);
and U7992 (N_7992,N_3438,N_4175);
nand U7993 (N_7993,N_3373,N_5199);
nand U7994 (N_7994,N_5214,N_4470);
and U7995 (N_7995,N_5209,N_5447);
nor U7996 (N_7996,N_4857,N_3196);
nor U7997 (N_7997,N_5676,N_4327);
or U7998 (N_7998,N_4143,N_5384);
or U7999 (N_7999,N_3257,N_5473);
xnor U8000 (N_8000,N_4203,N_3747);
xnor U8001 (N_8001,N_5568,N_5229);
or U8002 (N_8002,N_5021,N_3885);
nor U8003 (N_8003,N_5248,N_5846);
nand U8004 (N_8004,N_3257,N_3800);
nor U8005 (N_8005,N_4663,N_5591);
nand U8006 (N_8006,N_5514,N_5460);
nor U8007 (N_8007,N_5632,N_5055);
xor U8008 (N_8008,N_5395,N_5862);
nor U8009 (N_8009,N_3690,N_3307);
and U8010 (N_8010,N_3729,N_5830);
or U8011 (N_8011,N_5065,N_5425);
or U8012 (N_8012,N_5235,N_3779);
xnor U8013 (N_8013,N_3138,N_5556);
and U8014 (N_8014,N_5875,N_5831);
and U8015 (N_8015,N_5473,N_4071);
xnor U8016 (N_8016,N_4783,N_3275);
or U8017 (N_8017,N_3703,N_3038);
or U8018 (N_8018,N_5160,N_5401);
or U8019 (N_8019,N_5904,N_4704);
xnor U8020 (N_8020,N_3822,N_3769);
and U8021 (N_8021,N_3916,N_5974);
xnor U8022 (N_8022,N_3865,N_5923);
and U8023 (N_8023,N_3467,N_5907);
nor U8024 (N_8024,N_4428,N_3042);
xor U8025 (N_8025,N_4021,N_4595);
or U8026 (N_8026,N_4607,N_4102);
nand U8027 (N_8027,N_3599,N_5191);
and U8028 (N_8028,N_4053,N_4735);
nand U8029 (N_8029,N_3196,N_3970);
nor U8030 (N_8030,N_4991,N_5052);
or U8031 (N_8031,N_4952,N_4199);
nand U8032 (N_8032,N_5952,N_3070);
xor U8033 (N_8033,N_3941,N_5620);
nor U8034 (N_8034,N_3066,N_3160);
nand U8035 (N_8035,N_3081,N_3849);
nor U8036 (N_8036,N_3503,N_5793);
and U8037 (N_8037,N_5910,N_5723);
nor U8038 (N_8038,N_3888,N_4411);
nand U8039 (N_8039,N_4303,N_3789);
and U8040 (N_8040,N_5095,N_3006);
or U8041 (N_8041,N_3940,N_3560);
and U8042 (N_8042,N_4612,N_3987);
xnor U8043 (N_8043,N_4916,N_4944);
or U8044 (N_8044,N_4468,N_4049);
and U8045 (N_8045,N_3635,N_3542);
and U8046 (N_8046,N_5127,N_3476);
xor U8047 (N_8047,N_5920,N_4766);
xnor U8048 (N_8048,N_3349,N_4238);
or U8049 (N_8049,N_4851,N_4852);
xor U8050 (N_8050,N_5094,N_4892);
xnor U8051 (N_8051,N_3320,N_5289);
xnor U8052 (N_8052,N_5114,N_4018);
xor U8053 (N_8053,N_4417,N_4917);
and U8054 (N_8054,N_3332,N_5127);
or U8055 (N_8055,N_5585,N_4084);
nor U8056 (N_8056,N_4617,N_5895);
or U8057 (N_8057,N_5011,N_4795);
xnor U8058 (N_8058,N_5064,N_3565);
nand U8059 (N_8059,N_5388,N_5837);
nor U8060 (N_8060,N_4088,N_3089);
or U8061 (N_8061,N_3952,N_4360);
nand U8062 (N_8062,N_5870,N_4472);
or U8063 (N_8063,N_4413,N_5635);
or U8064 (N_8064,N_3303,N_4181);
nand U8065 (N_8065,N_5381,N_5532);
xor U8066 (N_8066,N_4237,N_3530);
nor U8067 (N_8067,N_5916,N_4236);
or U8068 (N_8068,N_4651,N_5737);
nor U8069 (N_8069,N_5207,N_4226);
xnor U8070 (N_8070,N_3371,N_4722);
xor U8071 (N_8071,N_5444,N_4517);
xnor U8072 (N_8072,N_4467,N_5815);
nand U8073 (N_8073,N_5153,N_5668);
xnor U8074 (N_8074,N_3402,N_4817);
nand U8075 (N_8075,N_5749,N_3989);
or U8076 (N_8076,N_4672,N_5491);
or U8077 (N_8077,N_5876,N_5715);
xor U8078 (N_8078,N_5967,N_4865);
or U8079 (N_8079,N_4581,N_3593);
xor U8080 (N_8080,N_3649,N_4541);
xnor U8081 (N_8081,N_3333,N_5863);
nor U8082 (N_8082,N_3997,N_5744);
xor U8083 (N_8083,N_5838,N_5333);
xnor U8084 (N_8084,N_5416,N_3689);
and U8085 (N_8085,N_4609,N_3188);
nor U8086 (N_8086,N_4119,N_3135);
xnor U8087 (N_8087,N_3442,N_4969);
nand U8088 (N_8088,N_3444,N_4149);
nand U8089 (N_8089,N_5655,N_3480);
nor U8090 (N_8090,N_5067,N_3553);
or U8091 (N_8091,N_5703,N_4300);
or U8092 (N_8092,N_3327,N_5908);
or U8093 (N_8093,N_5056,N_3082);
nand U8094 (N_8094,N_4063,N_4047);
nor U8095 (N_8095,N_3797,N_4661);
nor U8096 (N_8096,N_3639,N_4903);
xnor U8097 (N_8097,N_3556,N_3998);
or U8098 (N_8098,N_5835,N_5543);
nor U8099 (N_8099,N_5300,N_3902);
nand U8100 (N_8100,N_5343,N_4125);
nand U8101 (N_8101,N_5137,N_4809);
nand U8102 (N_8102,N_3152,N_5173);
xor U8103 (N_8103,N_4153,N_3328);
xnor U8104 (N_8104,N_5698,N_3703);
and U8105 (N_8105,N_3364,N_3108);
nor U8106 (N_8106,N_5841,N_3403);
nor U8107 (N_8107,N_3509,N_5934);
nor U8108 (N_8108,N_5908,N_4082);
xnor U8109 (N_8109,N_3042,N_4791);
xnor U8110 (N_8110,N_5098,N_4327);
nand U8111 (N_8111,N_4853,N_5550);
and U8112 (N_8112,N_5835,N_5968);
nor U8113 (N_8113,N_4669,N_3579);
xor U8114 (N_8114,N_4921,N_3411);
nand U8115 (N_8115,N_5028,N_3758);
nand U8116 (N_8116,N_4217,N_5045);
nor U8117 (N_8117,N_3421,N_5471);
xor U8118 (N_8118,N_5391,N_5118);
nor U8119 (N_8119,N_3990,N_5665);
nor U8120 (N_8120,N_4097,N_5376);
xor U8121 (N_8121,N_4175,N_3958);
nor U8122 (N_8122,N_4227,N_4668);
nor U8123 (N_8123,N_5312,N_4188);
xnor U8124 (N_8124,N_4986,N_4200);
nand U8125 (N_8125,N_4817,N_5712);
xor U8126 (N_8126,N_3418,N_3680);
xor U8127 (N_8127,N_3581,N_3834);
xor U8128 (N_8128,N_5869,N_5424);
nand U8129 (N_8129,N_4154,N_4476);
nor U8130 (N_8130,N_5226,N_4436);
xnor U8131 (N_8131,N_5990,N_4532);
nand U8132 (N_8132,N_3275,N_3319);
nand U8133 (N_8133,N_4998,N_4900);
nand U8134 (N_8134,N_4558,N_3051);
nand U8135 (N_8135,N_5588,N_3084);
and U8136 (N_8136,N_3880,N_3057);
xnor U8137 (N_8137,N_5870,N_5916);
nand U8138 (N_8138,N_3805,N_5530);
nor U8139 (N_8139,N_4894,N_5345);
xor U8140 (N_8140,N_5676,N_3677);
or U8141 (N_8141,N_4044,N_4208);
nand U8142 (N_8142,N_3942,N_3190);
nand U8143 (N_8143,N_4949,N_3444);
and U8144 (N_8144,N_3375,N_4157);
nor U8145 (N_8145,N_3529,N_5494);
nor U8146 (N_8146,N_4285,N_3813);
and U8147 (N_8147,N_5049,N_5667);
and U8148 (N_8148,N_5294,N_3832);
and U8149 (N_8149,N_4978,N_3588);
nand U8150 (N_8150,N_5772,N_4759);
xor U8151 (N_8151,N_5953,N_3852);
and U8152 (N_8152,N_3799,N_5651);
and U8153 (N_8153,N_4756,N_4046);
xnor U8154 (N_8154,N_3855,N_5000);
nor U8155 (N_8155,N_4265,N_5627);
nand U8156 (N_8156,N_3202,N_3957);
nor U8157 (N_8157,N_3214,N_4832);
or U8158 (N_8158,N_4173,N_4441);
xnor U8159 (N_8159,N_4801,N_5675);
and U8160 (N_8160,N_4593,N_4170);
or U8161 (N_8161,N_3195,N_5209);
nand U8162 (N_8162,N_5095,N_5730);
nand U8163 (N_8163,N_3489,N_5122);
or U8164 (N_8164,N_4817,N_4786);
nand U8165 (N_8165,N_4319,N_4714);
xor U8166 (N_8166,N_5794,N_4995);
or U8167 (N_8167,N_4708,N_4357);
or U8168 (N_8168,N_5478,N_3081);
nor U8169 (N_8169,N_4804,N_5184);
nand U8170 (N_8170,N_5780,N_5161);
nor U8171 (N_8171,N_5788,N_3790);
nand U8172 (N_8172,N_5337,N_4433);
nor U8173 (N_8173,N_4841,N_5731);
and U8174 (N_8174,N_5728,N_3170);
nor U8175 (N_8175,N_5908,N_3409);
and U8176 (N_8176,N_4135,N_4317);
xor U8177 (N_8177,N_3332,N_3133);
nor U8178 (N_8178,N_5854,N_4030);
nor U8179 (N_8179,N_5706,N_3540);
nand U8180 (N_8180,N_4413,N_3439);
xnor U8181 (N_8181,N_4095,N_3840);
nor U8182 (N_8182,N_3352,N_4623);
or U8183 (N_8183,N_5280,N_3363);
nor U8184 (N_8184,N_5923,N_4273);
or U8185 (N_8185,N_3223,N_5625);
nand U8186 (N_8186,N_4417,N_5620);
or U8187 (N_8187,N_4594,N_5187);
nand U8188 (N_8188,N_4196,N_4258);
nand U8189 (N_8189,N_4933,N_3009);
nand U8190 (N_8190,N_3641,N_3899);
nand U8191 (N_8191,N_3495,N_3542);
xnor U8192 (N_8192,N_3201,N_4534);
nand U8193 (N_8193,N_4458,N_5563);
nor U8194 (N_8194,N_3552,N_4368);
xnor U8195 (N_8195,N_4026,N_5013);
and U8196 (N_8196,N_3716,N_4079);
nand U8197 (N_8197,N_4016,N_3064);
xor U8198 (N_8198,N_3675,N_5481);
nor U8199 (N_8199,N_4265,N_3289);
and U8200 (N_8200,N_5154,N_4623);
nand U8201 (N_8201,N_3539,N_4747);
and U8202 (N_8202,N_5095,N_3044);
xor U8203 (N_8203,N_4442,N_3647);
or U8204 (N_8204,N_3609,N_5065);
nand U8205 (N_8205,N_4867,N_3217);
nand U8206 (N_8206,N_4609,N_4308);
nor U8207 (N_8207,N_5383,N_5293);
or U8208 (N_8208,N_3945,N_3936);
nor U8209 (N_8209,N_3960,N_3751);
nand U8210 (N_8210,N_3742,N_4404);
xnor U8211 (N_8211,N_5093,N_4346);
xor U8212 (N_8212,N_4669,N_5185);
or U8213 (N_8213,N_3477,N_3464);
or U8214 (N_8214,N_3973,N_3387);
nand U8215 (N_8215,N_4404,N_4498);
xor U8216 (N_8216,N_5847,N_4982);
nand U8217 (N_8217,N_4224,N_4183);
and U8218 (N_8218,N_3207,N_4491);
nand U8219 (N_8219,N_5940,N_5975);
and U8220 (N_8220,N_4556,N_4257);
or U8221 (N_8221,N_4138,N_3494);
nor U8222 (N_8222,N_4362,N_3228);
nand U8223 (N_8223,N_3281,N_5675);
or U8224 (N_8224,N_3230,N_5068);
and U8225 (N_8225,N_3963,N_4042);
and U8226 (N_8226,N_4669,N_5525);
nand U8227 (N_8227,N_5250,N_5506);
xnor U8228 (N_8228,N_5057,N_4036);
or U8229 (N_8229,N_3073,N_3888);
or U8230 (N_8230,N_4267,N_3673);
nand U8231 (N_8231,N_3747,N_3470);
xor U8232 (N_8232,N_4449,N_5461);
nand U8233 (N_8233,N_5632,N_5907);
nor U8234 (N_8234,N_4669,N_3308);
nand U8235 (N_8235,N_5044,N_3345);
or U8236 (N_8236,N_4369,N_5669);
and U8237 (N_8237,N_3034,N_5184);
or U8238 (N_8238,N_5460,N_5256);
nand U8239 (N_8239,N_3552,N_3675);
nand U8240 (N_8240,N_5339,N_3326);
and U8241 (N_8241,N_3400,N_3473);
and U8242 (N_8242,N_4703,N_4677);
nand U8243 (N_8243,N_3308,N_5917);
nand U8244 (N_8244,N_5666,N_3217);
or U8245 (N_8245,N_5356,N_4480);
and U8246 (N_8246,N_3918,N_5818);
nand U8247 (N_8247,N_5462,N_5363);
and U8248 (N_8248,N_3001,N_3417);
and U8249 (N_8249,N_3377,N_3738);
nand U8250 (N_8250,N_4572,N_3209);
nor U8251 (N_8251,N_3164,N_5677);
nand U8252 (N_8252,N_4421,N_5263);
and U8253 (N_8253,N_4940,N_4100);
nor U8254 (N_8254,N_5970,N_4606);
or U8255 (N_8255,N_3399,N_5440);
nand U8256 (N_8256,N_5504,N_5684);
nand U8257 (N_8257,N_4965,N_4295);
and U8258 (N_8258,N_4804,N_5015);
nor U8259 (N_8259,N_5521,N_5734);
nand U8260 (N_8260,N_4242,N_3917);
or U8261 (N_8261,N_5005,N_3479);
xnor U8262 (N_8262,N_3149,N_5145);
nand U8263 (N_8263,N_4171,N_4554);
xnor U8264 (N_8264,N_3892,N_5135);
or U8265 (N_8265,N_5600,N_5533);
nand U8266 (N_8266,N_4251,N_4816);
and U8267 (N_8267,N_5847,N_4187);
xor U8268 (N_8268,N_4153,N_4730);
xnor U8269 (N_8269,N_5676,N_5673);
xnor U8270 (N_8270,N_3637,N_5598);
xor U8271 (N_8271,N_3810,N_5537);
nor U8272 (N_8272,N_4831,N_3596);
xnor U8273 (N_8273,N_5117,N_5485);
or U8274 (N_8274,N_3281,N_5411);
nor U8275 (N_8275,N_4562,N_5657);
xor U8276 (N_8276,N_5850,N_3469);
xor U8277 (N_8277,N_3420,N_4359);
xnor U8278 (N_8278,N_3029,N_5513);
or U8279 (N_8279,N_3990,N_5403);
xnor U8280 (N_8280,N_4951,N_4231);
xor U8281 (N_8281,N_3497,N_3809);
and U8282 (N_8282,N_5136,N_4886);
nor U8283 (N_8283,N_3023,N_3533);
or U8284 (N_8284,N_5795,N_5365);
nand U8285 (N_8285,N_5204,N_5621);
nor U8286 (N_8286,N_3113,N_4620);
or U8287 (N_8287,N_3927,N_4937);
and U8288 (N_8288,N_4401,N_3534);
nand U8289 (N_8289,N_3068,N_4134);
and U8290 (N_8290,N_3210,N_3348);
nor U8291 (N_8291,N_5796,N_4050);
xor U8292 (N_8292,N_4457,N_5496);
nand U8293 (N_8293,N_4737,N_5953);
xor U8294 (N_8294,N_3802,N_4465);
nand U8295 (N_8295,N_3575,N_4904);
nand U8296 (N_8296,N_3036,N_4527);
xnor U8297 (N_8297,N_5059,N_5730);
xnor U8298 (N_8298,N_5559,N_3897);
or U8299 (N_8299,N_3903,N_4996);
and U8300 (N_8300,N_3366,N_3623);
nor U8301 (N_8301,N_3292,N_5104);
xnor U8302 (N_8302,N_4178,N_4409);
nor U8303 (N_8303,N_4485,N_3008);
and U8304 (N_8304,N_3116,N_5792);
and U8305 (N_8305,N_3382,N_3601);
nor U8306 (N_8306,N_3467,N_5380);
or U8307 (N_8307,N_3238,N_5404);
and U8308 (N_8308,N_3704,N_4384);
nor U8309 (N_8309,N_3270,N_3061);
nor U8310 (N_8310,N_5272,N_4980);
xnor U8311 (N_8311,N_5896,N_4842);
and U8312 (N_8312,N_5222,N_4509);
nor U8313 (N_8313,N_3947,N_5604);
xnor U8314 (N_8314,N_5786,N_3817);
and U8315 (N_8315,N_5875,N_3283);
nor U8316 (N_8316,N_4520,N_5795);
nand U8317 (N_8317,N_3636,N_3194);
and U8318 (N_8318,N_4055,N_4149);
nor U8319 (N_8319,N_4894,N_4869);
and U8320 (N_8320,N_5596,N_5062);
nor U8321 (N_8321,N_4097,N_3565);
and U8322 (N_8322,N_5415,N_4706);
nand U8323 (N_8323,N_3824,N_5326);
xor U8324 (N_8324,N_3891,N_3363);
xnor U8325 (N_8325,N_5223,N_5590);
nor U8326 (N_8326,N_3812,N_4857);
or U8327 (N_8327,N_5601,N_3597);
xor U8328 (N_8328,N_3002,N_4093);
xor U8329 (N_8329,N_5493,N_5933);
nand U8330 (N_8330,N_3835,N_5987);
nand U8331 (N_8331,N_4198,N_4752);
xnor U8332 (N_8332,N_5893,N_5667);
xnor U8333 (N_8333,N_3463,N_4911);
xor U8334 (N_8334,N_5436,N_5052);
nor U8335 (N_8335,N_4229,N_5713);
nor U8336 (N_8336,N_5242,N_5185);
xnor U8337 (N_8337,N_3571,N_5356);
or U8338 (N_8338,N_3250,N_3470);
and U8339 (N_8339,N_3349,N_5993);
or U8340 (N_8340,N_4831,N_3192);
or U8341 (N_8341,N_4521,N_4499);
nand U8342 (N_8342,N_5568,N_3261);
xor U8343 (N_8343,N_3705,N_5055);
nand U8344 (N_8344,N_4864,N_3378);
nor U8345 (N_8345,N_4168,N_3616);
and U8346 (N_8346,N_3656,N_3231);
or U8347 (N_8347,N_4614,N_5260);
or U8348 (N_8348,N_4340,N_5315);
xnor U8349 (N_8349,N_5339,N_3133);
xor U8350 (N_8350,N_4888,N_5510);
xor U8351 (N_8351,N_4633,N_3874);
nor U8352 (N_8352,N_3564,N_4036);
nand U8353 (N_8353,N_5101,N_3109);
xor U8354 (N_8354,N_3644,N_5472);
or U8355 (N_8355,N_3460,N_4364);
nand U8356 (N_8356,N_3634,N_5421);
or U8357 (N_8357,N_3372,N_3476);
nand U8358 (N_8358,N_4894,N_3561);
nand U8359 (N_8359,N_4825,N_3417);
and U8360 (N_8360,N_3424,N_4561);
nor U8361 (N_8361,N_5419,N_5201);
nor U8362 (N_8362,N_3198,N_3617);
xor U8363 (N_8363,N_5907,N_4268);
xor U8364 (N_8364,N_4720,N_4607);
nor U8365 (N_8365,N_3308,N_5657);
nor U8366 (N_8366,N_4908,N_5146);
or U8367 (N_8367,N_3292,N_5079);
or U8368 (N_8368,N_4491,N_4567);
nor U8369 (N_8369,N_4499,N_5253);
nand U8370 (N_8370,N_3120,N_4706);
nor U8371 (N_8371,N_5371,N_5051);
xnor U8372 (N_8372,N_4578,N_5314);
xor U8373 (N_8373,N_3074,N_3823);
nor U8374 (N_8374,N_4774,N_3842);
and U8375 (N_8375,N_3695,N_3597);
xor U8376 (N_8376,N_5830,N_3436);
nand U8377 (N_8377,N_3358,N_5524);
xnor U8378 (N_8378,N_3306,N_3777);
nand U8379 (N_8379,N_4024,N_4833);
xor U8380 (N_8380,N_4493,N_4323);
nor U8381 (N_8381,N_4052,N_4451);
or U8382 (N_8382,N_4375,N_3404);
and U8383 (N_8383,N_5614,N_3918);
xor U8384 (N_8384,N_3193,N_5024);
nor U8385 (N_8385,N_5825,N_3257);
or U8386 (N_8386,N_5939,N_3332);
and U8387 (N_8387,N_4333,N_3164);
nor U8388 (N_8388,N_4562,N_4356);
xor U8389 (N_8389,N_5436,N_3242);
nor U8390 (N_8390,N_5717,N_4523);
nand U8391 (N_8391,N_4168,N_4631);
or U8392 (N_8392,N_4190,N_3582);
nand U8393 (N_8393,N_3894,N_4343);
or U8394 (N_8394,N_4224,N_3913);
nor U8395 (N_8395,N_5667,N_3858);
or U8396 (N_8396,N_3680,N_3885);
nor U8397 (N_8397,N_4121,N_5075);
and U8398 (N_8398,N_3675,N_5461);
nand U8399 (N_8399,N_4420,N_5154);
and U8400 (N_8400,N_4272,N_3021);
nor U8401 (N_8401,N_4861,N_3926);
nand U8402 (N_8402,N_4595,N_4824);
xnor U8403 (N_8403,N_5084,N_5553);
or U8404 (N_8404,N_4443,N_5683);
nand U8405 (N_8405,N_4505,N_3277);
nand U8406 (N_8406,N_4983,N_3759);
nand U8407 (N_8407,N_4949,N_4247);
xnor U8408 (N_8408,N_4839,N_3317);
and U8409 (N_8409,N_5467,N_3798);
nand U8410 (N_8410,N_3099,N_5272);
nand U8411 (N_8411,N_3286,N_4433);
nand U8412 (N_8412,N_3135,N_3626);
xnor U8413 (N_8413,N_3725,N_4012);
and U8414 (N_8414,N_3965,N_5504);
nor U8415 (N_8415,N_4873,N_4674);
nor U8416 (N_8416,N_4218,N_5579);
nor U8417 (N_8417,N_3553,N_4295);
and U8418 (N_8418,N_5666,N_5095);
nand U8419 (N_8419,N_3071,N_4603);
and U8420 (N_8420,N_4829,N_4037);
or U8421 (N_8421,N_4941,N_3772);
nand U8422 (N_8422,N_4456,N_5216);
and U8423 (N_8423,N_3613,N_3628);
nand U8424 (N_8424,N_5747,N_4582);
nand U8425 (N_8425,N_4630,N_3723);
xnor U8426 (N_8426,N_4257,N_3853);
or U8427 (N_8427,N_3194,N_4935);
xnor U8428 (N_8428,N_3052,N_3805);
xor U8429 (N_8429,N_5811,N_5967);
nor U8430 (N_8430,N_5148,N_3596);
nand U8431 (N_8431,N_4790,N_3352);
or U8432 (N_8432,N_4161,N_5013);
nor U8433 (N_8433,N_3210,N_5646);
nor U8434 (N_8434,N_4510,N_4193);
nand U8435 (N_8435,N_5751,N_3395);
nand U8436 (N_8436,N_5282,N_3342);
and U8437 (N_8437,N_4990,N_4412);
nor U8438 (N_8438,N_3946,N_5552);
and U8439 (N_8439,N_3911,N_5251);
or U8440 (N_8440,N_4592,N_5730);
nand U8441 (N_8441,N_4775,N_3239);
and U8442 (N_8442,N_3717,N_3622);
or U8443 (N_8443,N_3939,N_5609);
xor U8444 (N_8444,N_3848,N_5770);
xor U8445 (N_8445,N_4529,N_5214);
and U8446 (N_8446,N_4053,N_4162);
nand U8447 (N_8447,N_3010,N_5614);
xor U8448 (N_8448,N_3550,N_3387);
or U8449 (N_8449,N_3809,N_3141);
nand U8450 (N_8450,N_3315,N_5848);
and U8451 (N_8451,N_5936,N_4298);
xor U8452 (N_8452,N_5068,N_4276);
and U8453 (N_8453,N_3006,N_5363);
nor U8454 (N_8454,N_3143,N_3844);
nor U8455 (N_8455,N_4232,N_3237);
or U8456 (N_8456,N_3363,N_4003);
nor U8457 (N_8457,N_5066,N_5222);
and U8458 (N_8458,N_3850,N_4411);
or U8459 (N_8459,N_4119,N_5546);
xor U8460 (N_8460,N_4714,N_3940);
or U8461 (N_8461,N_4731,N_4909);
and U8462 (N_8462,N_5454,N_5048);
and U8463 (N_8463,N_5466,N_5782);
or U8464 (N_8464,N_5018,N_3950);
xnor U8465 (N_8465,N_5095,N_4177);
nor U8466 (N_8466,N_3000,N_4873);
xnor U8467 (N_8467,N_3809,N_3828);
and U8468 (N_8468,N_5022,N_3430);
xnor U8469 (N_8469,N_3586,N_3858);
or U8470 (N_8470,N_4164,N_5829);
or U8471 (N_8471,N_3842,N_3721);
nand U8472 (N_8472,N_3661,N_5302);
nor U8473 (N_8473,N_4458,N_4016);
and U8474 (N_8474,N_4255,N_5754);
xnor U8475 (N_8475,N_3353,N_3220);
or U8476 (N_8476,N_4084,N_3158);
nor U8477 (N_8477,N_4645,N_3718);
and U8478 (N_8478,N_3892,N_5972);
and U8479 (N_8479,N_5442,N_3303);
nand U8480 (N_8480,N_5141,N_3898);
nand U8481 (N_8481,N_3499,N_5515);
nor U8482 (N_8482,N_4189,N_4689);
and U8483 (N_8483,N_3584,N_3849);
or U8484 (N_8484,N_3903,N_5445);
nand U8485 (N_8485,N_5882,N_4117);
xnor U8486 (N_8486,N_4344,N_5641);
xor U8487 (N_8487,N_4613,N_5125);
xnor U8488 (N_8488,N_3789,N_4897);
nor U8489 (N_8489,N_4181,N_5373);
and U8490 (N_8490,N_3492,N_4109);
nor U8491 (N_8491,N_4276,N_3148);
or U8492 (N_8492,N_3350,N_3863);
xnor U8493 (N_8493,N_3068,N_4808);
nor U8494 (N_8494,N_5631,N_5796);
nor U8495 (N_8495,N_3416,N_4440);
and U8496 (N_8496,N_5537,N_4022);
nand U8497 (N_8497,N_5867,N_3779);
and U8498 (N_8498,N_4039,N_3366);
xor U8499 (N_8499,N_5123,N_5843);
and U8500 (N_8500,N_4420,N_4919);
and U8501 (N_8501,N_5355,N_4068);
and U8502 (N_8502,N_4353,N_4883);
nor U8503 (N_8503,N_3789,N_4136);
nor U8504 (N_8504,N_3752,N_5720);
xor U8505 (N_8505,N_5649,N_3037);
nand U8506 (N_8506,N_4278,N_4632);
or U8507 (N_8507,N_3630,N_5001);
or U8508 (N_8508,N_4024,N_3698);
xnor U8509 (N_8509,N_3326,N_4468);
and U8510 (N_8510,N_3886,N_3553);
or U8511 (N_8511,N_3876,N_5419);
xnor U8512 (N_8512,N_4152,N_4989);
nand U8513 (N_8513,N_5993,N_4020);
or U8514 (N_8514,N_4626,N_3023);
nand U8515 (N_8515,N_5271,N_5817);
or U8516 (N_8516,N_5328,N_4704);
nor U8517 (N_8517,N_3029,N_5255);
or U8518 (N_8518,N_4574,N_5184);
nor U8519 (N_8519,N_5096,N_5054);
or U8520 (N_8520,N_4745,N_5206);
nand U8521 (N_8521,N_4737,N_5661);
and U8522 (N_8522,N_5589,N_5832);
nor U8523 (N_8523,N_4659,N_4683);
or U8524 (N_8524,N_3257,N_5003);
and U8525 (N_8525,N_4116,N_4615);
nand U8526 (N_8526,N_5763,N_3855);
xor U8527 (N_8527,N_5927,N_5638);
and U8528 (N_8528,N_4400,N_5417);
or U8529 (N_8529,N_4026,N_3587);
nand U8530 (N_8530,N_5698,N_3642);
xnor U8531 (N_8531,N_4073,N_4662);
and U8532 (N_8532,N_4585,N_5621);
and U8533 (N_8533,N_3248,N_3849);
xor U8534 (N_8534,N_4619,N_4545);
and U8535 (N_8535,N_4246,N_3101);
nand U8536 (N_8536,N_4559,N_5601);
nor U8537 (N_8537,N_5463,N_4511);
nor U8538 (N_8538,N_5824,N_5820);
nand U8539 (N_8539,N_4044,N_5637);
nor U8540 (N_8540,N_5551,N_3622);
and U8541 (N_8541,N_5454,N_5332);
or U8542 (N_8542,N_5602,N_3289);
nor U8543 (N_8543,N_3626,N_5885);
nand U8544 (N_8544,N_4011,N_5235);
and U8545 (N_8545,N_3231,N_5033);
xnor U8546 (N_8546,N_5219,N_4609);
xor U8547 (N_8547,N_4337,N_3556);
xor U8548 (N_8548,N_4947,N_3675);
and U8549 (N_8549,N_3053,N_3572);
xor U8550 (N_8550,N_5842,N_4738);
nand U8551 (N_8551,N_4939,N_3883);
nor U8552 (N_8552,N_4409,N_4072);
or U8553 (N_8553,N_5243,N_3685);
or U8554 (N_8554,N_5581,N_3398);
nand U8555 (N_8555,N_5953,N_5248);
or U8556 (N_8556,N_3866,N_5040);
xor U8557 (N_8557,N_5031,N_3011);
xnor U8558 (N_8558,N_3574,N_3991);
and U8559 (N_8559,N_4261,N_5854);
or U8560 (N_8560,N_4865,N_4395);
nand U8561 (N_8561,N_4682,N_4323);
or U8562 (N_8562,N_5580,N_4551);
xor U8563 (N_8563,N_4515,N_4703);
xnor U8564 (N_8564,N_5916,N_5947);
and U8565 (N_8565,N_4504,N_3023);
or U8566 (N_8566,N_4173,N_4118);
xor U8567 (N_8567,N_4355,N_5976);
xor U8568 (N_8568,N_5641,N_4820);
or U8569 (N_8569,N_3694,N_4592);
nand U8570 (N_8570,N_5453,N_3401);
nor U8571 (N_8571,N_3152,N_5981);
or U8572 (N_8572,N_4444,N_4063);
nand U8573 (N_8573,N_3262,N_5820);
xor U8574 (N_8574,N_4255,N_4246);
and U8575 (N_8575,N_4610,N_4893);
nor U8576 (N_8576,N_4425,N_3843);
nor U8577 (N_8577,N_5143,N_4084);
nor U8578 (N_8578,N_5353,N_3604);
or U8579 (N_8579,N_3429,N_4559);
or U8580 (N_8580,N_3902,N_3283);
or U8581 (N_8581,N_4880,N_3679);
nor U8582 (N_8582,N_5479,N_3775);
or U8583 (N_8583,N_5436,N_4088);
nand U8584 (N_8584,N_3791,N_5340);
and U8585 (N_8585,N_5887,N_4097);
or U8586 (N_8586,N_5872,N_3103);
nand U8587 (N_8587,N_4167,N_3369);
or U8588 (N_8588,N_4621,N_4743);
and U8589 (N_8589,N_4423,N_3628);
nor U8590 (N_8590,N_5626,N_5133);
nor U8591 (N_8591,N_4256,N_4645);
nand U8592 (N_8592,N_5370,N_3921);
or U8593 (N_8593,N_3767,N_3618);
and U8594 (N_8594,N_4087,N_3388);
or U8595 (N_8595,N_3499,N_3674);
or U8596 (N_8596,N_3334,N_4699);
nor U8597 (N_8597,N_4036,N_3698);
nor U8598 (N_8598,N_5849,N_4437);
or U8599 (N_8599,N_3903,N_4993);
or U8600 (N_8600,N_4018,N_4679);
nand U8601 (N_8601,N_5083,N_4324);
nor U8602 (N_8602,N_4881,N_3067);
xor U8603 (N_8603,N_3334,N_3968);
nand U8604 (N_8604,N_4182,N_3932);
nor U8605 (N_8605,N_5239,N_3460);
nand U8606 (N_8606,N_3419,N_5596);
nand U8607 (N_8607,N_5142,N_3003);
nor U8608 (N_8608,N_3646,N_4580);
and U8609 (N_8609,N_4737,N_3828);
or U8610 (N_8610,N_5605,N_3951);
nor U8611 (N_8611,N_5651,N_5600);
nor U8612 (N_8612,N_4143,N_5103);
nand U8613 (N_8613,N_3084,N_3466);
nand U8614 (N_8614,N_3181,N_4236);
xor U8615 (N_8615,N_5446,N_3899);
xnor U8616 (N_8616,N_3863,N_3724);
nor U8617 (N_8617,N_4056,N_4803);
nand U8618 (N_8618,N_5925,N_3338);
or U8619 (N_8619,N_3862,N_5030);
xnor U8620 (N_8620,N_4267,N_5271);
and U8621 (N_8621,N_4481,N_3705);
xnor U8622 (N_8622,N_3216,N_3148);
xor U8623 (N_8623,N_3060,N_4908);
nor U8624 (N_8624,N_5722,N_3273);
or U8625 (N_8625,N_5737,N_3333);
nand U8626 (N_8626,N_5743,N_3470);
xnor U8627 (N_8627,N_4243,N_3588);
and U8628 (N_8628,N_4292,N_5293);
xnor U8629 (N_8629,N_4370,N_4227);
xor U8630 (N_8630,N_3783,N_3704);
nand U8631 (N_8631,N_4745,N_5294);
or U8632 (N_8632,N_3878,N_5053);
and U8633 (N_8633,N_3890,N_5781);
and U8634 (N_8634,N_3232,N_4761);
xnor U8635 (N_8635,N_4478,N_3046);
and U8636 (N_8636,N_5438,N_3602);
or U8637 (N_8637,N_3033,N_4995);
nor U8638 (N_8638,N_4015,N_3944);
xnor U8639 (N_8639,N_3228,N_4571);
and U8640 (N_8640,N_5341,N_3039);
or U8641 (N_8641,N_3006,N_3046);
nand U8642 (N_8642,N_3672,N_4346);
or U8643 (N_8643,N_3842,N_5720);
nand U8644 (N_8644,N_3622,N_3381);
nand U8645 (N_8645,N_4161,N_3361);
or U8646 (N_8646,N_4195,N_5147);
nor U8647 (N_8647,N_5484,N_4500);
xor U8648 (N_8648,N_3706,N_4141);
nor U8649 (N_8649,N_4145,N_3194);
xor U8650 (N_8650,N_5953,N_5199);
and U8651 (N_8651,N_3619,N_4912);
nand U8652 (N_8652,N_5889,N_3560);
xor U8653 (N_8653,N_3671,N_5412);
nor U8654 (N_8654,N_3368,N_4026);
nor U8655 (N_8655,N_5176,N_5714);
nand U8656 (N_8656,N_4807,N_3918);
or U8657 (N_8657,N_5980,N_4196);
nor U8658 (N_8658,N_3842,N_5806);
nand U8659 (N_8659,N_5968,N_5127);
nor U8660 (N_8660,N_4953,N_4538);
nand U8661 (N_8661,N_5631,N_3099);
nand U8662 (N_8662,N_3055,N_5445);
or U8663 (N_8663,N_5888,N_5454);
nor U8664 (N_8664,N_4798,N_4811);
or U8665 (N_8665,N_3453,N_3328);
nor U8666 (N_8666,N_4374,N_3807);
and U8667 (N_8667,N_5712,N_4422);
and U8668 (N_8668,N_5807,N_5692);
xnor U8669 (N_8669,N_4003,N_4788);
nor U8670 (N_8670,N_3144,N_3990);
or U8671 (N_8671,N_4135,N_5397);
nand U8672 (N_8672,N_4417,N_5798);
or U8673 (N_8673,N_4211,N_3515);
xor U8674 (N_8674,N_4219,N_4812);
nor U8675 (N_8675,N_4883,N_4588);
nand U8676 (N_8676,N_5608,N_3438);
nand U8677 (N_8677,N_5654,N_5453);
and U8678 (N_8678,N_4919,N_3660);
nand U8679 (N_8679,N_5077,N_4827);
and U8680 (N_8680,N_3502,N_4201);
and U8681 (N_8681,N_4547,N_4021);
nor U8682 (N_8682,N_3769,N_4785);
nor U8683 (N_8683,N_4223,N_4238);
and U8684 (N_8684,N_5515,N_5265);
nand U8685 (N_8685,N_5650,N_3515);
nand U8686 (N_8686,N_5957,N_4014);
and U8687 (N_8687,N_4387,N_5526);
nand U8688 (N_8688,N_3455,N_3743);
nand U8689 (N_8689,N_5235,N_5308);
and U8690 (N_8690,N_3229,N_3466);
nand U8691 (N_8691,N_5831,N_5963);
nand U8692 (N_8692,N_3364,N_5049);
nor U8693 (N_8693,N_5288,N_4866);
xnor U8694 (N_8694,N_5791,N_5756);
nor U8695 (N_8695,N_4593,N_3320);
nand U8696 (N_8696,N_5482,N_5367);
nand U8697 (N_8697,N_4546,N_5782);
or U8698 (N_8698,N_4118,N_3038);
nand U8699 (N_8699,N_3278,N_5476);
and U8700 (N_8700,N_5274,N_3362);
and U8701 (N_8701,N_4495,N_4631);
nand U8702 (N_8702,N_5418,N_4843);
xnor U8703 (N_8703,N_3841,N_4487);
nor U8704 (N_8704,N_5845,N_5758);
nand U8705 (N_8705,N_5490,N_4021);
or U8706 (N_8706,N_3264,N_5970);
or U8707 (N_8707,N_5250,N_5400);
or U8708 (N_8708,N_4196,N_4839);
and U8709 (N_8709,N_3036,N_5139);
nand U8710 (N_8710,N_3132,N_5817);
nand U8711 (N_8711,N_3526,N_3123);
xnor U8712 (N_8712,N_3033,N_3827);
nand U8713 (N_8713,N_4995,N_4529);
and U8714 (N_8714,N_3956,N_4097);
or U8715 (N_8715,N_4974,N_4118);
and U8716 (N_8716,N_3519,N_3818);
and U8717 (N_8717,N_3106,N_4305);
and U8718 (N_8718,N_5732,N_5227);
xnor U8719 (N_8719,N_3805,N_3027);
nand U8720 (N_8720,N_5891,N_3246);
and U8721 (N_8721,N_5656,N_4877);
nor U8722 (N_8722,N_4005,N_4410);
nor U8723 (N_8723,N_5975,N_4456);
nand U8724 (N_8724,N_3014,N_4029);
nand U8725 (N_8725,N_5011,N_5186);
nand U8726 (N_8726,N_5296,N_3082);
xor U8727 (N_8727,N_4676,N_3545);
xnor U8728 (N_8728,N_3294,N_4107);
and U8729 (N_8729,N_4170,N_5987);
nand U8730 (N_8730,N_5687,N_4345);
and U8731 (N_8731,N_4379,N_3845);
nand U8732 (N_8732,N_3545,N_5044);
nand U8733 (N_8733,N_3035,N_5489);
nand U8734 (N_8734,N_4381,N_5854);
nand U8735 (N_8735,N_5242,N_3276);
and U8736 (N_8736,N_4323,N_3290);
or U8737 (N_8737,N_5073,N_3362);
nor U8738 (N_8738,N_4946,N_4796);
and U8739 (N_8739,N_4229,N_4045);
and U8740 (N_8740,N_3502,N_4946);
nand U8741 (N_8741,N_3552,N_3983);
nand U8742 (N_8742,N_4714,N_3882);
and U8743 (N_8743,N_3272,N_5462);
xor U8744 (N_8744,N_3944,N_3845);
nand U8745 (N_8745,N_5047,N_4468);
nand U8746 (N_8746,N_5531,N_5950);
nand U8747 (N_8747,N_3722,N_5412);
nand U8748 (N_8748,N_4249,N_4959);
and U8749 (N_8749,N_4574,N_3177);
and U8750 (N_8750,N_4784,N_5128);
and U8751 (N_8751,N_4189,N_4993);
nand U8752 (N_8752,N_5385,N_5880);
and U8753 (N_8753,N_4887,N_5158);
xnor U8754 (N_8754,N_4410,N_4330);
and U8755 (N_8755,N_3564,N_3380);
and U8756 (N_8756,N_3476,N_5743);
xnor U8757 (N_8757,N_4451,N_3855);
nor U8758 (N_8758,N_5572,N_5846);
and U8759 (N_8759,N_3231,N_4609);
xor U8760 (N_8760,N_3496,N_5358);
xnor U8761 (N_8761,N_5339,N_3518);
nand U8762 (N_8762,N_5407,N_3017);
nor U8763 (N_8763,N_3426,N_5875);
nand U8764 (N_8764,N_4536,N_5476);
nand U8765 (N_8765,N_3317,N_3017);
nor U8766 (N_8766,N_3059,N_3986);
and U8767 (N_8767,N_3103,N_3118);
or U8768 (N_8768,N_3768,N_3201);
or U8769 (N_8769,N_4556,N_5231);
xor U8770 (N_8770,N_5139,N_3757);
xor U8771 (N_8771,N_3622,N_3588);
nand U8772 (N_8772,N_3061,N_3990);
or U8773 (N_8773,N_4369,N_4497);
nand U8774 (N_8774,N_4338,N_3768);
nor U8775 (N_8775,N_4483,N_5164);
nor U8776 (N_8776,N_5802,N_5560);
or U8777 (N_8777,N_3466,N_5403);
nand U8778 (N_8778,N_4897,N_3198);
nand U8779 (N_8779,N_4755,N_5945);
or U8780 (N_8780,N_3718,N_5741);
or U8781 (N_8781,N_5998,N_4097);
xor U8782 (N_8782,N_5100,N_4690);
or U8783 (N_8783,N_3470,N_3427);
and U8784 (N_8784,N_3535,N_3636);
nand U8785 (N_8785,N_5779,N_5865);
xor U8786 (N_8786,N_5145,N_3785);
or U8787 (N_8787,N_4985,N_5694);
or U8788 (N_8788,N_4135,N_4323);
nand U8789 (N_8789,N_4132,N_5988);
nand U8790 (N_8790,N_3495,N_3880);
xor U8791 (N_8791,N_3686,N_5257);
xor U8792 (N_8792,N_5537,N_5022);
and U8793 (N_8793,N_3234,N_5019);
or U8794 (N_8794,N_5188,N_4217);
or U8795 (N_8795,N_3254,N_5105);
nand U8796 (N_8796,N_5467,N_4166);
xnor U8797 (N_8797,N_5462,N_5121);
nand U8798 (N_8798,N_3406,N_4674);
nand U8799 (N_8799,N_5390,N_5499);
or U8800 (N_8800,N_5676,N_5092);
and U8801 (N_8801,N_4670,N_5169);
xor U8802 (N_8802,N_4157,N_4651);
or U8803 (N_8803,N_4723,N_5299);
nor U8804 (N_8804,N_3757,N_3001);
or U8805 (N_8805,N_4525,N_5351);
or U8806 (N_8806,N_4236,N_3362);
nor U8807 (N_8807,N_4806,N_3004);
and U8808 (N_8808,N_3671,N_5842);
nor U8809 (N_8809,N_4025,N_3579);
nor U8810 (N_8810,N_4154,N_4951);
nand U8811 (N_8811,N_4560,N_3112);
or U8812 (N_8812,N_5926,N_5461);
and U8813 (N_8813,N_5169,N_3851);
and U8814 (N_8814,N_5599,N_4547);
nor U8815 (N_8815,N_3728,N_5181);
nand U8816 (N_8816,N_5944,N_3799);
nand U8817 (N_8817,N_3580,N_3893);
nor U8818 (N_8818,N_5796,N_3321);
or U8819 (N_8819,N_3722,N_5460);
nand U8820 (N_8820,N_5623,N_5526);
or U8821 (N_8821,N_4135,N_3328);
xnor U8822 (N_8822,N_5856,N_3688);
and U8823 (N_8823,N_5858,N_3115);
xor U8824 (N_8824,N_4173,N_4545);
xnor U8825 (N_8825,N_4663,N_4841);
nor U8826 (N_8826,N_4317,N_3977);
or U8827 (N_8827,N_3654,N_5010);
nor U8828 (N_8828,N_3593,N_5649);
xor U8829 (N_8829,N_3092,N_3674);
or U8830 (N_8830,N_4954,N_4302);
xor U8831 (N_8831,N_4740,N_5715);
and U8832 (N_8832,N_4729,N_4312);
nor U8833 (N_8833,N_4028,N_4510);
and U8834 (N_8834,N_4299,N_3082);
and U8835 (N_8835,N_3245,N_5947);
nand U8836 (N_8836,N_4210,N_4984);
xnor U8837 (N_8837,N_5815,N_3761);
xnor U8838 (N_8838,N_4466,N_3427);
nand U8839 (N_8839,N_5657,N_5621);
xnor U8840 (N_8840,N_3067,N_5034);
nand U8841 (N_8841,N_4610,N_5263);
and U8842 (N_8842,N_5754,N_5307);
and U8843 (N_8843,N_3100,N_3576);
or U8844 (N_8844,N_3720,N_4721);
xnor U8845 (N_8845,N_3758,N_4211);
and U8846 (N_8846,N_4890,N_3573);
nand U8847 (N_8847,N_4943,N_3061);
or U8848 (N_8848,N_3557,N_5606);
nand U8849 (N_8849,N_4504,N_5408);
and U8850 (N_8850,N_4015,N_3701);
xnor U8851 (N_8851,N_5478,N_3021);
nand U8852 (N_8852,N_5736,N_5959);
nand U8853 (N_8853,N_3819,N_5610);
or U8854 (N_8854,N_3351,N_4667);
or U8855 (N_8855,N_5602,N_4743);
and U8856 (N_8856,N_3821,N_3052);
nor U8857 (N_8857,N_4549,N_5658);
xnor U8858 (N_8858,N_5113,N_5259);
and U8859 (N_8859,N_4447,N_4838);
nor U8860 (N_8860,N_4791,N_4795);
nor U8861 (N_8861,N_3445,N_4423);
and U8862 (N_8862,N_5705,N_5959);
nor U8863 (N_8863,N_4410,N_3441);
nor U8864 (N_8864,N_3234,N_3339);
or U8865 (N_8865,N_5541,N_4929);
and U8866 (N_8866,N_4800,N_5347);
or U8867 (N_8867,N_3704,N_3248);
or U8868 (N_8868,N_4231,N_4092);
and U8869 (N_8869,N_4834,N_4598);
nor U8870 (N_8870,N_5489,N_4436);
xor U8871 (N_8871,N_4668,N_4726);
nor U8872 (N_8872,N_4102,N_4996);
nor U8873 (N_8873,N_5224,N_5951);
or U8874 (N_8874,N_5727,N_5971);
or U8875 (N_8875,N_4691,N_3455);
nor U8876 (N_8876,N_5352,N_5192);
nand U8877 (N_8877,N_4755,N_5091);
xnor U8878 (N_8878,N_5397,N_4448);
or U8879 (N_8879,N_5759,N_4529);
xnor U8880 (N_8880,N_5562,N_5001);
nor U8881 (N_8881,N_3298,N_3753);
and U8882 (N_8882,N_3286,N_5264);
nor U8883 (N_8883,N_5769,N_5222);
or U8884 (N_8884,N_5760,N_4130);
nor U8885 (N_8885,N_4960,N_4437);
or U8886 (N_8886,N_3434,N_4463);
and U8887 (N_8887,N_5165,N_3422);
nand U8888 (N_8888,N_5060,N_3518);
and U8889 (N_8889,N_5907,N_4266);
nand U8890 (N_8890,N_3458,N_3569);
or U8891 (N_8891,N_3194,N_5715);
xor U8892 (N_8892,N_4044,N_5540);
nand U8893 (N_8893,N_4877,N_3493);
nor U8894 (N_8894,N_3966,N_3180);
or U8895 (N_8895,N_3403,N_4761);
and U8896 (N_8896,N_5192,N_4094);
nor U8897 (N_8897,N_4372,N_4291);
xor U8898 (N_8898,N_4345,N_5559);
and U8899 (N_8899,N_5717,N_5889);
and U8900 (N_8900,N_4772,N_5342);
and U8901 (N_8901,N_5529,N_4570);
nand U8902 (N_8902,N_4267,N_5976);
xnor U8903 (N_8903,N_3041,N_5922);
nand U8904 (N_8904,N_3433,N_4369);
or U8905 (N_8905,N_3461,N_4089);
and U8906 (N_8906,N_5220,N_5326);
xor U8907 (N_8907,N_4438,N_3851);
nand U8908 (N_8908,N_4872,N_4599);
or U8909 (N_8909,N_5759,N_4944);
or U8910 (N_8910,N_3880,N_4847);
xnor U8911 (N_8911,N_5016,N_3156);
xor U8912 (N_8912,N_5258,N_4856);
nor U8913 (N_8913,N_5884,N_3141);
xnor U8914 (N_8914,N_5644,N_4784);
nor U8915 (N_8915,N_5437,N_5009);
nand U8916 (N_8916,N_5642,N_4440);
and U8917 (N_8917,N_4324,N_3049);
xnor U8918 (N_8918,N_4507,N_5437);
xor U8919 (N_8919,N_4497,N_5076);
or U8920 (N_8920,N_3741,N_3798);
or U8921 (N_8921,N_4786,N_5162);
nor U8922 (N_8922,N_3560,N_4358);
and U8923 (N_8923,N_3420,N_5240);
xor U8924 (N_8924,N_5451,N_4743);
xnor U8925 (N_8925,N_4537,N_5838);
or U8926 (N_8926,N_3792,N_3761);
and U8927 (N_8927,N_5893,N_4509);
xor U8928 (N_8928,N_3609,N_5669);
and U8929 (N_8929,N_5160,N_4330);
nand U8930 (N_8930,N_4911,N_5887);
nor U8931 (N_8931,N_4066,N_3702);
nor U8932 (N_8932,N_3692,N_3779);
or U8933 (N_8933,N_5862,N_3668);
nand U8934 (N_8934,N_4677,N_5562);
xnor U8935 (N_8935,N_3055,N_3353);
and U8936 (N_8936,N_5969,N_4174);
and U8937 (N_8937,N_4825,N_5913);
nor U8938 (N_8938,N_4058,N_3529);
nor U8939 (N_8939,N_4209,N_5053);
nor U8940 (N_8940,N_3805,N_3197);
and U8941 (N_8941,N_4124,N_3948);
nand U8942 (N_8942,N_5819,N_5958);
and U8943 (N_8943,N_4152,N_4010);
nor U8944 (N_8944,N_4331,N_5152);
nor U8945 (N_8945,N_3520,N_3758);
or U8946 (N_8946,N_4481,N_4056);
or U8947 (N_8947,N_5934,N_4290);
xor U8948 (N_8948,N_5126,N_3154);
nand U8949 (N_8949,N_3108,N_4147);
or U8950 (N_8950,N_4024,N_4792);
and U8951 (N_8951,N_5527,N_4482);
or U8952 (N_8952,N_5877,N_5038);
or U8953 (N_8953,N_3044,N_3210);
and U8954 (N_8954,N_4526,N_4775);
xnor U8955 (N_8955,N_3011,N_3839);
xor U8956 (N_8956,N_4007,N_5367);
and U8957 (N_8957,N_5665,N_4109);
and U8958 (N_8958,N_3934,N_5275);
nand U8959 (N_8959,N_3205,N_3834);
nor U8960 (N_8960,N_4348,N_3842);
nand U8961 (N_8961,N_5319,N_4434);
nor U8962 (N_8962,N_4338,N_3105);
nand U8963 (N_8963,N_5704,N_4218);
nor U8964 (N_8964,N_3641,N_3317);
nand U8965 (N_8965,N_3114,N_4341);
and U8966 (N_8966,N_3350,N_4674);
and U8967 (N_8967,N_3105,N_4622);
nand U8968 (N_8968,N_4565,N_4508);
or U8969 (N_8969,N_4392,N_4951);
nand U8970 (N_8970,N_4961,N_3214);
xor U8971 (N_8971,N_3685,N_5236);
nand U8972 (N_8972,N_4628,N_3499);
or U8973 (N_8973,N_4565,N_4839);
nor U8974 (N_8974,N_5667,N_3254);
and U8975 (N_8975,N_5687,N_5283);
nor U8976 (N_8976,N_5050,N_4244);
xor U8977 (N_8977,N_5713,N_4219);
nor U8978 (N_8978,N_4885,N_5747);
nand U8979 (N_8979,N_5729,N_5599);
xnor U8980 (N_8980,N_5557,N_5135);
or U8981 (N_8981,N_3091,N_4861);
nand U8982 (N_8982,N_3534,N_4262);
or U8983 (N_8983,N_5099,N_5544);
or U8984 (N_8984,N_3628,N_3706);
and U8985 (N_8985,N_3837,N_4699);
nor U8986 (N_8986,N_3799,N_4985);
nand U8987 (N_8987,N_4376,N_4220);
nand U8988 (N_8988,N_5515,N_4199);
nand U8989 (N_8989,N_4106,N_3553);
xor U8990 (N_8990,N_3327,N_5868);
xnor U8991 (N_8991,N_4528,N_4848);
nand U8992 (N_8992,N_5242,N_5740);
nor U8993 (N_8993,N_3152,N_3217);
xnor U8994 (N_8994,N_4394,N_4964);
or U8995 (N_8995,N_3165,N_5868);
xnor U8996 (N_8996,N_5351,N_3329);
xor U8997 (N_8997,N_3900,N_4739);
and U8998 (N_8998,N_3591,N_3204);
or U8999 (N_8999,N_5262,N_4733);
nand U9000 (N_9000,N_7784,N_7424);
nand U9001 (N_9001,N_6448,N_6779);
or U9002 (N_9002,N_8029,N_7243);
and U9003 (N_9003,N_7052,N_6966);
or U9004 (N_9004,N_7919,N_6756);
or U9005 (N_9005,N_6899,N_8759);
nor U9006 (N_9006,N_7217,N_8260);
and U9007 (N_9007,N_8669,N_7227);
xnor U9008 (N_9008,N_7530,N_7594);
nand U9009 (N_9009,N_6598,N_8082);
nor U9010 (N_9010,N_6040,N_8439);
nor U9011 (N_9011,N_6208,N_7178);
nand U9012 (N_9012,N_6695,N_7763);
nand U9013 (N_9013,N_6774,N_8915);
nor U9014 (N_9014,N_8844,N_8597);
nor U9015 (N_9015,N_8797,N_7023);
nand U9016 (N_9016,N_7629,N_7200);
xor U9017 (N_9017,N_7191,N_6801);
xor U9018 (N_9018,N_8688,N_6029);
or U9019 (N_9019,N_8776,N_6506);
or U9020 (N_9020,N_7244,N_8087);
nand U9021 (N_9021,N_6084,N_8754);
and U9022 (N_9022,N_7418,N_6873);
or U9023 (N_9023,N_7878,N_6898);
nand U9024 (N_9024,N_8244,N_8518);
xor U9025 (N_9025,N_6343,N_6999);
xnor U9026 (N_9026,N_6590,N_7745);
and U9027 (N_9027,N_6935,N_7376);
and U9028 (N_9028,N_8622,N_6349);
or U9029 (N_9029,N_6907,N_7326);
nor U9030 (N_9030,N_7478,N_7860);
and U9031 (N_9031,N_8895,N_6411);
nand U9032 (N_9032,N_6551,N_6422);
xnor U9033 (N_9033,N_7938,N_6521);
or U9034 (N_9034,N_8255,N_8629);
and U9035 (N_9035,N_8861,N_6215);
or U9036 (N_9036,N_7181,N_7519);
xor U9037 (N_9037,N_6891,N_8530);
nand U9038 (N_9038,N_8151,N_8001);
xor U9039 (N_9039,N_8616,N_7676);
nand U9040 (N_9040,N_7098,N_7902);
or U9041 (N_9041,N_6330,N_8654);
or U9042 (N_9042,N_7157,N_8003);
or U9043 (N_9043,N_7333,N_7672);
or U9044 (N_9044,N_6620,N_6870);
xor U9045 (N_9045,N_8474,N_7666);
xnor U9046 (N_9046,N_8345,N_6185);
nor U9047 (N_9047,N_8467,N_7287);
xor U9048 (N_9048,N_7348,N_6415);
nor U9049 (N_9049,N_6998,N_6202);
xor U9050 (N_9050,N_6361,N_8750);
or U9051 (N_9051,N_8918,N_7887);
and U9052 (N_9052,N_6304,N_6842);
xnor U9053 (N_9053,N_7083,N_8777);
nor U9054 (N_9054,N_8563,N_8090);
or U9055 (N_9055,N_6477,N_8224);
xor U9056 (N_9056,N_7759,N_7803);
nand U9057 (N_9057,N_7789,N_8453);
nand U9058 (N_9058,N_6922,N_8377);
xor U9059 (N_9059,N_8832,N_7673);
or U9060 (N_9060,N_8753,N_8781);
nand U9061 (N_9061,N_7103,N_8922);
and U9062 (N_9062,N_8725,N_7468);
xnor U9063 (N_9063,N_8322,N_8778);
or U9064 (N_9064,N_7029,N_7204);
or U9065 (N_9065,N_8280,N_8136);
nor U9066 (N_9066,N_7319,N_6570);
or U9067 (N_9067,N_7026,N_7202);
or U9068 (N_9068,N_6409,N_7393);
and U9069 (N_9069,N_8748,N_6048);
and U9070 (N_9070,N_8574,N_6589);
xnor U9071 (N_9071,N_7558,N_8408);
xnor U9072 (N_9072,N_6032,N_6007);
xnor U9073 (N_9073,N_6693,N_8925);
and U9074 (N_9074,N_7601,N_7667);
or U9075 (N_9075,N_8153,N_6802);
xor U9076 (N_9076,N_8806,N_7039);
and U9077 (N_9077,N_6763,N_8486);
nor U9078 (N_9078,N_6168,N_7271);
xor U9079 (N_9079,N_6161,N_6716);
and U9080 (N_9080,N_8773,N_8263);
xor U9081 (N_9081,N_8594,N_8638);
and U9082 (N_9082,N_6086,N_7552);
xor U9083 (N_9083,N_8580,N_7131);
nand U9084 (N_9084,N_8653,N_8994);
or U9085 (N_9085,N_6910,N_8975);
and U9086 (N_9086,N_7937,N_7008);
or U9087 (N_9087,N_7410,N_8651);
or U9088 (N_9088,N_8064,N_6162);
xor U9089 (N_9089,N_8902,N_6925);
and U9090 (N_9090,N_7416,N_6386);
nand U9091 (N_9091,N_6450,N_8191);
and U9092 (N_9092,N_8125,N_8936);
nand U9093 (N_9093,N_7078,N_6368);
nand U9094 (N_9094,N_8145,N_7034);
and U9095 (N_9095,N_8046,N_7733);
xnor U9096 (N_9096,N_6252,N_8928);
nand U9097 (N_9097,N_8893,N_8610);
nand U9098 (N_9098,N_8685,N_6292);
nand U9099 (N_9099,N_8156,N_8342);
or U9100 (N_9100,N_6788,N_6517);
or U9101 (N_9101,N_6243,N_7510);
xnor U9102 (N_9102,N_7305,N_7934);
nand U9103 (N_9103,N_6761,N_6491);
xor U9104 (N_9104,N_7038,N_6860);
xnor U9105 (N_9105,N_6698,N_8202);
nand U9106 (N_9106,N_8394,N_7250);
nor U9107 (N_9107,N_8572,N_8337);
or U9108 (N_9108,N_8398,N_6358);
xnor U9109 (N_9109,N_8127,N_8171);
nand U9110 (N_9110,N_7105,N_8708);
nand U9111 (N_9111,N_6047,N_6204);
nand U9112 (N_9112,N_6970,N_6837);
and U9113 (N_9113,N_7084,N_7089);
or U9114 (N_9114,N_6840,N_6535);
nand U9115 (N_9115,N_6081,N_6263);
nand U9116 (N_9116,N_8935,N_7586);
and U9117 (N_9117,N_8147,N_8901);
or U9118 (N_9118,N_6225,N_8547);
or U9119 (N_9119,N_7972,N_6518);
nand U9120 (N_9120,N_8746,N_7927);
nor U9121 (N_9121,N_8416,N_8025);
nand U9122 (N_9122,N_8236,N_7422);
or U9123 (N_9123,N_6890,N_8927);
xor U9124 (N_9124,N_6692,N_8076);
nand U9125 (N_9125,N_6500,N_7109);
nand U9126 (N_9126,N_7388,N_6128);
or U9127 (N_9127,N_7423,N_8612);
nor U9128 (N_9128,N_6496,N_6606);
nor U9129 (N_9129,N_8070,N_8630);
xor U9130 (N_9130,N_8045,N_8387);
or U9131 (N_9131,N_7566,N_6638);
nor U9132 (N_9132,N_8815,N_7709);
and U9133 (N_9133,N_6834,N_8048);
and U9134 (N_9134,N_6908,N_8189);
xnor U9135 (N_9135,N_7020,N_8799);
and U9136 (N_9136,N_7133,N_6015);
or U9137 (N_9137,N_7143,N_7992);
or U9138 (N_9138,N_8253,N_7500);
nor U9139 (N_9139,N_8699,N_6089);
or U9140 (N_9140,N_8016,N_7979);
nand U9141 (N_9141,N_8309,N_7520);
and U9142 (N_9142,N_6223,N_7978);
nand U9143 (N_9143,N_7785,N_8193);
nand U9144 (N_9144,N_8455,N_7627);
or U9145 (N_9145,N_6236,N_7555);
nand U9146 (N_9146,N_8917,N_6315);
or U9147 (N_9147,N_6845,N_7296);
nor U9148 (N_9148,N_6511,N_8664);
nor U9149 (N_9149,N_8535,N_8524);
xor U9150 (N_9150,N_6614,N_6778);
xnor U9151 (N_9151,N_6053,N_8110);
nand U9152 (N_9152,N_7955,N_8246);
nand U9153 (N_9153,N_6193,N_8174);
xnor U9154 (N_9154,N_7009,N_7342);
xor U9155 (N_9155,N_7230,N_8564);
nand U9156 (N_9156,N_7998,N_6163);
xnor U9157 (N_9157,N_6197,N_7572);
and U9158 (N_9158,N_8100,N_8912);
and U9159 (N_9159,N_7757,N_8143);
nor U9160 (N_9160,N_8876,N_8307);
xor U9161 (N_9161,N_8586,N_8198);
and U9162 (N_9162,N_7889,N_8814);
xor U9163 (N_9163,N_8060,N_6189);
nor U9164 (N_9164,N_7075,N_6749);
or U9165 (N_9165,N_6284,N_8468);
xor U9166 (N_9166,N_6699,N_8625);
and U9167 (N_9167,N_8479,N_6227);
xnor U9168 (N_9168,N_8656,N_6760);
nor U9169 (N_9169,N_7918,N_8865);
nor U9170 (N_9170,N_7716,N_7496);
xnor U9171 (N_9171,N_8511,N_7363);
nand U9172 (N_9172,N_7177,N_7433);
xor U9173 (N_9173,N_6482,N_8424);
nand U9174 (N_9174,N_7769,N_7207);
or U9175 (N_9175,N_6540,N_8554);
xor U9176 (N_9176,N_8437,N_7462);
nand U9177 (N_9177,N_6920,N_7474);
or U9178 (N_9178,N_6099,N_7808);
xor U9179 (N_9179,N_8691,N_8148);
nor U9180 (N_9180,N_8724,N_6525);
and U9181 (N_9181,N_8353,N_8386);
and U9182 (N_9182,N_6577,N_8780);
or U9183 (N_9183,N_8744,N_6444);
and U9184 (N_9184,N_6339,N_6293);
nand U9185 (N_9185,N_6461,N_7869);
and U9186 (N_9186,N_8376,N_7688);
nand U9187 (N_9187,N_8497,N_6078);
or U9188 (N_9188,N_6268,N_7206);
or U9189 (N_9189,N_7260,N_8954);
and U9190 (N_9190,N_6861,N_7527);
or U9191 (N_9191,N_6403,N_6667);
and U9192 (N_9192,N_8138,N_6855);
nor U9193 (N_9193,N_8545,N_8661);
and U9194 (N_9194,N_8821,N_7336);
nor U9195 (N_9195,N_7814,N_7324);
xnor U9196 (N_9196,N_7389,N_7349);
xnor U9197 (N_9197,N_7628,N_6331);
xor U9198 (N_9198,N_8624,N_8720);
or U9199 (N_9199,N_7135,N_6217);
nand U9200 (N_9200,N_6465,N_8932);
or U9201 (N_9201,N_6153,N_6641);
nand U9202 (N_9202,N_6270,N_8388);
or U9203 (N_9203,N_6932,N_6811);
xor U9204 (N_9204,N_6827,N_7382);
xnor U9205 (N_9205,N_8812,N_8719);
nor U9206 (N_9206,N_7471,N_6248);
xor U9207 (N_9207,N_7635,N_8733);
or U9208 (N_9208,N_7440,N_7561);
nand U9209 (N_9209,N_7925,N_6136);
nor U9210 (N_9210,N_8252,N_8351);
nor U9211 (N_9211,N_8571,N_7021);
nor U9212 (N_9212,N_7871,N_6279);
and U9213 (N_9213,N_8772,N_7354);
nor U9214 (N_9214,N_7697,N_6923);
or U9215 (N_9215,N_6785,N_6792);
nand U9216 (N_9216,N_7128,N_7618);
or U9217 (N_9217,N_8953,N_6637);
xor U9218 (N_9218,N_8347,N_8181);
and U9219 (N_9219,N_8751,N_7237);
nor U9220 (N_9220,N_6581,N_8283);
or U9221 (N_9221,N_7653,N_6242);
xnor U9222 (N_9222,N_6328,N_6245);
nand U9223 (N_9223,N_8568,N_6554);
nor U9224 (N_9224,N_7855,N_6362);
xnor U9225 (N_9225,N_6991,N_6406);
or U9226 (N_9226,N_7674,N_8331);
xor U9227 (N_9227,N_7080,N_6211);
nand U9228 (N_9228,N_6904,N_8695);
xor U9229 (N_9229,N_8275,N_7507);
nand U9230 (N_9230,N_6574,N_7812);
nor U9231 (N_9231,N_6902,N_6940);
xor U9232 (N_9232,N_7345,N_7239);
nor U9233 (N_9233,N_7715,N_6066);
or U9234 (N_9234,N_7751,N_6360);
and U9235 (N_9235,N_7266,N_6296);
nand U9236 (N_9236,N_8934,N_6661);
nor U9237 (N_9237,N_7100,N_8997);
and U9238 (N_9238,N_7509,N_6959);
or U9239 (N_9239,N_6416,N_8643);
nand U9240 (N_9240,N_7257,N_7567);
nor U9241 (N_9241,N_6659,N_7587);
nor U9242 (N_9242,N_8949,N_7735);
or U9243 (N_9243,N_6808,N_8475);
and U9244 (N_9244,N_6050,N_6370);
nand U9245 (N_9245,N_8820,N_7141);
nor U9246 (N_9246,N_7600,N_6192);
or U9247 (N_9247,N_8621,N_7174);
nor U9248 (N_9248,N_6673,N_8277);
nand U9249 (N_9249,N_7051,N_6658);
nand U9250 (N_9250,N_7828,N_7891);
xnor U9251 (N_9251,N_8598,N_6373);
or U9252 (N_9252,N_7799,N_8047);
xor U9253 (N_9253,N_8856,N_6196);
xnor U9254 (N_9254,N_7946,N_6240);
and U9255 (N_9255,N_6074,N_7280);
or U9256 (N_9256,N_8282,N_6526);
nor U9257 (N_9257,N_6390,N_7463);
xnor U9258 (N_9258,N_7439,N_8200);
xor U9259 (N_9259,N_8701,N_7291);
nand U9260 (N_9260,N_8271,N_7330);
or U9261 (N_9261,N_8058,N_7107);
or U9262 (N_9262,N_8817,N_6736);
and U9263 (N_9263,N_6076,N_6557);
and U9264 (N_9264,N_7169,N_6072);
nor U9265 (N_9265,N_6900,N_7398);
nand U9266 (N_9266,N_6119,N_8370);
nor U9267 (N_9267,N_8992,N_8159);
or U9268 (N_9268,N_6847,N_6665);
or U9269 (N_9269,N_6713,N_8019);
nand U9270 (N_9270,N_7882,N_6775);
nor U9271 (N_9271,N_8175,N_8783);
nand U9272 (N_9272,N_6501,N_6068);
xor U9273 (N_9273,N_7351,N_8752);
xnor U9274 (N_9274,N_7778,N_7525);
and U9275 (N_9275,N_8531,N_8526);
and U9276 (N_9276,N_6804,N_8577);
nor U9277 (N_9277,N_8482,N_7888);
xor U9278 (N_9278,N_6093,N_6660);
or U9279 (N_9279,N_7866,N_7685);
nand U9280 (N_9280,N_8581,N_6594);
nor U9281 (N_9281,N_7166,N_8466);
or U9282 (N_9282,N_7355,N_7328);
xnor U9283 (N_9283,N_8608,N_6332);
xnor U9284 (N_9284,N_8118,N_6744);
and U9285 (N_9285,N_7249,N_8083);
nand U9286 (N_9286,N_7314,N_8051);
nand U9287 (N_9287,N_8272,N_8465);
nand U9288 (N_9288,N_7153,N_8167);
xnor U9289 (N_9289,N_7677,N_8767);
or U9290 (N_9290,N_6051,N_8242);
or U9291 (N_9291,N_6680,N_6401);
nand U9292 (N_9292,N_8484,N_6681);
and U9293 (N_9293,N_6479,N_7288);
nand U9294 (N_9294,N_6138,N_6486);
nor U9295 (N_9295,N_6783,N_7449);
xnor U9296 (N_9296,N_8114,N_7329);
nor U9297 (N_9297,N_6466,N_8418);
nor U9298 (N_9298,N_6278,N_7989);
nor U9299 (N_9299,N_8160,N_6283);
or U9300 (N_9300,N_6709,N_8626);
nor U9301 (N_9301,N_7655,N_6038);
and U9302 (N_9302,N_7472,N_6033);
nor U9303 (N_9303,N_7589,N_8472);
xnor U9304 (N_9304,N_7861,N_8061);
nor U9305 (N_9305,N_6558,N_8130);
nor U9306 (N_9306,N_7366,N_8292);
and U9307 (N_9307,N_6275,N_8066);
nand U9308 (N_9308,N_7242,N_7603);
or U9309 (N_9309,N_7428,N_8600);
or U9310 (N_9310,N_8808,N_7403);
and U9311 (N_9311,N_7926,N_8254);
nor U9312 (N_9312,N_7438,N_7201);
or U9313 (N_9313,N_8596,N_6190);
xor U9314 (N_9314,N_8631,N_8328);
nor U9315 (N_9315,N_7779,N_8393);
nor U9316 (N_9316,N_8205,N_7486);
or U9317 (N_9317,N_6114,N_7359);
nand U9318 (N_9318,N_8286,N_6451);
nand U9319 (N_9319,N_8412,N_8150);
and U9320 (N_9320,N_8105,N_7695);
nor U9321 (N_9321,N_6126,N_7796);
nand U9322 (N_9322,N_6226,N_7450);
nand U9323 (N_9323,N_7172,N_8721);
nor U9324 (N_9324,N_6568,N_8022);
xor U9325 (N_9325,N_6460,N_8305);
nor U9326 (N_9326,N_8062,N_8711);
nor U9327 (N_9327,N_6648,N_8320);
nand U9328 (N_9328,N_8509,N_8988);
nand U9329 (N_9329,N_7331,N_7114);
or U9330 (N_9330,N_6421,N_6538);
nor U9331 (N_9331,N_6382,N_6941);
nand U9332 (N_9332,N_8903,N_6286);
and U9333 (N_9333,N_6791,N_6198);
nor U9334 (N_9334,N_8591,N_6928);
nor U9335 (N_9335,N_7737,N_6952);
xnor U9336 (N_9336,N_8566,N_6235);
and U9337 (N_9337,N_7731,N_7112);
nand U9338 (N_9338,N_7126,N_7658);
xnor U9339 (N_9339,N_7203,N_8015);
and U9340 (N_9340,N_7660,N_8553);
nand U9341 (N_9341,N_8262,N_8500);
or U9342 (N_9342,N_8976,N_6462);
nand U9343 (N_9343,N_8888,N_8120);
nor U9344 (N_9344,N_8668,N_6174);
or U9345 (N_9345,N_6201,N_7059);
xnor U9346 (N_9346,N_7180,N_8040);
xnor U9347 (N_9347,N_8335,N_7150);
or U9348 (N_9348,N_8537,N_8454);
nand U9349 (N_9349,N_7602,N_8505);
nor U9350 (N_9350,N_7831,N_6957);
xnor U9351 (N_9351,N_8312,N_8380);
nand U9352 (N_9352,N_8447,N_8095);
or U9353 (N_9353,N_7088,N_6915);
xor U9354 (N_9354,N_8214,N_6110);
and U9355 (N_9355,N_6261,N_8306);
nor U9356 (N_9356,N_8715,N_8117);
or U9357 (N_9357,N_7301,N_8161);
nor U9358 (N_9358,N_8540,N_6320);
xor U9359 (N_9359,N_8186,N_6397);
or U9360 (N_9360,N_7003,N_8614);
nor U9361 (N_9361,N_8055,N_6177);
nor U9362 (N_9362,N_8548,N_6008);
nor U9363 (N_9363,N_8887,N_7581);
or U9364 (N_9364,N_7962,N_8444);
or U9365 (N_9365,N_6572,N_8169);
nor U9366 (N_9366,N_7455,N_8080);
xnor U9367 (N_9367,N_7453,N_8067);
nand U9368 (N_9368,N_8894,N_7948);
or U9369 (N_9369,N_8765,N_8667);
and U9370 (N_9370,N_8704,N_6063);
nor U9371 (N_9371,N_6951,N_7770);
xnor U9372 (N_9372,N_8247,N_8421);
and U9373 (N_9373,N_6575,N_6524);
nor U9374 (N_9374,N_7849,N_6569);
and U9375 (N_9375,N_8199,N_7797);
nand U9376 (N_9376,N_6186,N_8538);
and U9377 (N_9377,N_6478,N_7848);
xor U9378 (N_9378,N_6254,N_6670);
nand U9379 (N_9379,N_8965,N_6702);
nand U9380 (N_9380,N_8536,N_6143);
or U9381 (N_9381,N_7536,N_8793);
nor U9382 (N_9382,N_8883,N_8227);
nand U9383 (N_9383,N_8495,N_7494);
nor U9384 (N_9384,N_6653,N_8796);
nand U9385 (N_9385,N_8483,N_8384);
nor U9386 (N_9386,N_6183,N_8492);
xor U9387 (N_9387,N_6821,N_6893);
xor U9388 (N_9388,N_7646,N_6430);
and U9389 (N_9389,N_7903,N_7727);
nor U9390 (N_9390,N_8769,N_8020);
nor U9391 (N_9391,N_7286,N_7215);
and U9392 (N_9392,N_8017,N_8038);
nor U9393 (N_9393,N_8411,N_7742);
nand U9394 (N_9394,N_6833,N_7338);
nand U9395 (N_9395,N_8768,N_6758);
or U9396 (N_9396,N_8462,N_7850);
xnor U9397 (N_9397,N_8502,N_7829);
nand U9398 (N_9398,N_7027,N_7661);
or U9399 (N_9399,N_6743,N_8555);
nand U9400 (N_9400,N_8297,N_8897);
nand U9401 (N_9401,N_6355,N_8684);
or U9402 (N_9402,N_7504,N_8809);
or U9403 (N_9403,N_6218,N_7935);
and U9404 (N_9404,N_8670,N_6070);
and U9405 (N_9405,N_7060,N_7617);
nor U9406 (N_9406,N_8542,N_8361);
nand U9407 (N_9407,N_7920,N_7991);
and U9408 (N_9408,N_6171,N_6534);
xnor U9409 (N_9409,N_8420,N_8094);
and U9410 (N_9410,N_6828,N_6629);
and U9411 (N_9411,N_8603,N_7068);
xnor U9412 (N_9412,N_7134,N_7495);
or U9413 (N_9413,N_7095,N_8871);
nand U9414 (N_9414,N_8923,N_8021);
xor U9415 (N_9415,N_6747,N_8556);
and U9416 (N_9416,N_6983,N_8517);
nor U9417 (N_9417,N_7939,N_6541);
and U9418 (N_9418,N_7758,N_7490);
or U9419 (N_9419,N_8513,N_8672);
nand U9420 (N_9420,N_7951,N_8284);
nor U9421 (N_9421,N_8298,N_6080);
nand U9422 (N_9422,N_6381,N_7642);
nand U9423 (N_9423,N_8694,N_7198);
or U9424 (N_9424,N_8033,N_8985);
and U9425 (N_9425,N_8811,N_7999);
xnor U9426 (N_9426,N_6117,N_7631);
nand U9427 (N_9427,N_6604,N_7826);
or U9428 (N_9428,N_6948,N_8978);
and U9429 (N_9429,N_6666,N_8613);
and U9430 (N_9430,N_8329,N_8269);
and U9431 (N_9431,N_7311,N_6872);
and U9432 (N_9432,N_8392,N_8233);
and U9433 (N_9433,N_7452,N_7115);
nand U9434 (N_9434,N_7657,N_6018);
nor U9435 (N_9435,N_7671,N_6230);
or U9436 (N_9436,N_7417,N_7212);
nor U9437 (N_9437,N_8921,N_7563);
nand U9438 (N_9438,N_6393,N_8757);
nand U9439 (N_9439,N_8889,N_6576);
nand U9440 (N_9440,N_6603,N_8627);
and U9441 (N_9441,N_7976,N_6071);
and U9442 (N_9442,N_7821,N_8357);
and U9443 (N_9443,N_7294,N_7235);
or U9444 (N_9444,N_8822,N_6650);
nand U9445 (N_9445,N_6023,N_6389);
nor U9446 (N_9446,N_8792,N_7892);
and U9447 (N_9447,N_6762,N_8012);
and U9448 (N_9448,N_6195,N_7419);
nor U9449 (N_9449,N_6400,N_7526);
xnor U9450 (N_9450,N_7531,N_8259);
or U9451 (N_9451,N_7997,N_7929);
or U9452 (N_9452,N_8770,N_7912);
nor U9453 (N_9453,N_6404,N_6046);
and U9454 (N_9454,N_8360,N_8550);
or U9455 (N_9455,N_7633,N_8606);
nor U9456 (N_9456,N_6733,N_8740);
nand U9457 (N_9457,N_7605,N_6676);
and U9458 (N_9458,N_8862,N_7046);
and U9459 (N_9459,N_6490,N_6618);
xnor U9460 (N_9460,N_6687,N_7016);
xnor U9461 (N_9461,N_7612,N_6327);
nand U9462 (N_9462,N_7216,N_7232);
and U9463 (N_9463,N_7122,N_7273);
and U9464 (N_9464,N_6992,N_6823);
xor U9465 (N_9465,N_7461,N_8683);
nor U9466 (N_9466,N_7401,N_7833);
and U9467 (N_9467,N_7263,N_7847);
nand U9468 (N_9468,N_6892,N_8476);
nand U9469 (N_9469,N_6273,N_6075);
or U9470 (N_9470,N_7322,N_6936);
nand U9471 (N_9471,N_7721,N_8354);
and U9472 (N_9472,N_7876,N_8703);
nor U9473 (N_9473,N_8679,N_7961);
and U9474 (N_9474,N_7321,N_8875);
nor U9475 (N_9475,N_7304,N_7337);
or U9476 (N_9476,N_7844,N_8023);
xor U9477 (N_9477,N_7868,N_7437);
nor U9478 (N_9478,N_7915,N_6799);
nand U9479 (N_9479,N_8558,N_6776);
xnor U9480 (N_9480,N_6357,N_8432);
nand U9481 (N_9481,N_6468,N_7024);
nor U9482 (N_9482,N_7993,N_7011);
nor U9483 (N_9483,N_7923,N_7158);
nor U9484 (N_9484,N_7819,N_6244);
or U9485 (N_9485,N_6635,N_6895);
nor U9486 (N_9486,N_8739,N_8135);
and U9487 (N_9487,N_7664,N_8587);
or U9488 (N_9488,N_7974,N_8009);
nor U9489 (N_9489,N_8706,N_8024);
nand U9490 (N_9490,N_7533,N_7082);
nor U9491 (N_9491,N_8267,N_7541);
and U9492 (N_9492,N_7343,N_8355);
nand U9493 (N_9493,N_7987,N_6825);
xnor U9494 (N_9494,N_8460,N_6566);
or U9495 (N_9495,N_7678,N_8201);
nand U9496 (N_9496,N_6232,N_6850);
and U9497 (N_9497,N_6605,N_7963);
nor U9498 (N_9498,N_6701,N_8313);
xnor U9499 (N_9499,N_7801,N_8841);
xnor U9500 (N_9500,N_6976,N_8842);
or U9501 (N_9501,N_7857,N_6246);
xor U9502 (N_9502,N_6287,N_7700);
and U9503 (N_9503,N_7765,N_7981);
nand U9504 (N_9504,N_8315,N_6337);
xnor U9505 (N_9505,N_7684,N_8162);
or U9506 (N_9506,N_6944,N_7076);
and U9507 (N_9507,N_6154,N_8212);
nand U9508 (N_9508,N_7371,N_8998);
nor U9509 (N_9509,N_6470,N_8219);
nand U9510 (N_9510,N_8787,N_8471);
or U9511 (N_9511,N_7795,N_7741);
xor U9512 (N_9512,N_6544,N_6249);
nor U9513 (N_9513,N_7863,N_7385);
or U9514 (N_9514,N_7632,N_6519);
or U9515 (N_9515,N_8636,N_7782);
nand U9516 (N_9516,N_6250,N_8726);
nand U9517 (N_9517,N_8823,N_7996);
nand U9518 (N_9518,N_8601,N_6786);
and U9519 (N_9519,N_6338,N_6257);
nand U9520 (N_9520,N_7692,N_6447);
or U9521 (N_9521,N_6098,N_7704);
and U9522 (N_9522,N_6067,N_8941);
or U9523 (N_9523,N_8018,N_8031);
and U9524 (N_9524,N_8123,N_7087);
nand U9525 (N_9525,N_6280,N_8419);
and U9526 (N_9526,N_7619,N_6159);
xor U9527 (N_9527,N_8177,N_6132);
and U9528 (N_9528,N_7163,N_7245);
or U9529 (N_9529,N_8266,N_7284);
nor U9530 (N_9530,N_6259,N_8137);
or U9531 (N_9531,N_6927,N_7448);
and U9532 (N_9532,N_7813,N_7256);
and U9533 (N_9533,N_6815,N_8011);
nand U9534 (N_9534,N_6251,N_7442);
nand U9535 (N_9535,N_7985,N_8052);
and U9536 (N_9536,N_6340,N_8857);
or U9537 (N_9537,N_7630,N_6065);
or U9538 (N_9538,N_7580,N_8044);
nor U9539 (N_9539,N_8851,N_6556);
xnor U9540 (N_9540,N_7002,N_7056);
nor U9541 (N_9541,N_7508,N_6025);
nand U9542 (N_9542,N_7295,N_7432);
nor U9543 (N_9543,N_6418,N_8766);
and U9544 (N_9544,N_8878,N_6265);
and U9545 (N_9545,N_6878,N_7641);
nor U9546 (N_9546,N_6125,N_6914);
or U9547 (N_9547,N_6609,N_6272);
nor U9548 (N_9548,N_7063,N_6642);
or U9549 (N_9549,N_6213,N_6711);
or U9550 (N_9550,N_6645,N_8290);
nor U9551 (N_9551,N_8204,N_8413);
and U9552 (N_9552,N_8406,N_6166);
xor U9553 (N_9553,N_7156,N_7576);
nor U9554 (N_9554,N_6313,N_8737);
nand U9555 (N_9555,N_8223,N_7125);
nor U9556 (N_9556,N_8884,N_6934);
nor U9557 (N_9557,N_6303,N_8617);
and U9558 (N_9558,N_6432,N_8506);
nand U9559 (N_9559,N_7261,N_6512);
or U9560 (N_9560,N_6322,N_7521);
xor U9561 (N_9561,N_8002,N_7537);
xor U9562 (N_9562,N_8677,N_6759);
and U9563 (N_9563,N_7044,N_8964);
nor U9564 (N_9564,N_6316,N_7179);
and U9565 (N_9565,N_8734,N_6423);
xor U9566 (N_9566,N_7072,N_7622);
and U9567 (N_9567,N_6777,N_6685);
nand U9568 (N_9568,N_7571,N_6147);
or U9569 (N_9569,N_8732,N_6580);
xnor U9570 (N_9570,N_8341,N_7540);
nand U9571 (N_9571,N_6854,N_7880);
and U9572 (N_9572,N_7189,N_7254);
or U9573 (N_9573,N_6011,N_7830);
or U9574 (N_9574,N_7139,N_8707);
xnor U9575 (N_9575,N_6896,N_7548);
nor U9576 (N_9576,N_7884,N_6090);
or U9577 (N_9577,N_7037,N_8623);
nand U9578 (N_9578,N_8035,N_6818);
nand U9579 (N_9579,N_6822,N_8404);
or U9580 (N_9580,N_8551,N_6180);
xnor U9581 (N_9581,N_7872,N_7396);
and U9582 (N_9582,N_6567,N_6104);
xnor U9583 (N_9583,N_7269,N_7771);
and U9584 (N_9584,N_7551,N_6930);
xor U9585 (N_9585,N_7292,N_7019);
and U9586 (N_9586,N_7917,N_7340);
nand U9587 (N_9587,N_7377,N_8967);
nor U9588 (N_9588,N_8265,N_6030);
nor U9589 (N_9589,N_6591,N_7381);
xor U9590 (N_9590,N_7665,N_6142);
xnor U9591 (N_9591,N_6323,N_6314);
nand U9592 (N_9592,N_8729,N_7092);
and U9593 (N_9593,N_8172,N_6173);
xor U9594 (N_9594,N_7547,N_7744);
nor U9595 (N_9595,N_8325,N_6919);
xnor U9596 (N_9596,N_7047,N_8755);
and U9597 (N_9597,N_6472,N_7289);
nand U9598 (N_9598,N_8069,N_6069);
nor U9599 (N_9599,N_6151,N_8180);
and U9600 (N_9600,N_6341,N_8559);
xnor U9601 (N_9601,N_6938,N_8234);
or U9602 (N_9602,N_7560,N_6954);
or U9603 (N_9603,N_7117,N_8635);
nand U9604 (N_9604,N_8527,N_6000);
nand U9605 (N_9605,N_8168,N_7147);
nor U9606 (N_9606,N_6017,N_6014);
or U9607 (N_9607,N_8727,N_6559);
and U9608 (N_9608,N_8660,N_7429);
or U9609 (N_9609,N_8141,N_6429);
nand U9610 (N_9610,N_6455,N_8804);
xor U9611 (N_9611,N_6597,N_6671);
xnor U9612 (N_9612,N_8079,N_6116);
xor U9613 (N_9613,N_8399,N_8364);
xnor U9614 (N_9614,N_7883,N_7932);
or U9615 (N_9615,N_6282,N_7870);
xnor U9616 (N_9616,N_7588,N_8702);
xnor U9617 (N_9617,N_6674,N_7413);
and U9618 (N_9618,N_7783,N_6144);
nor U9619 (N_9619,N_7030,N_7116);
nor U9620 (N_9620,N_6564,N_8334);
and U9621 (N_9621,N_6683,N_6579);
and U9622 (N_9622,N_6634,N_8774);
xnor U9623 (N_9623,N_6181,N_6961);
and U9624 (N_9624,N_6026,N_8963);
or U9625 (N_9625,N_8593,N_6717);
and U9626 (N_9626,N_8321,N_6347);
and U9627 (N_9627,N_7815,N_8116);
nand U9628 (N_9628,N_8000,N_7318);
xor U9629 (N_9629,N_6200,N_8228);
nand U9630 (N_9630,N_6956,N_8469);
nor U9631 (N_9631,N_7723,N_6057);
xor U9632 (N_9632,N_7766,N_8512);
nor U9633 (N_9633,N_6626,N_8560);
and U9634 (N_9634,N_8775,N_8779);
and U9635 (N_9635,N_7485,N_8640);
xnor U9636 (N_9636,N_8366,N_7190);
xnor U9637 (N_9637,N_8279,N_6990);
nand U9638 (N_9638,N_6929,N_7253);
and U9639 (N_9639,N_8642,N_6120);
and U9640 (N_9640,N_8858,N_7211);
xnor U9641 (N_9641,N_8385,N_8108);
nor U9642 (N_9642,N_7807,N_8389);
nor U9643 (N_9643,N_6109,N_7123);
or U9644 (N_9644,N_7748,N_8911);
nand U9645 (N_9645,N_6724,N_8788);
or U9646 (N_9646,N_6844,N_6346);
nand U9647 (N_9647,N_8245,N_8619);
or U9648 (N_9648,N_7310,N_7077);
or U9649 (N_9649,N_7859,N_7093);
and U9650 (N_9650,N_6981,N_8440);
or U9651 (N_9651,N_6795,N_6152);
or U9652 (N_9652,N_8155,N_8831);
nand U9653 (N_9653,N_7980,N_7055);
nor U9654 (N_9654,N_8872,N_8543);
nand U9655 (N_9655,N_8723,N_6843);
and U9656 (N_9656,N_6984,N_7446);
and U9657 (N_9657,N_7346,N_6971);
and U9658 (N_9658,N_6334,N_7248);
nand U9659 (N_9659,N_7032,N_8712);
xor U9660 (N_9660,N_8864,N_7689);
xor U9661 (N_9661,N_8582,N_8473);
or U9662 (N_9662,N_6742,N_8948);
nand U9663 (N_9663,N_8289,N_6738);
and U9664 (N_9664,N_8583,N_6056);
xor U9665 (N_9665,N_6157,N_8929);
and U9666 (N_9666,N_6751,N_8457);
or U9667 (N_9667,N_7501,N_8544);
xor U9668 (N_9668,N_6483,N_6396);
and U9669 (N_9669,N_8436,N_7793);
nor U9670 (N_9670,N_8824,N_7223);
nor U9671 (N_9671,N_8615,N_6677);
and U9672 (N_9672,N_6329,N_6917);
and U9673 (N_9673,N_8034,N_7543);
and U9674 (N_9674,N_7936,N_7773);
and U9675 (N_9675,N_7928,N_6527);
xor U9676 (N_9676,N_6514,N_8112);
and U9677 (N_9677,N_6371,N_7514);
xor U9678 (N_9678,N_6097,N_7764);
nor U9679 (N_9679,N_6796,N_6228);
xnor U9680 (N_9680,N_6100,N_6820);
xnor U9681 (N_9681,N_7220,N_6729);
xnor U9682 (N_9682,N_6721,N_8216);
xor U9683 (N_9683,N_6459,N_7910);
nand U9684 (N_9684,N_8026,N_8287);
and U9685 (N_9685,N_7822,N_6391);
xor U9686 (N_9686,N_8710,N_6819);
and U9687 (N_9687,N_7730,N_8868);
nand U9688 (N_9688,N_7183,N_8802);
xnor U9689 (N_9689,N_7550,N_7977);
or U9690 (N_9690,N_6877,N_7234);
and U9691 (N_9691,N_7298,N_7140);
nor U9692 (N_9692,N_7491,N_7693);
or U9693 (N_9693,N_6942,N_7197);
or U9694 (N_9694,N_7058,N_6652);
xor U9695 (N_9695,N_7497,N_8059);
nand U9696 (N_9696,N_7644,N_6616);
or U9697 (N_9697,N_6536,N_8299);
xnor U9698 (N_9698,N_8400,N_8485);
or U9699 (N_9699,N_8968,N_7170);
and U9700 (N_9700,N_8532,N_7898);
nor U9701 (N_9701,N_6385,N_6880);
nor U9702 (N_9702,N_8952,N_8987);
or U9703 (N_9703,N_6812,N_8520);
or U9704 (N_9704,N_7669,N_7534);
nor U9705 (N_9705,N_6306,N_7300);
xnor U9706 (N_9706,N_6587,N_8515);
and U9707 (N_9707,N_8316,N_6672);
nand U9708 (N_9708,N_7506,N_6407);
xnor U9709 (N_9709,N_7426,N_6004);
and U9710 (N_9710,N_7908,N_8652);
and U9711 (N_9711,N_7944,N_7431);
xor U9712 (N_9712,N_6867,N_8240);
nor U9713 (N_9713,N_6124,N_6019);
nand U9714 (N_9714,N_7668,N_7590);
and U9715 (N_9715,N_7986,N_8368);
and U9716 (N_9716,N_7516,N_7823);
or U9717 (N_9717,N_8166,N_7277);
xor U9718 (N_9718,N_6746,N_6207);
nor U9719 (N_9719,N_7940,N_8218);
nor U9720 (N_9720,N_6405,N_8369);
nor U9721 (N_9721,N_8434,N_8195);
or U9722 (N_9722,N_7802,N_7682);
nor U9723 (N_9723,N_6542,N_7896);
nor U9724 (N_9724,N_7707,N_8826);
nand U9725 (N_9725,N_8250,N_6498);
nand U9726 (N_9726,N_8647,N_8761);
xnor U9727 (N_9727,N_7853,N_7171);
nor U9728 (N_9728,N_6394,N_6964);
nor U9729 (N_9729,N_6264,N_8196);
or U9730 (N_9730,N_6584,N_8499);
nand U9731 (N_9731,N_6824,N_8170);
and U9732 (N_9732,N_6428,N_8960);
nor U9733 (N_9733,N_6027,N_8036);
xor U9734 (N_9734,N_7137,N_8365);
or U9735 (N_9735,N_7865,N_8588);
and U9736 (N_9736,N_6059,N_6533);
nand U9737 (N_9737,N_7930,N_8914);
or U9738 (N_9738,N_6798,N_8863);
nand U9739 (N_9739,N_8144,N_8281);
nand U9740 (N_9740,N_7054,N_7687);
and U9741 (N_9741,N_8333,N_8790);
nor U9742 (N_9742,N_6255,N_6102);
and U9743 (N_9743,N_6545,N_7625);
and U9744 (N_9744,N_7535,N_6253);
xnor U9745 (N_9745,N_8991,N_8573);
and U9746 (N_9746,N_7774,N_6436);
xnor U9747 (N_9747,N_8939,N_8230);
or U9748 (N_9748,N_6868,N_8931);
nor U9749 (N_9749,N_7767,N_8798);
nor U9750 (N_9750,N_6849,N_7283);
nor U9751 (N_9751,N_6176,N_7621);
nor U9752 (N_9752,N_8005,N_7846);
and U9753 (N_9753,N_6042,N_6456);
or U9754 (N_9754,N_6947,N_6573);
xor U9755 (N_9755,N_8860,N_6494);
or U9756 (N_9756,N_6419,N_6123);
or U9757 (N_9757,N_8698,N_7036);
nand U9758 (N_9758,N_6841,N_7113);
or U9759 (N_9759,N_6060,N_8576);
nand U9760 (N_9760,N_6112,N_6467);
nand U9761 (N_9761,N_8226,N_6184);
nor U9762 (N_9762,N_7460,N_8395);
nor U9763 (N_9763,N_8782,N_7854);
nand U9764 (N_9764,N_6413,N_7593);
nor U9765 (N_9765,N_8977,N_7893);
nand U9766 (N_9766,N_8104,N_8239);
xor U9767 (N_9767,N_7168,N_6203);
or U9768 (N_9768,N_7837,N_7699);
or U9769 (N_9769,N_8211,N_6438);
nor U9770 (N_9770,N_6767,N_7106);
and U9771 (N_9771,N_8742,N_6975);
and U9772 (N_9772,N_7144,N_8944);
and U9773 (N_9773,N_7573,N_7824);
nor U9774 (N_9774,N_6039,N_8187);
and U9775 (N_9775,N_6471,N_8122);
or U9776 (N_9776,N_6473,N_6463);
and U9777 (N_9777,N_7383,N_7221);
nand U9778 (N_9778,N_7862,N_7369);
nor U9779 (N_9779,N_6507,N_7626);
xnor U9780 (N_9780,N_7647,N_6592);
and U9781 (N_9781,N_7971,N_8655);
nor U9782 (N_9782,N_6291,N_6481);
or U9783 (N_9783,N_8716,N_6912);
nor U9784 (N_9784,N_7367,N_8641);
and U9785 (N_9785,N_7643,N_7164);
nor U9786 (N_9786,N_7231,N_8541);
or U9787 (N_9787,N_7913,N_7943);
nand U9788 (N_9788,N_8324,N_8032);
nand U9789 (N_9789,N_7701,N_8892);
or U9790 (N_9790,N_7499,N_8042);
nand U9791 (N_9791,N_6206,N_6838);
and U9792 (N_9792,N_8423,N_7065);
or U9793 (N_9793,N_8973,N_8470);
nand U9794 (N_9794,N_7240,N_7409);
and U9795 (N_9795,N_7279,N_8336);
nand U9796 (N_9796,N_6707,N_6344);
xnor U9797 (N_9797,N_7722,N_7362);
nand U9798 (N_9798,N_8014,N_8043);
or U9799 (N_9799,N_7062,N_8920);
or U9800 (N_9800,N_8238,N_8414);
or U9801 (N_9801,N_6835,N_8899);
nand U9802 (N_9802,N_7564,N_8133);
and U9803 (N_9803,N_7710,N_7005);
xor U9804 (N_9804,N_7464,N_7746);
nor U9805 (N_9805,N_6364,N_8791);
or U9806 (N_9806,N_7392,N_8693);
nand U9807 (N_9807,N_8873,N_8084);
nor U9808 (N_9808,N_7316,N_8605);
nand U9809 (N_9809,N_8176,N_6182);
xor U9810 (N_9810,N_7420,N_7390);
nand U9811 (N_9811,N_7400,N_6882);
nor U9812 (N_9812,N_7804,N_8374);
xnor U9813 (N_9813,N_6644,N_8718);
and U9814 (N_9814,N_6049,N_7467);
nand U9815 (N_9815,N_7155,N_6269);
xor U9816 (N_9816,N_6655,N_7465);
nor U9817 (N_9817,N_7881,N_6599);
xnor U9818 (N_9818,N_8107,N_6205);
nand U9819 (N_9819,N_6810,N_6499);
xor U9820 (N_9820,N_6164,N_7775);
nand U9821 (N_9821,N_7768,N_8681);
nand U9822 (N_9822,N_6475,N_6794);
and U9823 (N_9823,N_8498,N_7755);
nor U9824 (N_9824,N_8663,N_8743);
and U9825 (N_9825,N_8373,N_6022);
nor U9826 (N_9826,N_8958,N_7959);
xor U9827 (N_9827,N_7209,N_7193);
and U9828 (N_9828,N_8085,N_6170);
or U9829 (N_9829,N_6222,N_8229);
nand U9830 (N_9830,N_6866,N_6987);
and U9831 (N_9831,N_6869,N_7415);
or U9832 (N_9832,N_6503,N_8163);
nand U9833 (N_9833,N_7942,N_7965);
and U9834 (N_9834,N_7958,N_8456);
or U9835 (N_9835,N_7982,N_8763);
and U9836 (N_9836,N_8539,N_7726);
and U9837 (N_9837,N_8516,N_8349);
nor U9838 (N_9838,N_8081,N_6135);
and U9839 (N_9839,N_6427,N_7957);
nand U9840 (N_9840,N_7756,N_7205);
nand U9841 (N_9841,N_7832,N_8310);
or U9842 (N_9842,N_8119,N_7378);
nand U9843 (N_9843,N_6814,N_7427);
nand U9844 (N_9844,N_8478,N_6305);
or U9845 (N_9845,N_7358,N_8367);
nor U9846 (N_9846,N_8165,N_8291);
or U9847 (N_9847,N_6712,N_6865);
xnor U9848 (N_9848,N_7391,N_7734);
nand U9849 (N_9849,N_8441,N_6309);
xor U9850 (N_9850,N_6073,N_8907);
nand U9851 (N_9851,N_7405,N_8128);
xnor U9852 (N_9852,N_6354,N_7901);
nor U9853 (N_9853,N_8459,N_7827);
nand U9854 (N_9854,N_7320,N_8496);
xnor U9855 (N_9855,N_7161,N_7553);
or U9856 (N_9856,N_7136,N_7798);
nand U9857 (N_9857,N_7649,N_6764);
xnor U9858 (N_9858,N_6212,N_6613);
xor U9859 (N_9859,N_8338,N_7043);
nor U9860 (N_9860,N_8243,N_6826);
and U9861 (N_9861,N_7258,N_7042);
and U9862 (N_9862,N_7360,N_7399);
and U9863 (N_9863,N_8835,N_7867);
nand U9864 (N_9864,N_7761,N_7386);
nand U9865 (N_9865,N_8662,N_8425);
xor U9866 (N_9866,N_7781,N_6041);
or U9867 (N_9867,N_7545,N_8209);
xnor U9868 (N_9868,N_6884,N_6348);
xnor U9869 (N_9869,N_6994,N_6276);
nor U9870 (N_9870,N_7498,N_8208);
nand U9871 (N_9871,N_7323,N_6950);
or U9872 (N_9872,N_7228,N_6832);
xnor U9873 (N_9873,N_7794,N_6435);
nor U9874 (N_9874,N_7596,N_8371);
xnor U9875 (N_9875,N_7210,N_6563);
and U9876 (N_9876,N_8225,N_7841);
nand U9877 (N_9877,N_6317,N_8945);
xor U9878 (N_9878,N_8959,N_6931);
nor U9879 (N_9879,N_6901,N_8675);
xnor U9880 (N_9880,N_7947,N_6875);
or U9881 (N_9881,N_6752,N_6651);
and U9882 (N_9882,N_8319,N_6377);
nor U9883 (N_9883,N_6973,N_6636);
and U9884 (N_9884,N_8645,N_7578);
nand U9885 (N_9885,N_6342,N_7048);
xor U9886 (N_9886,N_7066,N_7656);
and U9887 (N_9887,N_6887,N_7236);
and U9888 (N_9888,N_7760,N_8595);
or U9889 (N_9889,N_7914,N_8609);
nand U9890 (N_9890,N_6734,N_6565);
nor U9891 (N_9891,N_7638,N_6532);
nand U9892 (N_9892,N_7090,N_6234);
nand U9893 (N_9893,N_8833,N_8332);
xor U9894 (N_9894,N_8213,N_7022);
nand U9895 (N_9895,N_6857,N_8129);
nor U9896 (N_9896,N_6839,N_8891);
nand U9897 (N_9897,N_8477,N_7001);
xnor U9898 (N_9898,N_8628,N_7456);
or U9899 (N_9899,N_8562,N_6537);
xnor U9900 (N_9900,N_6510,N_7028);
or U9901 (N_9901,N_6476,N_8448);
xor U9902 (N_9902,N_8993,N_6816);
or U9903 (N_9903,N_8758,N_7811);
nor U9904 (N_9904,N_7894,N_7108);
nor U9905 (N_9905,N_7636,N_8943);
and U9906 (N_9906,N_8311,N_8190);
or U9907 (N_9907,N_6630,N_6682);
or U9908 (N_9908,N_7546,N_7347);
or U9909 (N_9909,N_6092,N_6622);
nand U9910 (N_9910,N_8152,N_8445);
and U9911 (N_9911,N_8359,N_7609);
nand U9912 (N_9912,N_6686,N_6889);
xnor U9913 (N_9913,N_7208,N_8906);
nor U9914 (N_9914,N_6356,N_6772);
xnor U9915 (N_9915,N_8449,N_7339);
nor U9916 (N_9916,N_7511,N_8962);
and U9917 (N_9917,N_7040,N_7791);
nor U9918 (N_9918,N_7282,N_6924);
or U9919 (N_9919,N_8206,N_7469);
nand U9920 (N_9920,N_7599,N_6150);
or U9921 (N_9921,N_8274,N_8569);
nor U9922 (N_9922,N_8678,N_6719);
nor U9923 (N_9923,N_6392,N_7591);
xnor U9924 (N_9924,N_6684,N_6710);
nor U9925 (N_9925,N_6588,N_7057);
nor U9926 (N_9926,N_7683,N_6530);
nand U9927 (N_9927,N_6548,N_7712);
and U9928 (N_9928,N_6953,N_7950);
xnor U9929 (N_9929,N_7443,N_7035);
nor U9930 (N_9930,N_7079,N_6034);
and U9931 (N_9931,N_7274,N_7949);
nor U9932 (N_9932,N_7489,N_8521);
or U9933 (N_9933,N_7544,N_8845);
or U9934 (N_9934,N_6773,N_6384);
or U9935 (N_9935,N_7152,N_6797);
xor U9936 (N_9936,N_7364,N_8142);
xnor U9937 (N_9937,N_6696,N_8027);
and U9938 (N_9938,N_7916,N_6943);
nor U9939 (N_9939,N_6488,N_6036);
and U9940 (N_9940,N_6420,N_7875);
or U9941 (N_9941,N_6977,N_8528);
or U9942 (N_9942,N_7834,N_8602);
and U9943 (N_9943,N_6372,N_8680);
or U9944 (N_9944,N_6583,N_7696);
nand U9945 (N_9945,N_7121,N_8756);
nand U9946 (N_9946,N_8258,N_6480);
xor U9947 (N_9947,N_7162,N_7505);
nor U9948 (N_9948,N_7718,N_7241);
and U9949 (N_9949,N_8525,N_8146);
nor U9950 (N_9950,N_7278,N_7195);
nor U9951 (N_9951,N_8300,N_7694);
nor U9952 (N_9952,N_7691,N_6088);
nor U9953 (N_9953,N_7213,N_7568);
nor U9954 (N_9954,N_7006,N_7031);
nor U9955 (N_9955,N_6061,N_6469);
and U9956 (N_9956,N_6691,N_8762);
or U9957 (N_9957,N_7639,N_7858);
or U9958 (N_9958,N_7705,N_8288);
xor U9959 (N_9959,N_7435,N_8487);
nand U9960 (N_9960,N_8113,N_8346);
and U9961 (N_9961,N_7724,N_6529);
and U9962 (N_9962,N_6440,N_6631);
nor U9963 (N_9963,N_8950,N_6229);
nand U9964 (N_9964,N_6903,N_6561);
nand U9965 (N_9965,N_6700,N_8529);
xnor U9966 (N_9966,N_7975,N_8947);
nor U9967 (N_9967,N_7387,N_8840);
nand U9968 (N_9968,N_7167,N_8261);
and U9969 (N_9969,N_6546,N_7816);
nand U9970 (N_9970,N_7327,N_6487);
and U9971 (N_9971,N_6694,N_6395);
nor U9972 (N_9972,N_8730,N_6863);
nor U9973 (N_9973,N_7652,N_6290);
and U9974 (N_9974,N_7577,N_8158);
xnor U9975 (N_9975,N_6562,N_7651);
nand U9976 (N_9976,N_6725,N_6096);
xor U9977 (N_9977,N_6945,N_8657);
xor U9978 (N_9978,N_6402,N_8039);
xor U9979 (N_9979,N_8552,N_8403);
or U9980 (N_9980,N_8235,N_6375);
or U9981 (N_9981,N_8401,N_8049);
nand U9982 (N_9982,N_7421,N_8736);
or U9983 (N_9983,N_8430,N_8221);
nand U9984 (N_9984,N_6515,N_7702);
nand U9985 (N_9985,N_6353,N_7787);
or U9986 (N_9986,N_7897,N_6044);
nand U9987 (N_9987,N_6216,N_7013);
nor U9988 (N_9988,N_6439,N_6731);
nand U9989 (N_9989,N_8579,N_6474);
nor U9990 (N_9990,N_8426,N_8904);
xor U9991 (N_9991,N_8886,N_6087);
xor U9992 (N_9992,N_6664,N_8296);
or U9993 (N_9993,N_6426,N_7061);
xnor U9994 (N_9994,N_8686,N_6324);
xor U9995 (N_9995,N_7120,N_6005);
nor U9996 (N_9996,N_7281,N_6781);
nor U9997 (N_9997,N_8154,N_6441);
nand U9998 (N_9998,N_6210,N_8490);
nor U9999 (N_9999,N_7559,N_6351);
or U10000 (N_10000,N_6079,N_7907);
nor U10001 (N_10001,N_6485,N_7720);
nor U10002 (N_10002,N_8124,N_6445);
and U10003 (N_10003,N_6127,N_7595);
xnor U10004 (N_10004,N_8068,N_6058);
nor U10005 (N_10005,N_8905,N_6300);
or U10006 (N_10006,N_6993,N_7941);
or U10007 (N_10007,N_6094,N_6131);
xnor U10008 (N_10008,N_8356,N_7592);
nor U10009 (N_10009,N_6379,N_6663);
xnor U10010 (N_10010,N_7493,N_6160);
nor U10011 (N_10011,N_8909,N_6489);
nand U10012 (N_10012,N_7184,N_6378);
or U10013 (N_10013,N_8362,N_8885);
or U10014 (N_10014,N_6289,N_7457);
and U10015 (N_10015,N_6388,N_6301);
xor U10016 (N_10016,N_6130,N_6043);
xor U10017 (N_10017,N_8164,N_6452);
nor U10018 (N_10018,N_6732,N_8115);
nand U10019 (N_10019,N_7874,N_6607);
and U10020 (N_10020,N_8969,N_8093);
and U10021 (N_10021,N_8741,N_7488);
xor U10022 (N_10022,N_6188,N_6807);
xor U10023 (N_10023,N_7864,N_6016);
or U10024 (N_10024,N_6623,N_7104);
nor U10025 (N_10025,N_6274,N_6704);
nor U10026 (N_10026,N_6874,N_8986);
nand U10027 (N_10027,N_8344,N_8249);
nor U10028 (N_10028,N_7542,N_6539);
or U10029 (N_10029,N_8533,N_6111);
or U10030 (N_10030,N_7290,N_6888);
or U10031 (N_10031,N_8514,N_7297);
nand U10032 (N_10032,N_8828,N_7970);
nor U10033 (N_10033,N_7270,N_7749);
and U10034 (N_10034,N_8464,N_8933);
nand U10035 (N_10035,N_6697,N_7365);
xor U10036 (N_10036,N_6553,N_6013);
or U10037 (N_10037,N_8508,N_6757);
or U10038 (N_10038,N_8381,N_7945);
xnor U10039 (N_10039,N_6852,N_8390);
or U10040 (N_10040,N_6586,N_7332);
or U10041 (N_10041,N_6522,N_7073);
and U10042 (N_10042,N_6224,N_8818);
nor U10043 (N_10043,N_7272,N_7267);
nand U10044 (N_10044,N_8519,N_6982);
nor U10045 (N_10045,N_6003,N_8853);
xnor U10046 (N_10046,N_7306,N_7806);
xor U10047 (N_10047,N_8981,N_7640);
nand U10048 (N_10048,N_6457,N_8604);
xnor U10049 (N_10049,N_7663,N_6103);
nor U10050 (N_10050,N_7554,N_7900);
nor U10051 (N_10051,N_7251,N_7285);
xnor U10052 (N_10052,N_8348,N_8074);
nand U10053 (N_10053,N_8690,N_6939);
or U10054 (N_10054,N_8870,N_8050);
nor U10055 (N_10055,N_7549,N_7477);
nand U10056 (N_10056,N_7430,N_6369);
or U10057 (N_10057,N_8989,N_7611);
and U10058 (N_10058,N_7394,N_7074);
xnor U10059 (N_10059,N_8825,N_6266);
or U10060 (N_10060,N_6689,N_8713);
nor U10061 (N_10061,N_6675,N_8957);
xnor U10062 (N_10062,N_8053,N_6918);
xnor U10063 (N_10063,N_7582,N_7071);
xor U10064 (N_10064,N_6308,N_7247);
xnor U10065 (N_10065,N_6024,N_7659);
or U10066 (N_10066,N_8304,N_8658);
or U10067 (N_10067,N_6454,N_8270);
nor U10068 (N_10068,N_8940,N_6453);
xor U10069 (N_10069,N_8659,N_8273);
nand U10070 (N_10070,N_7800,N_6101);
and U10071 (N_10071,N_8966,N_8409);
or U10072 (N_10072,N_8382,N_8999);
or U10073 (N_10073,N_6417,N_7681);
and U10074 (N_10074,N_8882,N_8407);
xor U10075 (N_10075,N_7686,N_6656);
or U10076 (N_10076,N_8458,N_6158);
or U10077 (N_10077,N_8805,N_6258);
xor U10078 (N_10078,N_6179,N_6167);
nand U10079 (N_10079,N_7185,N_6679);
or U10080 (N_10080,N_8760,N_8910);
xor U10081 (N_10081,N_7522,N_7303);
and U10082 (N_10082,N_8056,N_8007);
nor U10083 (N_10083,N_6513,N_8971);
xor U10084 (N_10084,N_8131,N_8446);
nand U10085 (N_10085,N_8837,N_7650);
and U10086 (N_10086,N_8301,N_6113);
or U10087 (N_10087,N_6805,N_7373);
nand U10088 (N_10088,N_6425,N_6906);
and U10089 (N_10089,N_6446,N_7762);
nor U10090 (N_10090,N_8847,N_6813);
xnor U10091 (N_10091,N_7714,N_7402);
xor U10092 (N_10092,N_6508,N_6325);
nand U10093 (N_10093,N_7356,N_8132);
and U10094 (N_10094,N_7186,N_6593);
nor U10095 (N_10095,N_7307,N_7877);
and U10096 (N_10096,N_8961,N_8955);
and U10097 (N_10097,N_6741,N_8795);
nand U10098 (N_10098,N_8676,N_8534);
nor U10099 (N_10099,N_6739,N_7994);
or U10100 (N_10100,N_8480,N_6851);
xnor U10101 (N_10101,N_8589,N_7624);
or U10102 (N_10102,N_6333,N_6963);
and U10103 (N_10103,N_6769,N_8073);
or U10104 (N_10104,N_8326,N_7194);
and U10105 (N_10105,N_8488,N_7620);
or U10106 (N_10106,N_7302,N_7334);
xor U10107 (N_10107,N_8620,N_8700);
and U10108 (N_10108,N_7264,N_7097);
or U10109 (N_10109,N_7445,N_8111);
xor U10110 (N_10110,N_7218,N_8578);
xor U10111 (N_10111,N_6055,N_7335);
nor U10112 (N_10112,N_6862,N_6484);
nand U10113 (N_10113,N_8037,N_7899);
or U10114 (N_10114,N_6549,N_6376);
nand U10115 (N_10115,N_7614,N_8092);
and U10116 (N_10116,N_6028,N_8072);
nor U10117 (N_10117,N_7325,N_7124);
nor U10118 (N_10118,N_7532,N_8192);
nor U10119 (N_10119,N_7725,N_6608);
nand U10120 (N_10120,N_7648,N_7703);
xor U10121 (N_10121,N_8379,N_7466);
xor U10122 (N_10122,N_7952,N_7873);
nand U10123 (N_10123,N_7276,N_7129);
nor U10124 (N_10124,N_7317,N_8682);
and U10125 (N_10125,N_8650,N_8570);
nor U10126 (N_10126,N_8452,N_6829);
or U10127 (N_10127,N_8924,N_7597);
xnor U10128 (N_10128,N_7099,N_6765);
xor U10129 (N_10129,N_8937,N_6722);
or U10130 (N_10130,N_6367,N_8810);
nor U10131 (N_10131,N_6555,N_8256);
nor U10132 (N_10132,N_8302,N_6241);
and U10133 (N_10133,N_6398,N_7447);
xor U10134 (N_10134,N_8415,N_6083);
or U10135 (N_10135,N_6091,N_6516);
and U10136 (N_10136,N_8607,N_6237);
nand U10137 (N_10137,N_6336,N_7750);
nor U10138 (N_10138,N_8979,N_7397);
nand U10139 (N_10139,N_6911,N_6175);
nor U10140 (N_10140,N_6831,N_7810);
nor U10141 (N_10141,N_7598,N_6876);
and U10142 (N_10142,N_7451,N_8295);
or U10143 (N_10143,N_7406,N_8140);
or U10144 (N_10144,N_6106,N_6856);
and U10145 (N_10145,N_8303,N_6052);
nor U10146 (N_10146,N_6706,N_7119);
nor U10147 (N_10147,N_8634,N_8687);
or U10148 (N_10148,N_7613,N_8391);
xor U10149 (N_10149,N_6495,N_7473);
nor U10150 (N_10150,N_7680,N_6728);
nand U10151 (N_10151,N_8028,N_7728);
nor U10152 (N_10152,N_8438,N_8803);
or U10153 (N_10153,N_8006,N_8330);
nor U10154 (N_10154,N_6281,N_7523);
and U10155 (N_10155,N_8008,N_8089);
nand U10156 (N_10156,N_7852,N_6434);
nor U10157 (N_10157,N_8995,N_6965);
and U10158 (N_10158,N_8849,N_8378);
nand U10159 (N_10159,N_6705,N_7146);
or U10160 (N_10160,N_6858,N_8854);
or U10161 (N_10161,N_7481,N_8317);
nand U10162 (N_10162,N_6363,N_6913);
xor U10163 (N_10163,N_8507,N_6926);
nand U10164 (N_10164,N_8637,N_7954);
xor U10165 (N_10165,N_7479,N_6294);
and U10166 (N_10166,N_8880,N_8217);
xor U10167 (N_10167,N_7085,N_8565);
or U10168 (N_10168,N_7132,N_8522);
or U10169 (N_10169,N_8318,N_8103);
xnor U10170 (N_10170,N_7187,N_8184);
and U10171 (N_10171,N_6547,N_8241);
nor U10172 (N_10172,N_7425,N_8088);
nand U10173 (N_10173,N_6318,N_7482);
and U10174 (N_10174,N_6946,N_8557);
or U10175 (N_10175,N_7836,N_8785);
and U10176 (N_10176,N_7556,N_7151);
nor U10177 (N_10177,N_6780,N_6640);
xnor U10178 (N_10178,N_8749,N_6806);
and U10179 (N_10179,N_7313,N_8109);
nor U10180 (N_10180,N_6321,N_8461);
nor U10181 (N_10181,N_7226,N_6531);
nand U10182 (N_10182,N_8735,N_6718);
nor U10183 (N_10183,N_6155,N_8278);
or U10184 (N_10184,N_8590,N_8881);
and U10185 (N_10185,N_8951,N_8402);
or U10186 (N_10186,N_7246,N_8674);
and U10187 (N_10187,N_8896,N_6031);
nor U10188 (N_10188,N_6520,N_8942);
and U10189 (N_10189,N_6054,N_6082);
and U10190 (N_10190,N_6909,N_7067);
nand U10191 (N_10191,N_8869,N_8984);
xnor U10192 (N_10192,N_6064,N_6960);
and U10193 (N_10193,N_7698,N_6770);
nor U10194 (N_10194,N_8494,N_6596);
or U10195 (N_10195,N_6894,N_8575);
nor U10196 (N_10196,N_8908,N_8375);
and U10197 (N_10197,N_7353,N_7441);
nand U10198 (N_10198,N_6753,N_6690);
or U10199 (N_10199,N_6639,N_7513);
and U10200 (N_10200,N_6897,N_7370);
xnor U10201 (N_10201,N_8859,N_8843);
and U10202 (N_10202,N_6310,N_8086);
nor U10203 (N_10203,N_6632,N_8938);
nor U10204 (N_10204,N_6600,N_7729);
nor U10205 (N_10205,N_8188,N_7475);
nor U10206 (N_10206,N_6509,N_6504);
xnor U10207 (N_10207,N_8549,N_6662);
nor U10208 (N_10208,N_8648,N_7575);
or U10209 (N_10209,N_7739,N_6955);
nand U10210 (N_10210,N_8237,N_6297);
nor U10211 (N_10211,N_6319,N_8463);
and U10212 (N_10212,N_6881,N_8980);
and U10213 (N_10213,N_8523,N_7188);
nand U10214 (N_10214,N_8179,N_8705);
and U10215 (N_10215,N_7792,N_7255);
and U10216 (N_10216,N_7738,N_6149);
nor U10217 (N_10217,N_7753,N_6627);
xor U10218 (N_10218,N_6886,N_7229);
or U10219 (N_10219,N_8633,N_7856);
nand U10220 (N_10220,N_7719,N_6601);
xor U10221 (N_10221,N_7690,N_8096);
xnor U10222 (N_10222,N_7101,N_6260);
nor U10223 (N_10223,N_6262,N_8173);
xor U10224 (N_10224,N_6668,N_7102);
and U10225 (N_10225,N_6437,N_7007);
and U10226 (N_10226,N_8930,N_7524);
nand U10227 (N_10227,N_6740,N_7458);
or U10228 (N_10228,N_6431,N_6688);
xor U10229 (N_10229,N_8431,N_8350);
nor U10230 (N_10230,N_7118,N_6621);
or U10231 (N_10231,N_7293,N_7512);
xor U10232 (N_10232,N_8352,N_8850);
and U10233 (N_10233,N_6359,N_6714);
nand U10234 (N_10234,N_6295,N_6830);
or U10235 (N_10235,N_8077,N_6178);
nor U10236 (N_10236,N_7933,N_6209);
xnor U10237 (N_10237,N_6933,N_7111);
xor U10238 (N_10238,N_7890,N_6399);
or U10239 (N_10239,N_6649,N_6077);
nor U10240 (N_10240,N_8102,N_8819);
or U10241 (N_10241,N_8220,N_7983);
xor U10242 (N_10242,N_6134,N_8121);
or U10243 (N_10243,N_6239,N_6610);
nand U10244 (N_10244,N_7154,N_6133);
and U10245 (N_10245,N_8834,N_6708);
nor U10246 (N_10246,N_7840,N_7743);
nand U10247 (N_10247,N_8194,N_6006);
and U10248 (N_10248,N_6148,N_8916);
or U10249 (N_10249,N_8063,N_8276);
nor U10250 (N_10250,N_7015,N_6326);
nand U10251 (N_10251,N_7579,N_7214);
nor U10252 (N_10252,N_8285,N_8106);
nand U10253 (N_10253,N_8405,N_8185);
and U10254 (N_10254,N_6748,N_6615);
and U10255 (N_10255,N_8816,N_6169);
xnor U10256 (N_10256,N_6009,N_8972);
nand U10257 (N_10257,N_6853,N_6140);
xor U10258 (N_10258,N_6122,N_6001);
xor U10259 (N_10259,N_6410,N_7662);
nor U10260 (N_10260,N_7000,N_7777);
nand U10261 (N_10261,N_6974,N_6165);
and U10262 (N_10262,N_6299,N_6723);
nand U10263 (N_10263,N_6625,N_8618);
and U10264 (N_10264,N_6905,N_8293);
nand U10265 (N_10265,N_8065,N_6968);
and U10266 (N_10266,N_6619,N_6633);
nand U10267 (N_10267,N_7308,N_7820);
xor U10268 (N_10268,N_6267,N_8717);
or U10269 (N_10269,N_7130,N_8731);
or U10270 (N_10270,N_6045,N_8057);
nor U10271 (N_10271,N_7835,N_8098);
or U10272 (N_10272,N_8363,N_6219);
or U10273 (N_10273,N_6647,N_7518);
xnor U10274 (N_10274,N_8134,N_6194);
or U10275 (N_10275,N_7574,N_7921);
nor U10276 (N_10276,N_6787,N_6997);
and U10277 (N_10277,N_6012,N_8800);
or U10278 (N_10278,N_6864,N_6578);
nand U10279 (N_10279,N_6277,N_7315);
nand U10280 (N_10280,N_7096,N_6085);
nor U10281 (N_10281,N_8838,N_7747);
nor U10282 (N_10282,N_6643,N_8974);
xor U10283 (N_10283,N_7142,N_6335);
or U10284 (N_10284,N_8257,N_6311);
or U10285 (N_10285,N_7809,N_8839);
or U10286 (N_10286,N_8358,N_6220);
nand U10287 (N_10287,N_6628,N_7968);
xor U10288 (N_10288,N_7404,N_8671);
xor U10289 (N_10289,N_8599,N_6745);
nor U10290 (N_10290,N_6985,N_6543);
nand U10291 (N_10291,N_6793,N_6464);
and U10292 (N_10292,N_7817,N_7990);
xor U10293 (N_10293,N_8611,N_8855);
nor U10294 (N_10294,N_7740,N_7615);
and U10295 (N_10295,N_6095,N_8919);
nor U10296 (N_10296,N_6995,N_8867);
nand U10297 (N_10297,N_7196,N_7503);
or U10298 (N_10298,N_8004,N_6298);
xnor U10299 (N_10299,N_6768,N_7583);
or U10300 (N_10300,N_6105,N_8091);
nor U10301 (N_10301,N_7679,N_7967);
or U10302 (N_10302,N_6755,N_6414);
or U10303 (N_10303,N_6037,N_6972);
or U10304 (N_10304,N_7454,N_7222);
and U10305 (N_10305,N_8372,N_8714);
nor U10306 (N_10306,N_8794,N_7706);
or U10307 (N_10307,N_8232,N_7436);
and U10308 (N_10308,N_6062,N_7012);
and U10309 (N_10309,N_8231,N_8789);
or U10310 (N_10310,N_6424,N_8041);
or U10311 (N_10311,N_8874,N_7265);
or U10312 (N_10312,N_7515,N_6108);
and U10313 (N_10313,N_7752,N_7675);
nand U10314 (N_10314,N_6969,N_6782);
xor U10315 (N_10315,N_7312,N_8030);
nor U10316 (N_10316,N_6307,N_8327);
nand U10317 (N_10317,N_6836,N_8501);
or U10318 (N_10318,N_7786,N_7969);
nand U10319 (N_10319,N_6703,N_8830);
or U10320 (N_10320,N_6550,N_7953);
or U10321 (N_10321,N_8567,N_6238);
xor U10322 (N_10322,N_6789,N_6967);
xnor U10323 (N_10323,N_7886,N_6345);
nand U10324 (N_10324,N_6020,N_6552);
xnor U10325 (N_10325,N_8149,N_7182);
nand U10326 (N_10326,N_7344,N_7069);
or U10327 (N_10327,N_6809,N_6624);
xnor U10328 (N_10328,N_6669,N_7341);
and U10329 (N_10329,N_7379,N_6505);
nand U10330 (N_10330,N_8665,N_7538);
and U10331 (N_10331,N_8013,N_7127);
and U10332 (N_10332,N_7557,N_7262);
xor U10333 (N_10333,N_6449,N_7173);
or U10334 (N_10334,N_7309,N_7984);
xor U10335 (N_10335,N_7375,N_6602);
and U10336 (N_10336,N_6800,N_7895);
or U10337 (N_10337,N_7017,N_7086);
nor U10338 (N_10338,N_7352,N_8771);
nor U10339 (N_10339,N_6137,N_7732);
or U10340 (N_10340,N_6172,N_8071);
nor U10341 (N_10341,N_7492,N_7838);
or U10342 (N_10342,N_7470,N_8561);
nor U10343 (N_10343,N_8248,N_8427);
nor U10344 (N_10344,N_7014,N_6288);
nand U10345 (N_10345,N_8207,N_8343);
nor U10346 (N_10346,N_6949,N_7960);
xnor U10347 (N_10347,N_8900,N_7924);
nor U10348 (N_10348,N_7372,N_8383);
and U10349 (N_10349,N_7149,N_8970);
xor U10350 (N_10350,N_8877,N_7569);
xor U10351 (N_10351,N_6139,N_8410);
xnor U10352 (N_10352,N_8510,N_8848);
and U10353 (N_10353,N_8728,N_8481);
nor U10354 (N_10354,N_7091,N_7275);
nor U10355 (N_10355,N_8807,N_7788);
nor U10356 (N_10356,N_8644,N_8078);
and U10357 (N_10357,N_6387,N_6191);
xnor U10358 (N_10358,N_7148,N_7434);
xnor U10359 (N_10359,N_7041,N_6247);
nand U10360 (N_10360,N_6010,N_7233);
nand U10361 (N_10361,N_7053,N_8396);
and U10362 (N_10362,N_8323,N_8443);
and U10363 (N_10363,N_7480,N_7444);
nor U10364 (N_10364,N_8294,N_7711);
xnor U10365 (N_10365,N_6231,N_6916);
nor U10366 (N_10366,N_8422,N_8491);
nand U10367 (N_10367,N_8099,N_6156);
nor U10368 (N_10368,N_8745,N_7790);
nor U10369 (N_10369,N_7004,N_7528);
xor U10370 (N_10370,N_7736,N_8890);
nor U10371 (N_10371,N_8503,N_8829);
or U10372 (N_10372,N_7713,N_6141);
nand U10373 (N_10373,N_6107,N_8982);
or U10374 (N_10374,N_7110,N_6383);
or U10375 (N_10375,N_8183,N_8827);
nand U10376 (N_10376,N_7708,N_7754);
nor U10377 (N_10377,N_6118,N_8866);
nand U10378 (N_10378,N_8504,N_8926);
xor U10379 (N_10379,N_6771,N_8632);
nor U10380 (N_10380,N_7299,N_7964);
xor U10381 (N_10381,N_6352,N_7616);
nand U10382 (N_10382,N_7192,N_7160);
xor U10383 (N_10383,N_7585,N_6885);
and U10384 (N_10384,N_8251,N_6978);
xnor U10385 (N_10385,N_7911,N_7879);
xor U10386 (N_10386,N_7851,N_7606);
and U10387 (N_10387,N_7414,N_8722);
xor U10388 (N_10388,N_8649,N_7176);
nor U10389 (N_10389,N_8546,N_8101);
xnor U10390 (N_10390,N_6214,N_7219);
xnor U10391 (N_10391,N_7670,N_6921);
and U10392 (N_10392,N_8983,N_7484);
nor U10393 (N_10393,N_7843,N_7094);
and U10394 (N_10394,N_7374,N_6443);
nor U10395 (N_10395,N_6726,N_7805);
xor U10396 (N_10396,N_7839,N_6115);
xnor U10397 (N_10397,N_6988,N_6737);
nand U10398 (N_10398,N_8846,N_8898);
or U10399 (N_10399,N_7909,N_6146);
nand U10400 (N_10400,N_8493,N_6735);
or U10401 (N_10401,N_8139,N_7138);
xor U10402 (N_10402,N_7064,N_6996);
and U10403 (N_10403,N_7931,N_8157);
nor U10404 (N_10404,N_7818,N_6784);
xnor U10405 (N_10405,N_7905,N_7350);
or U10406 (N_10406,N_6958,N_8784);
and U10407 (N_10407,N_8697,N_7384);
or U10408 (N_10408,N_7357,N_7539);
nand U10409 (N_10409,N_8210,N_7238);
and U10410 (N_10410,N_6754,N_6582);
nor U10411 (N_10411,N_7050,N_6859);
and U10412 (N_10412,N_7483,N_6199);
or U10413 (N_10413,N_6129,N_6937);
nand U10414 (N_10414,N_8673,N_6380);
xnor U10415 (N_10415,N_6989,N_7973);
and U10416 (N_10416,N_8956,N_8738);
nor U10417 (N_10417,N_7634,N_7368);
xnor U10418 (N_10418,N_7584,N_7645);
nand U10419 (N_10419,N_6408,N_6528);
nor U10420 (N_10420,N_7623,N_8692);
or U10421 (N_10421,N_7780,N_6678);
nor U10422 (N_10422,N_6523,N_7018);
or U10423 (N_10423,N_6502,N_7565);
or U10424 (N_10424,N_8268,N_7361);
or U10425 (N_10425,N_6848,N_7049);
and U10426 (N_10426,N_7885,N_6271);
and U10427 (N_10427,N_6412,N_6145);
nand U10428 (N_10428,N_6846,N_8314);
and U10429 (N_10429,N_7904,N_8451);
nor U10430 (N_10430,N_6433,N_6750);
or U10431 (N_10431,N_8646,N_6979);
xor U10432 (N_10432,N_8126,N_7407);
nor U10433 (N_10433,N_7268,N_7772);
and U10434 (N_10434,N_7412,N_7159);
xnor U10435 (N_10435,N_7966,N_8222);
and U10436 (N_10436,N_7081,N_6962);
or U10437 (N_10437,N_8585,N_6256);
and U10438 (N_10438,N_6187,N_7570);
nand U10439 (N_10439,N_6617,N_8584);
xnor U10440 (N_10440,N_7411,N_7825);
and U10441 (N_10441,N_6002,N_6035);
nand U10442 (N_10442,N_6571,N_8489);
nor U10443 (N_10443,N_8836,N_6312);
or U10444 (N_10444,N_6879,N_8428);
xor U10445 (N_10445,N_7502,N_7610);
nand U10446 (N_10446,N_6497,N_6715);
nand U10447 (N_10447,N_7025,N_7145);
and U10448 (N_10448,N_7776,N_7717);
xnor U10449 (N_10449,N_6727,N_7199);
xor U10450 (N_10450,N_6986,N_8264);
nor U10451 (N_10451,N_8450,N_7637);
xnor U10452 (N_10452,N_6980,N_7224);
nor U10453 (N_10453,N_7033,N_8696);
or U10454 (N_10454,N_7175,N_7070);
or U10455 (N_10455,N_6021,N_8340);
nand U10456 (N_10456,N_8197,N_8417);
or U10457 (N_10457,N_8689,N_8178);
nand U10458 (N_10458,N_8666,N_6442);
nand U10459 (N_10459,N_6883,N_6595);
nor U10460 (N_10460,N_6233,N_7395);
and U10461 (N_10461,N_8433,N_8182);
and U10462 (N_10462,N_8801,N_7608);
nand U10463 (N_10463,N_6612,N_6458);
xnor U10464 (N_10464,N_6365,N_6493);
and U10465 (N_10465,N_6646,N_6803);
xor U10466 (N_10466,N_7380,N_6302);
xor U10467 (N_10467,N_7408,N_8747);
and U10468 (N_10468,N_6285,N_7988);
or U10469 (N_10469,N_8339,N_8990);
and U10470 (N_10470,N_7225,N_8442);
nand U10471 (N_10471,N_6766,N_8813);
or U10472 (N_10472,N_6611,N_7604);
nor U10473 (N_10473,N_8913,N_6730);
xnor U10474 (N_10474,N_8996,N_7529);
nand U10475 (N_10475,N_7517,N_7562);
and U10476 (N_10476,N_6585,N_8852);
nor U10477 (N_10477,N_7995,N_7956);
and U10478 (N_10478,N_7165,N_8010);
and U10479 (N_10479,N_8397,N_8215);
or U10480 (N_10480,N_8786,N_6654);
nand U10481 (N_10481,N_8429,N_8709);
nand U10482 (N_10482,N_8054,N_6492);
nand U10483 (N_10483,N_6560,N_8764);
and U10484 (N_10484,N_7010,N_6657);
nor U10485 (N_10485,N_7906,N_7252);
nor U10486 (N_10486,N_7607,N_7259);
nand U10487 (N_10487,N_7922,N_6121);
and U10488 (N_10488,N_6221,N_7459);
nand U10489 (N_10489,N_8946,N_6817);
xnor U10490 (N_10490,N_8435,N_8879);
and U10491 (N_10491,N_8097,N_8639);
nor U10492 (N_10492,N_6374,N_8203);
nand U10493 (N_10493,N_6871,N_6350);
or U10494 (N_10494,N_7487,N_6366);
or U10495 (N_10495,N_7654,N_8592);
and U10496 (N_10496,N_7845,N_6720);
nand U10497 (N_10497,N_6790,N_8308);
nor U10498 (N_10498,N_7045,N_8075);
nand U10499 (N_10499,N_7476,N_7842);
nor U10500 (N_10500,N_8808,N_6569);
nor U10501 (N_10501,N_7964,N_8820);
or U10502 (N_10502,N_8087,N_7756);
nor U10503 (N_10503,N_7235,N_6463);
xor U10504 (N_10504,N_8784,N_6196);
nor U10505 (N_10505,N_8834,N_6430);
nand U10506 (N_10506,N_6647,N_6900);
and U10507 (N_10507,N_8125,N_8607);
nand U10508 (N_10508,N_7674,N_8114);
nor U10509 (N_10509,N_7935,N_8981);
or U10510 (N_10510,N_7684,N_8832);
and U10511 (N_10511,N_6072,N_6262);
nand U10512 (N_10512,N_7403,N_6830);
xnor U10513 (N_10513,N_7452,N_6739);
nor U10514 (N_10514,N_8031,N_8985);
nor U10515 (N_10515,N_6494,N_7190);
xnor U10516 (N_10516,N_6845,N_6066);
nor U10517 (N_10517,N_8574,N_7499);
xnor U10518 (N_10518,N_8578,N_6441);
and U10519 (N_10519,N_8058,N_8481);
nor U10520 (N_10520,N_8926,N_8044);
or U10521 (N_10521,N_6454,N_8265);
or U10522 (N_10522,N_6703,N_6435);
and U10523 (N_10523,N_8538,N_6121);
nor U10524 (N_10524,N_8002,N_8024);
nand U10525 (N_10525,N_7146,N_8867);
nor U10526 (N_10526,N_8490,N_7689);
and U10527 (N_10527,N_6185,N_8041);
xnor U10528 (N_10528,N_7977,N_6576);
nor U10529 (N_10529,N_6496,N_7848);
or U10530 (N_10530,N_7462,N_8568);
nand U10531 (N_10531,N_7587,N_8441);
or U10532 (N_10532,N_8086,N_6508);
or U10533 (N_10533,N_7807,N_6208);
xor U10534 (N_10534,N_7364,N_6323);
and U10535 (N_10535,N_8759,N_8210);
xor U10536 (N_10536,N_6515,N_8801);
xnor U10537 (N_10537,N_7994,N_8465);
nand U10538 (N_10538,N_6651,N_7329);
nor U10539 (N_10539,N_8936,N_7806);
or U10540 (N_10540,N_7988,N_6713);
and U10541 (N_10541,N_8013,N_7335);
nand U10542 (N_10542,N_7645,N_8258);
nand U10543 (N_10543,N_7268,N_6324);
nor U10544 (N_10544,N_7645,N_8621);
or U10545 (N_10545,N_6995,N_8130);
xor U10546 (N_10546,N_8317,N_7988);
nand U10547 (N_10547,N_7388,N_7163);
nor U10548 (N_10548,N_7016,N_6567);
nand U10549 (N_10549,N_6614,N_6859);
xor U10550 (N_10550,N_6934,N_7897);
or U10551 (N_10551,N_6016,N_8375);
and U10552 (N_10552,N_7312,N_7808);
nand U10553 (N_10553,N_7497,N_7737);
nand U10554 (N_10554,N_6935,N_7318);
and U10555 (N_10555,N_6498,N_7169);
or U10556 (N_10556,N_6428,N_7989);
nand U10557 (N_10557,N_7822,N_8855);
or U10558 (N_10558,N_6634,N_8908);
nand U10559 (N_10559,N_6497,N_8823);
nor U10560 (N_10560,N_6668,N_7300);
and U10561 (N_10561,N_8308,N_7594);
or U10562 (N_10562,N_8843,N_7312);
nand U10563 (N_10563,N_6893,N_6327);
nand U10564 (N_10564,N_7248,N_8361);
nor U10565 (N_10565,N_8691,N_7404);
nor U10566 (N_10566,N_8312,N_6817);
nand U10567 (N_10567,N_6312,N_6597);
or U10568 (N_10568,N_7663,N_8028);
xnor U10569 (N_10569,N_7641,N_7818);
and U10570 (N_10570,N_8868,N_7709);
xor U10571 (N_10571,N_7726,N_8306);
xnor U10572 (N_10572,N_7119,N_6519);
xor U10573 (N_10573,N_6113,N_8219);
nor U10574 (N_10574,N_6222,N_8625);
xor U10575 (N_10575,N_6931,N_7533);
xor U10576 (N_10576,N_7117,N_6590);
nor U10577 (N_10577,N_6535,N_6747);
nor U10578 (N_10578,N_7576,N_7336);
and U10579 (N_10579,N_6054,N_8529);
and U10580 (N_10580,N_6981,N_8310);
nand U10581 (N_10581,N_7489,N_7424);
xor U10582 (N_10582,N_8323,N_7821);
nand U10583 (N_10583,N_7275,N_6608);
or U10584 (N_10584,N_8595,N_8348);
or U10585 (N_10585,N_6073,N_6868);
nand U10586 (N_10586,N_8552,N_8801);
or U10587 (N_10587,N_7426,N_8910);
nand U10588 (N_10588,N_6892,N_8763);
or U10589 (N_10589,N_6361,N_7368);
nor U10590 (N_10590,N_8541,N_8745);
nand U10591 (N_10591,N_6804,N_6802);
nand U10592 (N_10592,N_6666,N_7644);
or U10593 (N_10593,N_6995,N_7968);
and U10594 (N_10594,N_7639,N_7660);
nand U10595 (N_10595,N_7114,N_8929);
xnor U10596 (N_10596,N_8263,N_8216);
xnor U10597 (N_10597,N_7644,N_8840);
or U10598 (N_10598,N_6725,N_6469);
nand U10599 (N_10599,N_6078,N_7157);
and U10600 (N_10600,N_7203,N_6543);
and U10601 (N_10601,N_6874,N_8499);
xor U10602 (N_10602,N_7333,N_7995);
nor U10603 (N_10603,N_8427,N_8936);
or U10604 (N_10604,N_8519,N_7827);
or U10605 (N_10605,N_8345,N_7498);
nor U10606 (N_10606,N_7973,N_8741);
nand U10607 (N_10607,N_6320,N_8143);
and U10608 (N_10608,N_8075,N_8003);
xnor U10609 (N_10609,N_6268,N_8658);
nand U10610 (N_10610,N_8183,N_6227);
nor U10611 (N_10611,N_6752,N_8468);
and U10612 (N_10612,N_8317,N_6363);
or U10613 (N_10613,N_6114,N_8664);
nor U10614 (N_10614,N_6279,N_6119);
nor U10615 (N_10615,N_7993,N_8064);
nor U10616 (N_10616,N_8712,N_7392);
nor U10617 (N_10617,N_8908,N_8057);
or U10618 (N_10618,N_6086,N_6753);
nand U10619 (N_10619,N_7177,N_7996);
nor U10620 (N_10620,N_6977,N_6619);
or U10621 (N_10621,N_8363,N_6392);
and U10622 (N_10622,N_7220,N_6769);
xor U10623 (N_10623,N_7197,N_7741);
xor U10624 (N_10624,N_8578,N_8709);
or U10625 (N_10625,N_7222,N_7136);
xnor U10626 (N_10626,N_8631,N_7780);
nor U10627 (N_10627,N_6002,N_6007);
xnor U10628 (N_10628,N_7652,N_6548);
xor U10629 (N_10629,N_7605,N_7289);
nor U10630 (N_10630,N_8184,N_7745);
nand U10631 (N_10631,N_7061,N_8759);
and U10632 (N_10632,N_7694,N_8145);
nor U10633 (N_10633,N_7466,N_7930);
and U10634 (N_10634,N_8136,N_7588);
or U10635 (N_10635,N_7688,N_7677);
and U10636 (N_10636,N_8072,N_6303);
nor U10637 (N_10637,N_8302,N_7710);
and U10638 (N_10638,N_8713,N_6856);
nand U10639 (N_10639,N_6383,N_7929);
or U10640 (N_10640,N_8894,N_7875);
xor U10641 (N_10641,N_7851,N_7099);
or U10642 (N_10642,N_8565,N_8354);
xor U10643 (N_10643,N_6409,N_8061);
and U10644 (N_10644,N_7108,N_8599);
xnor U10645 (N_10645,N_6947,N_7915);
or U10646 (N_10646,N_7535,N_8162);
xor U10647 (N_10647,N_8544,N_7610);
nor U10648 (N_10648,N_7826,N_8045);
nand U10649 (N_10649,N_6071,N_8569);
or U10650 (N_10650,N_6633,N_7621);
and U10651 (N_10651,N_8355,N_7194);
and U10652 (N_10652,N_6078,N_8315);
nor U10653 (N_10653,N_8443,N_6424);
nor U10654 (N_10654,N_7283,N_7456);
nand U10655 (N_10655,N_8229,N_7656);
nand U10656 (N_10656,N_8282,N_6984);
nor U10657 (N_10657,N_8257,N_8476);
nor U10658 (N_10658,N_7967,N_6337);
xor U10659 (N_10659,N_6911,N_8009);
nor U10660 (N_10660,N_6602,N_7345);
or U10661 (N_10661,N_6435,N_7870);
nor U10662 (N_10662,N_8547,N_6926);
xor U10663 (N_10663,N_7693,N_8382);
and U10664 (N_10664,N_6755,N_8914);
and U10665 (N_10665,N_6863,N_6100);
or U10666 (N_10666,N_7739,N_8845);
nand U10667 (N_10667,N_8586,N_7938);
nor U10668 (N_10668,N_8440,N_8521);
nor U10669 (N_10669,N_8917,N_7600);
nor U10670 (N_10670,N_8781,N_8110);
xor U10671 (N_10671,N_7669,N_6141);
nor U10672 (N_10672,N_7476,N_6471);
or U10673 (N_10673,N_6723,N_7039);
nor U10674 (N_10674,N_6941,N_8691);
and U10675 (N_10675,N_6874,N_6148);
and U10676 (N_10676,N_7710,N_6370);
xor U10677 (N_10677,N_8855,N_8804);
nor U10678 (N_10678,N_8336,N_6059);
or U10679 (N_10679,N_6289,N_8696);
xnor U10680 (N_10680,N_7798,N_8211);
xnor U10681 (N_10681,N_8288,N_8282);
xor U10682 (N_10682,N_6597,N_8266);
nor U10683 (N_10683,N_6864,N_8339);
and U10684 (N_10684,N_6177,N_8717);
nor U10685 (N_10685,N_8679,N_6290);
nand U10686 (N_10686,N_8139,N_7345);
nor U10687 (N_10687,N_7097,N_8699);
and U10688 (N_10688,N_8130,N_8384);
or U10689 (N_10689,N_6433,N_7776);
and U10690 (N_10690,N_7666,N_8070);
or U10691 (N_10691,N_8336,N_6158);
and U10692 (N_10692,N_6318,N_6664);
xnor U10693 (N_10693,N_7270,N_6311);
nor U10694 (N_10694,N_6901,N_7167);
nand U10695 (N_10695,N_6327,N_7183);
or U10696 (N_10696,N_8792,N_7174);
nand U10697 (N_10697,N_6203,N_8941);
xnor U10698 (N_10698,N_8193,N_6265);
xor U10699 (N_10699,N_6739,N_7486);
nand U10700 (N_10700,N_7376,N_6657);
nand U10701 (N_10701,N_7473,N_7270);
nor U10702 (N_10702,N_8500,N_7940);
nor U10703 (N_10703,N_7897,N_8754);
nor U10704 (N_10704,N_7326,N_6761);
xor U10705 (N_10705,N_6414,N_7545);
and U10706 (N_10706,N_7573,N_8199);
and U10707 (N_10707,N_8848,N_6376);
or U10708 (N_10708,N_7682,N_8237);
or U10709 (N_10709,N_8870,N_8405);
nand U10710 (N_10710,N_6488,N_8981);
nor U10711 (N_10711,N_8502,N_8094);
nor U10712 (N_10712,N_7760,N_6823);
nand U10713 (N_10713,N_7980,N_8130);
xor U10714 (N_10714,N_8889,N_7749);
or U10715 (N_10715,N_6498,N_8901);
nor U10716 (N_10716,N_7341,N_6143);
nand U10717 (N_10717,N_8967,N_7496);
nand U10718 (N_10718,N_6766,N_6463);
or U10719 (N_10719,N_8694,N_6427);
nand U10720 (N_10720,N_7217,N_6353);
nand U10721 (N_10721,N_6483,N_6587);
nand U10722 (N_10722,N_7418,N_8804);
nor U10723 (N_10723,N_7951,N_6115);
nor U10724 (N_10724,N_6949,N_6770);
xnor U10725 (N_10725,N_8221,N_6788);
nand U10726 (N_10726,N_8248,N_7138);
nor U10727 (N_10727,N_8762,N_6648);
nor U10728 (N_10728,N_6042,N_8070);
and U10729 (N_10729,N_6202,N_8813);
and U10730 (N_10730,N_8773,N_8987);
xor U10731 (N_10731,N_6591,N_6738);
nor U10732 (N_10732,N_8538,N_6844);
and U10733 (N_10733,N_6546,N_7846);
xor U10734 (N_10734,N_7686,N_7727);
or U10735 (N_10735,N_6015,N_6175);
nand U10736 (N_10736,N_8801,N_8428);
nor U10737 (N_10737,N_7807,N_8335);
nand U10738 (N_10738,N_8317,N_7837);
and U10739 (N_10739,N_7244,N_7762);
or U10740 (N_10740,N_8834,N_8099);
nor U10741 (N_10741,N_6342,N_7428);
and U10742 (N_10742,N_7826,N_7873);
nand U10743 (N_10743,N_8033,N_8102);
or U10744 (N_10744,N_6288,N_8549);
or U10745 (N_10745,N_6235,N_8717);
and U10746 (N_10746,N_8683,N_7588);
or U10747 (N_10747,N_6422,N_8863);
and U10748 (N_10748,N_6569,N_6649);
or U10749 (N_10749,N_6754,N_6811);
xor U10750 (N_10750,N_8756,N_8371);
or U10751 (N_10751,N_7282,N_7899);
or U10752 (N_10752,N_8180,N_8509);
xnor U10753 (N_10753,N_6644,N_6009);
xnor U10754 (N_10754,N_6558,N_8223);
nand U10755 (N_10755,N_7939,N_6066);
nand U10756 (N_10756,N_8905,N_7683);
nor U10757 (N_10757,N_8768,N_6909);
xnor U10758 (N_10758,N_6229,N_8902);
or U10759 (N_10759,N_6763,N_7742);
nand U10760 (N_10760,N_6104,N_7588);
xnor U10761 (N_10761,N_6853,N_6113);
nand U10762 (N_10762,N_7825,N_6982);
and U10763 (N_10763,N_7747,N_6941);
nand U10764 (N_10764,N_7412,N_8726);
nand U10765 (N_10765,N_6415,N_8649);
nand U10766 (N_10766,N_8384,N_8339);
and U10767 (N_10767,N_7684,N_6974);
nor U10768 (N_10768,N_7922,N_8853);
or U10769 (N_10769,N_6005,N_6606);
or U10770 (N_10770,N_6424,N_8351);
and U10771 (N_10771,N_8865,N_7241);
xor U10772 (N_10772,N_7768,N_8547);
xnor U10773 (N_10773,N_7957,N_8696);
nand U10774 (N_10774,N_7336,N_6170);
or U10775 (N_10775,N_6742,N_8195);
nor U10776 (N_10776,N_8306,N_6324);
and U10777 (N_10777,N_6329,N_8600);
nor U10778 (N_10778,N_8623,N_8330);
nor U10779 (N_10779,N_7087,N_6617);
nor U10780 (N_10780,N_8558,N_7469);
or U10781 (N_10781,N_6072,N_8404);
and U10782 (N_10782,N_8549,N_6438);
nor U10783 (N_10783,N_6609,N_6808);
nand U10784 (N_10784,N_7490,N_7856);
xnor U10785 (N_10785,N_8852,N_6266);
or U10786 (N_10786,N_6514,N_6492);
or U10787 (N_10787,N_6189,N_8757);
and U10788 (N_10788,N_7186,N_7628);
xnor U10789 (N_10789,N_8689,N_7392);
xor U10790 (N_10790,N_6243,N_8523);
xnor U10791 (N_10791,N_6322,N_6906);
and U10792 (N_10792,N_8836,N_6158);
or U10793 (N_10793,N_6416,N_7306);
or U10794 (N_10794,N_8926,N_6275);
nand U10795 (N_10795,N_8102,N_7775);
nand U10796 (N_10796,N_8626,N_8998);
xor U10797 (N_10797,N_8510,N_8374);
nor U10798 (N_10798,N_7930,N_7483);
nand U10799 (N_10799,N_8925,N_8126);
and U10800 (N_10800,N_8342,N_7294);
nand U10801 (N_10801,N_8975,N_7108);
or U10802 (N_10802,N_6052,N_8057);
or U10803 (N_10803,N_6371,N_6540);
nand U10804 (N_10804,N_7927,N_8135);
nand U10805 (N_10805,N_6712,N_8280);
or U10806 (N_10806,N_6203,N_8497);
nand U10807 (N_10807,N_8443,N_8964);
nor U10808 (N_10808,N_8279,N_8229);
nand U10809 (N_10809,N_7299,N_8752);
or U10810 (N_10810,N_8109,N_8272);
nand U10811 (N_10811,N_8061,N_6333);
nand U10812 (N_10812,N_8812,N_8891);
nand U10813 (N_10813,N_7420,N_8000);
nor U10814 (N_10814,N_8859,N_8983);
nand U10815 (N_10815,N_6879,N_7779);
and U10816 (N_10816,N_7290,N_6492);
nor U10817 (N_10817,N_7077,N_7438);
xor U10818 (N_10818,N_6444,N_6003);
xor U10819 (N_10819,N_7303,N_8486);
nor U10820 (N_10820,N_8931,N_8859);
or U10821 (N_10821,N_6535,N_7683);
nor U10822 (N_10822,N_7859,N_7492);
nand U10823 (N_10823,N_7193,N_6025);
or U10824 (N_10824,N_7224,N_8408);
nand U10825 (N_10825,N_7158,N_7037);
or U10826 (N_10826,N_8920,N_7214);
and U10827 (N_10827,N_6081,N_6060);
nand U10828 (N_10828,N_6751,N_8252);
and U10829 (N_10829,N_8793,N_6638);
nor U10830 (N_10830,N_6742,N_7776);
or U10831 (N_10831,N_6598,N_8665);
xor U10832 (N_10832,N_8826,N_8925);
nand U10833 (N_10833,N_8280,N_8337);
nand U10834 (N_10834,N_7784,N_8152);
xor U10835 (N_10835,N_8027,N_6877);
or U10836 (N_10836,N_6271,N_6170);
xor U10837 (N_10837,N_8138,N_8294);
nand U10838 (N_10838,N_8357,N_7949);
xor U10839 (N_10839,N_8090,N_8181);
xor U10840 (N_10840,N_6103,N_7802);
and U10841 (N_10841,N_7507,N_6870);
nor U10842 (N_10842,N_7970,N_7540);
or U10843 (N_10843,N_7344,N_7841);
nor U10844 (N_10844,N_7998,N_7778);
nand U10845 (N_10845,N_6102,N_6643);
and U10846 (N_10846,N_7383,N_8842);
or U10847 (N_10847,N_6764,N_7425);
or U10848 (N_10848,N_6260,N_7849);
or U10849 (N_10849,N_8458,N_6613);
nor U10850 (N_10850,N_6232,N_7107);
nand U10851 (N_10851,N_8518,N_7801);
nor U10852 (N_10852,N_6516,N_6892);
or U10853 (N_10853,N_8004,N_6423);
and U10854 (N_10854,N_7230,N_8459);
or U10855 (N_10855,N_8685,N_7298);
nand U10856 (N_10856,N_7658,N_8941);
and U10857 (N_10857,N_6006,N_7749);
nor U10858 (N_10858,N_6500,N_7470);
and U10859 (N_10859,N_6063,N_6713);
or U10860 (N_10860,N_7783,N_6433);
nor U10861 (N_10861,N_6417,N_6916);
xnor U10862 (N_10862,N_6205,N_8811);
nand U10863 (N_10863,N_6185,N_7831);
nand U10864 (N_10864,N_8322,N_8128);
xnor U10865 (N_10865,N_6111,N_6629);
xor U10866 (N_10866,N_6914,N_8042);
nand U10867 (N_10867,N_8773,N_8920);
xor U10868 (N_10868,N_6306,N_6788);
and U10869 (N_10869,N_6726,N_6707);
and U10870 (N_10870,N_8230,N_7785);
nand U10871 (N_10871,N_8496,N_7385);
and U10872 (N_10872,N_8158,N_8434);
xor U10873 (N_10873,N_7116,N_7987);
or U10874 (N_10874,N_8101,N_8042);
or U10875 (N_10875,N_6020,N_6980);
nand U10876 (N_10876,N_7453,N_8356);
nand U10877 (N_10877,N_7747,N_7406);
and U10878 (N_10878,N_8228,N_6539);
and U10879 (N_10879,N_8228,N_7621);
xnor U10880 (N_10880,N_8487,N_6435);
or U10881 (N_10881,N_8928,N_8152);
and U10882 (N_10882,N_6902,N_6684);
nor U10883 (N_10883,N_7348,N_7612);
xor U10884 (N_10884,N_6549,N_8591);
and U10885 (N_10885,N_8569,N_7206);
nand U10886 (N_10886,N_6273,N_8241);
nor U10887 (N_10887,N_8700,N_7105);
or U10888 (N_10888,N_7615,N_6301);
or U10889 (N_10889,N_6510,N_6910);
or U10890 (N_10890,N_6739,N_7149);
nor U10891 (N_10891,N_8903,N_7059);
nor U10892 (N_10892,N_6333,N_8651);
xor U10893 (N_10893,N_8709,N_8246);
and U10894 (N_10894,N_6755,N_6302);
or U10895 (N_10895,N_8692,N_6512);
xor U10896 (N_10896,N_6296,N_8634);
and U10897 (N_10897,N_6200,N_6498);
nand U10898 (N_10898,N_6280,N_7978);
and U10899 (N_10899,N_7031,N_7720);
or U10900 (N_10900,N_7056,N_8625);
nand U10901 (N_10901,N_8686,N_6453);
and U10902 (N_10902,N_7076,N_8867);
xor U10903 (N_10903,N_7475,N_6538);
and U10904 (N_10904,N_7340,N_8364);
and U10905 (N_10905,N_6462,N_6640);
nor U10906 (N_10906,N_7625,N_7813);
and U10907 (N_10907,N_8454,N_7400);
nor U10908 (N_10908,N_6165,N_7202);
xnor U10909 (N_10909,N_8924,N_8504);
and U10910 (N_10910,N_8459,N_6209);
nand U10911 (N_10911,N_6164,N_7242);
nand U10912 (N_10912,N_7246,N_6618);
and U10913 (N_10913,N_8168,N_6073);
nor U10914 (N_10914,N_7759,N_7258);
or U10915 (N_10915,N_7099,N_8813);
or U10916 (N_10916,N_6919,N_8434);
xor U10917 (N_10917,N_8516,N_6783);
nand U10918 (N_10918,N_8989,N_8664);
nor U10919 (N_10919,N_6096,N_7615);
xnor U10920 (N_10920,N_7119,N_7297);
nor U10921 (N_10921,N_7192,N_6848);
xor U10922 (N_10922,N_8810,N_6666);
or U10923 (N_10923,N_6605,N_6574);
nor U10924 (N_10924,N_8946,N_6716);
or U10925 (N_10925,N_6333,N_8998);
nor U10926 (N_10926,N_7949,N_6309);
xor U10927 (N_10927,N_6706,N_6153);
nor U10928 (N_10928,N_8151,N_6250);
or U10929 (N_10929,N_7137,N_8979);
nor U10930 (N_10930,N_6041,N_7227);
nor U10931 (N_10931,N_8168,N_8147);
or U10932 (N_10932,N_8559,N_7274);
nor U10933 (N_10933,N_7277,N_8019);
nor U10934 (N_10934,N_8451,N_6378);
nand U10935 (N_10935,N_6645,N_6823);
nand U10936 (N_10936,N_6956,N_8001);
and U10937 (N_10937,N_7882,N_8658);
nand U10938 (N_10938,N_7394,N_8152);
nor U10939 (N_10939,N_8214,N_6883);
xnor U10940 (N_10940,N_6500,N_8247);
xor U10941 (N_10941,N_6931,N_6350);
nor U10942 (N_10942,N_6257,N_8444);
or U10943 (N_10943,N_6175,N_7272);
nor U10944 (N_10944,N_7874,N_7360);
nand U10945 (N_10945,N_6766,N_8131);
nand U10946 (N_10946,N_6029,N_6605);
nand U10947 (N_10947,N_6090,N_8868);
or U10948 (N_10948,N_8612,N_8735);
nand U10949 (N_10949,N_6416,N_7655);
nand U10950 (N_10950,N_8213,N_8583);
nor U10951 (N_10951,N_8984,N_8375);
or U10952 (N_10952,N_8664,N_7255);
xnor U10953 (N_10953,N_8261,N_8076);
and U10954 (N_10954,N_7319,N_7832);
or U10955 (N_10955,N_7695,N_8503);
and U10956 (N_10956,N_8237,N_8733);
nand U10957 (N_10957,N_7088,N_7773);
or U10958 (N_10958,N_8113,N_8699);
nand U10959 (N_10959,N_8972,N_6593);
and U10960 (N_10960,N_7593,N_7942);
nor U10961 (N_10961,N_8744,N_8820);
and U10962 (N_10962,N_6146,N_7713);
xor U10963 (N_10963,N_8406,N_8353);
xnor U10964 (N_10964,N_8982,N_8040);
nand U10965 (N_10965,N_8901,N_6053);
and U10966 (N_10966,N_7922,N_7656);
nor U10967 (N_10967,N_7730,N_6714);
xnor U10968 (N_10968,N_7151,N_8442);
nand U10969 (N_10969,N_8184,N_6946);
nand U10970 (N_10970,N_7482,N_6821);
nor U10971 (N_10971,N_6380,N_8112);
and U10972 (N_10972,N_7902,N_7958);
xor U10973 (N_10973,N_7478,N_7211);
nor U10974 (N_10974,N_7045,N_6913);
and U10975 (N_10975,N_7969,N_7127);
nor U10976 (N_10976,N_6611,N_6900);
nor U10977 (N_10977,N_8703,N_8592);
or U10978 (N_10978,N_7399,N_8777);
nor U10979 (N_10979,N_8511,N_8383);
nor U10980 (N_10980,N_7603,N_6646);
nor U10981 (N_10981,N_7193,N_6963);
xor U10982 (N_10982,N_8728,N_7125);
and U10983 (N_10983,N_7304,N_8560);
nand U10984 (N_10984,N_7191,N_8185);
nor U10985 (N_10985,N_8874,N_7051);
nor U10986 (N_10986,N_8040,N_7507);
or U10987 (N_10987,N_6295,N_6207);
xor U10988 (N_10988,N_8569,N_7806);
nor U10989 (N_10989,N_8634,N_8292);
nand U10990 (N_10990,N_6448,N_6225);
and U10991 (N_10991,N_6458,N_8774);
nor U10992 (N_10992,N_8299,N_7337);
or U10993 (N_10993,N_8228,N_6182);
or U10994 (N_10994,N_6891,N_7411);
nand U10995 (N_10995,N_6992,N_7214);
xnor U10996 (N_10996,N_8520,N_8326);
or U10997 (N_10997,N_7770,N_6029);
xor U10998 (N_10998,N_7704,N_7711);
or U10999 (N_10999,N_8411,N_7843);
or U11000 (N_11000,N_7056,N_6962);
or U11001 (N_11001,N_7098,N_7814);
nor U11002 (N_11002,N_6932,N_7611);
xor U11003 (N_11003,N_6158,N_6983);
xnor U11004 (N_11004,N_6719,N_7294);
xnor U11005 (N_11005,N_7283,N_7951);
xnor U11006 (N_11006,N_7773,N_8768);
and U11007 (N_11007,N_6783,N_6915);
and U11008 (N_11008,N_6546,N_6989);
xnor U11009 (N_11009,N_8605,N_7614);
and U11010 (N_11010,N_8017,N_6482);
nor U11011 (N_11011,N_8305,N_8606);
and U11012 (N_11012,N_8614,N_7673);
and U11013 (N_11013,N_6564,N_8510);
nor U11014 (N_11014,N_6409,N_7694);
or U11015 (N_11015,N_7146,N_6821);
nor U11016 (N_11016,N_8598,N_8249);
or U11017 (N_11017,N_6042,N_8038);
xor U11018 (N_11018,N_7387,N_7466);
nand U11019 (N_11019,N_7212,N_8668);
nand U11020 (N_11020,N_7686,N_6544);
nand U11021 (N_11021,N_6141,N_8961);
nand U11022 (N_11022,N_7441,N_8210);
xnor U11023 (N_11023,N_7855,N_6901);
and U11024 (N_11024,N_6972,N_6284);
nor U11025 (N_11025,N_6330,N_7247);
nand U11026 (N_11026,N_7257,N_8350);
or U11027 (N_11027,N_6007,N_8334);
nand U11028 (N_11028,N_7285,N_6500);
xnor U11029 (N_11029,N_6522,N_7632);
or U11030 (N_11030,N_7123,N_7239);
nand U11031 (N_11031,N_7791,N_6870);
and U11032 (N_11032,N_8892,N_6569);
nor U11033 (N_11033,N_6463,N_7482);
nand U11034 (N_11034,N_8930,N_7653);
xnor U11035 (N_11035,N_8754,N_8991);
xnor U11036 (N_11036,N_6610,N_8360);
nor U11037 (N_11037,N_8695,N_7605);
or U11038 (N_11038,N_8096,N_7831);
or U11039 (N_11039,N_8306,N_6335);
nor U11040 (N_11040,N_7103,N_6979);
or U11041 (N_11041,N_7416,N_7070);
and U11042 (N_11042,N_7927,N_8463);
and U11043 (N_11043,N_8644,N_8757);
nor U11044 (N_11044,N_8441,N_7324);
nand U11045 (N_11045,N_7832,N_6406);
xor U11046 (N_11046,N_6690,N_7093);
xnor U11047 (N_11047,N_7301,N_7909);
and U11048 (N_11048,N_6624,N_6938);
xnor U11049 (N_11049,N_6305,N_7377);
nor U11050 (N_11050,N_8642,N_6014);
nor U11051 (N_11051,N_8496,N_6260);
nor U11052 (N_11052,N_7329,N_8935);
and U11053 (N_11053,N_7662,N_6805);
and U11054 (N_11054,N_8356,N_8369);
and U11055 (N_11055,N_6341,N_7825);
or U11056 (N_11056,N_6585,N_8065);
nand U11057 (N_11057,N_7958,N_8996);
nor U11058 (N_11058,N_7557,N_7973);
xor U11059 (N_11059,N_8350,N_7511);
xor U11060 (N_11060,N_6358,N_7733);
nand U11061 (N_11061,N_7823,N_8283);
or U11062 (N_11062,N_6316,N_6622);
and U11063 (N_11063,N_7167,N_8641);
nor U11064 (N_11064,N_6436,N_7358);
and U11065 (N_11065,N_7399,N_8628);
xor U11066 (N_11066,N_6913,N_8744);
xnor U11067 (N_11067,N_7573,N_6678);
nor U11068 (N_11068,N_7867,N_8088);
nor U11069 (N_11069,N_7348,N_8223);
nor U11070 (N_11070,N_7253,N_6260);
nor U11071 (N_11071,N_8746,N_8578);
nor U11072 (N_11072,N_6752,N_6631);
nor U11073 (N_11073,N_7934,N_8414);
or U11074 (N_11074,N_7447,N_7894);
or U11075 (N_11075,N_7099,N_8961);
nand U11076 (N_11076,N_8995,N_7773);
or U11077 (N_11077,N_7691,N_7764);
or U11078 (N_11078,N_6253,N_6590);
or U11079 (N_11079,N_7817,N_6355);
nor U11080 (N_11080,N_6700,N_6730);
or U11081 (N_11081,N_7928,N_8198);
and U11082 (N_11082,N_7171,N_8222);
xnor U11083 (N_11083,N_7794,N_7220);
nor U11084 (N_11084,N_6599,N_7668);
xor U11085 (N_11085,N_6590,N_8505);
xor U11086 (N_11086,N_6757,N_7429);
and U11087 (N_11087,N_8145,N_7323);
xor U11088 (N_11088,N_7593,N_7684);
nor U11089 (N_11089,N_6786,N_7525);
and U11090 (N_11090,N_8199,N_6641);
nor U11091 (N_11091,N_6887,N_6572);
or U11092 (N_11092,N_8381,N_7515);
xnor U11093 (N_11093,N_8051,N_7783);
and U11094 (N_11094,N_8763,N_8967);
nand U11095 (N_11095,N_7879,N_6993);
nand U11096 (N_11096,N_6330,N_8071);
or U11097 (N_11097,N_6344,N_6215);
xor U11098 (N_11098,N_8945,N_6184);
or U11099 (N_11099,N_8114,N_6147);
xor U11100 (N_11100,N_6006,N_6721);
nor U11101 (N_11101,N_6368,N_7286);
nand U11102 (N_11102,N_6945,N_7248);
nor U11103 (N_11103,N_7370,N_8120);
and U11104 (N_11104,N_8016,N_8247);
and U11105 (N_11105,N_6952,N_8482);
and U11106 (N_11106,N_6261,N_8589);
or U11107 (N_11107,N_6556,N_6956);
nand U11108 (N_11108,N_8219,N_8164);
nor U11109 (N_11109,N_8199,N_6901);
nor U11110 (N_11110,N_7656,N_6688);
or U11111 (N_11111,N_7921,N_7307);
nand U11112 (N_11112,N_8453,N_8712);
or U11113 (N_11113,N_8037,N_7316);
nand U11114 (N_11114,N_6597,N_7903);
and U11115 (N_11115,N_6415,N_8540);
xor U11116 (N_11116,N_6670,N_7520);
nand U11117 (N_11117,N_8084,N_8353);
xnor U11118 (N_11118,N_8432,N_7108);
and U11119 (N_11119,N_6543,N_7208);
and U11120 (N_11120,N_7498,N_8174);
or U11121 (N_11121,N_6486,N_7016);
nor U11122 (N_11122,N_7675,N_7026);
or U11123 (N_11123,N_7284,N_6034);
nor U11124 (N_11124,N_6067,N_6262);
nor U11125 (N_11125,N_8938,N_7642);
nand U11126 (N_11126,N_8763,N_7032);
xor U11127 (N_11127,N_6928,N_6587);
nor U11128 (N_11128,N_6797,N_6500);
xor U11129 (N_11129,N_8717,N_8144);
or U11130 (N_11130,N_8800,N_8791);
xnor U11131 (N_11131,N_7226,N_7889);
nor U11132 (N_11132,N_6881,N_7600);
and U11133 (N_11133,N_8834,N_7424);
or U11134 (N_11134,N_7132,N_8747);
and U11135 (N_11135,N_8766,N_6074);
nand U11136 (N_11136,N_8383,N_8100);
nand U11137 (N_11137,N_8757,N_8428);
nand U11138 (N_11138,N_7524,N_6422);
nand U11139 (N_11139,N_8185,N_6866);
and U11140 (N_11140,N_8381,N_7115);
or U11141 (N_11141,N_7522,N_8883);
or U11142 (N_11142,N_8272,N_7516);
nor U11143 (N_11143,N_6801,N_8580);
or U11144 (N_11144,N_8324,N_6144);
xor U11145 (N_11145,N_7356,N_6264);
nand U11146 (N_11146,N_6657,N_6479);
nand U11147 (N_11147,N_6265,N_8129);
nor U11148 (N_11148,N_7629,N_6007);
or U11149 (N_11149,N_7381,N_7241);
and U11150 (N_11150,N_6298,N_6584);
nor U11151 (N_11151,N_7460,N_8519);
nand U11152 (N_11152,N_8604,N_6269);
xor U11153 (N_11153,N_6406,N_6189);
and U11154 (N_11154,N_8609,N_6661);
or U11155 (N_11155,N_6057,N_6623);
or U11156 (N_11156,N_7796,N_6717);
and U11157 (N_11157,N_6943,N_7059);
nor U11158 (N_11158,N_7239,N_7471);
or U11159 (N_11159,N_8126,N_6854);
nor U11160 (N_11160,N_8040,N_6733);
and U11161 (N_11161,N_6632,N_6929);
xor U11162 (N_11162,N_8271,N_8196);
or U11163 (N_11163,N_7195,N_8414);
xnor U11164 (N_11164,N_8522,N_8490);
nor U11165 (N_11165,N_8959,N_8498);
nand U11166 (N_11166,N_6996,N_7316);
nor U11167 (N_11167,N_8769,N_7941);
xnor U11168 (N_11168,N_7404,N_7439);
xor U11169 (N_11169,N_8064,N_6939);
or U11170 (N_11170,N_8159,N_6136);
or U11171 (N_11171,N_7082,N_7898);
and U11172 (N_11172,N_8378,N_7611);
nand U11173 (N_11173,N_6120,N_6798);
xnor U11174 (N_11174,N_7086,N_7091);
nand U11175 (N_11175,N_6811,N_7050);
nand U11176 (N_11176,N_8432,N_6971);
xor U11177 (N_11177,N_7444,N_8509);
xnor U11178 (N_11178,N_8101,N_8703);
or U11179 (N_11179,N_6446,N_8356);
xor U11180 (N_11180,N_8953,N_8674);
and U11181 (N_11181,N_7191,N_7965);
or U11182 (N_11182,N_7447,N_7996);
xnor U11183 (N_11183,N_6236,N_8852);
xnor U11184 (N_11184,N_8272,N_7371);
xor U11185 (N_11185,N_7488,N_8012);
xnor U11186 (N_11186,N_7462,N_6474);
nor U11187 (N_11187,N_8033,N_8888);
nor U11188 (N_11188,N_6650,N_8510);
nor U11189 (N_11189,N_8270,N_8444);
nor U11190 (N_11190,N_8034,N_7008);
nor U11191 (N_11191,N_7523,N_6862);
nor U11192 (N_11192,N_8294,N_6962);
nand U11193 (N_11193,N_8861,N_7435);
or U11194 (N_11194,N_7667,N_6016);
xnor U11195 (N_11195,N_7927,N_8227);
xor U11196 (N_11196,N_8251,N_6771);
and U11197 (N_11197,N_7525,N_7581);
and U11198 (N_11198,N_8179,N_8161);
xnor U11199 (N_11199,N_6957,N_7805);
or U11200 (N_11200,N_8428,N_6147);
and U11201 (N_11201,N_6780,N_6131);
and U11202 (N_11202,N_6936,N_6932);
nor U11203 (N_11203,N_7207,N_6959);
and U11204 (N_11204,N_7141,N_8202);
and U11205 (N_11205,N_6144,N_7015);
nand U11206 (N_11206,N_8073,N_8544);
and U11207 (N_11207,N_7896,N_6693);
nor U11208 (N_11208,N_6215,N_7404);
or U11209 (N_11209,N_7576,N_7573);
nor U11210 (N_11210,N_6796,N_6005);
nor U11211 (N_11211,N_8870,N_8633);
xnor U11212 (N_11212,N_7098,N_8283);
nor U11213 (N_11213,N_6134,N_7288);
nor U11214 (N_11214,N_7281,N_7252);
xnor U11215 (N_11215,N_8564,N_6633);
nand U11216 (N_11216,N_6491,N_7201);
and U11217 (N_11217,N_7339,N_7534);
nor U11218 (N_11218,N_6290,N_7325);
or U11219 (N_11219,N_7722,N_7948);
nand U11220 (N_11220,N_8054,N_7118);
and U11221 (N_11221,N_6741,N_7079);
nand U11222 (N_11222,N_8189,N_7837);
nor U11223 (N_11223,N_8492,N_8087);
nor U11224 (N_11224,N_7034,N_7003);
nor U11225 (N_11225,N_7114,N_8630);
nand U11226 (N_11226,N_8643,N_8676);
or U11227 (N_11227,N_8937,N_6587);
nor U11228 (N_11228,N_8393,N_7863);
and U11229 (N_11229,N_7332,N_7046);
xnor U11230 (N_11230,N_8590,N_8775);
and U11231 (N_11231,N_8891,N_7909);
xnor U11232 (N_11232,N_6335,N_6042);
nor U11233 (N_11233,N_6561,N_8967);
or U11234 (N_11234,N_8072,N_6058);
and U11235 (N_11235,N_6727,N_6334);
xnor U11236 (N_11236,N_7121,N_8299);
and U11237 (N_11237,N_6835,N_6348);
nor U11238 (N_11238,N_8812,N_6421);
nor U11239 (N_11239,N_8956,N_7631);
nor U11240 (N_11240,N_8787,N_8217);
and U11241 (N_11241,N_8171,N_7251);
and U11242 (N_11242,N_7471,N_7116);
nand U11243 (N_11243,N_7730,N_8563);
or U11244 (N_11244,N_6892,N_8165);
or U11245 (N_11245,N_6943,N_7105);
or U11246 (N_11246,N_6130,N_6653);
and U11247 (N_11247,N_8659,N_6952);
xnor U11248 (N_11248,N_6583,N_7733);
or U11249 (N_11249,N_8799,N_7885);
nand U11250 (N_11250,N_6227,N_6190);
nor U11251 (N_11251,N_6780,N_8421);
nor U11252 (N_11252,N_7100,N_8838);
xnor U11253 (N_11253,N_6565,N_6249);
xnor U11254 (N_11254,N_8747,N_6801);
nand U11255 (N_11255,N_6143,N_7246);
xor U11256 (N_11256,N_7371,N_6394);
and U11257 (N_11257,N_6405,N_8241);
and U11258 (N_11258,N_7355,N_8001);
nor U11259 (N_11259,N_6240,N_8504);
xor U11260 (N_11260,N_6738,N_6908);
xor U11261 (N_11261,N_8075,N_6470);
nand U11262 (N_11262,N_6627,N_7370);
xnor U11263 (N_11263,N_6752,N_8476);
nor U11264 (N_11264,N_6226,N_6622);
xor U11265 (N_11265,N_6527,N_6904);
xnor U11266 (N_11266,N_6578,N_7287);
nand U11267 (N_11267,N_8440,N_6704);
or U11268 (N_11268,N_7581,N_8456);
and U11269 (N_11269,N_7223,N_8729);
and U11270 (N_11270,N_7072,N_7933);
and U11271 (N_11271,N_6454,N_6200);
or U11272 (N_11272,N_6494,N_7088);
or U11273 (N_11273,N_8750,N_8664);
or U11274 (N_11274,N_6933,N_6668);
nor U11275 (N_11275,N_7834,N_6579);
nor U11276 (N_11276,N_7139,N_6591);
xnor U11277 (N_11277,N_7770,N_8334);
xnor U11278 (N_11278,N_6307,N_7708);
xnor U11279 (N_11279,N_6524,N_6619);
nand U11280 (N_11280,N_6409,N_8967);
xnor U11281 (N_11281,N_7284,N_8357);
nor U11282 (N_11282,N_8549,N_8579);
xor U11283 (N_11283,N_6056,N_7204);
or U11284 (N_11284,N_8102,N_6295);
or U11285 (N_11285,N_8367,N_6206);
nor U11286 (N_11286,N_8383,N_6812);
or U11287 (N_11287,N_7784,N_6561);
or U11288 (N_11288,N_7936,N_7602);
nand U11289 (N_11289,N_6630,N_8494);
xor U11290 (N_11290,N_6363,N_8655);
or U11291 (N_11291,N_6160,N_6355);
nor U11292 (N_11292,N_8286,N_7162);
and U11293 (N_11293,N_7057,N_6269);
nor U11294 (N_11294,N_7907,N_8389);
or U11295 (N_11295,N_7631,N_8252);
xnor U11296 (N_11296,N_7964,N_7870);
and U11297 (N_11297,N_6613,N_8884);
nor U11298 (N_11298,N_7674,N_7377);
nand U11299 (N_11299,N_7625,N_8460);
xor U11300 (N_11300,N_8502,N_7300);
or U11301 (N_11301,N_8278,N_8261);
or U11302 (N_11302,N_6663,N_8617);
and U11303 (N_11303,N_7509,N_7411);
xnor U11304 (N_11304,N_7892,N_6530);
and U11305 (N_11305,N_6182,N_6627);
nand U11306 (N_11306,N_7119,N_8314);
nor U11307 (N_11307,N_7371,N_6141);
xnor U11308 (N_11308,N_7871,N_8957);
or U11309 (N_11309,N_6211,N_8605);
nand U11310 (N_11310,N_8337,N_7791);
and U11311 (N_11311,N_7043,N_8515);
nor U11312 (N_11312,N_6652,N_8133);
and U11313 (N_11313,N_8955,N_7101);
and U11314 (N_11314,N_7188,N_7058);
xnor U11315 (N_11315,N_7929,N_8561);
or U11316 (N_11316,N_8538,N_7930);
and U11317 (N_11317,N_6928,N_8712);
nor U11318 (N_11318,N_6391,N_7576);
nand U11319 (N_11319,N_8535,N_8074);
or U11320 (N_11320,N_8596,N_7768);
and U11321 (N_11321,N_6353,N_7332);
or U11322 (N_11322,N_7833,N_7794);
nor U11323 (N_11323,N_6477,N_8173);
xor U11324 (N_11324,N_8991,N_6642);
xor U11325 (N_11325,N_6717,N_6408);
xor U11326 (N_11326,N_6938,N_6108);
or U11327 (N_11327,N_7469,N_7525);
and U11328 (N_11328,N_8475,N_6571);
nor U11329 (N_11329,N_6049,N_6738);
or U11330 (N_11330,N_7248,N_6840);
and U11331 (N_11331,N_8072,N_6721);
or U11332 (N_11332,N_8457,N_6591);
nand U11333 (N_11333,N_7366,N_7474);
nor U11334 (N_11334,N_7959,N_6048);
nor U11335 (N_11335,N_7554,N_8440);
xor U11336 (N_11336,N_7165,N_7350);
or U11337 (N_11337,N_7100,N_7993);
nand U11338 (N_11338,N_8890,N_8850);
xnor U11339 (N_11339,N_6920,N_6205);
nand U11340 (N_11340,N_8853,N_6665);
nand U11341 (N_11341,N_6996,N_7441);
nor U11342 (N_11342,N_8862,N_7905);
nand U11343 (N_11343,N_6369,N_8180);
and U11344 (N_11344,N_8373,N_8787);
and U11345 (N_11345,N_8865,N_7121);
nor U11346 (N_11346,N_6863,N_6038);
nand U11347 (N_11347,N_8326,N_6785);
nor U11348 (N_11348,N_6340,N_7058);
nor U11349 (N_11349,N_8348,N_8353);
nand U11350 (N_11350,N_8132,N_8471);
nor U11351 (N_11351,N_6038,N_7721);
or U11352 (N_11352,N_8531,N_7727);
nor U11353 (N_11353,N_8501,N_7190);
nor U11354 (N_11354,N_8438,N_8534);
xnor U11355 (N_11355,N_8394,N_6084);
nor U11356 (N_11356,N_7629,N_7695);
and U11357 (N_11357,N_7036,N_6527);
xnor U11358 (N_11358,N_8767,N_6729);
or U11359 (N_11359,N_8899,N_7595);
nor U11360 (N_11360,N_7891,N_7478);
nor U11361 (N_11361,N_8455,N_7899);
and U11362 (N_11362,N_8846,N_8877);
xnor U11363 (N_11363,N_8236,N_8239);
nand U11364 (N_11364,N_8832,N_8055);
and U11365 (N_11365,N_8916,N_8450);
nor U11366 (N_11366,N_6063,N_7563);
and U11367 (N_11367,N_8160,N_7872);
nand U11368 (N_11368,N_7517,N_6505);
xnor U11369 (N_11369,N_7621,N_7638);
xor U11370 (N_11370,N_7020,N_8140);
and U11371 (N_11371,N_8369,N_8049);
nor U11372 (N_11372,N_8786,N_7485);
and U11373 (N_11373,N_8590,N_8125);
nand U11374 (N_11374,N_8551,N_8315);
xor U11375 (N_11375,N_8820,N_6854);
and U11376 (N_11376,N_7160,N_6850);
or U11377 (N_11377,N_8426,N_8051);
or U11378 (N_11378,N_8793,N_8683);
xnor U11379 (N_11379,N_8613,N_8763);
and U11380 (N_11380,N_6490,N_7595);
or U11381 (N_11381,N_7093,N_8676);
nor U11382 (N_11382,N_6597,N_6611);
nand U11383 (N_11383,N_7858,N_7371);
xnor U11384 (N_11384,N_7858,N_8744);
or U11385 (N_11385,N_6204,N_7428);
nor U11386 (N_11386,N_6462,N_6409);
or U11387 (N_11387,N_8059,N_6370);
or U11388 (N_11388,N_7851,N_8268);
or U11389 (N_11389,N_7779,N_7285);
nand U11390 (N_11390,N_6710,N_7389);
and U11391 (N_11391,N_8139,N_7082);
nand U11392 (N_11392,N_7790,N_6701);
and U11393 (N_11393,N_7457,N_7297);
and U11394 (N_11394,N_8659,N_8122);
or U11395 (N_11395,N_8937,N_7863);
or U11396 (N_11396,N_7613,N_7645);
or U11397 (N_11397,N_8368,N_6079);
and U11398 (N_11398,N_6795,N_8717);
nand U11399 (N_11399,N_7601,N_8831);
or U11400 (N_11400,N_8246,N_7818);
or U11401 (N_11401,N_6643,N_7956);
nor U11402 (N_11402,N_8645,N_7812);
and U11403 (N_11403,N_8346,N_7859);
and U11404 (N_11404,N_7872,N_7063);
xor U11405 (N_11405,N_6986,N_7685);
nor U11406 (N_11406,N_7799,N_7723);
nand U11407 (N_11407,N_7200,N_7631);
nor U11408 (N_11408,N_6788,N_7362);
nand U11409 (N_11409,N_7426,N_7192);
or U11410 (N_11410,N_7397,N_8298);
or U11411 (N_11411,N_6038,N_7052);
and U11412 (N_11412,N_8995,N_6267);
nor U11413 (N_11413,N_7249,N_7357);
or U11414 (N_11414,N_6758,N_8008);
and U11415 (N_11415,N_7612,N_7184);
xor U11416 (N_11416,N_7571,N_8938);
nand U11417 (N_11417,N_7073,N_6966);
xor U11418 (N_11418,N_7697,N_7778);
nor U11419 (N_11419,N_6771,N_7024);
nand U11420 (N_11420,N_6855,N_6951);
and U11421 (N_11421,N_8947,N_6943);
or U11422 (N_11422,N_7277,N_8498);
nand U11423 (N_11423,N_8516,N_7811);
and U11424 (N_11424,N_6724,N_6593);
and U11425 (N_11425,N_6827,N_6218);
xor U11426 (N_11426,N_7129,N_6272);
nor U11427 (N_11427,N_6361,N_8097);
nand U11428 (N_11428,N_8456,N_6607);
nand U11429 (N_11429,N_8917,N_8290);
nand U11430 (N_11430,N_6266,N_7581);
nand U11431 (N_11431,N_6890,N_6981);
nor U11432 (N_11432,N_6917,N_6879);
or U11433 (N_11433,N_8663,N_8967);
nor U11434 (N_11434,N_7004,N_8704);
or U11435 (N_11435,N_8805,N_8621);
nand U11436 (N_11436,N_6320,N_6359);
nor U11437 (N_11437,N_7097,N_7252);
nor U11438 (N_11438,N_7312,N_6117);
nand U11439 (N_11439,N_7708,N_8310);
or U11440 (N_11440,N_7983,N_8376);
or U11441 (N_11441,N_6474,N_8543);
or U11442 (N_11442,N_7024,N_6365);
nand U11443 (N_11443,N_7484,N_8706);
nor U11444 (N_11444,N_8704,N_6350);
nor U11445 (N_11445,N_8476,N_8814);
or U11446 (N_11446,N_7091,N_6022);
xor U11447 (N_11447,N_7793,N_6912);
nor U11448 (N_11448,N_7578,N_7396);
and U11449 (N_11449,N_7871,N_8931);
nand U11450 (N_11450,N_7477,N_7877);
nor U11451 (N_11451,N_8038,N_7843);
xor U11452 (N_11452,N_7529,N_7640);
or U11453 (N_11453,N_6870,N_6046);
nor U11454 (N_11454,N_6548,N_8401);
and U11455 (N_11455,N_8437,N_7786);
xnor U11456 (N_11456,N_8511,N_7082);
nand U11457 (N_11457,N_8359,N_7631);
and U11458 (N_11458,N_8457,N_6180);
or U11459 (N_11459,N_8151,N_7087);
xnor U11460 (N_11460,N_8856,N_7919);
xor U11461 (N_11461,N_8469,N_8427);
and U11462 (N_11462,N_6535,N_8108);
nand U11463 (N_11463,N_6459,N_8415);
and U11464 (N_11464,N_6980,N_6889);
nand U11465 (N_11465,N_6024,N_7263);
and U11466 (N_11466,N_7239,N_8935);
or U11467 (N_11467,N_7580,N_8246);
nand U11468 (N_11468,N_7478,N_7971);
or U11469 (N_11469,N_8038,N_7289);
or U11470 (N_11470,N_8421,N_7416);
and U11471 (N_11471,N_7911,N_7230);
or U11472 (N_11472,N_8884,N_8911);
or U11473 (N_11473,N_7762,N_7923);
and U11474 (N_11474,N_6996,N_8162);
and U11475 (N_11475,N_7890,N_6083);
xnor U11476 (N_11476,N_7825,N_8947);
or U11477 (N_11477,N_8035,N_8990);
or U11478 (N_11478,N_6578,N_7602);
and U11479 (N_11479,N_7881,N_7447);
nand U11480 (N_11480,N_7048,N_8878);
nand U11481 (N_11481,N_7959,N_7203);
nand U11482 (N_11482,N_6537,N_6597);
xnor U11483 (N_11483,N_6982,N_8737);
nor U11484 (N_11484,N_7953,N_7471);
xnor U11485 (N_11485,N_6242,N_8469);
nand U11486 (N_11486,N_8455,N_7015);
or U11487 (N_11487,N_6690,N_8856);
nor U11488 (N_11488,N_6050,N_7661);
xnor U11489 (N_11489,N_8861,N_6097);
nand U11490 (N_11490,N_7630,N_8177);
and U11491 (N_11491,N_8628,N_7402);
xor U11492 (N_11492,N_8019,N_8627);
nor U11493 (N_11493,N_6404,N_8755);
and U11494 (N_11494,N_7867,N_8279);
and U11495 (N_11495,N_7962,N_8962);
nand U11496 (N_11496,N_6121,N_8129);
nor U11497 (N_11497,N_7238,N_8610);
nand U11498 (N_11498,N_6234,N_7201);
and U11499 (N_11499,N_6939,N_6270);
or U11500 (N_11500,N_7978,N_7933);
or U11501 (N_11501,N_6398,N_6764);
or U11502 (N_11502,N_6170,N_6495);
and U11503 (N_11503,N_6898,N_6336);
and U11504 (N_11504,N_8104,N_7189);
nand U11505 (N_11505,N_7967,N_8836);
or U11506 (N_11506,N_7995,N_6501);
nand U11507 (N_11507,N_7554,N_8152);
nor U11508 (N_11508,N_8286,N_8343);
or U11509 (N_11509,N_8837,N_7961);
nor U11510 (N_11510,N_7604,N_6411);
and U11511 (N_11511,N_7935,N_8912);
or U11512 (N_11512,N_8984,N_6781);
nand U11513 (N_11513,N_8793,N_7974);
or U11514 (N_11514,N_8783,N_7550);
or U11515 (N_11515,N_6128,N_6688);
or U11516 (N_11516,N_8599,N_6305);
nor U11517 (N_11517,N_8828,N_8587);
and U11518 (N_11518,N_7856,N_7528);
nor U11519 (N_11519,N_6101,N_8551);
nor U11520 (N_11520,N_6223,N_6213);
or U11521 (N_11521,N_8183,N_6597);
or U11522 (N_11522,N_8579,N_8046);
xnor U11523 (N_11523,N_6689,N_6873);
and U11524 (N_11524,N_8102,N_6626);
xnor U11525 (N_11525,N_6425,N_7893);
and U11526 (N_11526,N_7143,N_6658);
nor U11527 (N_11527,N_7730,N_7522);
and U11528 (N_11528,N_7015,N_6713);
xor U11529 (N_11529,N_7382,N_6269);
nor U11530 (N_11530,N_7609,N_8561);
and U11531 (N_11531,N_7371,N_8035);
or U11532 (N_11532,N_8543,N_7316);
and U11533 (N_11533,N_6201,N_7979);
and U11534 (N_11534,N_7576,N_6933);
nor U11535 (N_11535,N_8461,N_7143);
xor U11536 (N_11536,N_7625,N_8441);
or U11537 (N_11537,N_8239,N_7072);
and U11538 (N_11538,N_6043,N_6376);
nand U11539 (N_11539,N_8106,N_6381);
xnor U11540 (N_11540,N_6329,N_7670);
xor U11541 (N_11541,N_8424,N_8734);
xor U11542 (N_11542,N_7199,N_6701);
nand U11543 (N_11543,N_6636,N_6062);
xor U11544 (N_11544,N_8109,N_7747);
nor U11545 (N_11545,N_6822,N_8245);
or U11546 (N_11546,N_8165,N_7381);
xor U11547 (N_11547,N_7862,N_6176);
and U11548 (N_11548,N_7509,N_6018);
and U11549 (N_11549,N_8396,N_6780);
nor U11550 (N_11550,N_8380,N_6842);
and U11551 (N_11551,N_8923,N_7879);
nor U11552 (N_11552,N_6452,N_7084);
nand U11553 (N_11553,N_7229,N_8215);
xor U11554 (N_11554,N_7864,N_8173);
nor U11555 (N_11555,N_7818,N_8015);
nor U11556 (N_11556,N_8579,N_8578);
or U11557 (N_11557,N_6245,N_8939);
xnor U11558 (N_11558,N_6595,N_8705);
xor U11559 (N_11559,N_6599,N_8453);
nor U11560 (N_11560,N_7868,N_8478);
nand U11561 (N_11561,N_7298,N_8795);
nor U11562 (N_11562,N_6552,N_7516);
and U11563 (N_11563,N_7547,N_6687);
or U11564 (N_11564,N_7123,N_8709);
or U11565 (N_11565,N_6886,N_7294);
xnor U11566 (N_11566,N_6003,N_7029);
xnor U11567 (N_11567,N_7204,N_6118);
or U11568 (N_11568,N_7777,N_7699);
nor U11569 (N_11569,N_8150,N_7676);
nor U11570 (N_11570,N_6036,N_7021);
and U11571 (N_11571,N_8788,N_7357);
nor U11572 (N_11572,N_8238,N_8079);
or U11573 (N_11573,N_8289,N_6582);
xor U11574 (N_11574,N_7466,N_8735);
and U11575 (N_11575,N_8567,N_8047);
nor U11576 (N_11576,N_7434,N_7737);
and U11577 (N_11577,N_8623,N_7443);
nand U11578 (N_11578,N_8285,N_6905);
nor U11579 (N_11579,N_6478,N_8065);
nand U11580 (N_11580,N_7773,N_7342);
nor U11581 (N_11581,N_8082,N_8736);
xor U11582 (N_11582,N_8505,N_7710);
xor U11583 (N_11583,N_8040,N_7728);
and U11584 (N_11584,N_7170,N_7993);
or U11585 (N_11585,N_8587,N_7387);
nand U11586 (N_11586,N_7752,N_6141);
xnor U11587 (N_11587,N_8201,N_7149);
nand U11588 (N_11588,N_8995,N_7217);
xor U11589 (N_11589,N_8824,N_8444);
nand U11590 (N_11590,N_6666,N_8899);
xor U11591 (N_11591,N_7998,N_7768);
or U11592 (N_11592,N_8171,N_6329);
and U11593 (N_11593,N_6042,N_8102);
nand U11594 (N_11594,N_6653,N_8886);
nand U11595 (N_11595,N_6483,N_6484);
xor U11596 (N_11596,N_8912,N_8051);
or U11597 (N_11597,N_6054,N_8783);
or U11598 (N_11598,N_7106,N_8135);
xor U11599 (N_11599,N_6218,N_8975);
or U11600 (N_11600,N_7321,N_6393);
nand U11601 (N_11601,N_7654,N_8721);
nand U11602 (N_11602,N_8497,N_6185);
or U11603 (N_11603,N_6898,N_7738);
or U11604 (N_11604,N_8549,N_6666);
nor U11605 (N_11605,N_6194,N_7493);
or U11606 (N_11606,N_8039,N_7569);
xor U11607 (N_11607,N_7000,N_7787);
xnor U11608 (N_11608,N_7834,N_6070);
nor U11609 (N_11609,N_8950,N_7518);
nor U11610 (N_11610,N_7423,N_6493);
nor U11611 (N_11611,N_7401,N_7456);
nand U11612 (N_11612,N_8818,N_6189);
nor U11613 (N_11613,N_6421,N_7659);
and U11614 (N_11614,N_8419,N_8012);
xnor U11615 (N_11615,N_6664,N_6119);
nor U11616 (N_11616,N_7854,N_8906);
or U11617 (N_11617,N_7588,N_6867);
nor U11618 (N_11618,N_8147,N_8556);
nor U11619 (N_11619,N_7182,N_7496);
nand U11620 (N_11620,N_6076,N_8316);
nand U11621 (N_11621,N_7528,N_8253);
and U11622 (N_11622,N_6857,N_7879);
xnor U11623 (N_11623,N_7694,N_7390);
or U11624 (N_11624,N_6319,N_8496);
xor U11625 (N_11625,N_6394,N_6815);
nor U11626 (N_11626,N_8946,N_6321);
xor U11627 (N_11627,N_7777,N_6387);
nand U11628 (N_11628,N_7255,N_7431);
nor U11629 (N_11629,N_8300,N_6219);
nand U11630 (N_11630,N_6841,N_6260);
nor U11631 (N_11631,N_7328,N_8387);
nand U11632 (N_11632,N_8336,N_6693);
or U11633 (N_11633,N_6153,N_6607);
or U11634 (N_11634,N_6434,N_8724);
nand U11635 (N_11635,N_8741,N_8833);
or U11636 (N_11636,N_6097,N_6477);
and U11637 (N_11637,N_7219,N_8806);
nor U11638 (N_11638,N_6500,N_6242);
nor U11639 (N_11639,N_6615,N_7674);
and U11640 (N_11640,N_7951,N_7906);
or U11641 (N_11641,N_8321,N_8865);
xor U11642 (N_11642,N_7096,N_8384);
xor U11643 (N_11643,N_7400,N_6038);
or U11644 (N_11644,N_7460,N_7303);
or U11645 (N_11645,N_6667,N_8086);
or U11646 (N_11646,N_8800,N_8490);
or U11647 (N_11647,N_7118,N_8073);
nand U11648 (N_11648,N_6728,N_8897);
nand U11649 (N_11649,N_6311,N_8627);
nand U11650 (N_11650,N_6967,N_6121);
nand U11651 (N_11651,N_6553,N_8907);
nand U11652 (N_11652,N_7645,N_7350);
nand U11653 (N_11653,N_6782,N_7457);
and U11654 (N_11654,N_7198,N_8047);
or U11655 (N_11655,N_8193,N_8578);
or U11656 (N_11656,N_6760,N_6134);
or U11657 (N_11657,N_8456,N_8304);
nand U11658 (N_11658,N_6791,N_6607);
and U11659 (N_11659,N_6417,N_6680);
or U11660 (N_11660,N_7726,N_8207);
and U11661 (N_11661,N_8898,N_8563);
or U11662 (N_11662,N_8123,N_8576);
or U11663 (N_11663,N_8781,N_8907);
nor U11664 (N_11664,N_6900,N_7203);
xnor U11665 (N_11665,N_6349,N_8248);
and U11666 (N_11666,N_8453,N_8302);
nand U11667 (N_11667,N_6119,N_6415);
nor U11668 (N_11668,N_8693,N_6197);
nand U11669 (N_11669,N_6170,N_8316);
nand U11670 (N_11670,N_8037,N_7395);
or U11671 (N_11671,N_7713,N_8998);
and U11672 (N_11672,N_7588,N_6816);
or U11673 (N_11673,N_7658,N_7667);
and U11674 (N_11674,N_6579,N_7252);
nor U11675 (N_11675,N_8023,N_8028);
nor U11676 (N_11676,N_8385,N_7728);
or U11677 (N_11677,N_7863,N_7206);
xnor U11678 (N_11678,N_6405,N_6593);
xor U11679 (N_11679,N_8893,N_8845);
or U11680 (N_11680,N_7186,N_6963);
and U11681 (N_11681,N_7757,N_7355);
nand U11682 (N_11682,N_6680,N_8359);
and U11683 (N_11683,N_8058,N_7678);
nand U11684 (N_11684,N_8366,N_8245);
or U11685 (N_11685,N_6996,N_6631);
xor U11686 (N_11686,N_7169,N_8689);
xor U11687 (N_11687,N_6153,N_8751);
nor U11688 (N_11688,N_7678,N_6313);
xor U11689 (N_11689,N_7973,N_7235);
xor U11690 (N_11690,N_6247,N_7767);
nor U11691 (N_11691,N_7001,N_6983);
xnor U11692 (N_11692,N_6562,N_6122);
or U11693 (N_11693,N_6414,N_7129);
nor U11694 (N_11694,N_6268,N_8881);
xnor U11695 (N_11695,N_6345,N_7413);
xnor U11696 (N_11696,N_6162,N_7270);
xnor U11697 (N_11697,N_6814,N_7586);
nand U11698 (N_11698,N_6055,N_7457);
nand U11699 (N_11699,N_6962,N_6713);
and U11700 (N_11700,N_7077,N_7560);
and U11701 (N_11701,N_7045,N_6328);
and U11702 (N_11702,N_6916,N_6482);
nand U11703 (N_11703,N_8556,N_7296);
xor U11704 (N_11704,N_7322,N_6234);
nand U11705 (N_11705,N_6405,N_8345);
and U11706 (N_11706,N_6177,N_7294);
nand U11707 (N_11707,N_6178,N_6419);
and U11708 (N_11708,N_6564,N_7618);
and U11709 (N_11709,N_8850,N_6972);
or U11710 (N_11710,N_6851,N_8198);
nand U11711 (N_11711,N_7360,N_7253);
xnor U11712 (N_11712,N_6408,N_7769);
and U11713 (N_11713,N_7811,N_8155);
xor U11714 (N_11714,N_7035,N_6726);
nor U11715 (N_11715,N_7789,N_8888);
nand U11716 (N_11716,N_6956,N_7562);
xnor U11717 (N_11717,N_7680,N_6374);
nor U11718 (N_11718,N_7866,N_8214);
nand U11719 (N_11719,N_7657,N_8474);
and U11720 (N_11720,N_7745,N_8806);
nand U11721 (N_11721,N_7556,N_6323);
xnor U11722 (N_11722,N_6629,N_6236);
nor U11723 (N_11723,N_8842,N_6858);
nor U11724 (N_11724,N_6455,N_6951);
and U11725 (N_11725,N_6378,N_6283);
and U11726 (N_11726,N_6583,N_7680);
or U11727 (N_11727,N_7953,N_8596);
nor U11728 (N_11728,N_8514,N_7021);
and U11729 (N_11729,N_7430,N_6870);
and U11730 (N_11730,N_7702,N_7350);
nor U11731 (N_11731,N_6391,N_6620);
nand U11732 (N_11732,N_6849,N_8730);
nor U11733 (N_11733,N_8272,N_7241);
xor U11734 (N_11734,N_8104,N_7984);
nor U11735 (N_11735,N_8800,N_7560);
and U11736 (N_11736,N_6991,N_6348);
or U11737 (N_11737,N_6944,N_8576);
and U11738 (N_11738,N_6173,N_6022);
nand U11739 (N_11739,N_7572,N_7985);
nand U11740 (N_11740,N_6656,N_8950);
nand U11741 (N_11741,N_6338,N_6627);
xnor U11742 (N_11742,N_7243,N_7083);
nor U11743 (N_11743,N_6737,N_6728);
nor U11744 (N_11744,N_6040,N_7249);
or U11745 (N_11745,N_7798,N_7768);
xor U11746 (N_11746,N_8124,N_6042);
nor U11747 (N_11747,N_8586,N_8432);
or U11748 (N_11748,N_7593,N_8658);
xor U11749 (N_11749,N_7042,N_7895);
nand U11750 (N_11750,N_8881,N_7327);
and U11751 (N_11751,N_7839,N_8064);
nor U11752 (N_11752,N_7653,N_6444);
nand U11753 (N_11753,N_7425,N_8501);
nand U11754 (N_11754,N_8746,N_7403);
nand U11755 (N_11755,N_8640,N_6888);
and U11756 (N_11756,N_8350,N_8823);
nor U11757 (N_11757,N_8125,N_7779);
nor U11758 (N_11758,N_8165,N_6009);
xnor U11759 (N_11759,N_7254,N_8133);
nor U11760 (N_11760,N_7824,N_6675);
nand U11761 (N_11761,N_8224,N_8421);
nor U11762 (N_11762,N_7646,N_7474);
xnor U11763 (N_11763,N_8604,N_8740);
or U11764 (N_11764,N_6618,N_6293);
nor U11765 (N_11765,N_7188,N_6193);
and U11766 (N_11766,N_6962,N_7046);
nor U11767 (N_11767,N_7400,N_6142);
nand U11768 (N_11768,N_8440,N_7147);
or U11769 (N_11769,N_8773,N_8256);
nor U11770 (N_11770,N_8572,N_8699);
nand U11771 (N_11771,N_7846,N_6055);
nand U11772 (N_11772,N_6773,N_6858);
nor U11773 (N_11773,N_7018,N_7849);
or U11774 (N_11774,N_7040,N_7170);
and U11775 (N_11775,N_7452,N_8182);
and U11776 (N_11776,N_6752,N_6116);
nor U11777 (N_11777,N_8571,N_6628);
or U11778 (N_11778,N_6107,N_8090);
nor U11779 (N_11779,N_6291,N_7869);
and U11780 (N_11780,N_6962,N_6927);
or U11781 (N_11781,N_7101,N_6859);
xnor U11782 (N_11782,N_7103,N_6322);
or U11783 (N_11783,N_7871,N_6691);
nand U11784 (N_11784,N_8599,N_6621);
nand U11785 (N_11785,N_8260,N_6320);
and U11786 (N_11786,N_6113,N_7250);
nand U11787 (N_11787,N_7608,N_7911);
and U11788 (N_11788,N_7733,N_7051);
xnor U11789 (N_11789,N_6061,N_7462);
or U11790 (N_11790,N_7522,N_6600);
nand U11791 (N_11791,N_8951,N_8688);
nand U11792 (N_11792,N_6700,N_8832);
nand U11793 (N_11793,N_6807,N_8304);
xor U11794 (N_11794,N_7424,N_7296);
nor U11795 (N_11795,N_8410,N_8987);
xor U11796 (N_11796,N_6027,N_7949);
nand U11797 (N_11797,N_6325,N_6362);
nand U11798 (N_11798,N_6086,N_7000);
and U11799 (N_11799,N_7818,N_7634);
and U11800 (N_11800,N_6649,N_8895);
xnor U11801 (N_11801,N_7513,N_7335);
and U11802 (N_11802,N_8665,N_6086);
nor U11803 (N_11803,N_6707,N_8550);
or U11804 (N_11804,N_7652,N_8348);
nor U11805 (N_11805,N_7901,N_6107);
nand U11806 (N_11806,N_7098,N_6282);
or U11807 (N_11807,N_6616,N_6855);
nand U11808 (N_11808,N_6702,N_7118);
nor U11809 (N_11809,N_8585,N_8616);
nand U11810 (N_11810,N_7013,N_6885);
or U11811 (N_11811,N_7761,N_8580);
or U11812 (N_11812,N_6585,N_6996);
or U11813 (N_11813,N_8746,N_6715);
xor U11814 (N_11814,N_7468,N_7278);
xnor U11815 (N_11815,N_6931,N_6575);
and U11816 (N_11816,N_7025,N_8274);
nor U11817 (N_11817,N_6105,N_7489);
and U11818 (N_11818,N_6608,N_7249);
and U11819 (N_11819,N_8605,N_6725);
xnor U11820 (N_11820,N_8782,N_7824);
and U11821 (N_11821,N_6751,N_8828);
or U11822 (N_11822,N_8461,N_6606);
or U11823 (N_11823,N_8154,N_8610);
and U11824 (N_11824,N_7542,N_7166);
nor U11825 (N_11825,N_7360,N_8301);
nand U11826 (N_11826,N_8180,N_8394);
nand U11827 (N_11827,N_6374,N_8130);
and U11828 (N_11828,N_6961,N_6601);
nand U11829 (N_11829,N_7404,N_7376);
xnor U11830 (N_11830,N_7967,N_8683);
nor U11831 (N_11831,N_8579,N_7005);
xor U11832 (N_11832,N_8474,N_6164);
nand U11833 (N_11833,N_7803,N_7376);
and U11834 (N_11834,N_8524,N_7983);
nor U11835 (N_11835,N_8712,N_8485);
xor U11836 (N_11836,N_8312,N_8113);
xnor U11837 (N_11837,N_7614,N_6394);
and U11838 (N_11838,N_8286,N_7035);
and U11839 (N_11839,N_7278,N_8306);
and U11840 (N_11840,N_6113,N_6692);
xor U11841 (N_11841,N_8034,N_6545);
and U11842 (N_11842,N_7628,N_7824);
and U11843 (N_11843,N_6881,N_8337);
and U11844 (N_11844,N_7835,N_7765);
or U11845 (N_11845,N_7617,N_7449);
nor U11846 (N_11846,N_7835,N_7490);
and U11847 (N_11847,N_8769,N_8819);
and U11848 (N_11848,N_6439,N_7690);
and U11849 (N_11849,N_8143,N_6893);
and U11850 (N_11850,N_8857,N_7480);
nor U11851 (N_11851,N_8672,N_6125);
and U11852 (N_11852,N_6841,N_6012);
or U11853 (N_11853,N_6345,N_6348);
nand U11854 (N_11854,N_7317,N_6951);
xor U11855 (N_11855,N_8831,N_8055);
xor U11856 (N_11856,N_7579,N_7921);
or U11857 (N_11857,N_6699,N_7650);
or U11858 (N_11858,N_8327,N_8980);
or U11859 (N_11859,N_6906,N_7939);
xnor U11860 (N_11860,N_6055,N_7006);
or U11861 (N_11861,N_8787,N_6582);
nor U11862 (N_11862,N_8542,N_6210);
nor U11863 (N_11863,N_8289,N_8668);
or U11864 (N_11864,N_7374,N_7573);
and U11865 (N_11865,N_7718,N_7186);
and U11866 (N_11866,N_8009,N_6410);
nor U11867 (N_11867,N_7906,N_6939);
nor U11868 (N_11868,N_8584,N_8969);
nor U11869 (N_11869,N_7215,N_7812);
and U11870 (N_11870,N_7533,N_6867);
nand U11871 (N_11871,N_8162,N_6089);
nand U11872 (N_11872,N_7101,N_8323);
or U11873 (N_11873,N_7111,N_8023);
and U11874 (N_11874,N_6230,N_8440);
nand U11875 (N_11875,N_8522,N_7461);
and U11876 (N_11876,N_8729,N_6719);
or U11877 (N_11877,N_8403,N_7100);
or U11878 (N_11878,N_8098,N_7624);
and U11879 (N_11879,N_7740,N_8453);
nor U11880 (N_11880,N_8881,N_8343);
or U11881 (N_11881,N_7927,N_8842);
xnor U11882 (N_11882,N_6885,N_7123);
and U11883 (N_11883,N_6280,N_7899);
and U11884 (N_11884,N_6840,N_6934);
and U11885 (N_11885,N_8624,N_7695);
and U11886 (N_11886,N_7565,N_6685);
xnor U11887 (N_11887,N_8041,N_6390);
nand U11888 (N_11888,N_7606,N_8998);
nand U11889 (N_11889,N_8718,N_8800);
nor U11890 (N_11890,N_7736,N_7065);
nor U11891 (N_11891,N_8504,N_7584);
and U11892 (N_11892,N_6988,N_7158);
and U11893 (N_11893,N_7537,N_7151);
xor U11894 (N_11894,N_6182,N_8629);
and U11895 (N_11895,N_7665,N_7237);
and U11896 (N_11896,N_7649,N_7354);
nand U11897 (N_11897,N_6656,N_7447);
nor U11898 (N_11898,N_7372,N_8749);
and U11899 (N_11899,N_6360,N_7425);
nand U11900 (N_11900,N_8089,N_6183);
nor U11901 (N_11901,N_8850,N_6729);
xnor U11902 (N_11902,N_7463,N_6276);
and U11903 (N_11903,N_8505,N_8314);
or U11904 (N_11904,N_6686,N_7933);
or U11905 (N_11905,N_7964,N_7423);
xnor U11906 (N_11906,N_7544,N_6947);
and U11907 (N_11907,N_8078,N_8426);
or U11908 (N_11908,N_8240,N_8452);
and U11909 (N_11909,N_8608,N_6676);
nand U11910 (N_11910,N_8802,N_6648);
xnor U11911 (N_11911,N_6607,N_7267);
xnor U11912 (N_11912,N_8860,N_6054);
xor U11913 (N_11913,N_8207,N_7504);
nand U11914 (N_11914,N_8076,N_8550);
nor U11915 (N_11915,N_7507,N_8028);
or U11916 (N_11916,N_8760,N_8787);
and U11917 (N_11917,N_6264,N_8607);
nand U11918 (N_11918,N_7607,N_6606);
and U11919 (N_11919,N_6566,N_8768);
nand U11920 (N_11920,N_8375,N_6927);
nor U11921 (N_11921,N_8294,N_6282);
nor U11922 (N_11922,N_6607,N_6445);
nor U11923 (N_11923,N_7684,N_6774);
nand U11924 (N_11924,N_7441,N_6455);
or U11925 (N_11925,N_7012,N_7507);
or U11926 (N_11926,N_7988,N_8409);
nand U11927 (N_11927,N_6513,N_7978);
nor U11928 (N_11928,N_7155,N_6005);
and U11929 (N_11929,N_7902,N_6121);
and U11930 (N_11930,N_7967,N_7832);
xnor U11931 (N_11931,N_6697,N_8371);
nand U11932 (N_11932,N_6534,N_6317);
nand U11933 (N_11933,N_6516,N_8502);
nor U11934 (N_11934,N_6454,N_8064);
nand U11935 (N_11935,N_8459,N_7511);
xnor U11936 (N_11936,N_7183,N_6093);
nor U11937 (N_11937,N_7750,N_8844);
nand U11938 (N_11938,N_7753,N_7971);
nand U11939 (N_11939,N_7590,N_8871);
and U11940 (N_11940,N_8085,N_6595);
nor U11941 (N_11941,N_8312,N_7096);
nor U11942 (N_11942,N_6631,N_8703);
xor U11943 (N_11943,N_6538,N_6574);
nor U11944 (N_11944,N_6131,N_7909);
xor U11945 (N_11945,N_6784,N_6079);
xnor U11946 (N_11946,N_8451,N_8055);
or U11947 (N_11947,N_6754,N_7167);
or U11948 (N_11948,N_8160,N_8556);
nor U11949 (N_11949,N_7186,N_7561);
and U11950 (N_11950,N_7945,N_7783);
nor U11951 (N_11951,N_8006,N_8206);
and U11952 (N_11952,N_8217,N_8024);
xor U11953 (N_11953,N_6324,N_6257);
xor U11954 (N_11954,N_7437,N_7148);
nor U11955 (N_11955,N_7786,N_8739);
xnor U11956 (N_11956,N_8964,N_8113);
nor U11957 (N_11957,N_7511,N_6955);
xnor U11958 (N_11958,N_6987,N_6968);
nand U11959 (N_11959,N_7357,N_6091);
or U11960 (N_11960,N_8035,N_7615);
and U11961 (N_11961,N_6802,N_7984);
xor U11962 (N_11962,N_7809,N_8155);
nor U11963 (N_11963,N_7348,N_8885);
nand U11964 (N_11964,N_8568,N_7124);
xnor U11965 (N_11965,N_6651,N_8966);
nand U11966 (N_11966,N_8334,N_6157);
and U11967 (N_11967,N_8790,N_6152);
nor U11968 (N_11968,N_6152,N_8811);
and U11969 (N_11969,N_8072,N_6107);
nor U11970 (N_11970,N_7398,N_6551);
and U11971 (N_11971,N_6568,N_6899);
xor U11972 (N_11972,N_6543,N_7383);
nor U11973 (N_11973,N_7690,N_6487);
or U11974 (N_11974,N_6663,N_8645);
and U11975 (N_11975,N_6042,N_8014);
nor U11976 (N_11976,N_7174,N_7644);
and U11977 (N_11977,N_8284,N_6481);
xor U11978 (N_11978,N_8531,N_8723);
and U11979 (N_11979,N_6380,N_6376);
nand U11980 (N_11980,N_8669,N_6323);
nor U11981 (N_11981,N_6312,N_6437);
and U11982 (N_11982,N_6037,N_6982);
nand U11983 (N_11983,N_7642,N_7122);
nand U11984 (N_11984,N_7227,N_6789);
or U11985 (N_11985,N_8778,N_8639);
or U11986 (N_11986,N_8684,N_8746);
nor U11987 (N_11987,N_8026,N_8708);
or U11988 (N_11988,N_7925,N_7203);
xor U11989 (N_11989,N_7027,N_6265);
and U11990 (N_11990,N_8566,N_7187);
nand U11991 (N_11991,N_8197,N_6355);
nor U11992 (N_11992,N_6612,N_7413);
nand U11993 (N_11993,N_7780,N_8512);
nand U11994 (N_11994,N_8972,N_6185);
xnor U11995 (N_11995,N_7561,N_7562);
nor U11996 (N_11996,N_6130,N_6520);
xor U11997 (N_11997,N_8856,N_8189);
nand U11998 (N_11998,N_8589,N_7691);
nand U11999 (N_11999,N_7099,N_8669);
and U12000 (N_12000,N_11467,N_10015);
xnor U12001 (N_12001,N_9001,N_10372);
or U12002 (N_12002,N_10917,N_10859);
xnor U12003 (N_12003,N_9889,N_9990);
nand U12004 (N_12004,N_11834,N_10121);
and U12005 (N_12005,N_9378,N_9672);
and U12006 (N_12006,N_9955,N_9466);
xnor U12007 (N_12007,N_9345,N_10415);
xor U12008 (N_12008,N_11179,N_11968);
nand U12009 (N_12009,N_11570,N_11476);
and U12010 (N_12010,N_10804,N_9209);
nor U12011 (N_12011,N_11639,N_9047);
or U12012 (N_12012,N_10697,N_10484);
or U12013 (N_12013,N_9764,N_10167);
nor U12014 (N_12014,N_9381,N_9374);
nand U12015 (N_12015,N_10950,N_9389);
nand U12016 (N_12016,N_10647,N_9654);
nand U12017 (N_12017,N_10665,N_11816);
nor U12018 (N_12018,N_11805,N_11128);
nor U12019 (N_12019,N_10151,N_9807);
xnor U12020 (N_12020,N_9846,N_11122);
nand U12021 (N_12021,N_10906,N_10456);
nand U12022 (N_12022,N_10937,N_9835);
xnor U12023 (N_12023,N_9030,N_11607);
nand U12024 (N_12024,N_9340,N_9747);
nand U12025 (N_12025,N_10867,N_9973);
or U12026 (N_12026,N_11771,N_10518);
nand U12027 (N_12027,N_11546,N_9546);
and U12028 (N_12028,N_11407,N_10050);
xor U12029 (N_12029,N_11691,N_9981);
nor U12030 (N_12030,N_9800,N_9709);
nand U12031 (N_12031,N_10000,N_11398);
nor U12032 (N_12032,N_10754,N_11117);
nand U12033 (N_12033,N_10265,N_11431);
nor U12034 (N_12034,N_9786,N_9867);
nor U12035 (N_12035,N_9490,N_9772);
or U12036 (N_12036,N_10190,N_10694);
or U12037 (N_12037,N_9945,N_10542);
nor U12038 (N_12038,N_10721,N_9142);
xor U12039 (N_12039,N_11698,N_11384);
or U12040 (N_12040,N_11520,N_11049);
nor U12041 (N_12041,N_11202,N_9127);
and U12042 (N_12042,N_9149,N_9681);
nor U12043 (N_12043,N_9545,N_11770);
or U12044 (N_12044,N_11421,N_11291);
nor U12045 (N_12045,N_11809,N_11586);
nand U12046 (N_12046,N_11230,N_11264);
xor U12047 (N_12047,N_11674,N_10091);
xor U12048 (N_12048,N_11950,N_9716);
and U12049 (N_12049,N_9177,N_9458);
nand U12050 (N_12050,N_9925,N_10898);
or U12051 (N_12051,N_11859,N_9262);
xnor U12052 (N_12052,N_11455,N_9088);
nand U12053 (N_12053,N_10349,N_11211);
xnor U12054 (N_12054,N_9424,N_9985);
nand U12055 (N_12055,N_9691,N_10334);
nor U12056 (N_12056,N_11312,N_11944);
xor U12057 (N_12057,N_10954,N_9791);
nor U12058 (N_12058,N_11796,N_11763);
nor U12059 (N_12059,N_9794,N_11108);
nor U12060 (N_12060,N_9021,N_9937);
and U12061 (N_12061,N_9708,N_11166);
nor U12062 (N_12062,N_9726,N_9443);
or U12063 (N_12063,N_11051,N_9022);
nand U12064 (N_12064,N_10820,N_9168);
xnor U12065 (N_12065,N_11373,N_9805);
nor U12066 (N_12066,N_10703,N_10828);
and U12067 (N_12067,N_9926,N_11335);
nor U12068 (N_12068,N_9015,N_11995);
nand U12069 (N_12069,N_11572,N_9317);
and U12070 (N_12070,N_11256,N_10182);
and U12071 (N_12071,N_9983,N_9268);
or U12072 (N_12072,N_10180,N_9701);
xnor U12073 (N_12073,N_10538,N_9840);
nor U12074 (N_12074,N_9178,N_11651);
xor U12075 (N_12075,N_10245,N_9230);
or U12076 (N_12076,N_11487,N_11239);
nand U12077 (N_12077,N_11736,N_10511);
nand U12078 (N_12078,N_10037,N_10631);
or U12079 (N_12079,N_10900,N_10239);
xor U12080 (N_12080,N_11194,N_11890);
or U12081 (N_12081,N_11257,N_11189);
or U12082 (N_12082,N_9774,N_10499);
nor U12083 (N_12083,N_10939,N_9175);
and U12084 (N_12084,N_11134,N_10202);
and U12085 (N_12085,N_11743,N_9765);
xor U12086 (N_12086,N_10895,N_11503);
nand U12087 (N_12087,N_11186,N_11522);
xnor U12088 (N_12088,N_11083,N_10025);
xor U12089 (N_12089,N_11430,N_9660);
and U12090 (N_12090,N_10548,N_11088);
or U12091 (N_12091,N_11009,N_11196);
nor U12092 (N_12092,N_9481,N_10213);
nor U12093 (N_12093,N_9941,N_11368);
or U12094 (N_12094,N_11259,N_9834);
nand U12095 (N_12095,N_10248,N_11285);
and U12096 (N_12096,N_11434,N_9690);
nand U12097 (N_12097,N_11016,N_9287);
or U12098 (N_12098,N_11830,N_10640);
nand U12099 (N_12099,N_9721,N_10159);
and U12100 (N_12100,N_9161,N_11680);
nand U12101 (N_12101,N_9741,N_10814);
and U12102 (N_12102,N_9806,N_9913);
nand U12103 (N_12103,N_10191,N_11638);
nor U12104 (N_12104,N_9853,N_10892);
nor U12105 (N_12105,N_10930,N_11375);
or U12106 (N_12106,N_10108,N_10829);
or U12107 (N_12107,N_11634,N_11420);
nand U12108 (N_12108,N_9606,N_9563);
or U12109 (N_12109,N_9787,N_9705);
nand U12110 (N_12110,N_9566,N_9877);
and U12111 (N_12111,N_10018,N_10357);
xnor U12112 (N_12112,N_9244,N_10552);
and U12113 (N_12113,N_10735,N_11273);
and U12114 (N_12114,N_11404,N_11824);
and U12115 (N_12115,N_9583,N_9947);
nand U12116 (N_12116,N_11185,N_9938);
xnor U12117 (N_12117,N_11506,N_10581);
and U12118 (N_12118,N_11329,N_10212);
xnor U12119 (N_12119,N_9222,N_9608);
xor U12120 (N_12120,N_10510,N_9676);
nand U12121 (N_12121,N_9232,N_9811);
and U12122 (N_12122,N_11881,N_11443);
xnor U12123 (N_12123,N_11954,N_10064);
or U12124 (N_12124,N_9026,N_11820);
or U12125 (N_12125,N_9152,N_9748);
nand U12126 (N_12126,N_11249,N_10026);
xnor U12127 (N_12127,N_10772,N_10262);
and U12128 (N_12128,N_10641,N_9313);
or U12129 (N_12129,N_11136,N_11992);
and U12130 (N_12130,N_9193,N_9050);
nand U12131 (N_12131,N_10436,N_10681);
nor U12132 (N_12132,N_9402,N_11232);
nor U12133 (N_12133,N_10711,N_9707);
nor U12134 (N_12134,N_9343,N_11887);
or U12135 (N_12135,N_10059,N_10536);
and U12136 (N_12136,N_10880,N_10393);
or U12137 (N_12137,N_10057,N_11018);
or U12138 (N_12138,N_9668,N_10529);
xor U12139 (N_12139,N_9089,N_11269);
and U12140 (N_12140,N_10002,N_11507);
xor U12141 (N_12141,N_11246,N_10979);
or U12142 (N_12142,N_11153,N_9248);
xor U12143 (N_12143,N_9002,N_9548);
xnor U12144 (N_12144,N_10731,N_9214);
xnor U12145 (N_12145,N_9101,N_11164);
or U12146 (N_12146,N_9602,N_9126);
nand U12147 (N_12147,N_11429,N_9036);
nand U12148 (N_12148,N_9302,N_11080);
nand U12149 (N_12149,N_10001,N_11645);
nand U12150 (N_12150,N_9713,N_11920);
and U12151 (N_12151,N_10080,N_10340);
nor U12152 (N_12152,N_11217,N_9674);
and U12153 (N_12153,N_10116,N_11508);
and U12154 (N_12154,N_10620,N_10571);
nand U12155 (N_12155,N_11659,N_10593);
nand U12156 (N_12156,N_10757,N_10983);
xnor U12157 (N_12157,N_11760,N_9326);
or U12158 (N_12158,N_11849,N_10667);
or U12159 (N_12159,N_9189,N_10294);
nand U12160 (N_12160,N_9383,N_11896);
or U12161 (N_12161,N_9095,N_10570);
nand U12162 (N_12162,N_9100,N_9419);
xnor U12163 (N_12163,N_11727,N_11005);
xnor U12164 (N_12164,N_11728,N_9267);
or U12165 (N_12165,N_9964,N_10081);
nand U12166 (N_12166,N_9322,N_9014);
or U12167 (N_12167,N_9770,N_10765);
nor U12168 (N_12168,N_9554,N_10168);
and U12169 (N_12169,N_9011,N_10621);
and U12170 (N_12170,N_9825,N_10138);
nor U12171 (N_12171,N_11167,N_10474);
nand U12172 (N_12172,N_10259,N_9530);
nor U12173 (N_12173,N_9498,N_9645);
or U12174 (N_12174,N_10435,N_11819);
and U12175 (N_12175,N_10661,N_9873);
or U12176 (N_12176,N_10795,N_9156);
or U12177 (N_12177,N_9497,N_10160);
or U12178 (N_12178,N_9745,N_9636);
and U12179 (N_12179,N_9453,N_10346);
nor U12180 (N_12180,N_10228,N_11690);
xor U12181 (N_12181,N_11390,N_11408);
nand U12182 (N_12182,N_11280,N_10833);
or U12183 (N_12183,N_9012,N_10690);
or U12184 (N_12184,N_10036,N_9148);
nand U12185 (N_12185,N_11862,N_11582);
or U12186 (N_12186,N_11931,N_11826);
xnor U12187 (N_12187,N_9457,N_9040);
xor U12188 (N_12188,N_9266,N_10326);
nand U12189 (N_12189,N_11198,N_9220);
or U12190 (N_12190,N_11411,N_11878);
xnor U12191 (N_12191,N_9775,N_10263);
xnor U12192 (N_12192,N_11521,N_9420);
nand U12193 (N_12193,N_11868,N_9632);
or U12194 (N_12194,N_11441,N_9804);
nand U12195 (N_12195,N_9961,N_10085);
and U12196 (N_12196,N_10249,N_9143);
or U12197 (N_12197,N_10139,N_9412);
nand U12198 (N_12198,N_10654,N_11795);
and U12199 (N_12199,N_10236,N_9948);
and U12200 (N_12200,N_9896,N_10705);
or U12201 (N_12201,N_11338,N_10952);
or U12202 (N_12202,N_11699,N_9622);
nand U12203 (N_12203,N_9856,N_11649);
nor U12204 (N_12204,N_9400,N_10580);
xor U12205 (N_12205,N_9939,N_11165);
nand U12206 (N_12206,N_11981,N_11359);
or U12207 (N_12207,N_11081,N_9934);
nor U12208 (N_12208,N_9960,N_11401);
nor U12209 (N_12209,N_9544,N_9826);
nand U12210 (N_12210,N_11275,N_11474);
xnor U12211 (N_12211,N_11311,N_10708);
nand U12212 (N_12212,N_11372,N_10823);
and U12213 (N_12213,N_11841,N_11528);
nor U12214 (N_12214,N_11208,N_10127);
nor U12215 (N_12215,N_11904,N_9959);
and U12216 (N_12216,N_10383,N_9532);
or U12217 (N_12217,N_9844,N_9695);
nand U12218 (N_12218,N_11022,N_10938);
xor U12219 (N_12219,N_11481,N_10974);
or U12220 (N_12220,N_11609,N_9102);
nand U12221 (N_12221,N_9935,N_10662);
or U12222 (N_12222,N_9473,N_10736);
and U12223 (N_12223,N_11405,N_10238);
nand U12224 (N_12224,N_10503,N_10306);
nor U12225 (N_12225,N_10733,N_11116);
nand U12226 (N_12226,N_11410,N_10584);
nor U12227 (N_12227,N_9505,N_11511);
nor U12228 (N_12228,N_9442,N_11940);
nand U12229 (N_12229,N_11353,N_10046);
nand U12230 (N_12230,N_11432,N_10734);
nor U12231 (N_12231,N_10543,N_9449);
nor U12232 (N_12232,N_9866,N_10148);
nor U12233 (N_12233,N_9282,N_9330);
xor U12234 (N_12234,N_9769,N_11409);
nor U12235 (N_12235,N_11855,N_9474);
and U12236 (N_12236,N_10179,N_10286);
xnor U12237 (N_12237,N_10112,N_10501);
and U12238 (N_12238,N_10786,N_10448);
xnor U12239 (N_12239,N_11113,N_11066);
nand U12240 (N_12240,N_9179,N_9386);
and U12241 (N_12241,N_10848,N_9212);
and U12242 (N_12242,N_11378,N_10131);
xnor U12243 (N_12243,N_10412,N_10333);
and U12244 (N_12244,N_11293,N_10320);
nor U12245 (N_12245,N_11234,N_9656);
and U12246 (N_12246,N_11436,N_10663);
xnor U12247 (N_12247,N_10195,N_11006);
or U12248 (N_12248,N_9452,N_11021);
nand U12249 (N_12249,N_9346,N_10853);
and U12250 (N_12250,N_10989,N_11695);
xnor U12251 (N_12251,N_10125,N_10360);
nor U12252 (N_12252,N_10551,N_11499);
xor U12253 (N_12253,N_9117,N_9114);
nor U12254 (N_12254,N_9472,N_11281);
nand U12255 (N_12255,N_11745,N_10612);
xnor U12256 (N_12256,N_10758,N_11513);
or U12257 (N_12257,N_11309,N_10969);
and U12258 (N_12258,N_11936,N_10856);
and U12259 (N_12259,N_9203,N_10966);
nor U12260 (N_12260,N_11884,N_11631);
xnor U12261 (N_12261,N_9710,N_10578);
nor U12262 (N_12262,N_10682,N_11093);
xor U12263 (N_12263,N_10978,N_11714);
nor U12264 (N_12264,N_9516,N_10628);
xnor U12265 (N_12265,N_11288,N_10385);
xnor U12266 (N_12266,N_11952,N_10752);
or U12267 (N_12267,N_10216,N_11054);
and U12268 (N_12268,N_9824,N_11712);
and U12269 (N_12269,N_9683,N_11315);
and U12270 (N_12270,N_9693,N_10762);
or U12271 (N_12271,N_11702,N_9782);
or U12272 (N_12272,N_11077,N_11104);
or U12273 (N_12273,N_10211,N_10070);
xor U12274 (N_12274,N_11068,N_10636);
nor U12275 (N_12275,N_10693,N_11150);
or U12276 (N_12276,N_11563,N_11626);
xnor U12277 (N_12277,N_11808,N_9451);
or U12278 (N_12278,N_10936,N_10051);
or U12279 (N_12279,N_10006,N_9255);
or U12280 (N_12280,N_9573,N_9965);
nand U12281 (N_12281,N_11029,N_11350);
xor U12282 (N_12282,N_10388,N_10639);
or U12283 (N_12283,N_10058,N_11686);
nor U12284 (N_12284,N_11615,N_9297);
and U12285 (N_12285,N_11241,N_11534);
and U12286 (N_12286,N_9727,N_10205);
xor U12287 (N_12287,N_11073,N_9590);
or U12288 (N_12288,N_11254,N_9984);
xnor U12289 (N_12289,N_9480,N_10336);
nor U12290 (N_12290,N_10029,N_10229);
nand U12291 (N_12291,N_11915,N_9899);
nor U12292 (N_12292,N_9671,N_11561);
xor U12293 (N_12293,N_11750,N_11243);
nor U12294 (N_12294,N_11562,N_9288);
and U12295 (N_12295,N_10339,N_10083);
or U12296 (N_12296,N_10223,N_9550);
nor U12297 (N_12297,N_9279,N_9489);
or U12298 (N_12298,N_10405,N_11075);
and U12299 (N_12299,N_9665,N_9612);
xor U12300 (N_12300,N_11493,N_11601);
nor U12301 (N_12301,N_10218,N_9717);
nor U12302 (N_12302,N_11569,N_9565);
xor U12303 (N_12303,N_9974,N_11462);
nor U12304 (N_12304,N_11304,N_10111);
and U12305 (N_12305,N_11523,N_10364);
and U12306 (N_12306,N_11716,N_11240);
and U12307 (N_12307,N_9600,N_10676);
or U12308 (N_12308,N_10684,N_11705);
or U12309 (N_12309,N_9184,N_9325);
or U12310 (N_12310,N_10416,N_11625);
nor U12311 (N_12311,N_11061,N_10816);
or U12312 (N_12312,N_9060,N_10444);
or U12313 (N_12313,N_9893,N_9885);
xor U12314 (N_12314,N_10288,N_11780);
nand U12315 (N_12315,N_10153,N_11928);
and U12316 (N_12316,N_10502,N_9215);
nor U12317 (N_12317,N_10342,N_10556);
nor U12318 (N_12318,N_9658,N_11848);
and U12319 (N_12319,N_9843,N_10399);
and U12320 (N_12320,N_10314,N_10382);
xnor U12321 (N_12321,N_10021,N_11220);
xnor U12322 (N_12322,N_10445,N_11589);
and U12323 (N_12323,N_11115,N_11330);
or U12324 (N_12324,N_9483,N_11752);
xor U12325 (N_12325,N_11180,N_11793);
and U12326 (N_12326,N_10362,N_11152);
nand U12327 (N_12327,N_11482,N_10537);
or U12328 (N_12328,N_10617,N_9260);
nor U12329 (N_12329,N_9261,N_11148);
xor U12330 (N_12330,N_11125,N_9018);
or U12331 (N_12331,N_10062,N_10359);
and U12332 (N_12332,N_10019,N_10233);
nand U12333 (N_12333,N_10532,N_10224);
xnor U12334 (N_12334,N_11227,N_10129);
xor U12335 (N_12335,N_9615,N_10965);
and U12336 (N_12336,N_11658,N_11886);
xor U12337 (N_12337,N_9781,N_11685);
and U12338 (N_12338,N_10763,N_11127);
and U12339 (N_12339,N_9808,N_10177);
nand U12340 (N_12340,N_11987,N_11870);
or U12341 (N_12341,N_9977,N_11885);
or U12342 (N_12342,N_11883,N_10933);
and U12343 (N_12343,N_10573,N_10598);
and U12344 (N_12344,N_9124,N_11500);
xnor U12345 (N_12345,N_9032,N_9172);
nand U12346 (N_12346,N_11155,N_10794);
nand U12347 (N_12347,N_9598,N_9509);
xnor U12348 (N_12348,N_10919,N_11548);
nor U12349 (N_12349,N_11930,N_11531);
xnor U12350 (N_12350,N_11472,N_9872);
nor U12351 (N_12351,N_9056,N_10178);
or U12352 (N_12352,N_9139,N_11140);
nand U12353 (N_12353,N_11380,N_10068);
xnor U12354 (N_12354,N_10275,N_11903);
xnor U12355 (N_12355,N_9855,N_9596);
nor U12356 (N_12356,N_10798,N_9416);
and U12357 (N_12357,N_9041,N_9434);
nor U12358 (N_12358,N_9321,N_11932);
or U12359 (N_12359,N_11772,N_11847);
or U12360 (N_12360,N_10749,N_9868);
or U12361 (N_12361,N_11457,N_10204);
nand U12362 (N_12362,N_10822,N_9802);
nand U12363 (N_12363,N_11617,N_10540);
xor U12364 (N_12364,N_11509,N_10398);
or U12365 (N_12365,N_9123,N_9033);
xnor U12366 (N_12366,N_11559,N_9153);
xor U12367 (N_12367,N_9553,N_10683);
xnor U12368 (N_12368,N_11823,N_10313);
and U12369 (N_12369,N_9949,N_10633);
or U12370 (N_12370,N_11906,N_11806);
xor U12371 (N_12371,N_11305,N_9098);
nor U12372 (N_12372,N_10792,N_11838);
xor U12373 (N_12373,N_9371,N_10347);
nand U12374 (N_12374,N_9329,N_9759);
or U12375 (N_12375,N_10250,N_11488);
nor U12376 (N_12376,N_10361,N_11213);
or U12377 (N_12377,N_11205,N_10114);
nand U12378 (N_12378,N_9028,N_11485);
or U12379 (N_12379,N_10657,N_9657);
or U12380 (N_12380,N_9663,N_10561);
xor U12381 (N_12381,N_10387,N_10904);
and U12382 (N_12382,N_11040,N_10130);
xor U12383 (N_12383,N_9933,N_10464);
nand U12384 (N_12384,N_10185,N_11732);
and U12385 (N_12385,N_11997,N_10656);
nor U12386 (N_12386,N_9336,N_10935);
or U12387 (N_12387,N_10496,N_11846);
or U12388 (N_12388,N_11945,N_10541);
nand U12389 (N_12389,N_10433,N_9975);
nand U12390 (N_12390,N_10826,N_10165);
nor U12391 (N_12391,N_10810,N_11203);
nor U12392 (N_12392,N_11779,N_9294);
and U12393 (N_12393,N_10293,N_9391);
xor U12394 (N_12394,N_9678,N_10449);
nand U12395 (N_12395,N_10843,N_11832);
and U12396 (N_12396,N_9485,N_9538);
and U12397 (N_12397,N_10315,N_9425);
and U12398 (N_12398,N_11385,N_10109);
xnor U12399 (N_12399,N_11190,N_10533);
nor U12400 (N_12400,N_10396,N_11027);
and U12401 (N_12401,N_10990,N_11584);
nand U12402 (N_12402,N_11381,N_9023);
nor U12403 (N_12403,N_10220,N_9039);
xnor U12404 (N_12404,N_10926,N_9281);
xnor U12405 (N_12405,N_10692,N_11106);
nand U12406 (N_12406,N_9200,N_10497);
or U12407 (N_12407,N_10100,N_11843);
nor U12408 (N_12408,N_10999,N_10685);
or U12409 (N_12409,N_10514,N_10171);
nand U12410 (N_12410,N_10522,N_9813);
nor U12411 (N_12411,N_10874,N_9836);
or U12412 (N_12412,N_11766,N_11025);
xnor U12413 (N_12413,N_9046,N_11327);
nand U12414 (N_12414,N_11266,N_11811);
nand U12415 (N_12415,N_9228,N_11339);
and U12416 (N_12416,N_9909,N_11605);
and U12417 (N_12417,N_9679,N_9579);
xnor U12418 (N_12418,N_11790,N_11861);
xor U12419 (N_12419,N_10964,N_10891);
and U12420 (N_12420,N_10377,N_11218);
and U12421 (N_12421,N_10120,N_9165);
and U12422 (N_12422,N_11326,N_10603);
or U12423 (N_12423,N_10270,N_9439);
nand U12424 (N_12424,N_10658,N_10894);
or U12425 (N_12425,N_11191,N_11024);
nor U12426 (N_12426,N_10323,N_11199);
and U12427 (N_12427,N_10428,N_11542);
or U12428 (N_12428,N_9686,N_11892);
xnor U12429 (N_12429,N_11654,N_11447);
or U12430 (N_12430,N_9580,N_11316);
nor U12431 (N_12431,N_9403,N_11360);
nand U12432 (N_12432,N_11112,N_11967);
and U12433 (N_12433,N_9243,N_10266);
nand U12434 (N_12434,N_10358,N_11011);
or U12435 (N_12435,N_10328,N_9128);
or U12436 (N_12436,N_10729,N_11103);
xnor U12437 (N_12437,N_11971,N_9789);
xnor U12438 (N_12438,N_10834,N_9652);
xnor U12439 (N_12439,N_10796,N_9858);
xnor U12440 (N_12440,N_10666,N_10498);
or U12441 (N_12441,N_10473,N_10840);
nand U12442 (N_12442,N_10566,N_9922);
nor U12443 (N_12443,N_10353,N_10258);
xnor U12444 (N_12444,N_11169,N_10196);
xnor U12445 (N_12445,N_11979,N_9799);
or U12446 (N_12446,N_10901,N_11387);
and U12447 (N_12447,N_10482,N_11473);
nor U12448 (N_12448,N_11754,N_11056);
and U12449 (N_12449,N_9524,N_9547);
xor U12450 (N_12450,N_11026,N_11730);
nand U12451 (N_12451,N_11369,N_11320);
nor U12452 (N_12452,N_9838,N_9183);
xor U12453 (N_12453,N_10296,N_10553);
nand U12454 (N_12454,N_9845,N_10038);
xor U12455 (N_12455,N_11512,N_9447);
and U12456 (N_12456,N_11086,N_9436);
nor U12457 (N_12457,N_9038,N_9982);
and U12458 (N_12458,N_10929,N_10122);
nor U12459 (N_12459,N_9534,N_9971);
nor U12460 (N_12460,N_11057,N_9841);
nand U12461 (N_12461,N_11501,N_11969);
xor U12462 (N_12462,N_9700,N_10755);
and U12463 (N_12463,N_9584,N_11621);
nor U12464 (N_12464,N_9073,N_9162);
and U12465 (N_12465,N_10743,N_11893);
xor U12466 (N_12466,N_9931,N_9815);
and U12467 (N_12467,N_9166,N_11744);
nor U12468 (N_12468,N_10219,N_9496);
xnor U12469 (N_12469,N_9379,N_10748);
nor U12470 (N_12470,N_10193,N_10927);
or U12471 (N_12471,N_9418,N_10045);
or U12472 (N_12472,N_11554,N_10897);
and U12473 (N_12473,N_10877,N_9950);
and U12474 (N_12474,N_10425,N_10043);
nor U12475 (N_12475,N_10630,N_9529);
or U12476 (N_12476,N_11646,N_9749);
and U12477 (N_12477,N_11255,N_10642);
xor U12478 (N_12478,N_11450,N_11865);
xnor U12479 (N_12479,N_11545,N_9293);
or U12480 (N_12480,N_9842,N_11435);
and U12481 (N_12481,N_10215,N_10118);
and U12482 (N_12482,N_9380,N_11677);
and U12483 (N_12483,N_11367,N_10857);
and U12484 (N_12484,N_11090,N_10504);
nand U12485 (N_12485,N_10992,N_11424);
nor U12486 (N_12486,N_10659,N_10457);
xnor U12487 (N_12487,N_11934,N_11610);
xor U12488 (N_12488,N_9309,N_11395);
nand U12489 (N_12489,N_9827,N_10872);
nor U12490 (N_12490,N_9176,N_9662);
and U12491 (N_12491,N_11135,N_11701);
nand U12492 (N_12492,N_10896,N_9421);
or U12493 (N_12493,N_11850,N_11210);
nor U12494 (N_12494,N_10591,N_11839);
or U12495 (N_12495,N_10056,N_11748);
nor U12496 (N_12496,N_9239,N_10660);
nor U12497 (N_12497,N_11069,N_10044);
xor U12498 (N_12498,N_9092,N_11858);
xor U12499 (N_12499,N_10481,N_9476);
xnor U12500 (N_12500,N_11620,N_9024);
and U12501 (N_12501,N_9921,N_10977);
nor U12502 (N_12502,N_10065,N_11703);
and U12503 (N_12503,N_10401,N_10776);
xnor U12504 (N_12504,N_9504,N_9637);
or U12505 (N_12505,N_10980,N_10588);
or U12506 (N_12506,N_10618,N_11681);
nor U12507 (N_12507,N_9667,N_10851);
nor U12508 (N_12508,N_10367,N_11977);
xnor U12509 (N_12509,N_11813,N_11539);
nor U12510 (N_12510,N_10087,N_11265);
nor U12511 (N_12511,N_11863,N_9053);
xnor U12512 (N_12512,N_9324,N_9688);
nor U12513 (N_12513,N_10727,N_11916);
or U12514 (N_12514,N_11993,N_11888);
and U12515 (N_12515,N_10115,N_11252);
nor U12516 (N_12516,N_10023,N_9519);
or U12517 (N_12517,N_9930,N_11271);
nor U12518 (N_12518,N_11183,N_9455);
nand U12519 (N_12519,N_11297,N_10572);
xor U12520 (N_12520,N_9048,N_10549);
nor U12521 (N_12521,N_10420,N_11679);
nand U12522 (N_12522,N_9456,N_10400);
or U12523 (N_12523,N_10614,N_10528);
and U12524 (N_12524,N_9467,N_11798);
xor U12525 (N_12525,N_9029,N_11573);
xor U12526 (N_12526,N_10861,N_11707);
or U12527 (N_12527,N_10063,N_11591);
xor U12528 (N_12528,N_11613,N_10813);
xor U12529 (N_12529,N_9208,N_11963);
or U12530 (N_12530,N_10284,N_10356);
xnor U12531 (N_12531,N_9861,N_9465);
nor U12532 (N_12532,N_10599,N_11096);
xor U12533 (N_12533,N_10836,N_9894);
xnor U12534 (N_12534,N_11442,N_10291);
or U12535 (N_12535,N_9188,N_10764);
or U12536 (N_12536,N_9331,N_9837);
and U12537 (N_12537,N_10010,N_11423);
nand U12538 (N_12538,N_9560,N_11675);
xnor U12539 (N_12539,N_10517,N_11307);
nand U12540 (N_12540,N_9904,N_10232);
nand U12541 (N_12541,N_9394,N_10285);
nand U12542 (N_12542,N_10301,N_11010);
nor U12543 (N_12543,N_9328,N_10777);
or U12544 (N_12544,N_10076,N_9978);
nand U12545 (N_12545,N_9979,N_10141);
and U12546 (N_12546,N_10247,N_9355);
xor U12547 (N_12547,N_10365,N_11287);
nor U12548 (N_12548,N_11452,N_10986);
xnor U12549 (N_12549,N_9185,N_10688);
nand U12550 (N_12550,N_9360,N_9353);
xnor U12551 (N_12551,N_10079,N_10375);
or U12552 (N_12552,N_11851,N_10750);
nor U12553 (N_12553,N_9118,N_10072);
nand U12554 (N_12554,N_11120,N_10778);
or U12555 (N_12555,N_9591,N_11678);
and U12556 (N_12556,N_9199,N_9542);
nand U12557 (N_12557,N_9291,N_11682);
nor U12558 (N_12558,N_9742,N_11994);
nor U12559 (N_12559,N_9758,N_10489);
nor U12560 (N_12560,N_11323,N_9862);
nor U12561 (N_12561,N_11564,N_10865);
and U12562 (N_12562,N_9833,N_10720);
xnor U12563 (N_12563,N_11219,N_11556);
nor U12564 (N_12564,N_11557,N_10394);
nor U12565 (N_12565,N_10800,N_11786);
or U12566 (N_12566,N_10946,N_9626);
and U12567 (N_12567,N_11131,N_9613);
or U12568 (N_12568,N_9723,N_9953);
nand U12569 (N_12569,N_10557,N_9648);
nor U12570 (N_12570,N_9988,N_9170);
and U12571 (N_12571,N_9871,N_10217);
nand U12572 (N_12572,N_9138,N_9191);
or U12573 (N_12573,N_9160,N_10567);
or U12574 (N_12574,N_11391,N_9275);
or U12575 (N_12575,N_10040,N_11298);
xor U12576 (N_12576,N_11810,N_11337);
and U12577 (N_12577,N_9607,N_10819);
xnor U12578 (N_12578,N_9577,N_9414);
and U12579 (N_12579,N_9397,N_10106);
nor U12580 (N_12580,N_9429,N_11854);
xor U12581 (N_12581,N_10166,N_9552);
nand U12582 (N_12582,N_11738,N_11400);
nor U12583 (N_12583,N_9225,N_11486);
xnor U12584 (N_12584,N_9238,N_10760);
xor U12585 (N_12585,N_9461,N_10067);
or U12586 (N_12586,N_10710,N_10132);
nor U12587 (N_12587,N_9049,N_9936);
nand U12588 (N_12588,N_11550,N_9743);
and U12589 (N_12589,N_9898,N_11074);
and U12590 (N_12590,N_9863,N_11082);
nor U12591 (N_12591,N_10104,N_10941);
and U12592 (N_12592,N_11347,N_9237);
nand U12593 (N_12593,N_9880,N_11438);
and U12594 (N_12594,N_11612,N_9890);
xor U12595 (N_12595,N_9919,N_10815);
and U12596 (N_12596,N_11470,N_9213);
xor U12597 (N_12597,N_11334,N_10831);
or U12598 (N_12598,N_11842,N_11354);
or U12599 (N_12599,N_9718,N_10351);
nand U12600 (N_12600,N_11603,N_9173);
nand U12601 (N_12601,N_10921,N_11028);
and U12602 (N_12602,N_9557,N_10961);
nand U12603 (N_12603,N_11835,N_9370);
nor U12604 (N_12604,N_9756,N_9471);
nand U12605 (N_12605,N_11095,N_11130);
xor U12606 (N_12606,N_9433,N_11785);
or U12607 (N_12607,N_10910,N_11126);
nand U12608 (N_12608,N_9251,N_9903);
nor U12609 (N_12609,N_10970,N_10200);
and U12610 (N_12610,N_11480,N_9915);
and U12611 (N_12611,N_10525,N_9013);
and U12612 (N_12612,N_9618,N_9940);
xor U12613 (N_12613,N_9647,N_9006);
and U12614 (N_12614,N_9150,N_10558);
or U12615 (N_12615,N_10609,N_11803);
and U12616 (N_12616,N_11784,N_9318);
xor U12617 (N_12617,N_11245,N_9205);
nor U12618 (N_12618,N_11471,N_11160);
nand U12619 (N_12619,N_10920,N_10225);
nand U12620 (N_12620,N_10048,N_9354);
nand U12621 (N_12621,N_9372,N_11017);
and U12622 (N_12622,N_9164,N_11034);
xor U12623 (N_12623,N_11961,N_9740);
or U12624 (N_12624,N_9422,N_11007);
xnor U12625 (N_12625,N_9634,N_10931);
nor U12626 (N_12626,N_9484,N_10082);
xnor U12627 (N_12627,N_11238,N_11146);
or U12628 (N_12628,N_11379,N_10338);
or U12629 (N_12629,N_11268,N_11403);
and U12630 (N_12630,N_11433,N_11147);
xnor U12631 (N_12631,N_10746,N_10279);
xnor U12632 (N_12632,N_9486,N_10886);
or U12633 (N_12633,N_11917,N_11362);
and U12634 (N_12634,N_9630,N_11966);
nand U12635 (N_12635,N_10653,N_10390);
and U12636 (N_12636,N_10084,N_11064);
nor U12637 (N_12637,N_11723,N_11789);
and U12638 (N_12638,N_9044,N_9075);
nand U12639 (N_12639,N_11262,N_11003);
nand U12640 (N_12640,N_9257,N_10506);
nor U12641 (N_12641,N_10417,N_10706);
or U12642 (N_12642,N_11553,N_9065);
nand U12643 (N_12643,N_11321,N_10427);
nand U12644 (N_12644,N_10871,N_10300);
and U12645 (N_12645,N_9906,N_9592);
and U12646 (N_12646,N_10035,N_11549);
nand U12647 (N_12647,N_10370,N_10422);
xor U12648 (N_12648,N_10251,N_9761);
nor U12649 (N_12649,N_9768,N_11118);
nand U12650 (N_12650,N_9722,N_11399);
xnor U12651 (N_12651,N_9078,N_10325);
or U12652 (N_12652,N_10868,N_11492);
or U12653 (N_12653,N_10914,N_11817);
or U12654 (N_12654,N_11235,N_10672);
nand U12655 (N_12655,N_11735,N_11302);
xnor U12656 (N_12656,N_9994,N_9967);
or U12657 (N_12657,N_10234,N_9494);
nor U12658 (N_12658,N_9064,N_9495);
and U12659 (N_12659,N_11880,N_11900);
xnor U12660 (N_12660,N_9219,N_11355);
xor U12661 (N_12661,N_10086,N_10671);
or U12662 (N_12662,N_10909,N_10227);
or U12663 (N_12663,N_10221,N_9801);
nor U12664 (N_12664,N_9760,N_10411);
or U12665 (N_12665,N_11270,N_11800);
or U12666 (N_12666,N_9058,N_9246);
and U12667 (N_12667,N_11781,N_10260);
and U12668 (N_12668,N_11604,N_9586);
nand U12669 (N_12669,N_9986,N_9137);
xnor U12670 (N_12670,N_10870,N_9010);
nor U12671 (N_12671,N_9207,N_9962);
or U12672 (N_12672,N_10971,N_10960);
xor U12673 (N_12673,N_10189,N_11371);
xor U12674 (N_12674,N_10322,N_11299);
and U12675 (N_12675,N_9154,N_11102);
or U12676 (N_12676,N_9609,N_9392);
nand U12677 (N_12677,N_9111,N_10099);
nor U12678 (N_12678,N_11181,N_10544);
or U12679 (N_12679,N_11310,N_11541);
xor U12680 (N_12680,N_10718,N_10513);
nand U12681 (N_12681,N_9831,N_9406);
nand U12682 (N_12682,N_9067,N_9852);
or U12683 (N_12683,N_9830,N_9594);
nand U12684 (N_12684,N_11643,N_10174);
and U12685 (N_12685,N_10889,N_9888);
or U12686 (N_12686,N_11935,N_10117);
and U12687 (N_12687,N_10841,N_9655);
nor U12688 (N_12688,N_10344,N_10144);
nor U12689 (N_12689,N_11577,N_9068);
xnor U12690 (N_12690,N_9103,N_11031);
and U12691 (N_12691,N_10337,N_11568);
and U12692 (N_12692,N_11356,N_9847);
xnor U12693 (N_12693,N_9732,N_11193);
nor U12694 (N_12694,N_11296,N_10381);
nand U12695 (N_12695,N_10378,N_9670);
and U12696 (N_12696,N_10317,N_11346);
nand U12697 (N_12697,N_10345,N_10832);
nor U12698 (N_12698,N_11300,N_11277);
and U12699 (N_12699,N_9643,N_10429);
nor U12700 (N_12700,N_11877,N_10838);
xnor U12701 (N_12701,N_9298,N_10197);
and U12702 (N_12702,N_11593,N_11715);
or U12703 (N_12703,N_10866,N_9897);
nor U12704 (N_12704,N_10264,N_10441);
or U12705 (N_12705,N_9005,N_11475);
nor U12706 (N_12706,N_10878,N_9106);
nor U12707 (N_12707,N_11137,N_9290);
nor U12708 (N_12708,N_11425,N_9905);
nand U12709 (N_12709,N_9788,N_11396);
nor U12710 (N_12710,N_11592,N_9589);
or U12711 (N_12711,N_11821,N_11015);
xor U12712 (N_12712,N_10041,N_9595);
or U12713 (N_12713,N_11709,N_9327);
nor U12714 (N_12714,N_11891,N_11002);
nor U12715 (N_12715,N_9365,N_11163);
or U12716 (N_12716,N_10717,N_9942);
nand U12717 (N_12717,N_9859,N_11072);
xor U12718 (N_12718,N_9527,N_10253);
and U12719 (N_12719,N_9508,N_9525);
and U12720 (N_12720,N_9777,N_11107);
xnor U12721 (N_12721,N_11984,N_11261);
or U12722 (N_12722,N_10854,N_9076);
nand U12723 (N_12723,N_11059,N_10454);
xnor U12724 (N_12724,N_9883,N_9136);
and U12725 (N_12725,N_11247,N_9426);
nor U12726 (N_12726,N_9373,N_11869);
nand U12727 (N_12727,N_11985,N_10821);
or U12728 (N_12728,N_11947,N_11764);
nand U12729 (N_12729,N_9502,N_10110);
or U12730 (N_12730,N_9430,N_10839);
xnor U12731 (N_12731,N_10146,N_9954);
and U12732 (N_12732,N_11538,N_9464);
xnor U12733 (N_12733,N_10194,N_11201);
nor U12734 (N_12734,N_11889,N_9724);
xor U12735 (N_12735,N_11121,N_10101);
xor U12736 (N_12736,N_11683,N_9112);
nand U12737 (N_12737,N_11050,N_11149);
nor U12738 (N_12738,N_10137,N_9217);
or U12739 (N_12739,N_11099,N_9358);
nand U12740 (N_12740,N_11767,N_11721);
or U12741 (N_12741,N_9356,N_10744);
nor U12742 (N_12742,N_11207,N_11144);
nor U12743 (N_12743,N_10066,N_11114);
xnor U12744 (N_12744,N_11282,N_9851);
nand U12745 (N_12745,N_10781,N_10095);
and U12746 (N_12746,N_10702,N_9120);
nand U12747 (N_12747,N_11394,N_10017);
nor U12748 (N_12748,N_9694,N_11902);
and U12749 (N_12749,N_10913,N_11919);
nand U12750 (N_12750,N_10446,N_11807);
or U12751 (N_12751,N_9517,N_10876);
and U12752 (N_12752,N_11336,N_9357);
nand U12753 (N_12753,N_10560,N_10951);
xor U12754 (N_12754,N_9085,N_11802);
or U12755 (N_12755,N_10039,N_10374);
xnor U12756 (N_12756,N_9084,N_9440);
and U12757 (N_12757,N_11953,N_11294);
and U12758 (N_12758,N_9692,N_9348);
xnor U12759 (N_12759,N_10716,N_11386);
nor U12760 (N_12760,N_9578,N_10589);
nand U12761 (N_12761,N_10007,N_11319);
nor U12762 (N_12762,N_10545,N_9520);
and U12763 (N_12763,N_11156,N_11955);
nor U12764 (N_12764,N_10928,N_11225);
nor U12765 (N_12765,N_10574,N_11912);
xnor U12766 (N_12766,N_10472,N_10741);
xor U12767 (N_12767,N_10761,N_9052);
and U12768 (N_12768,N_11357,N_11204);
xnor U12769 (N_12769,N_11451,N_10140);
xnor U12770 (N_12770,N_9460,N_10410);
nand U12771 (N_12771,N_11585,N_11382);
nor U12772 (N_12772,N_10469,N_11172);
nand U12773 (N_12773,N_11428,N_9091);
nand U12774 (N_12774,N_11661,N_9969);
nor U12775 (N_12775,N_10475,N_9952);
xnor U12776 (N_12776,N_9130,N_11078);
or U12777 (N_12777,N_11560,N_9912);
nor U12778 (N_12778,N_10689,N_9240);
nor U12779 (N_12779,N_11922,N_11986);
and U12780 (N_12780,N_11925,N_9401);
or U12781 (N_12781,N_10281,N_10903);
xor U12782 (N_12782,N_11540,N_10825);
nand U12783 (N_12783,N_9146,N_10278);
nand U12784 (N_12784,N_10883,N_9980);
and U12785 (N_12785,N_11035,N_9687);
and U12786 (N_12786,N_11668,N_11170);
and U12787 (N_12787,N_9341,N_9797);
or U12788 (N_12788,N_11648,N_11667);
nor U12789 (N_12789,N_9019,N_10812);
nand U12790 (N_12790,N_9405,N_10576);
or U12791 (N_12791,N_9428,N_11415);
nor U12792 (N_12792,N_10431,N_11055);
nor U12793 (N_12793,N_9259,N_10713);
or U12794 (N_12794,N_10331,N_10379);
nand U12795 (N_12795,N_11231,N_9878);
xor U12796 (N_12796,N_9752,N_10973);
nor U12797 (N_12797,N_11943,N_10592);
and U12798 (N_12798,N_10699,N_11587);
xnor U12799 (N_12799,N_10255,N_10793);
and U12800 (N_12800,N_9650,N_9390);
xnor U12801 (N_12801,N_10948,N_10539);
or U12802 (N_12802,N_10908,N_11614);
and U12803 (N_12803,N_10987,N_10206);
nand U12804 (N_12804,N_10849,N_9167);
nor U12805 (N_12805,N_9233,N_11233);
nand U12806 (N_12806,N_10397,N_11636);
or U12807 (N_12807,N_9366,N_11182);
nor U12808 (N_12808,N_9236,N_10801);
xor U12809 (N_12809,N_11762,N_10962);
nand U12810 (N_12810,N_10932,N_11822);
nand U12811 (N_12811,N_11530,N_10624);
xor U12812 (N_12812,N_9043,N_9202);
or U12813 (N_12813,N_10030,N_9928);
and U12814 (N_12814,N_10466,N_11791);
and U12815 (N_12815,N_11089,N_11110);
nor U12816 (N_12816,N_9274,N_10032);
nand U12817 (N_12817,N_10508,N_11788);
and U12818 (N_12818,N_11544,N_9285);
xnor U12819 (N_12819,N_10487,N_11019);
xnor U12820 (N_12820,N_10069,N_10450);
or U12821 (N_12821,N_9066,N_11761);
xor U12822 (N_12822,N_11491,N_9812);
nand U12823 (N_12823,N_11414,N_10075);
nand U12824 (N_12824,N_11801,N_11416);
nor U12825 (N_12825,N_9574,N_11283);
nor U12826 (N_12826,N_9512,N_11739);
and U12827 (N_12827,N_9963,N_9069);
xnor U12828 (N_12828,N_9720,N_9737);
or U12829 (N_12829,N_9055,N_9362);
nor U12830 (N_12830,N_10797,N_9776);
nor U12831 (N_12831,N_10304,N_9093);
or U12832 (N_12832,N_9195,N_9575);
nand U12833 (N_12833,N_9009,N_9364);
xor U12834 (N_12834,N_11637,N_11741);
or U12835 (N_12835,N_9410,N_11001);
nor U12836 (N_12836,N_11173,N_11119);
nand U12837 (N_12837,N_11600,N_11815);
xor U12838 (N_12838,N_9427,N_9235);
or U12839 (N_12839,N_9848,N_11999);
nor U12840 (N_12840,N_10088,N_10535);
nor U12841 (N_12841,N_11960,N_9854);
or U12842 (N_12842,N_10991,N_11704);
or U12843 (N_12843,N_9099,N_10564);
or U12844 (N_12844,N_10462,N_11032);
or U12845 (N_12845,N_11157,N_10024);
nor U12846 (N_12846,N_9003,N_10078);
or U12847 (N_12847,N_10105,N_10077);
or U12848 (N_12848,N_9269,N_10134);
xnor U12849 (N_12849,N_9680,N_9646);
nor U12850 (N_12850,N_9385,N_10097);
and U12851 (N_12851,N_9487,N_10047);
nor U12852 (N_12852,N_11794,N_10629);
or U12853 (N_12853,N_11301,N_9635);
and U12854 (N_12854,N_11547,N_9300);
nand U12855 (N_12855,N_10811,N_10318);
nor U12856 (N_12856,N_11237,N_9129);
nor U12857 (N_12857,N_10622,N_10555);
or U12858 (N_12858,N_11427,N_9666);
xor U12859 (N_12859,N_10012,N_9223);
or U12860 (N_12860,N_11827,N_11123);
xor U12861 (N_12861,N_11595,N_11688);
or U12862 (N_12862,N_11664,N_9377);
or U12863 (N_12863,N_10483,N_9528);
xor U12864 (N_12864,N_10698,N_10845);
and U12865 (N_12865,N_9463,N_9477);
nor U12866 (N_12866,N_9673,N_9587);
and U12867 (N_12867,N_10209,N_10463);
or U12868 (N_12868,N_9499,N_10451);
nor U12869 (N_12869,N_10649,N_11030);
nand U12870 (N_12870,N_10864,N_10280);
xnor U12871 (N_12871,N_9541,N_11640);
xor U12872 (N_12872,N_10997,N_9728);
nor U12873 (N_12873,N_11159,N_9932);
nor U12874 (N_12874,N_11852,N_10728);
and U12875 (N_12875,N_9914,N_9526);
xnor U12876 (N_12876,N_11720,N_11599);
nor U12877 (N_12877,N_11973,N_10261);
xnor U12878 (N_12878,N_9689,N_9629);
xor U12879 (N_12879,N_9083,N_9675);
nand U12880 (N_12880,N_10695,N_9850);
xnor U12881 (N_12881,N_10579,N_11825);
and U12882 (N_12882,N_9042,N_11663);
or U12883 (N_12883,N_11913,N_9911);
xor U12884 (N_12884,N_9171,N_9860);
and U12885 (N_12885,N_10352,N_11751);
xnor U12886 (N_12886,N_11742,N_11178);
and U12887 (N_12887,N_11756,N_9376);
and U12888 (N_12888,N_11468,N_11657);
or U12889 (N_12889,N_10305,N_9163);
xnor U12890 (N_12890,N_11459,N_11836);
or U12891 (N_12891,N_10102,N_11901);
nor U12892 (N_12892,N_9363,N_9684);
nor U12893 (N_12893,N_9224,N_9432);
nor U12894 (N_12894,N_11552,N_10409);
or U12895 (N_12895,N_10949,N_10460);
nand U12896 (N_12896,N_10550,N_10176);
and U12897 (N_12897,N_10424,N_9711);
nor U12898 (N_12898,N_10638,N_10747);
and U12899 (N_12899,N_10967,N_10465);
xor U12900 (N_12900,N_11465,N_9337);
nor U12901 (N_12901,N_11133,N_10809);
nor U12902 (N_12902,N_11757,N_9900);
nand U12903 (N_12903,N_10715,N_11212);
nor U12904 (N_12904,N_11214,N_10606);
nand U12905 (N_12905,N_11991,N_11937);
nand U12906 (N_12906,N_9562,N_9187);
nor U12907 (N_12907,N_9623,N_9539);
nand U12908 (N_12908,N_10471,N_10214);
xor U12909 (N_12909,N_9027,N_9902);
and U12910 (N_12910,N_9198,N_9310);
nor U12911 (N_12911,N_10210,N_10726);
or U12912 (N_12912,N_9561,N_9134);
or U12913 (N_12913,N_11290,N_9729);
and U12914 (N_12914,N_11989,N_9437);
or U12915 (N_12915,N_10714,N_10341);
or U12916 (N_12916,N_9501,N_11644);
nor U12917 (N_12917,N_9669,N_9121);
nor U12918 (N_12918,N_9828,N_11023);
xnor U12919 (N_12919,N_10386,N_9631);
or U12920 (N_12920,N_10207,N_9617);
nor U12921 (N_12921,N_9169,N_11941);
nand U12922 (N_12922,N_9870,N_10028);
and U12923 (N_12923,N_10302,N_9533);
xor U12924 (N_12924,N_9482,N_10707);
and U12925 (N_12925,N_10994,N_9944);
nand U12926 (N_12926,N_9849,N_9576);
or U12927 (N_12927,N_11478,N_11532);
nand U12928 (N_12928,N_9314,N_9731);
xor U12929 (N_12929,N_10230,N_11627);
xor U12930 (N_12930,N_11684,N_11036);
nor U12931 (N_12931,N_10157,N_9446);
nand U12932 (N_12932,N_10003,N_9778);
or U12933 (N_12933,N_9649,N_11176);
or U12934 (N_12934,N_9638,N_10637);
or U12935 (N_12935,N_10686,N_10391);
or U12936 (N_12936,N_10873,N_10332);
and U12937 (N_12937,N_9757,N_9507);
nor U12938 (N_12938,N_9218,N_9303);
and U12939 (N_12939,N_9025,N_10175);
xnor U12940 (N_12940,N_10934,N_10277);
and U12941 (N_12941,N_11856,N_9500);
nand U12942 (N_12942,N_10407,N_10371);
or U12943 (N_12943,N_11708,N_10443);
nor U12944 (N_12944,N_10918,N_9308);
xnor U12945 (N_12945,N_9783,N_11044);
xnor U12946 (N_12946,N_9725,N_9549);
and U12947 (N_12947,N_10884,N_9151);
nand U12948 (N_12948,N_11331,N_9368);
nor U12949 (N_12949,N_11286,N_10521);
nor U12950 (N_12950,N_10350,N_10575);
or U12951 (N_12951,N_9133,N_10343);
and U12952 (N_12952,N_10655,N_10268);
nand U12953 (N_12953,N_11039,N_10808);
xnor U12954 (N_12954,N_11633,N_9619);
or U12955 (N_12955,N_10802,N_9784);
nor U12956 (N_12956,N_11038,N_11656);
nand U12957 (N_12957,N_9886,N_9823);
xor U12958 (N_12958,N_11711,N_11797);
or U12959 (N_12959,N_9829,N_9976);
xnor U12960 (N_12960,N_10126,N_11576);
nor U12961 (N_12961,N_9086,N_10267);
nor U12962 (N_12962,N_9253,N_10170);
and U12963 (N_12963,N_10646,N_10423);
and U12964 (N_12964,N_10756,N_11322);
or U12965 (N_12965,N_11141,N_9438);
or U12966 (N_12966,N_9206,N_9194);
xnor U12967 (N_12967,N_10869,N_10745);
and U12968 (N_12968,N_10492,N_11306);
and U12969 (N_12969,N_11581,N_9475);
and U12970 (N_12970,N_10321,N_11376);
and U12971 (N_12971,N_10881,N_9079);
xor U12972 (N_12972,N_11325,N_11871);
nand U12973 (N_12973,N_11590,N_10652);
xnor U12974 (N_12974,N_9907,N_11042);
xor U12975 (N_12975,N_10290,N_10453);
nor U12976 (N_12976,N_10587,N_9766);
and U12977 (N_12977,N_11665,N_10701);
nand U12978 (N_12978,N_10807,N_11694);
nand U12979 (N_12979,N_10467,N_9140);
xnor U12980 (N_12980,N_10307,N_9347);
and U12981 (N_12981,N_9231,N_9640);
nor U12982 (N_12982,N_9256,N_11162);
nand U12983 (N_12983,N_9923,N_10520);
and U12984 (N_12984,N_11228,N_10274);
nor U12985 (N_12985,N_9910,N_9082);
nand U12986 (N_12986,N_10945,N_10490);
or U12987 (N_12987,N_11188,N_10477);
xor U12988 (N_12988,N_11696,N_10269);
nand U12989 (N_12989,N_11975,N_9929);
and U12990 (N_12990,N_11875,N_11402);
nor U12991 (N_12991,N_9289,N_10742);
and U12992 (N_12992,N_10252,N_10687);
nor U12993 (N_12993,N_10128,N_10022);
and U12994 (N_12994,N_9785,N_9395);
xor U12995 (N_12995,N_11910,N_9407);
nand U12996 (N_12996,N_10319,N_10524);
nor U12997 (N_12997,N_10103,N_9144);
nor U12998 (N_12998,N_10256,N_10586);
or U12999 (N_12999,N_10244,N_11972);
xnor U13000 (N_13000,N_9221,N_11660);
nor U13001 (N_13001,N_11828,N_10604);
and U13002 (N_13002,N_9796,N_10297);
or U13003 (N_13003,N_10875,N_10569);
nor U13004 (N_13004,N_10093,N_11439);
xnor U13005 (N_13005,N_11921,N_9132);
nor U13006 (N_13006,N_10478,N_9306);
xor U13007 (N_13007,N_9943,N_10312);
and U13008 (N_13008,N_10470,N_11184);
nand U13009 (N_13009,N_10563,N_10354);
xor U13010 (N_13010,N_10958,N_9247);
and U13011 (N_13011,N_9283,N_9746);
and U13012 (N_13012,N_11109,N_10597);
or U13013 (N_13013,N_11948,N_10491);
nand U13014 (N_13014,N_11317,N_9884);
nor U13015 (N_13015,N_10133,N_10512);
nand U13016 (N_13016,N_9059,N_10619);
and U13017 (N_13017,N_9968,N_10452);
nand U13018 (N_13018,N_9459,N_11996);
nor U13019 (N_13019,N_9469,N_11653);
and U13020 (N_13020,N_9479,N_9273);
or U13021 (N_13021,N_10073,N_11505);
nor U13022 (N_13022,N_11062,N_11924);
or U13023 (N_13023,N_10972,N_10327);
xor U13024 (N_13024,N_10495,N_10147);
or U13025 (N_13025,N_10373,N_11449);
nor U13026 (N_13026,N_10094,N_11348);
and U13027 (N_13027,N_10500,N_9229);
and U13028 (N_13028,N_10071,N_11769);
nor U13029 (N_13029,N_9641,N_9515);
xnor U13030 (N_13030,N_9567,N_11143);
nor U13031 (N_13031,N_10055,N_10523);
nor U13032 (N_13032,N_11949,N_11366);
and U13033 (N_13033,N_9174,N_11942);
or U13034 (N_13034,N_11879,N_11951);
nor U13035 (N_13035,N_9627,N_11111);
xnor U13036 (N_13036,N_10152,N_9869);
nor U13037 (N_13037,N_9349,N_9411);
nand U13038 (N_13038,N_9771,N_10602);
nor U13039 (N_13039,N_9588,N_11731);
xor U13040 (N_13040,N_10421,N_11734);
xnor U13041 (N_13041,N_9523,N_9399);
nand U13042 (N_13042,N_11747,N_11787);
or U13043 (N_13043,N_9624,N_11224);
nand U13044 (N_13044,N_11717,N_9513);
xor U13045 (N_13045,N_9211,N_9057);
nand U13046 (N_13046,N_10192,N_11067);
nand U13047 (N_13047,N_11412,N_9625);
nand U13048 (N_13048,N_9115,N_11895);
xnor U13049 (N_13049,N_10527,N_11630);
and U13050 (N_13050,N_11124,N_10242);
or U13051 (N_13051,N_9531,N_10769);
nor U13052 (N_13052,N_10547,N_10827);
and U13053 (N_13053,N_9295,N_9987);
and U13054 (N_13054,N_9995,N_9569);
and U13055 (N_13055,N_11517,N_11192);
and U13056 (N_13056,N_11527,N_11168);
xnor U13057 (N_13057,N_10246,N_10863);
nor U13058 (N_13058,N_9369,N_9891);
xnor U13059 (N_13059,N_11333,N_11013);
or U13060 (N_13060,N_10799,N_11187);
nand U13061 (N_13061,N_11998,N_9263);
or U13062 (N_13062,N_10198,N_11267);
nor U13063 (N_13063,N_9998,N_9332);
nor U13064 (N_13064,N_10061,N_9822);
or U13065 (N_13065,N_9445,N_11012);
and U13066 (N_13066,N_10154,N_11079);
and U13067 (N_13067,N_10053,N_9417);
or U13068 (N_13068,N_11158,N_11594);
xor U13069 (N_13069,N_9661,N_9323);
and U13070 (N_13070,N_9037,N_10565);
xnor U13071 (N_13071,N_9581,N_9582);
xnor U13072 (N_13072,N_10054,N_10782);
nor U13073 (N_13073,N_11154,N_11774);
or U13074 (N_13074,N_11229,N_9004);
nor U13075 (N_13075,N_11706,N_9031);
nor U13076 (N_13076,N_9054,N_11223);
xnor U13077 (N_13077,N_9809,N_9946);
and U13078 (N_13078,N_9131,N_9585);
nand U13079 (N_13079,N_9396,N_9072);
and U13080 (N_13080,N_10384,N_11831);
nand U13081 (N_13081,N_11389,N_10027);
nor U13082 (N_13082,N_11272,N_10240);
nand U13083 (N_13083,N_9719,N_11897);
nand U13084 (N_13084,N_9999,N_11454);
xor U13085 (N_13085,N_11676,N_10890);
or U13086 (N_13086,N_10956,N_9972);
xor U13087 (N_13087,N_10493,N_9090);
or U13088 (N_13088,N_11713,N_11778);
and U13089 (N_13089,N_10768,N_9192);
xnor U13090 (N_13090,N_9450,N_9644);
or U13091 (N_13091,N_10846,N_9506);
xor U13092 (N_13092,N_9094,N_9970);
and U13093 (N_13093,N_10775,N_10674);
nor U13094 (N_13094,N_9468,N_9712);
or U13095 (N_13095,N_9818,N_11340);
xor U13096 (N_13096,N_9755,N_11014);
and U13097 (N_13097,N_10590,N_11145);
nor U13098 (N_13098,N_11242,N_11927);
and U13099 (N_13099,N_9087,N_11328);
or U13100 (N_13100,N_9780,N_10442);
and U13101 (N_13101,N_9196,N_9887);
nor U13102 (N_13102,N_11076,N_11020);
and U13103 (N_13103,N_10413,N_9779);
or U13104 (N_13104,N_11833,N_11982);
and U13105 (N_13105,N_11812,N_11956);
and U13106 (N_13106,N_10292,N_11236);
nand U13107 (N_13107,N_9201,N_11873);
nand U13108 (N_13108,N_9773,N_9611);
xor U13109 (N_13109,N_9182,N_11700);
or U13110 (N_13110,N_11866,N_9034);
or U13111 (N_13111,N_11551,N_10369);
nand U13112 (N_13112,N_9839,N_10879);
nor U13113 (N_13113,N_11422,N_11872);
xnor U13114 (N_13114,N_9956,N_9108);
xnor U13115 (N_13115,N_11692,N_10616);
nor U13116 (N_13116,N_11958,N_10494);
and U13117 (N_13117,N_11174,N_10887);
xor U13118 (N_13118,N_11033,N_10554);
or U13119 (N_13119,N_10096,N_9503);
and U13120 (N_13120,N_10774,N_10942);
nand U13121 (N_13121,N_10645,N_11853);
and U13122 (N_13122,N_11737,N_11318);
or U13123 (N_13123,N_10922,N_11776);
nor U13124 (N_13124,N_11899,N_10899);
and U13125 (N_13125,N_9116,N_10226);
nand U13126 (N_13126,N_9007,N_9435);
and U13127 (N_13127,N_10976,N_9875);
and U13128 (N_13128,N_10678,N_10310);
xor U13129 (N_13129,N_10596,N_9735);
or U13130 (N_13130,N_11905,N_9350);
xor U13131 (N_13131,N_11574,N_9762);
or U13132 (N_13132,N_11303,N_11251);
xor U13133 (N_13133,N_9338,N_10311);
xor U13134 (N_13134,N_9518,N_10679);
nand U13135 (N_13135,N_10626,N_9616);
and U13136 (N_13136,N_9559,N_10998);
nor U13137 (N_13137,N_9190,N_11383);
xor U13138 (N_13138,N_10722,N_9431);
and U13139 (N_13139,N_11221,N_11719);
and U13140 (N_13140,N_11226,N_10858);
nor U13141 (N_13141,N_9107,N_9280);
nor U13142 (N_13142,N_10824,N_9181);
or U13143 (N_13143,N_11641,N_9997);
nand U13144 (N_13144,N_10669,N_10785);
nand U13145 (N_13145,N_10060,N_9135);
xnor U13146 (N_13146,N_10142,N_11558);
or U13147 (N_13147,N_10368,N_11882);
xor U13148 (N_13148,N_9610,N_10725);
xnor U13149 (N_13149,N_9493,N_10751);
nor U13150 (N_13150,N_11138,N_10562);
xor U13151 (N_13151,N_10458,N_9651);
xnor U13152 (N_13152,N_11845,N_11578);
xnor U13153 (N_13153,N_10298,N_11710);
and U13154 (N_13154,N_11611,N_9664);
xnor U13155 (N_13155,N_10430,N_9744);
nand U13156 (N_13156,N_9832,N_11669);
xnor U13157 (N_13157,N_9535,N_11894);
xnor U13158 (N_13158,N_10161,N_10882);
nand U13159 (N_13159,N_10507,N_10408);
or U13160 (N_13160,N_11914,N_11799);
and U13161 (N_13161,N_11647,N_11463);
xnor U13162 (N_13162,N_9278,N_11543);
nand U13163 (N_13163,N_11768,N_11726);
or U13164 (N_13164,N_10613,N_10231);
nor U13165 (N_13165,N_9272,N_9119);
or U13166 (N_13166,N_11583,N_10605);
nand U13167 (N_13167,N_9597,N_10643);
or U13168 (N_13168,N_11105,N_9492);
or U13169 (N_13169,N_11392,N_11332);
or U13170 (N_13170,N_11343,N_9599);
xor U13171 (N_13171,N_10149,N_9819);
or U13172 (N_13172,N_10893,N_9210);
or U13173 (N_13173,N_10459,N_9537);
nor U13174 (N_13174,N_9408,N_11976);
and U13175 (N_13175,N_11215,N_10183);
or U13176 (N_13176,N_10468,N_11596);
or U13177 (N_13177,N_11063,N_10324);
or U13178 (N_13178,N_9958,N_9335);
or U13179 (N_13179,N_11342,N_10515);
xnor U13180 (N_13180,N_9270,N_11746);
xnor U13181 (N_13181,N_9522,N_11461);
nand U13182 (N_13182,N_9226,N_11345);
and U13183 (N_13183,N_9157,N_11200);
or U13184 (N_13184,N_9062,N_11597);
or U13185 (N_13185,N_11139,N_10308);
nor U13186 (N_13186,N_10650,N_10770);
xnor U13187 (N_13187,N_9398,N_9633);
nand U13188 (N_13188,N_11406,N_10615);
nand U13189 (N_13189,N_11263,N_11579);
xnor U13190 (N_13190,N_10724,N_10530);
nand U13191 (N_13191,N_11978,N_10912);
xnor U13192 (N_13192,N_10257,N_11628);
or U13193 (N_13193,N_10534,N_11535);
nor U13194 (N_13194,N_11497,N_9071);
and U13195 (N_13195,N_9614,N_10271);
nor U13196 (N_13196,N_9045,N_11516);
and U13197 (N_13197,N_9441,N_10862);
and U13198 (N_13198,N_11962,N_10739);
nor U13199 (N_13199,N_10780,N_10155);
xor U13200 (N_13200,N_10380,N_10052);
and U13201 (N_13201,N_9704,N_10447);
xor U13202 (N_13202,N_10842,N_9320);
xor U13203 (N_13203,N_9540,N_10476);
or U13204 (N_13204,N_10406,N_9470);
nor U13205 (N_13205,N_11575,N_10531);
nor U13206 (N_13206,N_9570,N_10486);
or U13207 (N_13207,N_9284,N_11504);
and U13208 (N_13208,N_11437,N_10020);
and U13209 (N_13209,N_10803,N_9991);
nand U13210 (N_13210,N_10601,N_9696);
nor U13211 (N_13211,N_9245,N_10237);
nand U13212 (N_13212,N_9307,N_10712);
nor U13213 (N_13213,N_9593,N_9312);
or U13214 (N_13214,N_11758,N_11818);
and U13215 (N_13215,N_10773,N_11775);
nor U13216 (N_13216,N_11753,N_10016);
nand U13217 (N_13217,N_11370,N_10241);
xnor U13218 (N_13218,N_11087,N_11417);
nand U13219 (N_13219,N_11571,N_11397);
xor U13220 (N_13220,N_9250,N_9296);
nor U13221 (N_13221,N_10199,N_9924);
nor U13222 (N_13222,N_9147,N_11495);
and U13223 (N_13223,N_9234,N_10704);
xor U13224 (N_13224,N_9125,N_10996);
or U13225 (N_13225,N_9754,N_10623);
and U13226 (N_13226,N_10402,N_11673);
nand U13227 (N_13227,N_10568,N_11092);
and U13228 (N_13228,N_10759,N_11253);
nand U13229 (N_13229,N_9070,N_11502);
xnor U13230 (N_13230,N_11324,N_11289);
nand U13231 (N_13231,N_9462,N_10136);
xor U13232 (N_13232,N_10163,N_11393);
nand U13233 (N_13233,N_11629,N_11258);
xor U13234 (N_13234,N_10953,N_11974);
or U13235 (N_13235,N_9895,N_9572);
xor U13236 (N_13236,N_10968,N_10033);
and U13237 (N_13237,N_10753,N_9352);
nand U13238 (N_13238,N_11477,N_10664);
or U13239 (N_13239,N_11361,N_11970);
xnor U13240 (N_13240,N_9351,N_9821);
nor U13241 (N_13241,N_11983,N_11466);
xor U13242 (N_13242,N_10509,N_9882);
nor U13243 (N_13243,N_9702,N_11687);
nor U13244 (N_13244,N_11598,N_10272);
nor U13245 (N_13245,N_10817,N_10418);
xor U13246 (N_13246,N_11365,N_11619);
or U13247 (N_13247,N_11418,N_9927);
and U13248 (N_13248,N_11722,N_10957);
nor U13249 (N_13249,N_11142,N_11483);
and U13250 (N_13250,N_9966,N_10632);
or U13251 (N_13251,N_11484,N_10984);
or U13252 (N_13252,N_10042,N_11048);
nand U13253 (N_13253,N_9061,N_10404);
and U13254 (N_13254,N_10439,N_9556);
or U13255 (N_13255,N_9568,N_11524);
xor U13256 (N_13256,N_11065,N_9276);
nand U13257 (N_13257,N_11045,N_11448);
nor U13258 (N_13258,N_11308,N_11374);
nand U13259 (N_13259,N_11498,N_11518);
nor U13260 (N_13260,N_9286,N_11606);
or U13261 (N_13261,N_11840,N_9817);
xor U13262 (N_13262,N_9077,N_9706);
nand U13263 (N_13263,N_10113,N_11782);
or U13264 (N_13264,N_9763,N_11632);
nor U13265 (N_13265,N_11740,N_9035);
nor U13266 (N_13266,N_10222,N_11085);
nor U13267 (N_13267,N_9110,N_11043);
nor U13268 (N_13268,N_9514,N_10916);
nand U13269 (N_13269,N_10844,N_10975);
and U13270 (N_13270,N_9382,N_10330);
nor U13271 (N_13271,N_11580,N_9361);
and U13272 (N_13272,N_10680,N_9074);
xor U13273 (N_13273,N_11844,N_9751);
nor U13274 (N_13274,N_10837,N_11314);
nor U13275 (N_13275,N_10719,N_9008);
xor U13276 (N_13276,N_10888,N_10610);
xnor U13277 (N_13277,N_11419,N_10049);
nand U13278 (N_13278,N_10031,N_10119);
xor U13279 (N_13279,N_9155,N_11313);
nand U13280 (N_13280,N_10627,N_10818);
and U13281 (N_13281,N_11529,N_10595);
nand U13282 (N_13282,N_11765,N_9750);
or U13283 (N_13283,N_10607,N_11697);
nand U13284 (N_13284,N_10282,N_11206);
or U13285 (N_13285,N_9384,N_10789);
nand U13286 (N_13286,N_10303,N_11388);
nand U13287 (N_13287,N_9603,N_9864);
and U13288 (N_13288,N_10737,N_11377);
xnor U13289 (N_13289,N_11814,N_11990);
and U13290 (N_13290,N_9620,N_10902);
xor U13291 (N_13291,N_10625,N_9342);
and U13292 (N_13292,N_11662,N_11094);
or U13293 (N_13293,N_9159,N_9876);
xnor U13294 (N_13294,N_9699,N_11671);
nor U13295 (N_13295,N_9739,N_10924);
nor U13296 (N_13296,N_11929,N_9252);
nand U13297 (N_13297,N_11295,N_10668);
nand U13298 (N_13298,N_10389,N_10201);
and U13299 (N_13299,N_9798,N_9413);
or U13300 (N_13300,N_9989,N_9454);
and U13301 (N_13301,N_11129,N_10376);
nor U13302 (N_13302,N_10651,N_11635);
xnor U13303 (N_13303,N_10675,N_9734);
and U13304 (N_13304,N_9730,N_11510);
nor U13305 (N_13305,N_10648,N_9865);
nand U13306 (N_13306,N_9682,N_11250);
and U13307 (N_13307,N_10287,N_11479);
or U13308 (N_13308,N_11759,N_9715);
nand U13309 (N_13309,N_10850,N_9653);
nor U13310 (N_13310,N_10158,N_10008);
or U13311 (N_13311,N_11908,N_9339);
and U13312 (N_13312,N_10526,N_10438);
nor U13313 (N_13313,N_9109,N_11724);
xnor U13314 (N_13314,N_11980,N_10348);
nor U13315 (N_13315,N_11037,N_9792);
nand U13316 (N_13316,N_9810,N_11008);
nand U13317 (N_13317,N_9478,N_11413);
or U13318 (N_13318,N_11777,N_9301);
nor U13319 (N_13319,N_11946,N_11177);
and U13320 (N_13320,N_10004,N_9793);
nor U13321 (N_13321,N_10723,N_9703);
xor U13322 (N_13322,N_11000,N_10329);
or U13323 (N_13323,N_9388,N_11898);
or U13324 (N_13324,N_9051,N_11058);
or U13325 (N_13325,N_10847,N_10790);
and U13326 (N_13326,N_11965,N_9993);
nand U13327 (N_13327,N_9277,N_11773);
nor U13328 (N_13328,N_10009,N_11876);
xor U13329 (N_13329,N_9677,N_9319);
nand U13330 (N_13330,N_11197,N_11514);
and U13331 (N_13331,N_9315,N_11100);
and U13332 (N_13332,N_9685,N_10788);
xnor U13333 (N_13333,N_10169,N_10295);
xnor U13334 (N_13334,N_10993,N_11084);
xor U13335 (N_13335,N_9145,N_10164);
and U13336 (N_13336,N_11608,N_11939);
nand U13337 (N_13337,N_9659,N_11783);
or U13338 (N_13338,N_10135,N_10779);
or U13339 (N_13339,N_10172,N_11171);
and U13340 (N_13340,N_10145,N_11867);
nand U13341 (N_13341,N_10355,N_11496);
and U13342 (N_13342,N_11729,N_11060);
xor U13343 (N_13343,N_10673,N_10995);
nand U13344 (N_13344,N_11098,N_9105);
xnor U13345 (N_13345,N_10289,N_10767);
or U13346 (N_13346,N_11672,N_10461);
or U13347 (N_13347,N_9698,N_9571);
nor U13348 (N_13348,N_10611,N_11363);
nand U13349 (N_13349,N_11588,N_10143);
or U13350 (N_13350,N_10123,N_10426);
nor U13351 (N_13351,N_10092,N_11364);
nor U13352 (N_13352,N_9918,N_11445);
xnor U13353 (N_13353,N_11460,N_9733);
nor U13354 (N_13354,N_10432,N_10419);
nand U13355 (N_13355,N_10730,N_10014);
xor U13356 (N_13356,N_9551,N_9264);
nand U13357 (N_13357,N_11555,N_10806);
or U13358 (N_13358,N_11624,N_11923);
or U13359 (N_13359,N_10732,N_11052);
and U13360 (N_13360,N_11426,N_10947);
xnor U13361 (N_13361,N_9448,N_10915);
and U13362 (N_13362,N_11515,N_9491);
nor U13363 (N_13363,N_9180,N_11864);
xnor U13364 (N_13364,N_10309,N_9409);
nor U13365 (N_13365,N_11733,N_11244);
xor U13366 (N_13366,N_9242,N_10254);
and U13367 (N_13367,N_11344,N_10905);
xnor U13368 (N_13368,N_10546,N_11274);
and U13369 (N_13369,N_10577,N_11091);
nand U13370 (N_13370,N_10985,N_10784);
nand U13371 (N_13371,N_9063,N_10982);
or U13372 (N_13372,N_11755,N_10855);
nor U13373 (N_13373,N_10479,N_10519);
xor U13374 (N_13374,N_11341,N_10107);
xnor U13375 (N_13375,N_10188,N_10335);
nor U13376 (N_13376,N_10392,N_10925);
and U13377 (N_13377,N_10608,N_11689);
nor U13378 (N_13378,N_11567,N_9816);
nand U13379 (N_13379,N_10787,N_11195);
and U13380 (N_13380,N_9564,N_9901);
and U13381 (N_13381,N_11464,N_10283);
nor U13382 (N_13382,N_9511,N_10594);
nor U13383 (N_13383,N_11494,N_11933);
xor U13384 (N_13384,N_9555,N_11041);
nor U13385 (N_13385,N_9197,N_11749);
nor U13386 (N_13386,N_9601,N_11964);
nor U13387 (N_13387,N_10644,N_11458);
nand U13388 (N_13388,N_10955,N_11857);
or U13389 (N_13389,N_11278,N_10963);
and U13390 (N_13390,N_9558,N_9992);
or U13391 (N_13391,N_9249,N_9393);
and U13392 (N_13392,N_11440,N_10923);
and U13393 (N_13393,N_10771,N_9299);
xnor U13394 (N_13394,N_9305,N_10740);
and U13395 (N_13395,N_9334,N_10162);
nor U13396 (N_13396,N_11642,N_11988);
xor U13397 (N_13397,N_10437,N_9543);
and U13398 (N_13398,N_9604,N_11666);
and U13399 (N_13399,N_10074,N_11536);
and U13400 (N_13400,N_9488,N_10181);
and U13401 (N_13401,N_9158,N_10089);
or U13402 (N_13402,N_9304,N_11209);
or U13403 (N_13403,N_9367,N_10480);
xor U13404 (N_13404,N_11444,N_10940);
nor U13405 (N_13405,N_9316,N_10805);
nand U13406 (N_13406,N_9096,N_10316);
nor U13407 (N_13407,N_11260,N_9444);
nor U13408 (N_13408,N_9097,N_11918);
xor U13409 (N_13409,N_10299,N_11248);
nand U13410 (N_13410,N_9415,N_9881);
nor U13411 (N_13411,N_9081,N_10635);
nand U13412 (N_13412,N_9227,N_11718);
nand U13413 (N_13413,N_9113,N_10208);
xor U13414 (N_13414,N_11874,N_11053);
or U13415 (N_13415,N_11670,N_10583);
and U13416 (N_13416,N_9736,N_11725);
and U13417 (N_13417,N_10440,N_10582);
xor U13418 (N_13418,N_9767,N_10363);
xor U13419 (N_13419,N_9271,N_11352);
xor U13420 (N_13420,N_10366,N_11938);
and U13421 (N_13421,N_10156,N_9080);
nand U13422 (N_13422,N_11161,N_10559);
nor U13423 (N_13423,N_9359,N_11566);
nor U13424 (N_13424,N_9738,N_11004);
nor U13425 (N_13425,N_9857,N_9344);
nand U13426 (N_13426,N_10005,N_10485);
nor U13427 (N_13427,N_10034,N_9387);
xnor U13428 (N_13428,N_10276,N_10395);
nand U13429 (N_13429,N_9141,N_11957);
nand U13430 (N_13430,N_11537,N_11655);
nor U13431 (N_13431,N_9186,N_11097);
and U13432 (N_13432,N_11175,N_11622);
xor U13433 (N_13433,N_11453,N_11804);
or U13434 (N_13434,N_10516,N_9017);
or U13435 (N_13435,N_9016,N_11911);
or U13436 (N_13436,N_9814,N_9892);
nand U13437 (N_13437,N_11490,N_11279);
or U13438 (N_13438,N_11151,N_9621);
or U13439 (N_13439,N_10691,N_9753);
nor U13440 (N_13440,N_11349,N_11526);
xor U13441 (N_13441,N_9292,N_11070);
nand U13442 (N_13442,N_11860,N_9820);
and U13443 (N_13443,N_9951,N_10907);
or U13444 (N_13444,N_10835,N_10273);
or U13445 (N_13445,N_9795,N_11792);
nand U13446 (N_13446,N_10911,N_11456);
or U13447 (N_13447,N_10944,N_9258);
and U13448 (N_13448,N_11959,N_11926);
and U13449 (N_13449,N_9404,N_9122);
nor U13450 (N_13450,N_11525,N_10184);
or U13451 (N_13451,N_11837,N_11047);
or U13452 (N_13452,N_9605,N_9311);
and U13453 (N_13453,N_10090,N_10791);
xor U13454 (N_13454,N_11519,N_10403);
or U13455 (N_13455,N_9639,N_9510);
or U13456 (N_13456,N_10235,N_10709);
or U13457 (N_13457,N_10585,N_11446);
nor U13458 (N_13458,N_10455,N_11101);
nand U13459 (N_13459,N_10959,N_11652);
nand U13460 (N_13460,N_10434,N_9216);
xnor U13461 (N_13461,N_10243,N_10981);
nand U13462 (N_13462,N_11907,N_11469);
and U13463 (N_13463,N_10943,N_10670);
xnor U13464 (N_13464,N_10677,N_9920);
and U13465 (N_13465,N_11358,N_9803);
or U13466 (N_13466,N_9879,N_10187);
and U13467 (N_13467,N_10124,N_11618);
xor U13468 (N_13468,N_9423,N_10150);
or U13469 (N_13469,N_10173,N_9265);
or U13470 (N_13470,N_10634,N_9521);
xor U13471 (N_13471,N_11489,N_9628);
nor U13472 (N_13472,N_10488,N_10860);
nand U13473 (N_13473,N_11132,N_10830);
or U13474 (N_13474,N_9204,N_10852);
or U13475 (N_13475,N_11351,N_11276);
nor U13476 (N_13476,N_9697,N_9908);
and U13477 (N_13477,N_10783,N_9957);
xor U13478 (N_13478,N_9000,N_11623);
or U13479 (N_13479,N_10600,N_10011);
xnor U13480 (N_13480,N_11533,N_9333);
nand U13481 (N_13481,N_11284,N_11829);
and U13482 (N_13482,N_9916,N_9375);
and U13483 (N_13483,N_9020,N_11616);
nor U13484 (N_13484,N_9874,N_9536);
nand U13485 (N_13485,N_10186,N_11216);
nor U13486 (N_13486,N_11071,N_10696);
xnor U13487 (N_13487,N_11222,N_9642);
nor U13488 (N_13488,N_11565,N_10013);
or U13489 (N_13489,N_10414,N_10505);
and U13490 (N_13490,N_10738,N_11292);
nor U13491 (N_13491,N_10203,N_11693);
or U13492 (N_13492,N_9996,N_10988);
or U13493 (N_13493,N_11602,N_9254);
or U13494 (N_13494,N_10766,N_9104);
nand U13495 (N_13495,N_9917,N_10700);
xor U13496 (N_13496,N_10098,N_9714);
and U13497 (N_13497,N_11650,N_9790);
and U13498 (N_13498,N_9241,N_10885);
nor U13499 (N_13499,N_11909,N_11046);
nor U13500 (N_13500,N_10305,N_10533);
xnor U13501 (N_13501,N_9870,N_9364);
or U13502 (N_13502,N_9133,N_9201);
nor U13503 (N_13503,N_10577,N_9925);
nor U13504 (N_13504,N_10166,N_9734);
xnor U13505 (N_13505,N_10693,N_10353);
nor U13506 (N_13506,N_10316,N_9409);
xnor U13507 (N_13507,N_9353,N_10886);
xor U13508 (N_13508,N_11286,N_10414);
nand U13509 (N_13509,N_11433,N_9446);
nand U13510 (N_13510,N_10926,N_9219);
xor U13511 (N_13511,N_9539,N_11711);
nand U13512 (N_13512,N_10984,N_11277);
nand U13513 (N_13513,N_10367,N_10314);
xnor U13514 (N_13514,N_10830,N_9942);
xor U13515 (N_13515,N_9009,N_11616);
xor U13516 (N_13516,N_9704,N_11197);
nand U13517 (N_13517,N_10424,N_11163);
or U13518 (N_13518,N_9965,N_10998);
nand U13519 (N_13519,N_9201,N_10710);
xor U13520 (N_13520,N_9421,N_9446);
and U13521 (N_13521,N_10654,N_10883);
nand U13522 (N_13522,N_10835,N_11768);
or U13523 (N_13523,N_10883,N_11618);
nor U13524 (N_13524,N_10188,N_11099);
xnor U13525 (N_13525,N_11798,N_10290);
and U13526 (N_13526,N_11996,N_11671);
nand U13527 (N_13527,N_10560,N_10544);
and U13528 (N_13528,N_10390,N_11202);
xnor U13529 (N_13529,N_10838,N_11408);
and U13530 (N_13530,N_10660,N_10617);
or U13531 (N_13531,N_9681,N_11362);
nor U13532 (N_13532,N_11828,N_10721);
or U13533 (N_13533,N_10948,N_9883);
nor U13534 (N_13534,N_11137,N_11478);
nor U13535 (N_13535,N_10471,N_10361);
or U13536 (N_13536,N_9628,N_10274);
and U13537 (N_13537,N_10289,N_11969);
xor U13538 (N_13538,N_9405,N_11985);
nand U13539 (N_13539,N_10334,N_10843);
nor U13540 (N_13540,N_11843,N_10774);
and U13541 (N_13541,N_10763,N_9319);
xor U13542 (N_13542,N_11074,N_9127);
xor U13543 (N_13543,N_9772,N_10338);
nand U13544 (N_13544,N_10852,N_9786);
xor U13545 (N_13545,N_9904,N_9130);
nand U13546 (N_13546,N_11349,N_10156);
nand U13547 (N_13547,N_9923,N_11352);
or U13548 (N_13548,N_11082,N_9098);
xnor U13549 (N_13549,N_10047,N_9500);
xnor U13550 (N_13550,N_9699,N_10379);
nor U13551 (N_13551,N_10617,N_9565);
xnor U13552 (N_13552,N_9630,N_9027);
nand U13553 (N_13553,N_11391,N_11453);
or U13554 (N_13554,N_11664,N_10906);
nor U13555 (N_13555,N_10751,N_11623);
or U13556 (N_13556,N_9939,N_9301);
nor U13557 (N_13557,N_11920,N_11577);
and U13558 (N_13558,N_9067,N_11189);
and U13559 (N_13559,N_10240,N_10340);
nor U13560 (N_13560,N_10800,N_11365);
xnor U13561 (N_13561,N_9441,N_9596);
xnor U13562 (N_13562,N_9815,N_11854);
nand U13563 (N_13563,N_9917,N_11187);
or U13564 (N_13564,N_9196,N_9527);
nor U13565 (N_13565,N_11616,N_11338);
nand U13566 (N_13566,N_10176,N_11814);
or U13567 (N_13567,N_9969,N_9525);
xnor U13568 (N_13568,N_11190,N_9550);
or U13569 (N_13569,N_10441,N_11832);
nor U13570 (N_13570,N_11333,N_10679);
and U13571 (N_13571,N_11796,N_9904);
nand U13572 (N_13572,N_10371,N_9081);
nand U13573 (N_13573,N_9530,N_10023);
xor U13574 (N_13574,N_10778,N_9511);
nor U13575 (N_13575,N_11149,N_9696);
nor U13576 (N_13576,N_9049,N_9359);
xor U13577 (N_13577,N_9037,N_9926);
xnor U13578 (N_13578,N_10722,N_10360);
xor U13579 (N_13579,N_10138,N_10019);
nor U13580 (N_13580,N_11860,N_9788);
and U13581 (N_13581,N_11283,N_10978);
or U13582 (N_13582,N_10767,N_10532);
and U13583 (N_13583,N_10560,N_9801);
nor U13584 (N_13584,N_9481,N_10603);
xnor U13585 (N_13585,N_11694,N_10707);
or U13586 (N_13586,N_9115,N_11663);
nor U13587 (N_13587,N_10297,N_9996);
or U13588 (N_13588,N_11513,N_9024);
xor U13589 (N_13589,N_10149,N_9933);
nor U13590 (N_13590,N_10825,N_11489);
or U13591 (N_13591,N_11883,N_9701);
and U13592 (N_13592,N_10924,N_10808);
nand U13593 (N_13593,N_9306,N_10954);
and U13594 (N_13594,N_11055,N_11726);
xnor U13595 (N_13595,N_9497,N_9171);
xor U13596 (N_13596,N_10851,N_11944);
nor U13597 (N_13597,N_9515,N_10991);
nand U13598 (N_13598,N_10857,N_9622);
nor U13599 (N_13599,N_9945,N_10025);
nand U13600 (N_13600,N_9572,N_10665);
or U13601 (N_13601,N_9727,N_11420);
or U13602 (N_13602,N_11202,N_9654);
nor U13603 (N_13603,N_11823,N_9852);
nor U13604 (N_13604,N_9903,N_9936);
or U13605 (N_13605,N_10539,N_9185);
xor U13606 (N_13606,N_9376,N_10218);
nor U13607 (N_13607,N_11769,N_9335);
nor U13608 (N_13608,N_10609,N_9389);
nor U13609 (N_13609,N_11426,N_9224);
or U13610 (N_13610,N_11557,N_10434);
and U13611 (N_13611,N_11862,N_9475);
and U13612 (N_13612,N_9351,N_10210);
and U13613 (N_13613,N_11154,N_10196);
or U13614 (N_13614,N_10290,N_9207);
nor U13615 (N_13615,N_10905,N_11267);
nand U13616 (N_13616,N_10625,N_11981);
nor U13617 (N_13617,N_9395,N_9739);
and U13618 (N_13618,N_10719,N_11858);
nand U13619 (N_13619,N_10420,N_11823);
or U13620 (N_13620,N_9611,N_11508);
nand U13621 (N_13621,N_11272,N_9382);
or U13622 (N_13622,N_10208,N_9812);
or U13623 (N_13623,N_11914,N_10888);
and U13624 (N_13624,N_10050,N_11447);
nand U13625 (N_13625,N_11387,N_10842);
nor U13626 (N_13626,N_10743,N_9991);
or U13627 (N_13627,N_10652,N_10315);
nand U13628 (N_13628,N_11007,N_9316);
and U13629 (N_13629,N_9585,N_10151);
nor U13630 (N_13630,N_11863,N_9892);
nand U13631 (N_13631,N_11062,N_11899);
and U13632 (N_13632,N_10831,N_11564);
and U13633 (N_13633,N_11753,N_10113);
and U13634 (N_13634,N_11312,N_11810);
xnor U13635 (N_13635,N_9189,N_11978);
xor U13636 (N_13636,N_9677,N_10136);
or U13637 (N_13637,N_10985,N_10240);
or U13638 (N_13638,N_11118,N_11571);
nand U13639 (N_13639,N_10993,N_10280);
nand U13640 (N_13640,N_11314,N_11495);
nand U13641 (N_13641,N_9457,N_10847);
xor U13642 (N_13642,N_9713,N_10101);
nor U13643 (N_13643,N_9160,N_9391);
and U13644 (N_13644,N_9380,N_9678);
nor U13645 (N_13645,N_9963,N_11859);
xor U13646 (N_13646,N_10014,N_9035);
nor U13647 (N_13647,N_10325,N_11374);
xnor U13648 (N_13648,N_10774,N_9987);
nand U13649 (N_13649,N_10525,N_11109);
and U13650 (N_13650,N_10720,N_9272);
nor U13651 (N_13651,N_10659,N_11731);
nor U13652 (N_13652,N_9024,N_11200);
nand U13653 (N_13653,N_9939,N_10563);
nor U13654 (N_13654,N_10955,N_11177);
or U13655 (N_13655,N_10589,N_10022);
nand U13656 (N_13656,N_10828,N_9857);
nor U13657 (N_13657,N_9622,N_10344);
and U13658 (N_13658,N_11579,N_10365);
or U13659 (N_13659,N_9748,N_10823);
and U13660 (N_13660,N_11924,N_9106);
xor U13661 (N_13661,N_9194,N_10802);
xnor U13662 (N_13662,N_10014,N_11124);
nor U13663 (N_13663,N_9397,N_9347);
or U13664 (N_13664,N_9719,N_11312);
or U13665 (N_13665,N_9072,N_10157);
nor U13666 (N_13666,N_9171,N_10812);
nor U13667 (N_13667,N_10696,N_11956);
and U13668 (N_13668,N_10857,N_11813);
nand U13669 (N_13669,N_11158,N_9011);
or U13670 (N_13670,N_9913,N_9245);
and U13671 (N_13671,N_11170,N_11749);
and U13672 (N_13672,N_10201,N_11196);
xnor U13673 (N_13673,N_9580,N_11423);
xor U13674 (N_13674,N_11343,N_10842);
xor U13675 (N_13675,N_10289,N_10197);
and U13676 (N_13676,N_10688,N_11610);
xnor U13677 (N_13677,N_9235,N_10037);
and U13678 (N_13678,N_11521,N_10638);
and U13679 (N_13679,N_9236,N_10374);
nand U13680 (N_13680,N_11466,N_9791);
nor U13681 (N_13681,N_10230,N_9294);
nor U13682 (N_13682,N_10918,N_11028);
nor U13683 (N_13683,N_10800,N_9596);
and U13684 (N_13684,N_10887,N_9371);
nand U13685 (N_13685,N_10830,N_9653);
and U13686 (N_13686,N_10297,N_10924);
nor U13687 (N_13687,N_11150,N_9808);
or U13688 (N_13688,N_9438,N_11987);
or U13689 (N_13689,N_10268,N_11190);
xnor U13690 (N_13690,N_11633,N_9586);
nand U13691 (N_13691,N_11391,N_9295);
or U13692 (N_13692,N_10348,N_11759);
and U13693 (N_13693,N_10892,N_9339);
or U13694 (N_13694,N_10613,N_9042);
nand U13695 (N_13695,N_9032,N_10880);
and U13696 (N_13696,N_11417,N_9296);
and U13697 (N_13697,N_11326,N_11110);
and U13698 (N_13698,N_11633,N_11003);
xnor U13699 (N_13699,N_9073,N_10441);
or U13700 (N_13700,N_11517,N_9417);
or U13701 (N_13701,N_9814,N_9808);
nor U13702 (N_13702,N_11260,N_10970);
nor U13703 (N_13703,N_10587,N_11106);
nor U13704 (N_13704,N_10262,N_11453);
or U13705 (N_13705,N_11280,N_10804);
xor U13706 (N_13706,N_11676,N_11983);
nor U13707 (N_13707,N_11405,N_10029);
or U13708 (N_13708,N_11722,N_9878);
or U13709 (N_13709,N_9953,N_10350);
and U13710 (N_13710,N_10854,N_10029);
nand U13711 (N_13711,N_10474,N_9123);
xor U13712 (N_13712,N_10528,N_9662);
or U13713 (N_13713,N_11950,N_11299);
xnor U13714 (N_13714,N_11597,N_11818);
xnor U13715 (N_13715,N_11169,N_10353);
nor U13716 (N_13716,N_11256,N_11511);
and U13717 (N_13717,N_11225,N_10950);
and U13718 (N_13718,N_11650,N_9709);
nor U13719 (N_13719,N_11444,N_11348);
nand U13720 (N_13720,N_10169,N_9486);
nor U13721 (N_13721,N_10003,N_9641);
and U13722 (N_13722,N_11860,N_10289);
nor U13723 (N_13723,N_9787,N_9855);
or U13724 (N_13724,N_11491,N_10340);
or U13725 (N_13725,N_10825,N_11514);
or U13726 (N_13726,N_10732,N_11432);
or U13727 (N_13727,N_10008,N_10099);
or U13728 (N_13728,N_11337,N_9536);
or U13729 (N_13729,N_10917,N_10107);
nor U13730 (N_13730,N_9901,N_10621);
nand U13731 (N_13731,N_10131,N_10298);
xnor U13732 (N_13732,N_9271,N_9712);
and U13733 (N_13733,N_10679,N_9688);
and U13734 (N_13734,N_11444,N_9055);
and U13735 (N_13735,N_9431,N_11306);
nor U13736 (N_13736,N_11256,N_9846);
nand U13737 (N_13737,N_11094,N_10400);
xnor U13738 (N_13738,N_10695,N_11500);
and U13739 (N_13739,N_10504,N_10828);
nor U13740 (N_13740,N_9534,N_10586);
nor U13741 (N_13741,N_11424,N_9260);
and U13742 (N_13742,N_9925,N_9133);
nor U13743 (N_13743,N_9557,N_11624);
nand U13744 (N_13744,N_9344,N_9998);
nor U13745 (N_13745,N_9353,N_10513);
nand U13746 (N_13746,N_11564,N_10187);
nand U13747 (N_13747,N_9501,N_10396);
xnor U13748 (N_13748,N_10238,N_11649);
xnor U13749 (N_13749,N_9919,N_10432);
xor U13750 (N_13750,N_10670,N_10987);
nand U13751 (N_13751,N_11512,N_11830);
and U13752 (N_13752,N_9878,N_11377);
nand U13753 (N_13753,N_10161,N_9562);
nor U13754 (N_13754,N_9259,N_10499);
and U13755 (N_13755,N_11366,N_9996);
nand U13756 (N_13756,N_11334,N_10379);
and U13757 (N_13757,N_9565,N_11238);
xnor U13758 (N_13758,N_9641,N_9203);
xnor U13759 (N_13759,N_9288,N_9046);
xnor U13760 (N_13760,N_9787,N_9043);
xor U13761 (N_13761,N_10646,N_9618);
nand U13762 (N_13762,N_10368,N_11914);
or U13763 (N_13763,N_11615,N_10093);
and U13764 (N_13764,N_9658,N_9299);
or U13765 (N_13765,N_11284,N_9088);
or U13766 (N_13766,N_9556,N_11186);
nor U13767 (N_13767,N_11039,N_9946);
or U13768 (N_13768,N_9737,N_10062);
xor U13769 (N_13769,N_9067,N_10244);
nor U13770 (N_13770,N_9915,N_10421);
or U13771 (N_13771,N_9903,N_9247);
xnor U13772 (N_13772,N_9898,N_11223);
xnor U13773 (N_13773,N_11789,N_11094);
xor U13774 (N_13774,N_9445,N_9919);
nor U13775 (N_13775,N_11973,N_10139);
xnor U13776 (N_13776,N_10922,N_10084);
or U13777 (N_13777,N_10194,N_11024);
xor U13778 (N_13778,N_10042,N_9043);
or U13779 (N_13779,N_11933,N_9605);
nand U13780 (N_13780,N_9668,N_9246);
nand U13781 (N_13781,N_10020,N_9150);
nand U13782 (N_13782,N_11995,N_11274);
or U13783 (N_13783,N_9508,N_10442);
or U13784 (N_13784,N_11915,N_10857);
xor U13785 (N_13785,N_10711,N_11730);
nand U13786 (N_13786,N_11646,N_11497);
or U13787 (N_13787,N_11032,N_10798);
xor U13788 (N_13788,N_10048,N_11051);
nand U13789 (N_13789,N_10772,N_10415);
or U13790 (N_13790,N_11706,N_11635);
and U13791 (N_13791,N_10975,N_9701);
or U13792 (N_13792,N_9734,N_9750);
xnor U13793 (N_13793,N_10536,N_9582);
nand U13794 (N_13794,N_10411,N_9030);
and U13795 (N_13795,N_10740,N_11248);
or U13796 (N_13796,N_10934,N_10503);
or U13797 (N_13797,N_9975,N_9754);
and U13798 (N_13798,N_10561,N_9485);
nand U13799 (N_13799,N_10565,N_11182);
nor U13800 (N_13800,N_10462,N_9834);
and U13801 (N_13801,N_10731,N_10148);
and U13802 (N_13802,N_10504,N_9649);
or U13803 (N_13803,N_11767,N_11917);
xnor U13804 (N_13804,N_11344,N_11293);
xor U13805 (N_13805,N_9505,N_10662);
nand U13806 (N_13806,N_9748,N_10333);
or U13807 (N_13807,N_9154,N_11897);
nor U13808 (N_13808,N_10134,N_9760);
or U13809 (N_13809,N_10878,N_10624);
xor U13810 (N_13810,N_11123,N_11623);
and U13811 (N_13811,N_10444,N_9473);
nor U13812 (N_13812,N_9578,N_11385);
xnor U13813 (N_13813,N_10177,N_10534);
nor U13814 (N_13814,N_9381,N_10764);
nor U13815 (N_13815,N_10304,N_9078);
nor U13816 (N_13816,N_9645,N_10517);
xor U13817 (N_13817,N_10565,N_10403);
nor U13818 (N_13818,N_11143,N_9588);
nand U13819 (N_13819,N_9808,N_10224);
or U13820 (N_13820,N_11639,N_9094);
xnor U13821 (N_13821,N_10390,N_10108);
nor U13822 (N_13822,N_11429,N_9175);
nor U13823 (N_13823,N_9891,N_10597);
nor U13824 (N_13824,N_9331,N_9152);
nand U13825 (N_13825,N_10260,N_10689);
nor U13826 (N_13826,N_11841,N_11274);
and U13827 (N_13827,N_9880,N_10888);
nor U13828 (N_13828,N_11239,N_9054);
nand U13829 (N_13829,N_9066,N_10516);
or U13830 (N_13830,N_10157,N_10580);
nor U13831 (N_13831,N_9855,N_9466);
nor U13832 (N_13832,N_9612,N_9497);
nor U13833 (N_13833,N_9920,N_11968);
xor U13834 (N_13834,N_11113,N_11667);
xor U13835 (N_13835,N_10802,N_10468);
nand U13836 (N_13836,N_10148,N_9835);
or U13837 (N_13837,N_9059,N_9815);
and U13838 (N_13838,N_9687,N_11004);
nand U13839 (N_13839,N_9679,N_9084);
nor U13840 (N_13840,N_11757,N_9390);
nand U13841 (N_13841,N_9082,N_11851);
nand U13842 (N_13842,N_10672,N_10879);
nor U13843 (N_13843,N_11038,N_10514);
and U13844 (N_13844,N_9652,N_10952);
nor U13845 (N_13845,N_10607,N_10526);
xor U13846 (N_13846,N_9015,N_9804);
or U13847 (N_13847,N_10140,N_11875);
xor U13848 (N_13848,N_9807,N_11178);
nand U13849 (N_13849,N_10805,N_11618);
nor U13850 (N_13850,N_9581,N_10808);
xor U13851 (N_13851,N_9013,N_11191);
or U13852 (N_13852,N_11412,N_11220);
nand U13853 (N_13853,N_9222,N_9111);
xor U13854 (N_13854,N_9143,N_10077);
or U13855 (N_13855,N_10587,N_11229);
nand U13856 (N_13856,N_11677,N_9292);
nand U13857 (N_13857,N_9407,N_11222);
nor U13858 (N_13858,N_10247,N_9707);
xor U13859 (N_13859,N_11286,N_9563);
nor U13860 (N_13860,N_9940,N_11844);
and U13861 (N_13861,N_11054,N_11308);
or U13862 (N_13862,N_9320,N_10576);
or U13863 (N_13863,N_9333,N_9692);
nor U13864 (N_13864,N_11973,N_9376);
nor U13865 (N_13865,N_9519,N_9143);
or U13866 (N_13866,N_9298,N_10575);
xnor U13867 (N_13867,N_11545,N_11707);
and U13868 (N_13868,N_11538,N_11292);
nor U13869 (N_13869,N_11603,N_11459);
nor U13870 (N_13870,N_9806,N_9454);
xnor U13871 (N_13871,N_9980,N_10284);
or U13872 (N_13872,N_9950,N_10808);
or U13873 (N_13873,N_11797,N_11387);
or U13874 (N_13874,N_10895,N_11850);
xnor U13875 (N_13875,N_10327,N_10918);
xor U13876 (N_13876,N_10960,N_9913);
nand U13877 (N_13877,N_9519,N_11232);
nand U13878 (N_13878,N_9850,N_10739);
nor U13879 (N_13879,N_9939,N_10585);
or U13880 (N_13880,N_11714,N_11927);
and U13881 (N_13881,N_11477,N_11480);
nand U13882 (N_13882,N_11007,N_10597);
nor U13883 (N_13883,N_11167,N_10975);
or U13884 (N_13884,N_10253,N_10752);
nand U13885 (N_13885,N_11529,N_9812);
and U13886 (N_13886,N_11212,N_10012);
nand U13887 (N_13887,N_9872,N_11673);
nor U13888 (N_13888,N_10301,N_11574);
and U13889 (N_13889,N_9838,N_9291);
xor U13890 (N_13890,N_10571,N_9264);
nand U13891 (N_13891,N_9244,N_11245);
xor U13892 (N_13892,N_10999,N_10966);
nor U13893 (N_13893,N_11904,N_9183);
and U13894 (N_13894,N_9253,N_10748);
nor U13895 (N_13895,N_11941,N_10729);
nand U13896 (N_13896,N_11710,N_11120);
and U13897 (N_13897,N_10984,N_10341);
xor U13898 (N_13898,N_11503,N_10530);
nor U13899 (N_13899,N_9008,N_10650);
and U13900 (N_13900,N_9465,N_11494);
xnor U13901 (N_13901,N_9469,N_11445);
nand U13902 (N_13902,N_10096,N_10278);
and U13903 (N_13903,N_9420,N_9038);
nor U13904 (N_13904,N_11035,N_11360);
nand U13905 (N_13905,N_9197,N_10007);
nand U13906 (N_13906,N_10813,N_10693);
and U13907 (N_13907,N_10720,N_11924);
nor U13908 (N_13908,N_10668,N_10498);
xor U13909 (N_13909,N_9564,N_11786);
and U13910 (N_13910,N_11898,N_9502);
xnor U13911 (N_13911,N_11799,N_9842);
and U13912 (N_13912,N_10172,N_11088);
nand U13913 (N_13913,N_11527,N_10317);
nor U13914 (N_13914,N_11830,N_9658);
and U13915 (N_13915,N_11755,N_9862);
nand U13916 (N_13916,N_9782,N_10461);
nand U13917 (N_13917,N_11721,N_9576);
xor U13918 (N_13918,N_9866,N_9511);
and U13919 (N_13919,N_9164,N_10539);
nand U13920 (N_13920,N_10548,N_10060);
nand U13921 (N_13921,N_11366,N_9632);
nand U13922 (N_13922,N_11110,N_10071);
and U13923 (N_13923,N_9190,N_11154);
and U13924 (N_13924,N_10079,N_11494);
and U13925 (N_13925,N_10449,N_10129);
nand U13926 (N_13926,N_10779,N_11091);
and U13927 (N_13927,N_9877,N_9053);
and U13928 (N_13928,N_9126,N_9831);
and U13929 (N_13929,N_11260,N_10224);
or U13930 (N_13930,N_11439,N_10275);
or U13931 (N_13931,N_10870,N_9726);
nand U13932 (N_13932,N_11413,N_11415);
xor U13933 (N_13933,N_10033,N_10703);
nand U13934 (N_13934,N_9470,N_10379);
or U13935 (N_13935,N_10622,N_10423);
and U13936 (N_13936,N_9118,N_9615);
nor U13937 (N_13937,N_10938,N_11307);
xnor U13938 (N_13938,N_11175,N_11502);
and U13939 (N_13939,N_9438,N_9444);
or U13940 (N_13940,N_11526,N_11067);
nand U13941 (N_13941,N_9850,N_9654);
xnor U13942 (N_13942,N_10582,N_9774);
xor U13943 (N_13943,N_10371,N_11578);
nor U13944 (N_13944,N_11923,N_9470);
xor U13945 (N_13945,N_11907,N_9657);
or U13946 (N_13946,N_9698,N_11755);
nor U13947 (N_13947,N_9772,N_9581);
nor U13948 (N_13948,N_9722,N_11768);
nor U13949 (N_13949,N_11633,N_9461);
nor U13950 (N_13950,N_10416,N_11260);
xor U13951 (N_13951,N_9003,N_10470);
nor U13952 (N_13952,N_9328,N_11456);
xnor U13953 (N_13953,N_11083,N_9416);
xor U13954 (N_13954,N_10403,N_10349);
xor U13955 (N_13955,N_10227,N_11901);
nand U13956 (N_13956,N_10454,N_11931);
nand U13957 (N_13957,N_10527,N_11273);
xnor U13958 (N_13958,N_9525,N_11029);
or U13959 (N_13959,N_10793,N_9283);
nor U13960 (N_13960,N_11310,N_9185);
nand U13961 (N_13961,N_10525,N_10301);
xnor U13962 (N_13962,N_10727,N_10739);
xor U13963 (N_13963,N_11513,N_11906);
nor U13964 (N_13964,N_9338,N_9368);
and U13965 (N_13965,N_11058,N_9432);
xor U13966 (N_13966,N_11348,N_11813);
xor U13967 (N_13967,N_10203,N_11849);
nand U13968 (N_13968,N_10471,N_10661);
or U13969 (N_13969,N_11730,N_9413);
and U13970 (N_13970,N_9231,N_11394);
or U13971 (N_13971,N_11216,N_10772);
nor U13972 (N_13972,N_9868,N_11698);
nand U13973 (N_13973,N_11271,N_9288);
or U13974 (N_13974,N_10219,N_9668);
or U13975 (N_13975,N_11182,N_10893);
or U13976 (N_13976,N_10784,N_9852);
and U13977 (N_13977,N_9161,N_11611);
or U13978 (N_13978,N_9731,N_10824);
and U13979 (N_13979,N_10687,N_11034);
nand U13980 (N_13980,N_10435,N_10187);
and U13981 (N_13981,N_9906,N_11169);
nor U13982 (N_13982,N_11980,N_11326);
and U13983 (N_13983,N_9089,N_11349);
or U13984 (N_13984,N_9637,N_11039);
nand U13985 (N_13985,N_11114,N_9329);
and U13986 (N_13986,N_10238,N_11962);
and U13987 (N_13987,N_10652,N_11409);
nand U13988 (N_13988,N_9027,N_9183);
or U13989 (N_13989,N_11322,N_11948);
nor U13990 (N_13990,N_10622,N_10595);
or U13991 (N_13991,N_10247,N_11506);
nor U13992 (N_13992,N_10380,N_10635);
and U13993 (N_13993,N_11789,N_11822);
and U13994 (N_13994,N_11749,N_9631);
or U13995 (N_13995,N_9938,N_11819);
xor U13996 (N_13996,N_11063,N_9526);
xnor U13997 (N_13997,N_10493,N_9304);
and U13998 (N_13998,N_11669,N_11434);
xor U13999 (N_13999,N_11177,N_11814);
nor U14000 (N_14000,N_10542,N_11283);
nand U14001 (N_14001,N_11291,N_11261);
nand U14002 (N_14002,N_11168,N_11342);
or U14003 (N_14003,N_11641,N_11999);
nand U14004 (N_14004,N_11515,N_11022);
nand U14005 (N_14005,N_10018,N_11012);
nor U14006 (N_14006,N_11522,N_11491);
or U14007 (N_14007,N_10664,N_9934);
and U14008 (N_14008,N_10125,N_9334);
xnor U14009 (N_14009,N_9442,N_10923);
nor U14010 (N_14010,N_9415,N_11894);
nand U14011 (N_14011,N_10135,N_10862);
nand U14012 (N_14012,N_10250,N_11694);
nor U14013 (N_14013,N_10866,N_10505);
nand U14014 (N_14014,N_9922,N_9568);
or U14015 (N_14015,N_10339,N_10927);
or U14016 (N_14016,N_9989,N_10902);
and U14017 (N_14017,N_9201,N_10989);
nor U14018 (N_14018,N_11345,N_11221);
xor U14019 (N_14019,N_11775,N_10437);
or U14020 (N_14020,N_11836,N_11710);
or U14021 (N_14021,N_10844,N_10880);
nand U14022 (N_14022,N_10774,N_11509);
or U14023 (N_14023,N_11570,N_9895);
nor U14024 (N_14024,N_10851,N_9278);
or U14025 (N_14025,N_11603,N_11831);
xnor U14026 (N_14026,N_10889,N_10550);
xor U14027 (N_14027,N_9927,N_11443);
nand U14028 (N_14028,N_9828,N_11458);
or U14029 (N_14029,N_11213,N_9449);
xnor U14030 (N_14030,N_10164,N_10277);
xor U14031 (N_14031,N_10047,N_9898);
or U14032 (N_14032,N_9194,N_11108);
nand U14033 (N_14033,N_11565,N_9777);
xor U14034 (N_14034,N_9280,N_10749);
xor U14035 (N_14035,N_9041,N_10908);
and U14036 (N_14036,N_10502,N_11895);
xor U14037 (N_14037,N_9307,N_9823);
xor U14038 (N_14038,N_10910,N_11406);
xor U14039 (N_14039,N_10652,N_11343);
and U14040 (N_14040,N_11145,N_10970);
nor U14041 (N_14041,N_10009,N_11271);
nor U14042 (N_14042,N_10366,N_9987);
or U14043 (N_14043,N_10297,N_11404);
nand U14044 (N_14044,N_11351,N_11058);
nor U14045 (N_14045,N_11259,N_11814);
and U14046 (N_14046,N_11302,N_9673);
and U14047 (N_14047,N_11925,N_10038);
nor U14048 (N_14048,N_10963,N_11153);
xor U14049 (N_14049,N_9796,N_9527);
nor U14050 (N_14050,N_11496,N_9344);
nand U14051 (N_14051,N_11359,N_9745);
and U14052 (N_14052,N_10283,N_11595);
xnor U14053 (N_14053,N_10496,N_10185);
xor U14054 (N_14054,N_10678,N_9912);
nand U14055 (N_14055,N_9338,N_9522);
nor U14056 (N_14056,N_10232,N_10967);
nand U14057 (N_14057,N_9058,N_11708);
or U14058 (N_14058,N_10836,N_11169);
or U14059 (N_14059,N_11926,N_9791);
nor U14060 (N_14060,N_11637,N_10749);
or U14061 (N_14061,N_9176,N_11566);
and U14062 (N_14062,N_9549,N_10489);
nand U14063 (N_14063,N_9847,N_11279);
xnor U14064 (N_14064,N_10597,N_9583);
nor U14065 (N_14065,N_10022,N_9326);
nand U14066 (N_14066,N_11702,N_9000);
nor U14067 (N_14067,N_9994,N_9416);
xnor U14068 (N_14068,N_9952,N_9597);
or U14069 (N_14069,N_10266,N_9950);
xnor U14070 (N_14070,N_11306,N_10188);
or U14071 (N_14071,N_10160,N_10166);
and U14072 (N_14072,N_9203,N_9348);
nor U14073 (N_14073,N_11334,N_11410);
and U14074 (N_14074,N_11340,N_9754);
or U14075 (N_14075,N_11505,N_9359);
nor U14076 (N_14076,N_9287,N_11292);
or U14077 (N_14077,N_11972,N_9438);
and U14078 (N_14078,N_10704,N_11236);
xnor U14079 (N_14079,N_9015,N_11653);
nand U14080 (N_14080,N_10037,N_11040);
nand U14081 (N_14081,N_11968,N_10769);
and U14082 (N_14082,N_10510,N_10362);
nand U14083 (N_14083,N_9126,N_9587);
xor U14084 (N_14084,N_10801,N_11688);
and U14085 (N_14085,N_11278,N_9533);
or U14086 (N_14086,N_9643,N_10787);
and U14087 (N_14087,N_11119,N_11208);
and U14088 (N_14088,N_9329,N_10085);
xor U14089 (N_14089,N_9212,N_11677);
nor U14090 (N_14090,N_9965,N_9621);
or U14091 (N_14091,N_9007,N_10641);
and U14092 (N_14092,N_11000,N_9218);
xnor U14093 (N_14093,N_10369,N_9573);
nor U14094 (N_14094,N_11850,N_10995);
or U14095 (N_14095,N_9371,N_9428);
xnor U14096 (N_14096,N_11925,N_11639);
xor U14097 (N_14097,N_10591,N_10647);
nor U14098 (N_14098,N_9566,N_11851);
nand U14099 (N_14099,N_10473,N_9803);
xor U14100 (N_14100,N_10495,N_10660);
nor U14101 (N_14101,N_9155,N_9978);
nand U14102 (N_14102,N_11264,N_9669);
xnor U14103 (N_14103,N_10993,N_9074);
and U14104 (N_14104,N_9703,N_11140);
nor U14105 (N_14105,N_10380,N_9970);
nand U14106 (N_14106,N_11667,N_10601);
xor U14107 (N_14107,N_9784,N_9008);
xnor U14108 (N_14108,N_11587,N_9658);
xor U14109 (N_14109,N_9892,N_9999);
or U14110 (N_14110,N_9754,N_11629);
or U14111 (N_14111,N_11029,N_10592);
or U14112 (N_14112,N_9664,N_10777);
nor U14113 (N_14113,N_11180,N_10886);
nand U14114 (N_14114,N_9316,N_11580);
nor U14115 (N_14115,N_11228,N_10484);
xnor U14116 (N_14116,N_10971,N_9163);
nand U14117 (N_14117,N_9923,N_9656);
nor U14118 (N_14118,N_10534,N_9132);
or U14119 (N_14119,N_10482,N_9645);
and U14120 (N_14120,N_11489,N_10105);
xnor U14121 (N_14121,N_10883,N_10523);
nor U14122 (N_14122,N_11621,N_10656);
nand U14123 (N_14123,N_10833,N_11170);
or U14124 (N_14124,N_11164,N_11696);
or U14125 (N_14125,N_10286,N_9499);
nand U14126 (N_14126,N_10117,N_10395);
or U14127 (N_14127,N_11424,N_11836);
nor U14128 (N_14128,N_9914,N_9313);
or U14129 (N_14129,N_11350,N_11484);
nand U14130 (N_14130,N_11236,N_10699);
xor U14131 (N_14131,N_11535,N_9452);
nor U14132 (N_14132,N_9347,N_11264);
and U14133 (N_14133,N_11444,N_10852);
and U14134 (N_14134,N_11065,N_9317);
nor U14135 (N_14135,N_10177,N_11769);
xor U14136 (N_14136,N_11005,N_9223);
nor U14137 (N_14137,N_11708,N_11170);
xnor U14138 (N_14138,N_10639,N_11505);
nand U14139 (N_14139,N_11226,N_9121);
nor U14140 (N_14140,N_9058,N_10947);
nand U14141 (N_14141,N_11157,N_10962);
and U14142 (N_14142,N_10704,N_10856);
nand U14143 (N_14143,N_9423,N_11511);
xor U14144 (N_14144,N_10445,N_11923);
nand U14145 (N_14145,N_9095,N_9047);
nor U14146 (N_14146,N_11714,N_11691);
and U14147 (N_14147,N_9660,N_9347);
or U14148 (N_14148,N_11974,N_10242);
or U14149 (N_14149,N_11154,N_9735);
nor U14150 (N_14150,N_9832,N_11530);
nor U14151 (N_14151,N_9158,N_11656);
xnor U14152 (N_14152,N_11230,N_11870);
xor U14153 (N_14153,N_9002,N_9234);
nor U14154 (N_14154,N_10023,N_10101);
nand U14155 (N_14155,N_11830,N_9595);
and U14156 (N_14156,N_11675,N_10921);
and U14157 (N_14157,N_10538,N_11605);
nand U14158 (N_14158,N_9359,N_11700);
nor U14159 (N_14159,N_10807,N_10866);
nand U14160 (N_14160,N_9478,N_10794);
xnor U14161 (N_14161,N_11017,N_10328);
nor U14162 (N_14162,N_9001,N_9004);
or U14163 (N_14163,N_10211,N_9010);
nand U14164 (N_14164,N_11860,N_10253);
and U14165 (N_14165,N_9955,N_9103);
xor U14166 (N_14166,N_10892,N_9471);
or U14167 (N_14167,N_9761,N_10084);
xor U14168 (N_14168,N_10110,N_11536);
nor U14169 (N_14169,N_11791,N_10850);
xor U14170 (N_14170,N_9923,N_9569);
or U14171 (N_14171,N_11647,N_10687);
nand U14172 (N_14172,N_10285,N_10282);
nand U14173 (N_14173,N_9510,N_9384);
nor U14174 (N_14174,N_11272,N_10482);
or U14175 (N_14175,N_11155,N_9703);
and U14176 (N_14176,N_10108,N_9577);
nand U14177 (N_14177,N_9722,N_10985);
xor U14178 (N_14178,N_11928,N_11229);
nor U14179 (N_14179,N_9968,N_9703);
or U14180 (N_14180,N_9229,N_10289);
or U14181 (N_14181,N_10746,N_11542);
nand U14182 (N_14182,N_9786,N_10229);
nand U14183 (N_14183,N_10723,N_9618);
nand U14184 (N_14184,N_9689,N_11771);
nor U14185 (N_14185,N_9860,N_9722);
or U14186 (N_14186,N_11189,N_10227);
xor U14187 (N_14187,N_10517,N_11290);
or U14188 (N_14188,N_11243,N_10055);
nand U14189 (N_14189,N_9585,N_11321);
nor U14190 (N_14190,N_9799,N_9243);
nor U14191 (N_14191,N_10877,N_11940);
nand U14192 (N_14192,N_11112,N_11272);
and U14193 (N_14193,N_11342,N_11862);
and U14194 (N_14194,N_11021,N_11925);
or U14195 (N_14195,N_9338,N_11860);
and U14196 (N_14196,N_11870,N_10532);
nor U14197 (N_14197,N_9980,N_10585);
nand U14198 (N_14198,N_9248,N_10593);
nor U14199 (N_14199,N_11153,N_10522);
nand U14200 (N_14200,N_11605,N_10964);
or U14201 (N_14201,N_9902,N_11133);
and U14202 (N_14202,N_9878,N_11228);
and U14203 (N_14203,N_11675,N_11486);
nand U14204 (N_14204,N_10615,N_9853);
and U14205 (N_14205,N_11077,N_10046);
xnor U14206 (N_14206,N_11856,N_9879);
and U14207 (N_14207,N_9674,N_10198);
xnor U14208 (N_14208,N_9089,N_11970);
xor U14209 (N_14209,N_10770,N_10455);
and U14210 (N_14210,N_10847,N_10112);
xnor U14211 (N_14211,N_11337,N_11931);
nor U14212 (N_14212,N_10261,N_9278);
xor U14213 (N_14213,N_11544,N_10307);
and U14214 (N_14214,N_11905,N_10446);
and U14215 (N_14215,N_9592,N_10298);
or U14216 (N_14216,N_11034,N_11944);
nand U14217 (N_14217,N_10979,N_11937);
and U14218 (N_14218,N_9482,N_11893);
nand U14219 (N_14219,N_11816,N_9871);
or U14220 (N_14220,N_9593,N_9432);
or U14221 (N_14221,N_11333,N_10497);
or U14222 (N_14222,N_10825,N_9424);
xor U14223 (N_14223,N_9917,N_11521);
and U14224 (N_14224,N_9794,N_9638);
nor U14225 (N_14225,N_9990,N_9936);
nor U14226 (N_14226,N_9802,N_11417);
nand U14227 (N_14227,N_10921,N_10465);
nor U14228 (N_14228,N_10488,N_9955);
nor U14229 (N_14229,N_10095,N_10442);
nor U14230 (N_14230,N_11299,N_11162);
nor U14231 (N_14231,N_9900,N_11953);
xnor U14232 (N_14232,N_10281,N_10361);
or U14233 (N_14233,N_11414,N_11804);
nand U14234 (N_14234,N_9875,N_9682);
nand U14235 (N_14235,N_10587,N_9524);
and U14236 (N_14236,N_11087,N_11493);
xor U14237 (N_14237,N_10487,N_10459);
nand U14238 (N_14238,N_11984,N_9396);
and U14239 (N_14239,N_10145,N_10276);
or U14240 (N_14240,N_10186,N_10124);
xor U14241 (N_14241,N_10535,N_11482);
nor U14242 (N_14242,N_9723,N_11529);
xnor U14243 (N_14243,N_9374,N_11511);
or U14244 (N_14244,N_10082,N_11468);
or U14245 (N_14245,N_10605,N_9403);
or U14246 (N_14246,N_9237,N_10363);
nand U14247 (N_14247,N_9080,N_11433);
nand U14248 (N_14248,N_10364,N_10092);
nand U14249 (N_14249,N_11542,N_9399);
or U14250 (N_14250,N_11087,N_9802);
nand U14251 (N_14251,N_9380,N_11644);
or U14252 (N_14252,N_10529,N_9504);
nor U14253 (N_14253,N_9296,N_10136);
nand U14254 (N_14254,N_10269,N_10611);
nor U14255 (N_14255,N_11021,N_10276);
nand U14256 (N_14256,N_9680,N_11506);
or U14257 (N_14257,N_11070,N_9158);
nor U14258 (N_14258,N_9626,N_9658);
xor U14259 (N_14259,N_10446,N_9420);
nand U14260 (N_14260,N_9687,N_11328);
and U14261 (N_14261,N_10350,N_10308);
nor U14262 (N_14262,N_9757,N_9057);
nand U14263 (N_14263,N_11021,N_9872);
nor U14264 (N_14264,N_10056,N_9778);
xor U14265 (N_14265,N_10073,N_11377);
xnor U14266 (N_14266,N_10596,N_9583);
nor U14267 (N_14267,N_11776,N_10030);
nor U14268 (N_14268,N_9885,N_11769);
nand U14269 (N_14269,N_10598,N_11553);
xor U14270 (N_14270,N_11044,N_9257);
nor U14271 (N_14271,N_10379,N_9996);
xnor U14272 (N_14272,N_9517,N_10950);
nand U14273 (N_14273,N_9941,N_9566);
nor U14274 (N_14274,N_10306,N_10429);
nor U14275 (N_14275,N_10144,N_9905);
nor U14276 (N_14276,N_11814,N_10359);
and U14277 (N_14277,N_10558,N_9559);
xor U14278 (N_14278,N_11506,N_11421);
or U14279 (N_14279,N_9810,N_11159);
nor U14280 (N_14280,N_10894,N_10803);
and U14281 (N_14281,N_9617,N_9241);
xnor U14282 (N_14282,N_11573,N_9913);
or U14283 (N_14283,N_10204,N_10405);
xor U14284 (N_14284,N_11250,N_9755);
xnor U14285 (N_14285,N_11531,N_9781);
nand U14286 (N_14286,N_10545,N_10701);
or U14287 (N_14287,N_9244,N_9089);
or U14288 (N_14288,N_9739,N_11424);
nand U14289 (N_14289,N_11126,N_10007);
or U14290 (N_14290,N_10127,N_9519);
nand U14291 (N_14291,N_10531,N_10984);
or U14292 (N_14292,N_11048,N_11514);
xnor U14293 (N_14293,N_10638,N_9791);
nor U14294 (N_14294,N_11092,N_10810);
and U14295 (N_14295,N_11533,N_11835);
xnor U14296 (N_14296,N_11020,N_10596);
xnor U14297 (N_14297,N_9858,N_10453);
nor U14298 (N_14298,N_10574,N_9586);
and U14299 (N_14299,N_11576,N_9971);
xor U14300 (N_14300,N_10055,N_11234);
and U14301 (N_14301,N_9793,N_9001);
xnor U14302 (N_14302,N_11528,N_9427);
nor U14303 (N_14303,N_11193,N_9478);
nand U14304 (N_14304,N_11060,N_9162);
and U14305 (N_14305,N_10759,N_9089);
nor U14306 (N_14306,N_10787,N_9960);
nand U14307 (N_14307,N_11877,N_10086);
or U14308 (N_14308,N_9385,N_10972);
or U14309 (N_14309,N_10543,N_10038);
or U14310 (N_14310,N_9956,N_9699);
and U14311 (N_14311,N_11471,N_11232);
or U14312 (N_14312,N_9285,N_10560);
and U14313 (N_14313,N_9095,N_11106);
xnor U14314 (N_14314,N_9806,N_9271);
xor U14315 (N_14315,N_11293,N_11013);
or U14316 (N_14316,N_11365,N_9560);
nand U14317 (N_14317,N_9249,N_10501);
xor U14318 (N_14318,N_11042,N_10580);
or U14319 (N_14319,N_10963,N_10678);
xnor U14320 (N_14320,N_10264,N_9820);
or U14321 (N_14321,N_10457,N_11132);
xor U14322 (N_14322,N_9879,N_9866);
nand U14323 (N_14323,N_10446,N_9040);
nor U14324 (N_14324,N_9470,N_11919);
and U14325 (N_14325,N_10578,N_11272);
nand U14326 (N_14326,N_10309,N_9918);
and U14327 (N_14327,N_11213,N_10123);
and U14328 (N_14328,N_10375,N_9890);
xnor U14329 (N_14329,N_11121,N_11734);
and U14330 (N_14330,N_11025,N_10192);
nand U14331 (N_14331,N_10805,N_11022);
nor U14332 (N_14332,N_10641,N_9841);
and U14333 (N_14333,N_11323,N_11465);
nand U14334 (N_14334,N_10176,N_9390);
and U14335 (N_14335,N_11420,N_10035);
or U14336 (N_14336,N_10420,N_11102);
or U14337 (N_14337,N_10705,N_9673);
nor U14338 (N_14338,N_10257,N_10624);
or U14339 (N_14339,N_9736,N_11933);
or U14340 (N_14340,N_11882,N_9288);
or U14341 (N_14341,N_10268,N_10534);
or U14342 (N_14342,N_9898,N_9384);
nor U14343 (N_14343,N_10355,N_10952);
nand U14344 (N_14344,N_9815,N_9192);
xnor U14345 (N_14345,N_10044,N_10999);
or U14346 (N_14346,N_9200,N_10623);
nor U14347 (N_14347,N_9918,N_10400);
or U14348 (N_14348,N_10597,N_11550);
xor U14349 (N_14349,N_9932,N_9002);
nand U14350 (N_14350,N_11564,N_9982);
and U14351 (N_14351,N_10559,N_10696);
nor U14352 (N_14352,N_11722,N_9957);
nor U14353 (N_14353,N_9462,N_9387);
xor U14354 (N_14354,N_9744,N_11580);
nand U14355 (N_14355,N_10981,N_9415);
or U14356 (N_14356,N_11256,N_9591);
nand U14357 (N_14357,N_11147,N_11732);
nand U14358 (N_14358,N_9197,N_9640);
xnor U14359 (N_14359,N_10844,N_10409);
and U14360 (N_14360,N_10277,N_11393);
nand U14361 (N_14361,N_11892,N_10909);
and U14362 (N_14362,N_11520,N_11906);
or U14363 (N_14363,N_9285,N_11737);
nor U14364 (N_14364,N_10781,N_11116);
xor U14365 (N_14365,N_10053,N_11238);
nand U14366 (N_14366,N_11401,N_10867);
or U14367 (N_14367,N_9103,N_11977);
nor U14368 (N_14368,N_11973,N_11676);
nor U14369 (N_14369,N_9589,N_9400);
and U14370 (N_14370,N_9072,N_10428);
nor U14371 (N_14371,N_10426,N_11885);
xnor U14372 (N_14372,N_10806,N_11638);
xor U14373 (N_14373,N_10717,N_9097);
or U14374 (N_14374,N_10974,N_9574);
or U14375 (N_14375,N_9634,N_9190);
or U14376 (N_14376,N_11661,N_11226);
nor U14377 (N_14377,N_11191,N_10471);
nand U14378 (N_14378,N_10036,N_11303);
xnor U14379 (N_14379,N_10626,N_11535);
nand U14380 (N_14380,N_9786,N_11861);
nand U14381 (N_14381,N_9709,N_9318);
or U14382 (N_14382,N_9770,N_11240);
and U14383 (N_14383,N_9534,N_9076);
and U14384 (N_14384,N_9945,N_9786);
nor U14385 (N_14385,N_11734,N_10526);
or U14386 (N_14386,N_10482,N_10984);
nor U14387 (N_14387,N_10257,N_9127);
nor U14388 (N_14388,N_9219,N_11926);
xnor U14389 (N_14389,N_9445,N_11252);
or U14390 (N_14390,N_9819,N_10274);
xnor U14391 (N_14391,N_11264,N_10991);
nor U14392 (N_14392,N_9104,N_11214);
or U14393 (N_14393,N_9476,N_11152);
xor U14394 (N_14394,N_10367,N_10131);
nor U14395 (N_14395,N_9413,N_10613);
or U14396 (N_14396,N_9281,N_9238);
and U14397 (N_14397,N_10238,N_11402);
xor U14398 (N_14398,N_9316,N_10255);
and U14399 (N_14399,N_11602,N_11648);
nand U14400 (N_14400,N_10495,N_10579);
nor U14401 (N_14401,N_11591,N_10654);
and U14402 (N_14402,N_11912,N_11199);
and U14403 (N_14403,N_11663,N_9335);
xor U14404 (N_14404,N_10394,N_10900);
xor U14405 (N_14405,N_11269,N_9365);
and U14406 (N_14406,N_9725,N_11110);
xnor U14407 (N_14407,N_10244,N_11910);
nor U14408 (N_14408,N_10081,N_9858);
or U14409 (N_14409,N_9779,N_11926);
nor U14410 (N_14410,N_10976,N_9128);
xnor U14411 (N_14411,N_10148,N_11189);
xnor U14412 (N_14412,N_10080,N_9621);
nand U14413 (N_14413,N_10579,N_9323);
nor U14414 (N_14414,N_11048,N_10066);
xor U14415 (N_14415,N_11351,N_10351);
or U14416 (N_14416,N_10626,N_11152);
nand U14417 (N_14417,N_10992,N_11674);
nand U14418 (N_14418,N_9496,N_9246);
and U14419 (N_14419,N_10286,N_11345);
xnor U14420 (N_14420,N_9363,N_10100);
xnor U14421 (N_14421,N_11659,N_9931);
nor U14422 (N_14422,N_10516,N_11448);
and U14423 (N_14423,N_9141,N_9407);
nand U14424 (N_14424,N_9040,N_10846);
xnor U14425 (N_14425,N_9459,N_9052);
or U14426 (N_14426,N_11370,N_11363);
xor U14427 (N_14427,N_11855,N_10782);
or U14428 (N_14428,N_9127,N_10373);
xnor U14429 (N_14429,N_11548,N_10794);
xor U14430 (N_14430,N_10265,N_9347);
nor U14431 (N_14431,N_9751,N_11716);
or U14432 (N_14432,N_9908,N_10423);
nand U14433 (N_14433,N_10181,N_10430);
or U14434 (N_14434,N_10985,N_9425);
and U14435 (N_14435,N_9416,N_9494);
or U14436 (N_14436,N_11175,N_11947);
and U14437 (N_14437,N_10210,N_9152);
or U14438 (N_14438,N_10010,N_9263);
and U14439 (N_14439,N_10886,N_11365);
and U14440 (N_14440,N_11471,N_10569);
or U14441 (N_14441,N_10030,N_10703);
and U14442 (N_14442,N_11332,N_9401);
or U14443 (N_14443,N_9340,N_9213);
nor U14444 (N_14444,N_10167,N_9115);
nor U14445 (N_14445,N_11949,N_11110);
nor U14446 (N_14446,N_9956,N_11892);
xnor U14447 (N_14447,N_11770,N_9216);
nand U14448 (N_14448,N_11152,N_10391);
nand U14449 (N_14449,N_10705,N_9010);
and U14450 (N_14450,N_10105,N_11776);
xor U14451 (N_14451,N_9655,N_10133);
nor U14452 (N_14452,N_10898,N_11172);
or U14453 (N_14453,N_9082,N_11652);
nand U14454 (N_14454,N_9958,N_9818);
and U14455 (N_14455,N_9801,N_11682);
nor U14456 (N_14456,N_9011,N_9541);
and U14457 (N_14457,N_9782,N_11968);
and U14458 (N_14458,N_9584,N_9988);
nor U14459 (N_14459,N_11593,N_9169);
or U14460 (N_14460,N_11852,N_10483);
and U14461 (N_14461,N_10674,N_11093);
and U14462 (N_14462,N_10419,N_9277);
nand U14463 (N_14463,N_10207,N_10463);
or U14464 (N_14464,N_10801,N_11267);
and U14465 (N_14465,N_11568,N_9251);
xor U14466 (N_14466,N_9554,N_9791);
nor U14467 (N_14467,N_11580,N_11890);
or U14468 (N_14468,N_11138,N_11710);
or U14469 (N_14469,N_11522,N_11673);
nor U14470 (N_14470,N_11519,N_9950);
or U14471 (N_14471,N_10501,N_11652);
nor U14472 (N_14472,N_9870,N_11846);
nand U14473 (N_14473,N_9712,N_9587);
or U14474 (N_14474,N_10718,N_11594);
nand U14475 (N_14475,N_9797,N_9269);
xor U14476 (N_14476,N_9820,N_10769);
nor U14477 (N_14477,N_9892,N_11802);
nor U14478 (N_14478,N_11073,N_10651);
or U14479 (N_14479,N_11061,N_11219);
nor U14480 (N_14480,N_11048,N_9486);
and U14481 (N_14481,N_10786,N_10535);
or U14482 (N_14482,N_11120,N_11826);
nand U14483 (N_14483,N_9967,N_11042);
and U14484 (N_14484,N_10699,N_9844);
and U14485 (N_14485,N_11670,N_11691);
and U14486 (N_14486,N_10765,N_10145);
and U14487 (N_14487,N_11551,N_9095);
nor U14488 (N_14488,N_11250,N_11344);
nand U14489 (N_14489,N_10209,N_10995);
nand U14490 (N_14490,N_11737,N_10147);
xnor U14491 (N_14491,N_11407,N_9347);
or U14492 (N_14492,N_11299,N_11119);
xor U14493 (N_14493,N_10474,N_10441);
and U14494 (N_14494,N_9035,N_10324);
nand U14495 (N_14495,N_10874,N_11484);
or U14496 (N_14496,N_11509,N_9902);
nand U14497 (N_14497,N_11134,N_11688);
and U14498 (N_14498,N_10890,N_10859);
xor U14499 (N_14499,N_11326,N_10202);
nor U14500 (N_14500,N_10578,N_11047);
or U14501 (N_14501,N_9112,N_10886);
xnor U14502 (N_14502,N_9596,N_11232);
and U14503 (N_14503,N_9846,N_10248);
xnor U14504 (N_14504,N_10395,N_9556);
xnor U14505 (N_14505,N_9320,N_9257);
nand U14506 (N_14506,N_10697,N_11759);
or U14507 (N_14507,N_11223,N_9726);
nor U14508 (N_14508,N_11822,N_9811);
xnor U14509 (N_14509,N_11374,N_11725);
nor U14510 (N_14510,N_9360,N_10669);
and U14511 (N_14511,N_10598,N_10575);
xnor U14512 (N_14512,N_11125,N_9750);
nor U14513 (N_14513,N_10190,N_11064);
nand U14514 (N_14514,N_9610,N_9714);
nand U14515 (N_14515,N_11141,N_10077);
nor U14516 (N_14516,N_10915,N_9416);
or U14517 (N_14517,N_9661,N_11856);
nand U14518 (N_14518,N_9512,N_11990);
or U14519 (N_14519,N_11483,N_10712);
and U14520 (N_14520,N_11947,N_9760);
nand U14521 (N_14521,N_11266,N_9240);
or U14522 (N_14522,N_10063,N_9120);
or U14523 (N_14523,N_9045,N_10853);
nor U14524 (N_14524,N_11107,N_9019);
nand U14525 (N_14525,N_11593,N_11103);
or U14526 (N_14526,N_11250,N_11908);
and U14527 (N_14527,N_9513,N_10083);
nor U14528 (N_14528,N_11206,N_10211);
nor U14529 (N_14529,N_11251,N_10746);
and U14530 (N_14530,N_9571,N_9972);
and U14531 (N_14531,N_10592,N_10217);
nand U14532 (N_14532,N_11969,N_10841);
or U14533 (N_14533,N_10447,N_11821);
or U14534 (N_14534,N_10367,N_11944);
nand U14535 (N_14535,N_11879,N_11396);
or U14536 (N_14536,N_9067,N_10990);
nand U14537 (N_14537,N_11783,N_11613);
and U14538 (N_14538,N_10349,N_10404);
or U14539 (N_14539,N_9889,N_11036);
nor U14540 (N_14540,N_10801,N_10382);
and U14541 (N_14541,N_9008,N_10641);
nor U14542 (N_14542,N_11149,N_10889);
nor U14543 (N_14543,N_10770,N_11025);
xor U14544 (N_14544,N_10550,N_9609);
nand U14545 (N_14545,N_10790,N_10308);
nor U14546 (N_14546,N_11640,N_11013);
nand U14547 (N_14547,N_9182,N_11965);
nand U14548 (N_14548,N_11054,N_10418);
and U14549 (N_14549,N_11281,N_9863);
nand U14550 (N_14550,N_10392,N_9073);
nand U14551 (N_14551,N_11285,N_9850);
xor U14552 (N_14552,N_11331,N_9115);
or U14553 (N_14553,N_9468,N_9362);
nor U14554 (N_14554,N_11615,N_11401);
or U14555 (N_14555,N_10879,N_9287);
xor U14556 (N_14556,N_11345,N_10593);
nor U14557 (N_14557,N_10882,N_9909);
or U14558 (N_14558,N_9086,N_9143);
xnor U14559 (N_14559,N_10251,N_9929);
nor U14560 (N_14560,N_9620,N_9661);
nor U14561 (N_14561,N_10399,N_11936);
nand U14562 (N_14562,N_10542,N_11208);
nand U14563 (N_14563,N_10937,N_10557);
nand U14564 (N_14564,N_10653,N_11159);
nor U14565 (N_14565,N_9346,N_9088);
nor U14566 (N_14566,N_11972,N_9184);
or U14567 (N_14567,N_10236,N_9624);
nor U14568 (N_14568,N_10784,N_9987);
and U14569 (N_14569,N_10381,N_11586);
xnor U14570 (N_14570,N_9625,N_11168);
and U14571 (N_14571,N_10447,N_9348);
and U14572 (N_14572,N_10626,N_9737);
nand U14573 (N_14573,N_9538,N_9000);
nor U14574 (N_14574,N_10643,N_9534);
nand U14575 (N_14575,N_9187,N_11449);
and U14576 (N_14576,N_9961,N_11039);
xnor U14577 (N_14577,N_11330,N_10801);
and U14578 (N_14578,N_9595,N_10146);
and U14579 (N_14579,N_10835,N_9062);
nor U14580 (N_14580,N_9239,N_10374);
nor U14581 (N_14581,N_10804,N_10673);
xnor U14582 (N_14582,N_9185,N_11726);
and U14583 (N_14583,N_10698,N_10300);
or U14584 (N_14584,N_9801,N_11684);
xor U14585 (N_14585,N_11499,N_11473);
and U14586 (N_14586,N_11123,N_11365);
or U14587 (N_14587,N_9397,N_11436);
nor U14588 (N_14588,N_11554,N_11069);
xnor U14589 (N_14589,N_9037,N_11080);
nor U14590 (N_14590,N_9699,N_10894);
and U14591 (N_14591,N_11265,N_10573);
nand U14592 (N_14592,N_10624,N_9894);
and U14593 (N_14593,N_9715,N_9252);
and U14594 (N_14594,N_11510,N_10334);
and U14595 (N_14595,N_11523,N_9018);
or U14596 (N_14596,N_10537,N_10733);
xnor U14597 (N_14597,N_9450,N_11303);
and U14598 (N_14598,N_10747,N_11367);
and U14599 (N_14599,N_10099,N_10774);
and U14600 (N_14600,N_9052,N_10979);
and U14601 (N_14601,N_11382,N_10514);
nand U14602 (N_14602,N_9904,N_9846);
nand U14603 (N_14603,N_11586,N_11714);
xor U14604 (N_14604,N_11894,N_10057);
and U14605 (N_14605,N_11671,N_11692);
nand U14606 (N_14606,N_11268,N_11724);
nor U14607 (N_14607,N_9930,N_11380);
xnor U14608 (N_14608,N_9367,N_11927);
and U14609 (N_14609,N_9724,N_9712);
and U14610 (N_14610,N_11687,N_11649);
nand U14611 (N_14611,N_9379,N_11657);
nor U14612 (N_14612,N_11320,N_10688);
xor U14613 (N_14613,N_10464,N_11654);
and U14614 (N_14614,N_11450,N_9760);
nor U14615 (N_14615,N_11762,N_11075);
and U14616 (N_14616,N_11265,N_10519);
xor U14617 (N_14617,N_11130,N_10222);
or U14618 (N_14618,N_11282,N_11311);
and U14619 (N_14619,N_11776,N_9763);
and U14620 (N_14620,N_11815,N_11853);
or U14621 (N_14621,N_9703,N_10057);
or U14622 (N_14622,N_10080,N_10307);
xor U14623 (N_14623,N_11761,N_10968);
and U14624 (N_14624,N_11713,N_9630);
or U14625 (N_14625,N_11421,N_9476);
nand U14626 (N_14626,N_11141,N_9045);
nand U14627 (N_14627,N_9604,N_9018);
nand U14628 (N_14628,N_9088,N_11559);
xnor U14629 (N_14629,N_11091,N_9315);
nand U14630 (N_14630,N_9394,N_11422);
nand U14631 (N_14631,N_10047,N_10716);
and U14632 (N_14632,N_11797,N_10029);
nor U14633 (N_14633,N_10012,N_9496);
or U14634 (N_14634,N_10650,N_10784);
nor U14635 (N_14635,N_11348,N_11900);
or U14636 (N_14636,N_9969,N_10915);
xor U14637 (N_14637,N_10905,N_9890);
nor U14638 (N_14638,N_10533,N_10263);
nor U14639 (N_14639,N_10227,N_10771);
nand U14640 (N_14640,N_10002,N_9296);
nor U14641 (N_14641,N_11694,N_11825);
xor U14642 (N_14642,N_9485,N_11237);
and U14643 (N_14643,N_11889,N_9833);
xnor U14644 (N_14644,N_9749,N_11801);
xnor U14645 (N_14645,N_10868,N_9439);
and U14646 (N_14646,N_11046,N_11926);
xnor U14647 (N_14647,N_9440,N_11305);
nand U14648 (N_14648,N_10281,N_10079);
xnor U14649 (N_14649,N_11388,N_10314);
nor U14650 (N_14650,N_11630,N_9791);
or U14651 (N_14651,N_10907,N_10335);
and U14652 (N_14652,N_10193,N_10571);
and U14653 (N_14653,N_10918,N_9721);
or U14654 (N_14654,N_11032,N_9732);
and U14655 (N_14655,N_11281,N_9938);
or U14656 (N_14656,N_11598,N_10425);
xnor U14657 (N_14657,N_10437,N_10650);
xnor U14658 (N_14658,N_9089,N_11156);
and U14659 (N_14659,N_10566,N_9614);
xor U14660 (N_14660,N_9385,N_9259);
nand U14661 (N_14661,N_11932,N_10692);
xnor U14662 (N_14662,N_9200,N_9451);
nand U14663 (N_14663,N_11119,N_9272);
nor U14664 (N_14664,N_10878,N_10889);
xnor U14665 (N_14665,N_9845,N_10858);
and U14666 (N_14666,N_11038,N_10788);
and U14667 (N_14667,N_10279,N_10934);
nor U14668 (N_14668,N_11952,N_11651);
or U14669 (N_14669,N_9797,N_10347);
xor U14670 (N_14670,N_9115,N_9670);
nor U14671 (N_14671,N_11403,N_10734);
or U14672 (N_14672,N_10544,N_10157);
nand U14673 (N_14673,N_11551,N_10667);
or U14674 (N_14674,N_11131,N_9782);
nand U14675 (N_14675,N_11413,N_9234);
nor U14676 (N_14676,N_9733,N_11718);
or U14677 (N_14677,N_11124,N_11311);
xnor U14678 (N_14678,N_9114,N_9233);
xnor U14679 (N_14679,N_11473,N_9832);
or U14680 (N_14680,N_11511,N_10400);
or U14681 (N_14681,N_11626,N_9566);
nand U14682 (N_14682,N_9387,N_11864);
or U14683 (N_14683,N_11948,N_10646);
or U14684 (N_14684,N_11047,N_9840);
or U14685 (N_14685,N_11578,N_9585);
nand U14686 (N_14686,N_10420,N_10381);
nand U14687 (N_14687,N_9680,N_9579);
and U14688 (N_14688,N_9209,N_10681);
or U14689 (N_14689,N_10526,N_11525);
nand U14690 (N_14690,N_11372,N_11121);
or U14691 (N_14691,N_10698,N_11248);
or U14692 (N_14692,N_11369,N_10725);
xnor U14693 (N_14693,N_9232,N_11438);
and U14694 (N_14694,N_11912,N_9449);
and U14695 (N_14695,N_11042,N_10309);
nor U14696 (N_14696,N_11781,N_10443);
nor U14697 (N_14697,N_11550,N_9520);
and U14698 (N_14698,N_9107,N_11318);
xnor U14699 (N_14699,N_10214,N_10146);
nor U14700 (N_14700,N_10499,N_10321);
and U14701 (N_14701,N_11300,N_11721);
or U14702 (N_14702,N_9934,N_10994);
nor U14703 (N_14703,N_10139,N_10087);
xnor U14704 (N_14704,N_10752,N_10238);
nor U14705 (N_14705,N_9057,N_11414);
nor U14706 (N_14706,N_11172,N_11995);
nor U14707 (N_14707,N_10833,N_10029);
nor U14708 (N_14708,N_9081,N_11297);
or U14709 (N_14709,N_9111,N_11568);
xnor U14710 (N_14710,N_9159,N_11358);
or U14711 (N_14711,N_10825,N_10354);
nor U14712 (N_14712,N_10285,N_11431);
and U14713 (N_14713,N_9232,N_11434);
or U14714 (N_14714,N_10415,N_10461);
or U14715 (N_14715,N_9679,N_11961);
and U14716 (N_14716,N_9008,N_10361);
nand U14717 (N_14717,N_10480,N_9414);
and U14718 (N_14718,N_11358,N_11634);
xnor U14719 (N_14719,N_11696,N_9908);
nand U14720 (N_14720,N_11459,N_9204);
and U14721 (N_14721,N_9173,N_11949);
or U14722 (N_14722,N_10678,N_11843);
xnor U14723 (N_14723,N_10587,N_10905);
nor U14724 (N_14724,N_9398,N_11223);
or U14725 (N_14725,N_11478,N_9161);
or U14726 (N_14726,N_10759,N_11881);
xor U14727 (N_14727,N_9598,N_9879);
and U14728 (N_14728,N_11010,N_11401);
xor U14729 (N_14729,N_11615,N_10538);
and U14730 (N_14730,N_9807,N_11496);
and U14731 (N_14731,N_10288,N_10135);
and U14732 (N_14732,N_9953,N_11533);
nand U14733 (N_14733,N_10354,N_9925);
and U14734 (N_14734,N_10454,N_11260);
xnor U14735 (N_14735,N_10646,N_9881);
xor U14736 (N_14736,N_9914,N_10965);
and U14737 (N_14737,N_9732,N_9150);
nor U14738 (N_14738,N_11036,N_9644);
nand U14739 (N_14739,N_11023,N_9208);
xor U14740 (N_14740,N_11173,N_9191);
nor U14741 (N_14741,N_11985,N_10286);
or U14742 (N_14742,N_10880,N_11341);
xnor U14743 (N_14743,N_9901,N_9435);
or U14744 (N_14744,N_9844,N_11044);
or U14745 (N_14745,N_11654,N_11197);
nor U14746 (N_14746,N_9068,N_9161);
nand U14747 (N_14747,N_10832,N_10274);
nand U14748 (N_14748,N_11359,N_11155);
xnor U14749 (N_14749,N_9994,N_10751);
and U14750 (N_14750,N_11212,N_10308);
nand U14751 (N_14751,N_9225,N_11500);
nor U14752 (N_14752,N_11664,N_11420);
xor U14753 (N_14753,N_10742,N_10228);
nand U14754 (N_14754,N_11671,N_11133);
nor U14755 (N_14755,N_9339,N_9098);
or U14756 (N_14756,N_11970,N_9022);
nor U14757 (N_14757,N_9842,N_9768);
or U14758 (N_14758,N_10300,N_9839);
or U14759 (N_14759,N_10789,N_9851);
xor U14760 (N_14760,N_11357,N_10008);
and U14761 (N_14761,N_11341,N_11418);
or U14762 (N_14762,N_11254,N_9679);
xnor U14763 (N_14763,N_11104,N_11108);
xor U14764 (N_14764,N_9712,N_10948);
nor U14765 (N_14765,N_10034,N_10938);
xnor U14766 (N_14766,N_9961,N_11405);
or U14767 (N_14767,N_11591,N_11937);
or U14768 (N_14768,N_11194,N_9967);
nand U14769 (N_14769,N_10751,N_11073);
nor U14770 (N_14770,N_11401,N_10561);
xor U14771 (N_14771,N_10298,N_11405);
nor U14772 (N_14772,N_10160,N_10734);
nand U14773 (N_14773,N_11946,N_9539);
nor U14774 (N_14774,N_9264,N_10020);
and U14775 (N_14775,N_11115,N_11873);
nand U14776 (N_14776,N_10406,N_11269);
and U14777 (N_14777,N_9977,N_11071);
nor U14778 (N_14778,N_9268,N_9692);
or U14779 (N_14779,N_11023,N_9770);
nor U14780 (N_14780,N_10402,N_9199);
nor U14781 (N_14781,N_9493,N_10173);
xnor U14782 (N_14782,N_11863,N_10347);
xnor U14783 (N_14783,N_11489,N_10002);
and U14784 (N_14784,N_9041,N_9209);
nor U14785 (N_14785,N_11212,N_11628);
xor U14786 (N_14786,N_11724,N_10706);
nand U14787 (N_14787,N_9305,N_11583);
and U14788 (N_14788,N_10421,N_11001);
or U14789 (N_14789,N_11320,N_11676);
or U14790 (N_14790,N_9962,N_9048);
nand U14791 (N_14791,N_11069,N_11537);
nor U14792 (N_14792,N_10744,N_9141);
nand U14793 (N_14793,N_9627,N_11362);
and U14794 (N_14794,N_9637,N_9442);
nand U14795 (N_14795,N_11607,N_11220);
nand U14796 (N_14796,N_10785,N_10827);
nand U14797 (N_14797,N_11587,N_9166);
or U14798 (N_14798,N_9456,N_9355);
and U14799 (N_14799,N_10457,N_11963);
or U14800 (N_14800,N_9575,N_11200);
or U14801 (N_14801,N_10477,N_9415);
and U14802 (N_14802,N_10936,N_10344);
nand U14803 (N_14803,N_10939,N_11651);
and U14804 (N_14804,N_10763,N_9073);
or U14805 (N_14805,N_11750,N_10697);
xor U14806 (N_14806,N_9666,N_10050);
nor U14807 (N_14807,N_9841,N_9047);
xnor U14808 (N_14808,N_10556,N_11237);
or U14809 (N_14809,N_10020,N_11305);
nand U14810 (N_14810,N_10589,N_10620);
or U14811 (N_14811,N_9181,N_10024);
xnor U14812 (N_14812,N_10822,N_10064);
xnor U14813 (N_14813,N_11609,N_9929);
xor U14814 (N_14814,N_11979,N_11142);
nor U14815 (N_14815,N_10455,N_9609);
xnor U14816 (N_14816,N_9987,N_11988);
and U14817 (N_14817,N_11802,N_11857);
nor U14818 (N_14818,N_9346,N_11164);
nor U14819 (N_14819,N_11886,N_10995);
nand U14820 (N_14820,N_9939,N_11164);
nand U14821 (N_14821,N_9240,N_11475);
or U14822 (N_14822,N_9884,N_11334);
xnor U14823 (N_14823,N_9550,N_9609);
nand U14824 (N_14824,N_11872,N_9531);
nor U14825 (N_14825,N_9188,N_10428);
nor U14826 (N_14826,N_10096,N_11712);
and U14827 (N_14827,N_11304,N_11263);
and U14828 (N_14828,N_11279,N_10473);
nand U14829 (N_14829,N_9960,N_9025);
and U14830 (N_14830,N_11404,N_11049);
or U14831 (N_14831,N_9893,N_11532);
nor U14832 (N_14832,N_9223,N_11243);
and U14833 (N_14833,N_11507,N_11350);
nor U14834 (N_14834,N_9192,N_11644);
xor U14835 (N_14835,N_10993,N_10864);
or U14836 (N_14836,N_9323,N_11457);
xor U14837 (N_14837,N_10247,N_9560);
and U14838 (N_14838,N_10299,N_10625);
xnor U14839 (N_14839,N_10792,N_10891);
nand U14840 (N_14840,N_9460,N_11632);
or U14841 (N_14841,N_11816,N_10542);
and U14842 (N_14842,N_9330,N_9302);
xnor U14843 (N_14843,N_9452,N_10350);
xnor U14844 (N_14844,N_11000,N_10904);
xnor U14845 (N_14845,N_9898,N_9192);
or U14846 (N_14846,N_10536,N_11322);
and U14847 (N_14847,N_11286,N_9568);
nand U14848 (N_14848,N_11060,N_11360);
xnor U14849 (N_14849,N_11736,N_9688);
or U14850 (N_14850,N_9484,N_9151);
xor U14851 (N_14851,N_10113,N_10931);
and U14852 (N_14852,N_9579,N_10747);
xor U14853 (N_14853,N_11013,N_9541);
nand U14854 (N_14854,N_10571,N_9086);
xor U14855 (N_14855,N_9353,N_11369);
xor U14856 (N_14856,N_10201,N_10365);
xnor U14857 (N_14857,N_11529,N_9239);
xnor U14858 (N_14858,N_10788,N_9454);
or U14859 (N_14859,N_10857,N_11139);
nor U14860 (N_14860,N_11797,N_10863);
nand U14861 (N_14861,N_10654,N_9314);
and U14862 (N_14862,N_11371,N_9670);
and U14863 (N_14863,N_10058,N_9008);
and U14864 (N_14864,N_11846,N_11844);
xnor U14865 (N_14865,N_9934,N_11173);
and U14866 (N_14866,N_9312,N_9459);
and U14867 (N_14867,N_9715,N_11637);
and U14868 (N_14868,N_10944,N_10924);
xor U14869 (N_14869,N_11005,N_11955);
or U14870 (N_14870,N_10889,N_10153);
or U14871 (N_14871,N_11584,N_11863);
xor U14872 (N_14872,N_9957,N_9086);
nand U14873 (N_14873,N_11951,N_10091);
nand U14874 (N_14874,N_11953,N_10395);
xor U14875 (N_14875,N_11652,N_10710);
xor U14876 (N_14876,N_9083,N_10941);
nor U14877 (N_14877,N_9747,N_9463);
and U14878 (N_14878,N_10928,N_10105);
nor U14879 (N_14879,N_9087,N_10913);
or U14880 (N_14880,N_10350,N_11285);
nor U14881 (N_14881,N_11880,N_11988);
and U14882 (N_14882,N_10759,N_9587);
and U14883 (N_14883,N_10027,N_9800);
nor U14884 (N_14884,N_10873,N_11106);
xnor U14885 (N_14885,N_10516,N_10807);
and U14886 (N_14886,N_11864,N_10861);
nor U14887 (N_14887,N_10460,N_11856);
or U14888 (N_14888,N_10851,N_9634);
nor U14889 (N_14889,N_9481,N_11370);
nor U14890 (N_14890,N_10465,N_11053);
nor U14891 (N_14891,N_10096,N_9270);
and U14892 (N_14892,N_10796,N_9434);
xor U14893 (N_14893,N_10405,N_10347);
nor U14894 (N_14894,N_10010,N_9557);
xor U14895 (N_14895,N_9757,N_9138);
xor U14896 (N_14896,N_11602,N_9478);
nor U14897 (N_14897,N_11264,N_10334);
or U14898 (N_14898,N_11282,N_9259);
or U14899 (N_14899,N_10890,N_11982);
nor U14900 (N_14900,N_10775,N_9537);
nand U14901 (N_14901,N_11258,N_10924);
or U14902 (N_14902,N_11953,N_9094);
nand U14903 (N_14903,N_10460,N_10662);
or U14904 (N_14904,N_10165,N_11703);
xnor U14905 (N_14905,N_9058,N_11447);
and U14906 (N_14906,N_9785,N_11374);
nand U14907 (N_14907,N_10952,N_11967);
or U14908 (N_14908,N_11006,N_11531);
nor U14909 (N_14909,N_9027,N_10383);
xor U14910 (N_14910,N_9023,N_10610);
and U14911 (N_14911,N_9715,N_11342);
nand U14912 (N_14912,N_10803,N_11803);
xnor U14913 (N_14913,N_10662,N_10894);
or U14914 (N_14914,N_11191,N_9805);
nand U14915 (N_14915,N_9208,N_11460);
nor U14916 (N_14916,N_9991,N_11328);
xnor U14917 (N_14917,N_11159,N_10908);
nor U14918 (N_14918,N_9571,N_9404);
nor U14919 (N_14919,N_11693,N_11935);
and U14920 (N_14920,N_11196,N_11818);
nand U14921 (N_14921,N_9020,N_10609);
and U14922 (N_14922,N_10739,N_9162);
nor U14923 (N_14923,N_11170,N_9608);
or U14924 (N_14924,N_9367,N_11594);
nor U14925 (N_14925,N_10351,N_10545);
or U14926 (N_14926,N_9191,N_11566);
xor U14927 (N_14927,N_9726,N_11673);
and U14928 (N_14928,N_10574,N_9535);
nand U14929 (N_14929,N_9952,N_10675);
nor U14930 (N_14930,N_11918,N_11260);
or U14931 (N_14931,N_9296,N_9706);
or U14932 (N_14932,N_11185,N_10948);
xnor U14933 (N_14933,N_11922,N_9499);
xor U14934 (N_14934,N_10043,N_10731);
or U14935 (N_14935,N_10155,N_11704);
nand U14936 (N_14936,N_10079,N_11731);
nand U14937 (N_14937,N_10411,N_11846);
and U14938 (N_14938,N_11540,N_10764);
nand U14939 (N_14939,N_10382,N_11177);
nand U14940 (N_14940,N_10823,N_10524);
nor U14941 (N_14941,N_10012,N_11721);
nand U14942 (N_14942,N_10720,N_9478);
xor U14943 (N_14943,N_10902,N_10483);
xnor U14944 (N_14944,N_10479,N_10847);
and U14945 (N_14945,N_10218,N_10139);
xor U14946 (N_14946,N_11562,N_10102);
or U14947 (N_14947,N_9201,N_11370);
or U14948 (N_14948,N_11242,N_10694);
nor U14949 (N_14949,N_10168,N_10805);
or U14950 (N_14950,N_10380,N_10149);
xnor U14951 (N_14951,N_9297,N_10019);
nand U14952 (N_14952,N_11550,N_10916);
and U14953 (N_14953,N_9484,N_9589);
or U14954 (N_14954,N_10033,N_11964);
nand U14955 (N_14955,N_11788,N_9605);
nand U14956 (N_14956,N_10863,N_10721);
nor U14957 (N_14957,N_11714,N_10948);
or U14958 (N_14958,N_10366,N_11093);
xor U14959 (N_14959,N_11657,N_10708);
and U14960 (N_14960,N_9290,N_10418);
nor U14961 (N_14961,N_10572,N_11355);
nor U14962 (N_14962,N_11528,N_11526);
nand U14963 (N_14963,N_9936,N_10329);
nand U14964 (N_14964,N_10896,N_11542);
xnor U14965 (N_14965,N_10632,N_9554);
or U14966 (N_14966,N_9177,N_9608);
or U14967 (N_14967,N_10249,N_11279);
nor U14968 (N_14968,N_11064,N_10696);
nand U14969 (N_14969,N_11727,N_11429);
nand U14970 (N_14970,N_10585,N_10919);
nor U14971 (N_14971,N_9892,N_11904);
nor U14972 (N_14972,N_10685,N_9825);
and U14973 (N_14973,N_9725,N_9825);
nand U14974 (N_14974,N_10350,N_10357);
xnor U14975 (N_14975,N_11482,N_11906);
and U14976 (N_14976,N_11130,N_9638);
xnor U14977 (N_14977,N_10692,N_11926);
and U14978 (N_14978,N_9706,N_10250);
and U14979 (N_14979,N_11589,N_11508);
nand U14980 (N_14980,N_10409,N_9718);
nand U14981 (N_14981,N_10163,N_10961);
nand U14982 (N_14982,N_9224,N_10011);
nand U14983 (N_14983,N_11731,N_9903);
and U14984 (N_14984,N_11427,N_9298);
nor U14985 (N_14985,N_9424,N_9669);
xor U14986 (N_14986,N_11170,N_9769);
nor U14987 (N_14987,N_9330,N_11322);
nand U14988 (N_14988,N_9752,N_9933);
and U14989 (N_14989,N_11370,N_11751);
xor U14990 (N_14990,N_11042,N_10549);
and U14991 (N_14991,N_10794,N_10229);
nor U14992 (N_14992,N_9469,N_9967);
nand U14993 (N_14993,N_10338,N_10222);
or U14994 (N_14994,N_9512,N_11732);
and U14995 (N_14995,N_9316,N_9411);
nor U14996 (N_14996,N_11754,N_11729);
and U14997 (N_14997,N_11282,N_11802);
nand U14998 (N_14998,N_11251,N_10462);
nand U14999 (N_14999,N_10170,N_10127);
nor U15000 (N_15000,N_12213,N_13439);
nand U15001 (N_15001,N_14007,N_14803);
xnor U15002 (N_15002,N_13524,N_12391);
or U15003 (N_15003,N_12680,N_13019);
xor U15004 (N_15004,N_12199,N_14793);
nand U15005 (N_15005,N_12422,N_14097);
and U15006 (N_15006,N_13667,N_13168);
and U15007 (N_15007,N_12989,N_14268);
and U15008 (N_15008,N_14246,N_13386);
and U15009 (N_15009,N_13937,N_14281);
and U15010 (N_15010,N_14758,N_14127);
nor U15011 (N_15011,N_14006,N_14103);
or U15012 (N_15012,N_13410,N_14371);
nand U15013 (N_15013,N_14972,N_12664);
nor U15014 (N_15014,N_13921,N_14947);
or U15015 (N_15015,N_13281,N_12816);
nor U15016 (N_15016,N_12076,N_13871);
and U15017 (N_15017,N_13986,N_14798);
xor U15018 (N_15018,N_12911,N_14068);
nand U15019 (N_15019,N_13167,N_14225);
or U15020 (N_15020,N_13969,N_13887);
or U15021 (N_15021,N_12333,N_12539);
nor U15022 (N_15022,N_13749,N_12345);
and U15023 (N_15023,N_14495,N_12166);
or U15024 (N_15024,N_13957,N_12194);
xor U15025 (N_15025,N_12088,N_14681);
nand U15026 (N_15026,N_13790,N_14792);
nand U15027 (N_15027,N_14005,N_14915);
nor U15028 (N_15028,N_13106,N_14756);
or U15029 (N_15029,N_12926,N_13214);
nor U15030 (N_15030,N_12826,N_14902);
xnor U15031 (N_15031,N_14968,N_14417);
nor U15032 (N_15032,N_12454,N_13597);
nand U15033 (N_15033,N_13358,N_12905);
nor U15034 (N_15034,N_12251,N_12398);
nor U15035 (N_15035,N_12399,N_14532);
or U15036 (N_15036,N_13825,N_13913);
xor U15037 (N_15037,N_12669,N_12739);
or U15038 (N_15038,N_14464,N_14847);
and U15039 (N_15039,N_14046,N_13072);
and U15040 (N_15040,N_14509,N_12029);
or U15041 (N_15041,N_14842,N_13351);
or U15042 (N_15042,N_14381,N_14908);
and U15043 (N_15043,N_12998,N_13459);
xor U15044 (N_15044,N_14649,N_12322);
or U15045 (N_15045,N_13136,N_12219);
nor U15046 (N_15046,N_13710,N_12512);
and U15047 (N_15047,N_14916,N_13763);
xnor U15048 (N_15048,N_13947,N_14468);
xor U15049 (N_15049,N_14304,N_12495);
xnor U15050 (N_15050,N_14351,N_14440);
xnor U15051 (N_15051,N_14493,N_13146);
nand U15052 (N_15052,N_14675,N_12145);
or U15053 (N_15053,N_12556,N_12176);
or U15054 (N_15054,N_12589,N_14372);
or U15055 (N_15055,N_13276,N_12943);
nand U15056 (N_15056,N_14621,N_12690);
or U15057 (N_15057,N_12853,N_14358);
nor U15058 (N_15058,N_12524,N_13850);
and U15059 (N_15059,N_13722,N_14602);
nand U15060 (N_15060,N_14737,N_12515);
or U15061 (N_15061,N_13251,N_12749);
or U15062 (N_15062,N_12559,N_13062);
nor U15063 (N_15063,N_14749,N_13028);
or U15064 (N_15064,N_12864,N_12000);
nor U15065 (N_15065,N_13772,N_14739);
and U15066 (N_15066,N_13200,N_13538);
xor U15067 (N_15067,N_12658,N_12234);
or U15068 (N_15068,N_14456,N_13342);
or U15069 (N_15069,N_13513,N_12041);
nor U15070 (N_15070,N_14134,N_13354);
xor U15071 (N_15071,N_12829,N_13254);
nand U15072 (N_15072,N_13783,N_13615);
and U15073 (N_15073,N_13040,N_12462);
or U15074 (N_15074,N_14132,N_12736);
and U15075 (N_15075,N_13693,N_13944);
nand U15076 (N_15076,N_12184,N_14364);
nor U15077 (N_15077,N_13742,N_14411);
and U15078 (N_15078,N_14685,N_14011);
xor U15079 (N_15079,N_14540,N_13553);
or U15080 (N_15080,N_12206,N_13719);
nor U15081 (N_15081,N_12730,N_14526);
nand U15082 (N_15082,N_12476,N_13976);
or U15083 (N_15083,N_12057,N_12668);
nor U15084 (N_15084,N_13148,N_13343);
and U15085 (N_15085,N_13467,N_14563);
xor U15086 (N_15086,N_12175,N_12483);
or U15087 (N_15087,N_14484,N_14565);
xnor U15088 (N_15088,N_12726,N_12182);
xor U15089 (N_15089,N_14619,N_14555);
nand U15090 (N_15090,N_12337,N_13882);
nand U15091 (N_15091,N_12205,N_14652);
xnor U15092 (N_15092,N_13177,N_13569);
and U15093 (N_15093,N_14929,N_13543);
and U15094 (N_15094,N_14935,N_14818);
and U15095 (N_15095,N_14766,N_14956);
nor U15096 (N_15096,N_13641,N_12044);
or U15097 (N_15097,N_13367,N_12456);
xor U15098 (N_15098,N_13691,N_12858);
xor U15099 (N_15099,N_13020,N_12444);
xor U15100 (N_15100,N_14668,N_13567);
xor U15101 (N_15101,N_12441,N_13816);
nand U15102 (N_15102,N_14030,N_13753);
nor U15103 (N_15103,N_12046,N_12949);
and U15104 (N_15104,N_14163,N_12033);
nor U15105 (N_15105,N_13007,N_13789);
or U15106 (N_15106,N_14362,N_12494);
and U15107 (N_15107,N_12626,N_13462);
xnor U15108 (N_15108,N_14850,N_14400);
xor U15109 (N_15109,N_14500,N_13156);
or U15110 (N_15110,N_14461,N_13978);
nor U15111 (N_15111,N_14707,N_12171);
nand U15112 (N_15112,N_12484,N_14794);
nor U15113 (N_15113,N_14193,N_14647);
nand U15114 (N_15114,N_13610,N_13003);
nor U15115 (N_15115,N_13183,N_13397);
nor U15116 (N_15116,N_14187,N_12957);
xor U15117 (N_15117,N_13135,N_13744);
nor U15118 (N_15118,N_14004,N_12112);
xnor U15119 (N_15119,N_14407,N_13891);
or U15120 (N_15120,N_12245,N_12226);
xor U15121 (N_15121,N_13005,N_14379);
xnor U15122 (N_15122,N_13406,N_14892);
and U15123 (N_15123,N_14871,N_14595);
nand U15124 (N_15124,N_14895,N_13356);
xnor U15125 (N_15125,N_14999,N_12884);
or U15126 (N_15126,N_14042,N_12636);
nand U15127 (N_15127,N_13290,N_13124);
nand U15128 (N_15128,N_12080,N_12666);
or U15129 (N_15129,N_12734,N_13131);
nor U15130 (N_15130,N_13961,N_13242);
or U15131 (N_15131,N_13466,N_12147);
or U15132 (N_15132,N_13125,N_12971);
and U15133 (N_15133,N_12903,N_12623);
xnor U15134 (N_15134,N_12603,N_12792);
nor U15135 (N_15135,N_14688,N_14917);
or U15136 (N_15136,N_12237,N_14251);
xnor U15137 (N_15137,N_14615,N_13048);
and U15138 (N_15138,N_14213,N_14995);
nor U15139 (N_15139,N_14264,N_13333);
and U15140 (N_15140,N_14777,N_14541);
nand U15141 (N_15141,N_13872,N_14611);
or U15142 (N_15142,N_13626,N_14087);
nor U15143 (N_15143,N_13540,N_14171);
and U15144 (N_15144,N_14853,N_14912);
nor U15145 (N_15145,N_14963,N_12093);
nor U15146 (N_15146,N_13927,N_12577);
xor U15147 (N_15147,N_13883,N_13951);
nor U15148 (N_15148,N_12125,N_14879);
and U15149 (N_15149,N_12875,N_14120);
and U15150 (N_15150,N_14763,N_12915);
nor U15151 (N_15151,N_12413,N_13192);
nand U15152 (N_15152,N_12394,N_12329);
xnor U15153 (N_15153,N_13987,N_14455);
xor U15154 (N_15154,N_13274,N_13534);
or U15155 (N_15155,N_12780,N_12448);
nor U15156 (N_15156,N_13811,N_14557);
xnor U15157 (N_15157,N_12975,N_12563);
nor U15158 (N_15158,N_12617,N_12340);
or U15159 (N_15159,N_12540,N_13181);
and U15160 (N_15160,N_12131,N_14476);
or U15161 (N_15161,N_12350,N_12066);
nand U15162 (N_15162,N_14978,N_13039);
and U15163 (N_15163,N_14144,N_12477);
nor U15164 (N_15164,N_13585,N_14740);
and U15165 (N_15165,N_14123,N_13703);
nor U15166 (N_15166,N_14458,N_13983);
xor U15167 (N_15167,N_13948,N_12202);
nor U15168 (N_15168,N_12355,N_12286);
and U15169 (N_15169,N_12635,N_13770);
nor U15170 (N_15170,N_13522,N_14599);
xor U15171 (N_15171,N_13227,N_14781);
nor U15172 (N_15172,N_13884,N_12160);
xor U15173 (N_15173,N_13328,N_13592);
and U15174 (N_15174,N_12745,N_13133);
nand U15175 (N_15175,N_13403,N_14911);
nor U15176 (N_15176,N_12607,N_14833);
and U15177 (N_15177,N_13207,N_13633);
nor U15178 (N_15178,N_12373,N_13849);
nand U15179 (N_15179,N_13088,N_14229);
nand U15180 (N_15180,N_12082,N_13676);
and U15181 (N_15181,N_14823,N_12279);
and U15182 (N_15182,N_14930,N_13739);
nand U15183 (N_15183,N_12002,N_14848);
or U15184 (N_15184,N_14319,N_13025);
or U15185 (N_15185,N_13143,N_12114);
xnor U15186 (N_15186,N_14328,N_13226);
xor U15187 (N_15187,N_13490,N_12438);
nor U15188 (N_15188,N_13249,N_14349);
and U15189 (N_15189,N_14648,N_12225);
and U15190 (N_15190,N_14657,N_13715);
xor U15191 (N_15191,N_13940,N_12302);
and U15192 (N_15192,N_14320,N_12528);
xnor U15193 (N_15193,N_13886,N_12346);
or U15194 (N_15194,N_14589,N_13400);
nand U15195 (N_15195,N_13260,N_13660);
nand U15196 (N_15196,N_12580,N_14402);
and U15197 (N_15197,N_13984,N_14782);
or U15198 (N_15198,N_13210,N_13321);
nand U15199 (N_15199,N_13711,N_14701);
and U15200 (N_15200,N_12595,N_14726);
xor U15201 (N_15201,N_12897,N_12283);
or U15202 (N_15202,N_14141,N_12157);
xnor U15203 (N_15203,N_12600,N_12096);
and U15204 (N_15204,N_14906,N_12017);
and U15205 (N_15205,N_12847,N_12833);
nand U15206 (N_15206,N_12011,N_13436);
nand U15207 (N_15207,N_13875,N_12244);
and U15208 (N_15208,N_14918,N_13587);
or U15209 (N_15209,N_14061,N_12266);
nor U15210 (N_15210,N_13701,N_12689);
and U15211 (N_15211,N_12253,N_12755);
nand U15212 (N_15212,N_14603,N_13113);
or U15213 (N_15213,N_12781,N_12168);
xor U15214 (N_15214,N_12397,N_12738);
and U15215 (N_15215,N_13175,N_13155);
and U15216 (N_15216,N_14969,N_12813);
nand U15217 (N_15217,N_12910,N_13578);
or U15218 (N_15218,N_13994,N_14815);
or U15219 (N_15219,N_14812,N_13809);
or U15220 (N_15220,N_13129,N_14125);
nor U15221 (N_15221,N_13182,N_13221);
or U15222 (N_15222,N_12697,N_12613);
nand U15223 (N_15223,N_13493,N_14583);
or U15224 (N_15224,N_13187,N_13097);
or U15225 (N_15225,N_14716,N_12652);
xnor U15226 (N_15226,N_14183,N_13824);
and U15227 (N_15227,N_12830,N_12846);
or U15228 (N_15228,N_14222,N_14462);
and U15229 (N_15229,N_14425,N_13017);
and U15230 (N_15230,N_13591,N_12174);
and U15231 (N_15231,N_13119,N_12047);
xor U15232 (N_15232,N_13154,N_13669);
nor U15233 (N_15233,N_12103,N_14430);
nor U15234 (N_15234,N_13504,N_13705);
xor U15235 (N_15235,N_13305,N_12179);
and U15236 (N_15236,N_12966,N_13902);
xor U15237 (N_15237,N_14830,N_13552);
xor U15238 (N_15238,N_12498,N_13781);
and U15239 (N_15239,N_14478,N_14406);
nor U15240 (N_15240,N_13145,N_14780);
or U15241 (N_15241,N_12775,N_14333);
xor U15242 (N_15242,N_12224,N_12463);
nor U15243 (N_15243,N_13974,N_13924);
or U15244 (N_15244,N_12542,N_14070);
or U15245 (N_15245,N_12885,N_12642);
and U15246 (N_15246,N_13029,N_12744);
xnor U15247 (N_15247,N_13943,N_12034);
nand U15248 (N_15248,N_12371,N_14426);
and U15249 (N_15249,N_14962,N_13796);
and U15250 (N_15250,N_14142,N_12190);
xor U15251 (N_15251,N_12963,N_13302);
and U15252 (N_15252,N_13688,N_13053);
or U15253 (N_15253,N_13928,N_12758);
nor U15254 (N_15254,N_13223,N_12920);
and U15255 (N_15255,N_13413,N_13656);
xor U15256 (N_15256,N_13117,N_13134);
xor U15257 (N_15257,N_13399,N_13383);
xor U15258 (N_15258,N_12056,N_13568);
nor U15259 (N_15259,N_12356,N_14475);
or U15260 (N_15260,N_14301,N_12369);
and U15261 (N_15261,N_14938,N_12578);
xor U15262 (N_15262,N_14308,N_12122);
or U15263 (N_15263,N_14022,N_14861);
xor U15264 (N_15264,N_12300,N_12774);
xor U15265 (N_15265,N_13162,N_14888);
xnor U15266 (N_15266,N_12250,N_13271);
or U15267 (N_15267,N_12073,N_12126);
or U15268 (N_15268,N_14044,N_14785);
nand U15269 (N_15269,N_13959,N_13191);
xnor U15270 (N_15270,N_12714,N_13843);
or U15271 (N_15271,N_14682,N_13714);
nand U15272 (N_15272,N_14762,N_13205);
nand U15273 (N_15273,N_12376,N_14883);
xor U15274 (N_15274,N_14829,N_12788);
and U15275 (N_15275,N_13692,N_13074);
xor U15276 (N_15276,N_14345,N_13139);
nor U15277 (N_15277,N_14985,N_14241);
nand U15278 (N_15278,N_14161,N_12660);
nor U15279 (N_15279,N_13889,N_12104);
xnor U15280 (N_15280,N_14029,N_13069);
or U15281 (N_15281,N_12328,N_14677);
nand U15282 (N_15282,N_14961,N_12985);
xnor U15283 (N_15283,N_14288,N_14531);
or U15284 (N_15284,N_12465,N_14421);
xnor U15285 (N_15285,N_13225,N_14820);
or U15286 (N_15286,N_13479,N_14567);
xnor U15287 (N_15287,N_14728,N_12220);
nand U15288 (N_15288,N_12261,N_12021);
nor U15289 (N_15289,N_13679,N_13516);
nor U15290 (N_15290,N_14428,N_14491);
and U15291 (N_15291,N_12880,N_14365);
or U15292 (N_15292,N_14732,N_12229);
xor U15293 (N_15293,N_14223,N_12865);
and U15294 (N_15294,N_13093,N_12488);
or U15295 (N_15295,N_12363,N_12639);
and U15296 (N_15296,N_13560,N_12027);
or U15297 (N_15297,N_14401,N_13417);
and U15298 (N_15298,N_13846,N_14653);
nand U15299 (N_15299,N_12348,N_13474);
nand U15300 (N_15300,N_12933,N_12522);
nand U15301 (N_15301,N_13502,N_12952);
nand U15302 (N_15302,N_12516,N_12324);
nand U15303 (N_15303,N_12361,N_14723);
xor U15304 (N_15304,N_14039,N_13256);
xor U15305 (N_15305,N_12485,N_13078);
and U15306 (N_15306,N_14506,N_14561);
nor U15307 (N_15307,N_14822,N_13378);
xor U15308 (N_15308,N_14524,N_14954);
and U15309 (N_15309,N_12930,N_14152);
nor U15310 (N_15310,N_14233,N_13863);
or U15311 (N_15311,N_12007,N_13021);
or U15312 (N_15312,N_12272,N_14252);
xnor U15313 (N_15313,N_12703,N_14078);
nor U15314 (N_15314,N_14897,N_12567);
nand U15315 (N_15315,N_13385,N_12979);
nand U15316 (N_15316,N_14274,N_12873);
or U15317 (N_15317,N_13334,N_14443);
xnor U15318 (N_15318,N_14130,N_12616);
nand U15319 (N_15319,N_13949,N_14975);
and U15320 (N_15320,N_13868,N_13603);
and U15321 (N_15321,N_12298,N_14368);
or U15322 (N_15322,N_14922,N_14247);
xnor U15323 (N_15323,N_12866,N_14654);
xor U15324 (N_15324,N_12503,N_12432);
nor U15325 (N_15325,N_14040,N_13644);
and U15326 (N_15326,N_13694,N_12746);
nand U15327 (N_15327,N_13391,N_14549);
or U15328 (N_15328,N_14587,N_12051);
nor U15329 (N_15329,N_12152,N_12845);
and U15330 (N_15330,N_13392,N_12777);
nor U15331 (N_15331,N_12657,N_13440);
xnor U15332 (N_15332,N_13132,N_12579);
xnor U15333 (N_15333,N_13726,N_12821);
nor U15334 (N_15334,N_12215,N_12216);
and U15335 (N_15335,N_14439,N_13509);
or U15336 (N_15336,N_14987,N_13277);
and U15337 (N_15337,N_12238,N_14361);
and U15338 (N_15338,N_14457,N_14168);
nand U15339 (N_15339,N_14138,N_14091);
and U15340 (N_15340,N_12869,N_13602);
nand U15341 (N_15341,N_12115,N_12951);
xnor U15342 (N_15342,N_14318,N_12505);
or U15343 (N_15343,N_14121,N_13613);
nand U15344 (N_15344,N_12123,N_13527);
and U15345 (N_15345,N_13776,N_14422);
xnor U15346 (N_15346,N_14750,N_12791);
nand U15347 (N_15347,N_12709,N_13185);
nand U15348 (N_15348,N_13962,N_13120);
nand U15349 (N_15349,N_14547,N_14660);
nand U15350 (N_15350,N_14979,N_13609);
xnor U15351 (N_15351,N_14859,N_14394);
nand U15352 (N_15352,N_13506,N_12451);
or U15353 (N_15353,N_13993,N_13465);
xnor U15354 (N_15354,N_13661,N_12466);
nand U15355 (N_15355,N_13443,N_13166);
xor U15356 (N_15356,N_14169,N_12135);
nand U15357 (N_15357,N_13786,N_12053);
xor U15358 (N_15358,N_14083,N_12936);
or U15359 (N_15359,N_14271,N_13275);
or U15360 (N_15360,N_13011,N_12545);
nand U15361 (N_15361,N_14625,N_13903);
and U15362 (N_15362,N_14207,N_13680);
nand U15363 (N_15363,N_13265,N_14092);
and U15364 (N_15364,N_13586,N_12043);
and U15365 (N_15365,N_12091,N_14463);
xor U15366 (N_15366,N_13027,N_14612);
and U15367 (N_15367,N_14810,N_13532);
nor U15368 (N_15368,N_12955,N_12392);
and U15369 (N_15369,N_12544,N_12032);
and U15370 (N_15370,N_13101,N_14018);
and U15371 (N_15371,N_12415,N_14118);
nand U15372 (N_15372,N_14324,N_12111);
xnor U15373 (N_15373,N_12785,N_14096);
or U15374 (N_15374,N_14727,N_12994);
xnor U15375 (N_15375,N_14572,N_14736);
or U15376 (N_15376,N_14444,N_14661);
and U15377 (N_15377,N_14951,N_13267);
nor U15378 (N_15378,N_12416,N_12139);
xor U15379 (N_15379,N_12059,N_14700);
or U15380 (N_15380,N_13252,N_12349);
nor U15381 (N_15381,N_13582,N_12177);
nor U15382 (N_15382,N_13057,N_14715);
and U15383 (N_15383,N_14131,N_14380);
and U15384 (N_15384,N_13463,N_13870);
xor U15385 (N_15385,N_14986,N_14576);
nor U15386 (N_15386,N_14585,N_14388);
nand U15387 (N_15387,N_12410,N_13127);
or U15388 (N_15388,N_14202,N_13831);
or U15389 (N_15389,N_12042,N_14913);
nand U15390 (N_15390,N_14841,N_12264);
nor U15391 (N_15391,N_13662,N_12742);
nand U15392 (N_15392,N_14721,N_14195);
xnor U15393 (N_15393,N_13398,N_13898);
xor U15394 (N_15394,N_12519,N_13310);
and U15395 (N_15395,N_14627,N_14082);
or U15396 (N_15396,N_14206,N_13890);
or U15397 (N_15397,N_12314,N_12321);
or U15398 (N_15398,N_12651,N_13222);
nand U15399 (N_15399,N_13013,N_12881);
nand U15400 (N_15400,N_14139,N_12638);
nor U15401 (N_15401,N_14694,N_12417);
or U15402 (N_15402,N_13738,N_12712);
xnor U15403 (N_15403,N_13432,N_12260);
xor U15404 (N_15404,N_14024,N_12601);
xor U15405 (N_15405,N_12079,N_13211);
nor U15406 (N_15406,N_13897,N_14373);
and U15407 (N_15407,N_14423,N_13515);
and U15408 (N_15408,N_12854,N_12271);
xnor U15409 (N_15409,N_13032,N_13652);
and U15410 (N_15410,N_14335,N_14340);
and U15411 (N_15411,N_12270,N_12497);
or U15412 (N_15412,N_14573,N_14086);
nor U15413 (N_15413,N_13253,N_13216);
nor U15414 (N_15414,N_12729,N_14544);
and U15415 (N_15415,N_14940,N_12307);
nand U15416 (N_15416,N_12287,N_13488);
nor U15417 (N_15417,N_14575,N_14215);
and U15418 (N_15418,N_12561,N_12453);
or U15419 (N_15419,N_14946,N_13838);
or U15420 (N_15420,N_13307,N_13409);
and U15421 (N_15421,N_12900,N_14391);
xor U15422 (N_15422,N_14899,N_14941);
xnor U15423 (N_15423,N_14058,N_14260);
or U15424 (N_15424,N_13499,N_12870);
xnor U15425 (N_15425,N_14480,N_13681);
nor U15426 (N_15426,N_14415,N_13746);
and U15427 (N_15427,N_14932,N_12455);
nand U15428 (N_15428,N_13584,N_13699);
or U15429 (N_15429,N_12388,N_14639);
nand U15430 (N_15430,N_13985,N_14560);
xnor U15431 (N_15431,N_13034,N_12811);
nand U15432 (N_15432,N_12895,N_12209);
and U15433 (N_15433,N_13230,N_14197);
nor U15434 (N_15434,N_14891,N_12183);
xnor U15435 (N_15435,N_14662,N_12711);
xor U15436 (N_15436,N_14433,N_13238);
nand U15437 (N_15437,N_14966,N_13458);
and U15438 (N_15438,N_12201,N_14176);
and U15439 (N_15439,N_14997,N_12045);
nand U15440 (N_15440,N_14671,N_13123);
xor U15441 (N_15441,N_14937,N_14343);
nand U15442 (N_15442,N_14106,N_12193);
nor U15443 (N_15443,N_13353,N_12670);
xnor U15444 (N_15444,N_13282,N_13394);
nor U15445 (N_15445,N_14242,N_13655);
nand U15446 (N_15446,N_12850,N_14538);
or U15447 (N_15447,N_12269,N_14837);
nand U15448 (N_15448,N_13745,N_12360);
nor U15449 (N_15449,N_13817,N_12396);
xor U15450 (N_15450,N_12095,N_12169);
nor U15451 (N_15451,N_13379,N_14684);
and U15452 (N_15452,N_13115,N_12604);
xor U15453 (N_15453,N_13009,N_12486);
or U15454 (N_15454,N_12647,N_12482);
and U15455 (N_15455,N_12297,N_14977);
or U15456 (N_15456,N_12984,N_13659);
or U15457 (N_15457,N_14360,N_13654);
xor U15458 (N_15458,N_13931,N_14839);
and U15459 (N_15459,N_12493,N_12764);
nand U15460 (N_15460,N_14105,N_12819);
or U15461 (N_15461,N_14175,N_13452);
or U15462 (N_15462,N_14156,N_12335);
xnor U15463 (N_15463,N_14693,N_13451);
nand U15464 (N_15464,N_12236,N_13808);
nor U15465 (N_15465,N_13186,N_12389);
and U15466 (N_15466,N_13064,N_13503);
or U15467 (N_15467,N_12980,N_14137);
and U15468 (N_15468,N_12167,N_14026);
xor U15469 (N_15469,N_14702,N_14814);
or U15470 (N_15470,N_13218,N_13634);
and U15471 (N_15471,N_13345,N_12706);
and U15472 (N_15472,N_12402,N_12150);
xnor U15473 (N_15473,N_14552,N_13043);
nand U15474 (N_15474,N_13593,N_12390);
nor U15475 (N_15475,N_12084,N_13730);
nor U15476 (N_15476,N_14746,N_14687);
or U15477 (N_15477,N_12976,N_14590);
nor U15478 (N_15478,N_13401,N_14043);
or U15479 (N_15479,N_13472,N_14686);
nor U15480 (N_15480,N_14192,N_12221);
xor U15481 (N_15481,N_13579,N_13911);
nor U15482 (N_15482,N_14133,N_13901);
nor U15483 (N_15483,N_13565,N_13718);
nor U15484 (N_15484,N_13247,N_12228);
nor U15485 (N_15485,N_12204,N_12377);
or U15486 (N_15486,N_14704,N_13338);
or U15487 (N_15487,N_14285,N_12550);
nand U15488 (N_15488,N_14370,N_14224);
or U15489 (N_15489,N_12208,N_13648);
nor U15490 (N_15490,N_12421,N_13697);
and U15491 (N_15491,N_14438,N_14632);
and U15492 (N_15492,N_13341,N_14243);
xnor U15493 (N_15493,N_13623,N_14479);
or U15494 (N_15494,N_14220,N_13500);
and U15495 (N_15495,N_13165,N_12937);
or U15496 (N_15496,N_13955,N_14331);
nand U15497 (N_15497,N_12254,N_13300);
nand U15498 (N_15498,N_12916,N_13541);
or U15499 (N_15499,N_12630,N_13456);
xnor U15500 (N_15500,N_12078,N_13036);
xor U15501 (N_15501,N_12502,N_12207);
and U15502 (N_15502,N_13598,N_13232);
nand U15503 (N_15503,N_13248,N_13314);
nor U15504 (N_15504,N_12248,N_13332);
or U15505 (N_15505,N_13087,N_13349);
and U15506 (N_15506,N_12479,N_13941);
or U15507 (N_15507,N_12268,N_12518);
xnor U15508 (N_15508,N_14804,N_12013);
nor U15509 (N_15509,N_14519,N_13766);
and U15510 (N_15510,N_13787,N_12981);
nand U15511 (N_15511,N_13449,N_12958);
nand U15512 (N_15512,N_13874,N_13651);
nor U15513 (N_15513,N_12301,N_12585);
and U15514 (N_15514,N_14258,N_13665);
nor U15515 (N_15515,N_14332,N_13303);
nand U15516 (N_15516,N_13429,N_14352);
xor U15517 (N_15517,N_12655,N_13357);
nor U15518 (N_15518,N_13382,N_14846);
or U15519 (N_15519,N_14870,N_14582);
and U15520 (N_15520,N_13990,N_13860);
xnor U15521 (N_15521,N_12077,N_12852);
or U15522 (N_15522,N_14214,N_13885);
and U15523 (N_15523,N_13589,N_12089);
nand U15524 (N_15524,N_13638,N_12424);
or U15525 (N_15525,N_12433,N_12312);
xor U15526 (N_15526,N_12794,N_14038);
nor U15527 (N_15527,N_13995,N_12673);
nand U15528 (N_15528,N_13759,N_13687);
xnor U15529 (N_15529,N_13239,N_12818);
xor U15530 (N_15530,N_12565,N_14828);
xnor U15531 (N_15531,N_14805,N_14237);
nand U15532 (N_15532,N_12318,N_12538);
xnor U15533 (N_15533,N_14754,N_12927);
nand U15534 (N_15534,N_14813,N_12754);
or U15535 (N_15535,N_12347,N_13630);
xnor U15536 (N_15536,N_12282,N_13294);
or U15537 (N_15537,N_12569,N_14273);
and U15538 (N_15538,N_13373,N_13805);
or U15539 (N_15539,N_13258,N_12747);
nand U15540 (N_15540,N_13208,N_12717);
xnor U15541 (N_15541,N_12748,N_13460);
or U15542 (N_15542,N_14178,N_14672);
nand U15543 (N_15543,N_14016,N_13798);
or U15544 (N_15544,N_13704,N_13428);
and U15545 (N_15545,N_12624,N_13363);
nor U15546 (N_15546,N_14445,N_14012);
nor U15547 (N_15547,N_14277,N_13727);
nor U15548 (N_15548,N_14236,N_13301);
nand U15549 (N_15549,N_13979,N_13150);
and U15550 (N_15550,N_12891,N_14460);
nand U15551 (N_15551,N_12768,N_14635);
or U15552 (N_15552,N_12908,N_13769);
or U15553 (N_15553,N_14036,N_14412);
nor U15554 (N_15554,N_13331,N_13147);
xor U15555 (N_15555,N_13108,N_13537);
nor U15556 (N_15556,N_12574,N_14337);
nor U15557 (N_15557,N_14586,N_12072);
nor U15558 (N_15558,N_12315,N_14387);
or U15559 (N_15559,N_12809,N_13973);
and U15560 (N_15560,N_14622,N_14184);
nor U15561 (N_15561,N_13604,N_13671);
and U15562 (N_15562,N_12196,N_13573);
xnor U15563 (N_15563,N_13720,N_12532);
xnor U15564 (N_15564,N_12531,N_14071);
and U15565 (N_15565,N_12716,N_12888);
or U15566 (N_15566,N_12804,N_13658);
or U15567 (N_15567,N_13981,N_14720);
xor U15568 (N_15568,N_14626,N_14907);
or U15569 (N_15569,N_14341,N_13561);
and U15570 (N_15570,N_12319,N_13220);
xor U15571 (N_15571,N_12299,N_12537);
or U15572 (N_15572,N_14298,N_14605);
nor U15573 (N_15573,N_13529,N_14579);
nor U15574 (N_15574,N_14607,N_14928);
xor U15575 (N_15575,N_13475,N_14384);
nand U15576 (N_15576,N_12688,N_12501);
xor U15577 (N_15577,N_13476,N_13337);
nor U15578 (N_15578,N_13355,N_14090);
and U15579 (N_15579,N_14316,N_12751);
nand U15580 (N_15580,N_12143,N_14459);
or U15581 (N_15581,N_13764,N_14312);
xor U15582 (N_15582,N_12987,N_13640);
and U15583 (N_15583,N_14201,N_12119);
nor U15584 (N_15584,N_14329,N_13105);
or U15585 (N_15585,N_14588,N_13768);
nor U15586 (N_15586,N_12530,N_13618);
nor U15587 (N_15587,N_13574,N_12163);
nand U15588 (N_15588,N_13231,N_13130);
xnor U15589 (N_15589,N_12899,N_13695);
nor U15590 (N_15590,N_14390,N_12267);
nor U15591 (N_15591,N_13404,N_14027);
or U15592 (N_15592,N_13563,N_14744);
or U15593 (N_15593,N_14310,N_13137);
xnor U15594 (N_15594,N_14054,N_14179);
and U15595 (N_15595,N_12724,N_14789);
nor U15596 (N_15596,N_14747,N_12074);
and U15597 (N_15597,N_14267,N_14295);
and U15598 (N_15598,N_14146,N_14293);
and U15599 (N_15599,N_12442,N_13668);
and U15600 (N_15600,N_12434,N_12786);
or U15601 (N_15601,N_13180,N_12814);
xor U15602 (N_15602,N_13163,N_12406);
or U15603 (N_15603,N_13457,N_14494);
nand U15604 (N_15604,N_14238,N_13765);
or U15605 (N_15605,N_13508,N_13468);
and U15606 (N_15606,N_13698,N_13347);
nand U15607 (N_15607,N_13086,N_14658);
nand U15608 (N_15608,N_13169,N_13804);
nand U15609 (N_15609,N_14010,N_13754);
nand U15610 (N_15610,N_13895,N_12929);
nor U15611 (N_15611,N_12142,N_14717);
nor U15612 (N_15612,N_12700,N_13492);
nor U15613 (N_15613,N_12140,N_13862);
and U15614 (N_15614,N_12619,N_14832);
or U15615 (N_15615,N_13645,N_13344);
xnor U15616 (N_15616,N_14949,N_13395);
xnor U15617 (N_15617,N_14507,N_12148);
and U15618 (N_15618,N_13411,N_14283);
nand U15619 (N_15619,N_14550,N_13844);
xnor U15620 (N_15620,N_12507,N_14235);
nand U15621 (N_15621,N_13380,N_14286);
nor U15622 (N_15622,N_12622,N_13322);
or U15623 (N_15623,N_12491,N_13748);
nor U15624 (N_15624,N_12036,N_12065);
nor U15625 (N_15625,N_12239,N_13972);
xnor U15626 (N_15626,N_14713,N_12917);
nand U15627 (N_15627,N_12086,N_14449);
nand U15628 (N_15628,N_12120,N_13126);
nor U15629 (N_15629,N_12732,N_14976);
or U15630 (N_15630,N_14398,N_14250);
or U15631 (N_15631,N_14725,N_14350);
nand U15632 (N_15632,N_12863,N_14009);
nand U15633 (N_15633,N_13518,N_14482);
and U15634 (N_15634,N_12474,N_12364);
nand U15635 (N_15635,N_12610,N_13867);
or U15636 (N_15636,N_13551,N_12621);
nor U15637 (N_15637,N_12292,N_13173);
nor U15638 (N_15638,N_13455,N_12099);
xor U15639 (N_15639,N_12129,N_12698);
and U15640 (N_15640,N_13487,N_14473);
nor U15641 (N_15641,N_13992,N_14160);
or U15642 (N_15642,N_13496,N_13352);
and U15643 (N_15643,N_14551,N_14014);
and U15644 (N_15644,N_12628,N_14342);
nor U15645 (N_15645,N_12411,N_13159);
or U15646 (N_15646,N_12993,N_12939);
xor U15647 (N_15647,N_14769,N_14546);
xor U15648 (N_15648,N_12961,N_14499);
or U15649 (N_15649,N_14974,N_13721);
nor U15650 (N_15650,N_13674,N_13308);
nor U15651 (N_15651,N_12592,N_13607);
and U15652 (N_15652,N_14363,N_13856);
xor U15653 (N_15653,N_13828,N_12534);
nor U15654 (N_15654,N_13077,N_12886);
nand U15655 (N_15655,N_12978,N_12257);
nor U15656 (N_15656,N_14767,N_12274);
nor U15657 (N_15657,N_14843,N_13953);
and U15658 (N_15658,N_14367,N_14489);
nor U15659 (N_15659,N_14548,N_13435);
xnor U15660 (N_15660,N_12343,N_13172);
and U15661 (N_15661,N_14052,N_14019);
or U15662 (N_15662,N_13736,N_14189);
nor U15663 (N_15663,N_12997,N_13707);
xor U15664 (N_15664,N_13149,N_13619);
xor U15665 (N_15665,N_12988,N_14768);
and U15666 (N_15666,N_13631,N_12566);
nand U15667 (N_15667,N_14165,N_14601);
nor U15668 (N_15668,N_13284,N_14697);
xnor U15669 (N_15669,N_14511,N_13076);
xor U15670 (N_15670,N_14306,N_14354);
xor U15671 (N_15671,N_12334,N_14510);
nor U15672 (N_15672,N_14673,N_13624);
or U15673 (N_15673,N_13283,N_14033);
and U15674 (N_15674,N_12068,N_14276);
nor U15675 (N_15675,N_14957,N_14199);
nand U15676 (N_15676,N_13908,N_12517);
xor U15677 (N_15677,N_13204,N_13988);
or U15678 (N_15678,N_13092,N_14450);
xnor U15679 (N_15679,N_14255,N_12907);
nand U15680 (N_15680,N_12656,N_14710);
nand U15681 (N_15681,N_14441,N_13755);
and U15682 (N_15682,N_14637,N_12707);
or U15683 (N_15683,N_13533,N_12313);
nand U15684 (N_15684,N_12330,N_14655);
nor U15685 (N_15685,N_14050,N_13326);
and U15686 (N_15686,N_13045,N_13740);
nand U15687 (N_15687,N_12436,N_14858);
nor U15688 (N_15688,N_13184,N_14613);
and U15689 (N_15689,N_14521,N_12778);
xnor U15690 (N_15690,N_13635,N_13683);
and U15691 (N_15691,N_12395,N_13477);
and U15692 (N_15692,N_13649,N_12473);
and U15693 (N_15693,N_14309,N_12817);
or U15694 (N_15694,N_13295,N_13390);
xnor U15695 (N_15695,N_13237,N_12982);
nor U15696 (N_15696,N_12510,N_13910);
or U15697 (N_15697,N_13642,N_12555);
xnor U15698 (N_15698,N_12403,N_12440);
nand U15699 (N_15699,N_13121,N_12472);
xor U15700 (N_15700,N_12405,N_14656);
nor U15701 (N_15701,N_12052,N_14170);
and U15702 (N_15702,N_12558,N_13815);
and U15703 (N_15703,N_12925,N_13833);
nor U15704 (N_15704,N_12625,N_13494);
nor U15705 (N_15705,N_14960,N_12450);
xor U15706 (N_15706,N_14167,N_13255);
nor U15707 (N_15707,N_13531,N_14706);
xnor U15708 (N_15708,N_14323,N_13311);
nand U15709 (N_15709,N_12648,N_13936);
xnor U15710 (N_15710,N_12155,N_14616);
xnor U15711 (N_15711,N_13008,N_13780);
nand U15712 (N_15712,N_14446,N_12584);
xor U15713 (N_15713,N_13639,N_14256);
nor U15714 (N_15714,N_12280,N_13408);
and U15715 (N_15715,N_14875,N_12048);
nor U15716 (N_15716,N_12022,N_13313);
nor U15717 (N_15717,N_13234,N_12211);
nand U15718 (N_15718,N_14429,N_13193);
nand U15719 (N_15719,N_12289,N_13082);
or U15720 (N_15720,N_14920,N_13595);
xor U15721 (N_15721,N_14745,N_12109);
or U15722 (N_15722,N_12291,N_14795);
xnor U15723 (N_15723,N_12727,N_14887);
nand U15724 (N_15724,N_13002,N_14474);
nand U15725 (N_15725,N_14289,N_13835);
or U15726 (N_15726,N_13461,N_14053);
nand U15727 (N_15727,N_14844,N_13061);
or U15728 (N_15728,N_13547,N_13520);
or U15729 (N_15729,N_14296,N_12180);
nor U15730 (N_15730,N_13090,N_14177);
xnor U15731 (N_15731,N_13576,N_14724);
nand U15732 (N_15732,N_13521,N_14290);
and U15733 (N_15733,N_14104,N_13000);
nor U15734 (N_15734,N_13279,N_12341);
nor U15735 (N_15735,N_12083,N_14403);
nand U15736 (N_15736,N_12842,N_14664);
xor U15737 (N_15737,N_12935,N_13643);
and U15738 (N_15738,N_13778,N_14084);
nand U15739 (N_15739,N_14593,N_14530);
or U15740 (N_15740,N_13767,N_14451);
xnor U15741 (N_15741,N_12081,N_12799);
nor U15742 (N_15742,N_14799,N_12797);
nor U15743 (N_15743,N_12667,N_13544);
or U15744 (N_15744,N_13171,N_12446);
nor U15745 (N_15745,N_12633,N_13206);
nor U15746 (N_15746,N_12117,N_14734);
or U15747 (N_15747,N_13842,N_13559);
and U15748 (N_15748,N_14527,N_14149);
nand U15749 (N_15749,N_13919,N_14630);
or U15750 (N_15750,N_14757,N_13056);
nor U15751 (N_15751,N_13892,N_14874);
xnor U15752 (N_15752,N_14709,N_13219);
or U15753 (N_15753,N_14037,N_14925);
and U15754 (N_15754,N_14369,N_12659);
or U15755 (N_15755,N_13427,N_13483);
and U15756 (N_15756,N_13806,N_14145);
and U15757 (N_15757,N_13329,N_14158);
nand U15758 (N_15758,N_12789,N_13388);
xnor U15759 (N_15759,N_14890,N_13601);
xnor U15760 (N_15760,N_12469,N_13195);
xnor U15761 (N_15761,N_12597,N_14136);
nand U15762 (N_15762,N_12602,N_13696);
xor U15763 (N_15763,N_14366,N_13810);
xnor U15764 (N_15764,N_14109,N_12904);
xor U15765 (N_15765,N_14307,N_13580);
and U15766 (N_15766,N_13514,N_12197);
and U15767 (N_15767,N_14924,N_13528);
xor U15768 (N_15768,N_14047,N_14013);
xnor U15769 (N_15769,N_12243,N_12825);
nand U15770 (N_15770,N_14392,N_14827);
or U15771 (N_15771,N_12685,N_14397);
nor U15772 (N_15772,N_12172,N_12387);
nor U15773 (N_15773,N_14182,N_12470);
or U15774 (N_15774,N_13080,N_14028);
and U15775 (N_15775,N_14851,N_12743);
nand U15776 (N_15776,N_13670,N_14099);
xor U15777 (N_15777,N_13377,N_14934);
xor U15778 (N_15778,N_14356,N_14325);
nand U15779 (N_15779,N_14515,N_13702);
nor U15780 (N_15780,N_14571,N_14676);
and U15781 (N_15781,N_12674,N_12110);
and U15782 (N_15782,N_14536,N_12807);
nor U15783 (N_15783,N_12576,N_14140);
and U15784 (N_15784,N_14857,N_12230);
nand U15785 (N_15785,N_12969,N_14452);
nor U15786 (N_15786,N_14069,N_14542);
or U15787 (N_15787,N_13421,N_14095);
or U15788 (N_15788,N_12831,N_14761);
or U15789 (N_15789,N_13030,N_12800);
or U15790 (N_15790,N_13554,N_14263);
or U15791 (N_15791,N_14074,N_12222);
nand U15792 (N_15792,N_13369,N_13616);
or U15793 (N_15793,N_13140,N_13058);
and U15794 (N_15794,N_14347,N_14797);
nor U15795 (N_15795,N_14869,N_13734);
and U15796 (N_15796,N_14523,N_12185);
and U15797 (N_15797,N_14926,N_14498);
and U15798 (N_15798,N_13319,N_12367);
xnor U15799 (N_15799,N_14437,N_12070);
and U15800 (N_15800,N_12504,N_13620);
nor U15801 (N_15801,N_14981,N_13558);
and U15802 (N_15802,N_12306,N_14989);
nand U15803 (N_15803,N_12461,N_14868);
and U15804 (N_15804,N_12351,N_12678);
nand U15805 (N_15805,N_12249,N_14651);
xor U15806 (N_15806,N_14950,N_13706);
xnor U15807 (N_15807,N_14191,N_14705);
and U15808 (N_15808,N_13419,N_12478);
nand U15809 (N_15809,N_12368,N_13564);
nor U15810 (N_15810,N_13916,N_14825);
or U15811 (N_15811,N_13723,N_13539);
and U15812 (N_15812,N_14631,N_13963);
nand U15813 (N_15813,N_12841,N_13826);
nor U15814 (N_15814,N_14205,N_12753);
nand U15815 (N_15815,N_13548,N_14817);
or U15816 (N_15816,N_14893,N_12384);
nand U15817 (N_15817,N_13713,N_13224);
nand U15818 (N_15818,N_13272,N_13758);
nand U15819 (N_15819,N_13004,N_12323);
or U15820 (N_15820,N_12662,N_12009);
and U15821 (N_15821,N_14819,N_13821);
nand U15822 (N_15822,N_13361,N_14886);
and U15823 (N_15823,N_12554,N_14759);
nor U15824 (N_15824,N_13330,N_13104);
xor U15825 (N_15825,N_13550,N_14045);
nand U15826 (N_15826,N_14719,N_12427);
nor U15827 (N_15827,N_14147,N_14481);
nor U15828 (N_15828,N_12594,N_13930);
nand U15829 (N_15829,N_12296,N_14900);
or U15830 (N_15830,N_13741,N_14678);
nand U15831 (N_15831,N_12898,N_12587);
and U15832 (N_15832,N_12118,N_14089);
nand U15833 (N_15833,N_14487,N_13965);
nor U15834 (N_15834,N_12731,N_12901);
nor U15835 (N_15835,N_13588,N_13160);
nand U15836 (N_15836,N_14570,N_13023);
nor U15837 (N_15837,N_12316,N_13315);
xor U15838 (N_15838,N_14079,N_12188);
or U15839 (N_15839,N_14410,N_12430);
or U15840 (N_15840,N_12443,N_12879);
xor U15841 (N_15841,N_12339,N_13934);
nand U15842 (N_15842,N_14330,N_14670);
xor U15843 (N_15843,N_13414,N_13438);
or U15844 (N_15844,N_13605,N_14558);
nand U15845 (N_15845,N_12896,N_12161);
nand U15846 (N_15846,N_13103,N_13203);
or U15847 (N_15847,N_13264,N_12154);
xor U15848 (N_15848,N_14378,N_12294);
xnor U15849 (N_15849,N_14982,N_12862);
nand U15850 (N_15850,N_12564,N_12481);
xnor U15851 (N_15851,N_13760,N_13033);
nor U15852 (N_15852,N_12851,N_13485);
or U15853 (N_15853,N_14419,N_14608);
nor U15854 (N_15854,N_14077,N_12092);
and U15855 (N_15855,N_12144,N_14778);
xnor U15856 (N_15856,N_13708,N_12964);
and U15857 (N_15857,N_12499,N_14181);
or U15858 (N_15858,N_12990,N_13259);
xor U15859 (N_15859,N_13999,N_13546);
xnor U15860 (N_15860,N_14865,N_14994);
xor U15861 (N_15861,N_12856,N_12100);
and U15862 (N_15862,N_14122,N_13299);
and U15863 (N_15863,N_13774,N_13111);
and U15864 (N_15864,N_14881,N_13241);
xor U15865 (N_15865,N_12889,N_13881);
xnor U15866 (N_15866,N_14302,N_14598);
and U15867 (N_15867,N_13562,N_13244);
and U15868 (N_15868,N_14909,N_12420);
or U15869 (N_15869,N_14703,N_12137);
and U15870 (N_15870,N_12634,N_12784);
nor U15871 (N_15871,N_14023,N_13453);
nand U15872 (N_15872,N_14409,N_14098);
nor U15873 (N_15873,N_14945,N_14303);
or U15874 (N_15874,N_13762,N_13682);
or U15875 (N_15875,N_12967,N_14518);
or U15876 (N_15876,N_14217,N_13266);
xnor U15877 (N_15877,N_13519,N_14666);
and U15878 (N_15878,N_14824,N_12354);
nand U15879 (N_15879,N_14674,N_13535);
or U15880 (N_15880,N_12040,N_14116);
xnor U15881 (N_15881,N_13368,N_12187);
nand U15882 (N_15882,N_12378,N_13278);
and U15883 (N_15883,N_13926,N_13100);
or U15884 (N_15884,N_12247,N_14101);
nand U15885 (N_15885,N_12087,N_12383);
nor U15886 (N_15886,N_14617,N_14162);
and U15887 (N_15887,N_14279,N_13637);
nor U15888 (N_15888,N_14564,N_12492);
nand U15889 (N_15889,N_14334,N_13712);
nor U15890 (N_15890,N_13814,N_13794);
nand U15891 (N_15891,N_12520,N_13851);
nor U15892 (N_15892,N_13996,N_14353);
or U15893 (N_15893,N_14245,N_12276);
and U15894 (N_15894,N_12526,N_12295);
or U15895 (N_15895,N_12192,N_12687);
nor U15896 (N_15896,N_14771,N_13906);
nor U15897 (N_15897,N_13059,N_13731);
xor U15898 (N_15898,N_14114,N_13606);
and U15899 (N_15899,N_12820,N_14374);
or U15900 (N_15900,N_13393,N_13426);
and U15901 (N_15901,N_12404,N_13375);
or U15902 (N_15902,N_14965,N_12722);
and U15903 (N_15903,N_14395,N_12049);
nor U15904 (N_15904,N_12810,N_12599);
xor U15905 (N_15905,N_14190,N_14240);
nand U15906 (N_15906,N_13864,N_13402);
or U15907 (N_15907,N_12010,N_12546);
nand U15908 (N_15908,N_12705,N_12151);
and U15909 (N_15909,N_12733,N_13022);
nor U15910 (N_15910,N_14610,N_12665);
nand U15911 (N_15911,N_12026,N_13257);
nor U15912 (N_15912,N_12614,N_13571);
and U15913 (N_15913,N_14955,N_13818);
xor U15914 (N_15914,N_12445,N_14107);
nor U15915 (N_15915,N_12787,N_14432);
and U15916 (N_15916,N_12227,N_13430);
or U15917 (N_15917,N_12996,N_14174);
nor U15918 (N_15918,N_14816,N_14669);
or U15919 (N_15919,N_13454,N_14266);
nand U15920 (N_15920,N_14017,N_12106);
and U15921 (N_15921,N_13900,N_12543);
or U15922 (N_15922,N_13085,N_12750);
xnor U15923 (N_15923,N_14076,N_13091);
nor U15924 (N_15924,N_13424,N_13950);
nand U15925 (N_15925,N_14072,N_13024);
nand U15926 (N_15926,N_13396,N_12246);
xor U15927 (N_15927,N_13549,N_13262);
xor U15928 (N_15928,N_14921,N_12812);
and U15929 (N_15929,N_12124,N_14852);
and U15930 (N_15930,N_12803,N_14618);
nand U15931 (N_15931,N_14836,N_14275);
nor U15932 (N_15932,N_12308,N_14566);
xor U15933 (N_15933,N_14322,N_12798);
and U15934 (N_15934,N_14787,N_14970);
and U15935 (N_15935,N_12790,N_14194);
xnor U15936 (N_15936,N_13823,N_14219);
or U15937 (N_15937,N_12113,N_13035);
nor U15938 (N_15938,N_14093,N_12288);
or U15939 (N_15939,N_13556,N_12382);
or U15940 (N_15940,N_14786,N_13423);
nand U15941 (N_15941,N_14645,N_13939);
xnor U15942 (N_15942,N_13664,N_12553);
nand U15943 (N_15943,N_13757,N_13050);
and U15944 (N_15944,N_12263,N_13015);
and U15945 (N_15945,N_14059,N_12773);
nor U15946 (N_15946,N_12275,N_13971);
nor U15947 (N_15947,N_14000,N_13196);
nor U15948 (N_15948,N_13636,N_12372);
and U15949 (N_15949,N_13109,N_13107);
nand U15950 (N_15950,N_12181,N_14434);
or U15951 (N_15951,N_12258,N_13346);
or U15952 (N_15952,N_12548,N_12407);
nand U15953 (N_15953,N_13795,N_14903);
nor U15954 (N_15954,N_12766,N_14983);
and U15955 (N_15955,N_12713,N_14594);
nor U15956 (N_15956,N_12159,N_12217);
and U15957 (N_15957,N_12018,N_14735);
xnor U15958 (N_15958,N_14427,N_14485);
or U15959 (N_15959,N_14692,N_12883);
xor U15960 (N_15960,N_13899,N_14003);
nand U15961 (N_15961,N_13829,N_12836);
and U15962 (N_15962,N_12590,N_12490);
and U15963 (N_15963,N_13689,N_14959);
nand U15964 (N_15964,N_12525,N_12704);
or U15965 (N_15965,N_12972,N_14944);
and U15966 (N_15966,N_13628,N_14773);
and U15967 (N_15967,N_14764,N_13599);
xor U15968 (N_15968,N_12942,N_12837);
and U15969 (N_15969,N_12233,N_14483);
nand U15970 (N_15970,N_12806,N_13188);
or U15971 (N_15971,N_14624,N_13381);
and U15972 (N_15972,N_13732,N_12401);
and U15973 (N_15973,N_13202,N_13174);
nand U15974 (N_15974,N_14866,N_13360);
nor U15975 (N_15975,N_14600,N_12940);
and U15976 (N_15976,N_12582,N_12598);
nand U15977 (N_15977,N_14939,N_14765);
nand U15978 (N_15978,N_13066,N_13837);
or U15979 (N_15979,N_14015,N_14261);
nand U15980 (N_15980,N_14466,N_14377);
nand U15981 (N_15981,N_14775,N_14150);
xor U15982 (N_15982,N_13339,N_12956);
nor U15983 (N_15983,N_14416,N_14063);
nor U15984 (N_15984,N_13415,N_14698);
and U15985 (N_15985,N_12344,N_12795);
nand U15986 (N_15986,N_13788,N_14772);
and U15987 (N_15987,N_14722,N_14287);
and U15988 (N_15988,N_14239,N_13387);
and U15989 (N_15989,N_12452,N_13942);
and U15990 (N_15990,N_12693,N_13791);
and U15991 (N_15991,N_12593,N_14313);
and U15992 (N_15992,N_14227,N_12393);
nor U15993 (N_15993,N_12893,N_14514);
nand U15994 (N_15994,N_13444,N_13611);
nand U15995 (N_15995,N_14435,N_12311);
nand U15996 (N_15996,N_14386,N_14508);
and U15997 (N_15997,N_12178,N_13878);
nor U15998 (N_15998,N_14714,N_13116);
nor U15999 (N_15999,N_12902,N_14872);
nor U16000 (N_16000,N_14683,N_12400);
xnor U16001 (N_16001,N_13512,N_12320);
or U16002 (N_16002,N_12695,N_14894);
xor U16003 (N_16003,N_14234,N_13933);
and U16004 (N_16004,N_12136,N_12098);
nor U16005 (N_16005,N_14522,N_14270);
nand U16006 (N_16006,N_12632,N_12186);
nor U16007 (N_16007,N_12849,N_13909);
nor U16008 (N_16008,N_13366,N_12960);
xor U16009 (N_16009,N_13037,N_12877);
nand U16010 (N_16010,N_13250,N_14788);
xnor U16011 (N_16011,N_14873,N_12629);
and U16012 (N_16012,N_12020,N_13923);
or U16013 (N_16013,N_13407,N_13170);
nor U16014 (N_16014,N_14025,N_14973);
and U16015 (N_16015,N_12547,N_12871);
or U16016 (N_16016,N_13505,N_12992);
or U16017 (N_16017,N_14991,N_13070);
xnor U16018 (N_16018,N_14760,N_13717);
and U16019 (N_16019,N_12631,N_12663);
xor U16020 (N_16020,N_13629,N_14953);
nor U16021 (N_16021,N_13873,N_13956);
or U16022 (N_16022,N_13751,N_13834);
nor U16023 (N_16023,N_12386,N_12922);
and U16024 (N_16024,N_12646,N_12691);
nand U16025 (N_16025,N_12977,N_14642);
and U16026 (N_16026,N_14385,N_14336);
xnor U16027 (N_16027,N_12608,N_12412);
nor U16028 (N_16028,N_13491,N_13775);
nor U16029 (N_16029,N_12968,N_12031);
and U16030 (N_16030,N_13245,N_12793);
and U16031 (N_16031,N_12067,N_12805);
and U16032 (N_16032,N_14115,N_13729);
xnor U16033 (N_16033,N_13917,N_12060);
and U16034 (N_16034,N_14186,N_12116);
nor U16035 (N_16035,N_12769,N_12235);
or U16036 (N_16036,N_14862,N_12262);
or U16037 (N_16037,N_14784,N_13672);
xor U16038 (N_16038,N_14933,N_13982);
or U16039 (N_16039,N_14151,N_12708);
and U16040 (N_16040,N_14988,N_13213);
nand U16041 (N_16041,N_14643,N_14128);
nor U16042 (N_16042,N_12189,N_13049);
xor U16043 (N_16043,N_13627,N_12839);
and U16044 (N_16044,N_14856,N_14806);
and U16045 (N_16045,N_13989,N_12611);
nor U16046 (N_16046,N_14854,N_13122);
or U16047 (N_16047,N_13577,N_12890);
nor U16048 (N_16048,N_13876,N_14904);
nor U16049 (N_16049,N_14638,N_13317);
nor U16050 (N_16050,N_12094,N_13298);
and U16051 (N_16051,N_12062,N_14231);
xor U16052 (N_16052,N_13293,N_13797);
or U16053 (N_16053,N_14512,N_12676);
xor U16054 (N_16054,N_12834,N_12409);
and U16055 (N_16055,N_13880,N_12281);
and U16056 (N_16056,N_13684,N_14282);
xor U16057 (N_16057,N_14111,N_13510);
nor U16058 (N_16058,N_14477,N_12684);
nand U16059 (N_16059,N_14936,N_14821);
or U16060 (N_16060,N_12919,N_12867);
nand U16061 (N_16061,N_12741,N_13617);
and U16062 (N_16062,N_14357,N_12710);
xnor U16063 (N_16063,N_12947,N_14321);
or U16064 (N_16064,N_14562,N_12770);
and U16065 (N_16065,N_13523,N_12357);
nor U16066 (N_16066,N_13289,N_14905);
nor U16067 (N_16067,N_14393,N_12725);
nand U16068 (N_16068,N_13888,N_13820);
and U16069 (N_16069,N_13801,N_12838);
xnor U16070 (N_16070,N_14155,N_13420);
nor U16071 (N_16071,N_13977,N_13907);
and U16072 (N_16072,N_12366,N_14591);
or U16073 (N_16073,N_13389,N_13968);
or U16074 (N_16074,N_13233,N_13083);
nor U16075 (N_16075,N_13784,N_14100);
nor U16076 (N_16076,N_12737,N_12682);
nand U16077 (N_16077,N_13594,N_12102);
nor U16078 (N_16078,N_13583,N_13422);
or U16079 (N_16079,N_14259,N_14265);
or U16080 (N_16080,N_14317,N_13306);
or U16081 (N_16081,N_13118,N_12331);
or U16082 (N_16082,N_12533,N_12428);
and U16083 (N_16083,N_13678,N_14399);
nor U16084 (N_16084,N_14748,N_14031);
xnor U16085 (N_16085,N_14634,N_12761);
nor U16086 (N_16086,N_14472,N_13481);
or U16087 (N_16087,N_14596,N_12868);
and U16088 (N_16088,N_12618,N_14173);
and U16089 (N_16089,N_12523,N_14269);
and U16090 (N_16090,N_14801,N_12914);
nor U16091 (N_16091,N_14790,N_13142);
nor U16092 (N_16092,N_12861,N_14209);
nor U16093 (N_16093,N_12304,N_13114);
xnor U16094 (N_16094,N_12557,N_14073);
and U16095 (N_16095,N_14898,N_12620);
or U16096 (N_16096,N_13437,N_12855);
or U16097 (N_16097,N_14971,N_13197);
xnor U16098 (N_16098,N_13012,N_14253);
and U16099 (N_16099,N_13840,N_14041);
nor U16100 (N_16100,N_13071,N_12001);
and U16101 (N_16101,N_14396,N_12859);
nand U16102 (N_16102,N_14326,N_12195);
and U16103 (N_16103,N_13663,N_12326);
or U16104 (N_16104,N_14471,N_13287);
and U16105 (N_16105,N_13325,N_14980);
xor U16106 (N_16106,N_14348,N_12783);
nor U16107 (N_16107,N_13046,N_12918);
and U16108 (N_16108,N_13484,N_12822);
or U16109 (N_16109,N_14210,N_14623);
nor U16110 (N_16110,N_12637,N_13647);
nand U16111 (N_16111,N_14129,N_13010);
nor U16112 (N_16112,N_14876,N_13433);
nand U16113 (N_16113,N_13464,N_13600);
xor U16114 (N_16114,N_12039,N_14581);
nand U16115 (N_16115,N_14826,N_12575);
nor U16116 (N_16116,N_13364,N_12061);
nand U16117 (N_16117,N_13416,N_12458);
nor U16118 (N_16118,N_13964,N_13189);
nor U16119 (N_16119,N_13517,N_12835);
xor U16120 (N_16120,N_12735,N_13296);
xnor U16121 (N_16121,N_14525,N_14154);
and U16122 (N_16122,N_13566,N_12284);
xnor U16123 (N_16123,N_14262,N_12570);
or U16124 (N_16124,N_13802,N_12132);
nor U16125 (N_16125,N_13075,N_12273);
or U16126 (N_16126,N_12037,N_12815);
and U16127 (N_16127,N_12643,N_14650);
nor U16128 (N_16128,N_13052,N_12572);
nor U16129 (N_16129,N_12277,N_12256);
nor U16130 (N_16130,N_13975,N_14604);
nand U16131 (N_16131,N_13309,N_14102);
and U16132 (N_16132,N_12508,N_12459);
nor U16133 (N_16133,N_13026,N_13065);
nor U16134 (N_16134,N_14517,N_12765);
nor U16135 (N_16135,N_12467,N_12058);
xor U16136 (N_16136,N_14609,N_14504);
xnor U16137 (N_16137,N_12198,N_13782);
xnor U16138 (N_16138,N_13199,N_12005);
nor U16139 (N_16139,N_14157,N_13280);
and U16140 (N_16140,N_14088,N_14204);
and U16141 (N_16141,N_13073,N_13473);
xor U16142 (N_16142,N_12085,N_13501);
nor U16143 (N_16143,N_13089,N_14284);
and U16144 (N_16144,N_12259,N_12134);
nand U16145 (N_16145,N_14064,N_12857);
or U16146 (N_16146,N_14143,N_14338);
or U16147 (N_16147,N_12941,N_12374);
or U16148 (N_16148,N_12808,N_14840);
or U16149 (N_16149,N_12771,N_13042);
or U16150 (N_16150,N_12358,N_13323);
nand U16151 (N_16151,N_13067,N_12848);
and U16152 (N_16152,N_12426,N_14327);
or U16153 (N_16153,N_12931,N_12551);
nor U16154 (N_16154,N_12882,N_13756);
or U16155 (N_16155,N_13268,N_12562);
or U16156 (N_16156,N_12353,N_13590);
nor U16157 (N_16157,N_13932,N_13904);
or U16158 (N_16158,N_14447,N_13151);
nand U16159 (N_16159,N_12723,N_14008);
xor U16160 (N_16160,N_13536,N_13632);
nand U16161 (N_16161,N_14166,N_14942);
and U16162 (N_16162,N_12772,N_13447);
nand U16163 (N_16163,N_13263,N_12591);
or U16164 (N_16164,N_14383,N_13318);
nor U16165 (N_16165,N_13827,N_12265);
nand U16166 (N_16166,N_14931,N_12719);
nand U16167 (N_16167,N_12752,N_12305);
nor U16168 (N_16168,N_12419,N_14057);
and U16169 (N_16169,N_12645,N_12757);
xor U16170 (N_16170,N_14807,N_12457);
or U16171 (N_16171,N_12156,N_12740);
and U16172 (N_16172,N_13614,N_13384);
nor U16173 (N_16173,N_14034,N_13153);
and U16174 (N_16174,N_13209,N_12671);
or U16175 (N_16175,N_13055,N_14731);
or U16176 (N_16176,N_12165,N_14200);
xor U16177 (N_16177,N_14730,N_14465);
nand U16178 (N_16178,N_14075,N_14055);
xnor U16179 (N_16179,N_12232,N_12973);
nand U16180 (N_16180,N_13482,N_13743);
xor U16181 (N_16181,N_12649,N_13157);
or U16182 (N_16182,N_13084,N_12012);
xor U16183 (N_16183,N_12923,N_12153);
and U16184 (N_16184,N_13952,N_12762);
xor U16185 (N_16185,N_14539,N_12173);
and U16186 (N_16186,N_12164,N_14470);
xnor U16187 (N_16187,N_13469,N_12075);
or U16188 (N_16188,N_12974,N_12827);
nor U16189 (N_16189,N_14831,N_14696);
nor U16190 (N_16190,N_14389,N_13724);
xor U16191 (N_16191,N_12721,N_13261);
xor U16192 (N_16192,N_13905,N_12529);
or U16193 (N_16193,N_12776,N_13677);
and U16194 (N_16194,N_12310,N_12874);
nand U16195 (N_16195,N_14578,N_14592);
xnor U16196 (N_16196,N_13967,N_14770);
xnor U16197 (N_16197,N_14280,N_12677);
or U16198 (N_16198,N_14849,N_14984);
and U16199 (N_16199,N_14641,N_12878);
nand U16200 (N_16200,N_13350,N_13894);
xnor U16201 (N_16201,N_14503,N_14992);
xor U16202 (N_16202,N_12571,N_14742);
nor U16203 (N_16203,N_14901,N_14467);
nand U16204 (N_16204,N_14249,N_14783);
nand U16205 (N_16205,N_12796,N_13970);
and U16206 (N_16206,N_14743,N_14196);
or U16207 (N_16207,N_14418,N_14776);
xor U16208 (N_16208,N_12359,N_14689);
nand U16209 (N_16209,N_12945,N_13495);
and U16210 (N_16210,N_12050,N_14711);
xor U16211 (N_16211,N_13690,N_14221);
xnor U16212 (N_16212,N_14584,N_13094);
or U16213 (N_16213,N_13812,N_14529);
and U16214 (N_16214,N_13198,N_12934);
nor U16215 (N_16215,N_13286,N_12514);
xnor U16216 (N_16216,N_13480,N_12991);
nand U16217 (N_16217,N_12309,N_12763);
and U16218 (N_16218,N_14257,N_13434);
nor U16219 (N_16219,N_14153,N_12912);
or U16220 (N_16220,N_12609,N_13855);
nor U16221 (N_16221,N_12108,N_13229);
nor U16222 (N_16222,N_12894,N_12028);
nand U16223 (N_16223,N_12962,N_12379);
and U16224 (N_16224,N_13112,N_12679);
xor U16225 (N_16225,N_13675,N_12782);
and U16226 (N_16226,N_14085,N_13803);
xor U16227 (N_16227,N_12995,N_13418);
nand U16228 (N_16228,N_14545,N_14535);
xnor U16229 (N_16229,N_12953,N_12489);
or U16230 (N_16230,N_13653,N_12468);
xnor U16231 (N_16231,N_13312,N_14835);
or U16232 (N_16232,N_14020,N_13946);
nor U16233 (N_16233,N_13486,N_12200);
or U16234 (N_16234,N_12605,N_13442);
nor U16235 (N_16235,N_14180,N_14032);
nor U16236 (N_16236,N_12715,N_14533);
or U16237 (N_16237,N_14659,N_14469);
xnor U16238 (N_16238,N_12661,N_13852);
nand U16239 (N_16239,N_12030,N_14135);
or U16240 (N_16240,N_13866,N_13800);
nand U16241 (N_16241,N_12370,N_14112);
nor U16242 (N_16242,N_12983,N_14679);
or U16243 (N_16243,N_12844,N_12675);
nor U16244 (N_16244,N_13525,N_14628);
nor U16245 (N_16245,N_12921,N_13138);
xnor U16246 (N_16246,N_12191,N_13596);
nor U16247 (N_16247,N_13161,N_14272);
nand U16248 (N_16248,N_12999,N_12004);
nor U16249 (N_16249,N_12338,N_13215);
nor U16250 (N_16250,N_14492,N_12336);
or U16251 (N_16251,N_12431,N_14958);
xor U16252 (N_16252,N_12107,N_14375);
or U16253 (N_16253,N_14597,N_12365);
and U16254 (N_16254,N_14580,N_14952);
nand U16255 (N_16255,N_14448,N_13848);
nor U16256 (N_16256,N_13998,N_13448);
nand U16257 (N_16257,N_14998,N_12425);
nand U16258 (N_16258,N_14292,N_14108);
or U16259 (N_16259,N_12924,N_14741);
nand U16260 (N_16260,N_13270,N_12101);
nor U16261 (N_16261,N_14291,N_12105);
nor U16262 (N_16262,N_13929,N_14640);
and U16263 (N_16263,N_13445,N_13966);
xor U16264 (N_16264,N_12801,N_14690);
and U16265 (N_16265,N_12986,N_13832);
nand U16266 (N_16266,N_14497,N_14382);
and U16267 (N_16267,N_13728,N_14910);
and U16268 (N_16268,N_13405,N_12824);
nand U16269 (N_16269,N_12681,N_14923);
xor U16270 (N_16270,N_12699,N_13285);
xnor U16271 (N_16271,N_13288,N_14035);
and U16272 (N_16272,N_14203,N_14081);
or U16273 (N_16273,N_13621,N_12293);
nand U16274 (N_16274,N_13666,N_13896);
or U16275 (N_16275,N_12008,N_13526);
and U16276 (N_16276,N_14574,N_14553);
xor U16277 (N_16277,N_12054,N_12203);
xor U16278 (N_16278,N_13938,N_13246);
xnor U16279 (N_16279,N_12928,N_12325);
nor U16280 (N_16280,N_12756,N_14486);
nor U16281 (N_16281,N_12003,N_13152);
nand U16282 (N_16282,N_14051,N_13374);
nand U16283 (N_16283,N_13102,N_13178);
or U16284 (N_16284,N_12696,N_13799);
xor U16285 (N_16285,N_12025,N_14208);
nand U16286 (N_16286,N_12586,N_12913);
xnor U16287 (N_16287,N_12948,N_13179);
nor U16288 (N_16288,N_13857,N_13236);
nor U16289 (N_16289,N_14896,N_12255);
nand U16290 (N_16290,N_12024,N_14513);
or U16291 (N_16291,N_12640,N_12887);
nor U16292 (N_16292,N_12612,N_14405);
nand U16293 (N_16293,N_14990,N_14845);
nand U16294 (N_16294,N_14712,N_12418);
nand U16295 (N_16295,N_13737,N_14699);
xor U16296 (N_16296,N_13709,N_13068);
and U16297 (N_16297,N_14644,N_14113);
and U16298 (N_16298,N_12146,N_14056);
nor U16299 (N_16299,N_14708,N_13031);
xnor U16300 (N_16300,N_13316,N_14884);
or U16301 (N_16301,N_12290,N_14967);
or U16302 (N_16302,N_13176,N_14060);
and U16303 (N_16303,N_12460,N_12876);
nor U16304 (N_16304,N_14680,N_14914);
nor U16305 (N_16305,N_12285,N_12437);
xnor U16306 (N_16306,N_14882,N_13016);
or U16307 (N_16307,N_13657,N_13725);
nand U16308 (N_16308,N_12641,N_13372);
and U16309 (N_16309,N_12615,N_12149);
nand U16310 (N_16310,N_12513,N_12938);
and U16311 (N_16311,N_12317,N_12023);
or U16312 (N_16312,N_13958,N_14413);
or U16313 (N_16313,N_13841,N_14568);
nand U16314 (N_16314,N_13575,N_12552);
and U16315 (N_16315,N_13859,N_12138);
xnor U16316 (N_16316,N_14636,N_12536);
and U16317 (N_16317,N_14620,N_12423);
nor U16318 (N_16318,N_14614,N_13646);
xnor U16319 (N_16319,N_12596,N_12686);
xor U16320 (N_16320,N_14733,N_12128);
and U16321 (N_16321,N_14516,N_14148);
xor U16322 (N_16322,N_14414,N_14729);
and U16323 (N_16323,N_13348,N_14629);
and U16324 (N_16324,N_12946,N_13997);
and U16325 (N_16325,N_14339,N_13320);
or U16326 (N_16326,N_14212,N_14646);
xor U16327 (N_16327,N_12718,N_14948);
nor U16328 (N_16328,N_12055,N_13194);
xor U16329 (N_16329,N_13054,N_14755);
xnor U16330 (N_16330,N_13839,N_14501);
and U16331 (N_16331,N_14889,N_13412);
nor U16332 (N_16332,N_12509,N_13376);
nand U16333 (N_16333,N_13793,N_13991);
nor U16334 (N_16334,N_13612,N_13498);
nor U16335 (N_16335,N_13608,N_12121);
or U16336 (N_16336,N_13650,N_14110);
nor U16337 (N_16337,N_12549,N_13622);
xnor U16338 (N_16338,N_14943,N_13044);
nor U16339 (N_16339,N_13041,N_12527);
nor U16340 (N_16340,N_14218,N_12141);
xor U16341 (N_16341,N_13297,N_13700);
nor U16342 (N_16342,N_13861,N_14346);
nand U16343 (N_16343,N_14066,N_13141);
nor U16344 (N_16344,N_13813,N_14067);
nand U16345 (N_16345,N_13853,N_13099);
and U16346 (N_16346,N_12362,N_13371);
and U16347 (N_16347,N_13370,N_13750);
nor U16348 (N_16348,N_14254,N_12521);
and U16349 (N_16349,N_12583,N_14294);
nor U16350 (N_16350,N_13819,N_12581);
xor U16351 (N_16351,N_14404,N_13925);
and U16352 (N_16352,N_12158,N_13779);
nand U16353 (N_16353,N_14117,N_13201);
and U16354 (N_16354,N_13240,N_13470);
xor U16355 (N_16355,N_14299,N_13096);
or U16356 (N_16356,N_14502,N_13935);
or U16357 (N_16357,N_14226,N_14453);
nor U16358 (N_16358,N_12500,N_12541);
nand U16359 (N_16359,N_14811,N_14751);
xnor U16360 (N_16360,N_12932,N_13006);
or U16361 (N_16361,N_12303,N_14211);
nand U16362 (N_16362,N_12016,N_12252);
and U16363 (N_16363,N_14919,N_12385);
xor U16364 (N_16364,N_12487,N_12560);
xnor U16365 (N_16365,N_13014,N_12653);
nand U16366 (N_16366,N_12439,N_12464);
and U16367 (N_16367,N_12380,N_12014);
xor U16368 (N_16368,N_14490,N_12909);
or U16369 (N_16369,N_12130,N_14667);
nand U16370 (N_16370,N_12480,N_14297);
or U16371 (N_16371,N_12694,N_13038);
nand U16372 (N_16372,N_14877,N_14126);
or U16373 (N_16373,N_12535,N_12231);
and U16374 (N_16374,N_14048,N_12843);
nor U16375 (N_16375,N_12475,N_13555);
nand U16376 (N_16376,N_12038,N_13869);
and U16377 (N_16377,N_12872,N_12728);
xor U16378 (N_16378,N_14528,N_14376);
xor U16379 (N_16379,N_12506,N_14021);
xnor U16380 (N_16380,N_14880,N_14878);
xor U16381 (N_16381,N_12242,N_14752);
xnor U16382 (N_16382,N_12720,N_13915);
or U16383 (N_16383,N_13018,N_13865);
xnor U16384 (N_16384,N_14124,N_14695);
xor U16385 (N_16385,N_12906,N_13190);
or U16386 (N_16386,N_14314,N_14867);
nor U16387 (N_16387,N_14927,N_13572);
nand U16388 (N_16388,N_12759,N_12496);
nand U16389 (N_16389,N_14718,N_14774);
nor U16390 (N_16390,N_13327,N_13324);
nand U16391 (N_16391,N_13292,N_12954);
or U16392 (N_16392,N_12959,N_14232);
xnor U16393 (N_16393,N_13581,N_12511);
nand U16394 (N_16394,N_13847,N_12892);
nor U16395 (N_16395,N_12573,N_12654);
nor U16396 (N_16396,N_13530,N_14420);
xor U16397 (N_16397,N_12210,N_14454);
and U16398 (N_16398,N_12683,N_12278);
and U16399 (N_16399,N_12950,N_14964);
xor U16400 (N_16400,N_12035,N_14442);
or U16401 (N_16401,N_13098,N_14505);
or U16402 (N_16402,N_14278,N_12429);
nor U16403 (N_16403,N_13685,N_13735);
nand U16404 (N_16404,N_14834,N_13060);
xnor U16405 (N_16405,N_12701,N_14606);
and U16406 (N_16406,N_12435,N_12327);
and U16407 (N_16407,N_14554,N_14359);
xnor U16408 (N_16408,N_13545,N_12970);
or U16409 (N_16409,N_12006,N_13570);
nand U16410 (N_16410,N_14062,N_12223);
xnor U16411 (N_16411,N_12965,N_13359);
or U16412 (N_16412,N_14800,N_12071);
nand U16413 (N_16413,N_14864,N_13079);
or U16414 (N_16414,N_14172,N_14791);
xnor U16415 (N_16415,N_14002,N_13110);
or U16416 (N_16416,N_12606,N_13752);
nand U16417 (N_16417,N_13471,N_13128);
nand U16418 (N_16418,N_14119,N_13960);
or U16419 (N_16419,N_12408,N_12767);
nand U16420 (N_16420,N_14520,N_14248);
nor U16421 (N_16421,N_14537,N_13792);
xor U16422 (N_16422,N_12692,N_12644);
xnor U16423 (N_16423,N_12241,N_13336);
xnor U16424 (N_16424,N_14863,N_14198);
nand U16425 (N_16425,N_13893,N_13557);
or U16426 (N_16426,N_13291,N_13489);
xor U16427 (N_16427,N_14244,N_14488);
xnor U16428 (N_16428,N_13733,N_12352);
or U16429 (N_16429,N_13914,N_13761);
xnor U16430 (N_16430,N_12840,N_12212);
xor U16431 (N_16431,N_14188,N_12090);
or U16432 (N_16432,N_13980,N_12414);
nand U16433 (N_16433,N_13777,N_12588);
nand U16434 (N_16434,N_13478,N_12828);
nand U16435 (N_16435,N_12568,N_14753);
xnor U16436 (N_16436,N_13507,N_13747);
xor U16437 (N_16437,N_12944,N_13673);
or U16438 (N_16438,N_12214,N_12471);
nand U16439 (N_16439,N_14534,N_14809);
and U16440 (N_16440,N_13340,N_13920);
nand U16441 (N_16441,N_14080,N_12832);
xnor U16442 (N_16442,N_14885,N_14796);
nand U16443 (N_16443,N_13822,N_12064);
nand U16444 (N_16444,N_13335,N_14556);
and U16445 (N_16445,N_13158,N_13095);
or U16446 (N_16446,N_12672,N_14185);
nor U16447 (N_16447,N_13954,N_12069);
or U16448 (N_16448,N_14431,N_12627);
and U16449 (N_16449,N_13243,N_12240);
nor U16450 (N_16450,N_12015,N_13362);
nor U16451 (N_16451,N_13001,N_14164);
xnor U16452 (N_16452,N_14094,N_13425);
nand U16453 (N_16453,N_13273,N_14663);
nand U16454 (N_16454,N_12449,N_14001);
nand U16455 (N_16455,N_14315,N_14838);
nand U16456 (N_16456,N_14577,N_13918);
nand U16457 (N_16457,N_14305,N_14691);
and U16458 (N_16458,N_14569,N_13686);
and U16459 (N_16459,N_14300,N_14408);
and U16460 (N_16460,N_12650,N_14802);
nor U16461 (N_16461,N_13945,N_13625);
or U16462 (N_16462,N_13365,N_12802);
nand U16463 (N_16463,N_14436,N_13807);
or U16464 (N_16464,N_14424,N_13877);
or U16465 (N_16465,N_13773,N_12127);
xnor U16466 (N_16466,N_13879,N_13212);
and U16467 (N_16467,N_13497,N_12170);
and U16468 (N_16468,N_14159,N_13228);
nand U16469 (N_16469,N_13771,N_13785);
nand U16470 (N_16470,N_14808,N_12332);
or U16471 (N_16471,N_14230,N_12063);
nand U16472 (N_16472,N_13051,N_13164);
xnor U16473 (N_16473,N_13858,N_12860);
and U16474 (N_16474,N_12702,N_12375);
nand U16475 (N_16475,N_14355,N_14543);
xor U16476 (N_16476,N_13063,N_13511);
nand U16477 (N_16477,N_12779,N_13854);
nand U16478 (N_16478,N_13431,N_14496);
or U16479 (N_16479,N_14633,N_14216);
nand U16480 (N_16480,N_13081,N_13450);
nor U16481 (N_16481,N_13304,N_14559);
and U16482 (N_16482,N_13922,N_14779);
nand U16483 (N_16483,N_14228,N_12760);
nor U16484 (N_16484,N_13235,N_14344);
and U16485 (N_16485,N_12019,N_13845);
nand U16486 (N_16486,N_12162,N_14311);
and U16487 (N_16487,N_12447,N_12381);
nand U16488 (N_16488,N_13446,N_14665);
nand U16489 (N_16489,N_13830,N_13269);
xor U16490 (N_16490,N_13716,N_14049);
and U16491 (N_16491,N_13441,N_12133);
xnor U16492 (N_16492,N_13836,N_12218);
nand U16493 (N_16493,N_12823,N_12342);
or U16494 (N_16494,N_14993,N_14996);
or U16495 (N_16495,N_12097,N_14738);
xor U16496 (N_16496,N_13912,N_14855);
and U16497 (N_16497,N_13542,N_13144);
nand U16498 (N_16498,N_14860,N_13217);
or U16499 (N_16499,N_14065,N_13047);
nor U16500 (N_16500,N_13216,N_12923);
xor U16501 (N_16501,N_14134,N_13907);
nor U16502 (N_16502,N_14183,N_13788);
and U16503 (N_16503,N_14222,N_14078);
xor U16504 (N_16504,N_14784,N_13473);
and U16505 (N_16505,N_14244,N_14609);
nor U16506 (N_16506,N_14064,N_12114);
nand U16507 (N_16507,N_12604,N_12055);
or U16508 (N_16508,N_12579,N_12492);
xnor U16509 (N_16509,N_12242,N_14940);
and U16510 (N_16510,N_13662,N_13325);
or U16511 (N_16511,N_13408,N_12955);
nor U16512 (N_16512,N_13104,N_13080);
or U16513 (N_16513,N_12722,N_13695);
or U16514 (N_16514,N_12402,N_14457);
or U16515 (N_16515,N_14445,N_14607);
or U16516 (N_16516,N_13915,N_13283);
and U16517 (N_16517,N_13367,N_13883);
nand U16518 (N_16518,N_12332,N_14501);
nor U16519 (N_16519,N_12862,N_12526);
and U16520 (N_16520,N_14220,N_14281);
nor U16521 (N_16521,N_12192,N_13468);
or U16522 (N_16522,N_13114,N_12573);
nor U16523 (N_16523,N_13772,N_13471);
and U16524 (N_16524,N_14393,N_12458);
nor U16525 (N_16525,N_14823,N_12347);
or U16526 (N_16526,N_12124,N_14455);
and U16527 (N_16527,N_13352,N_13966);
and U16528 (N_16528,N_14174,N_14552);
nand U16529 (N_16529,N_12495,N_14477);
nor U16530 (N_16530,N_14138,N_14702);
or U16531 (N_16531,N_13037,N_12393);
or U16532 (N_16532,N_14952,N_12084);
or U16533 (N_16533,N_12029,N_12514);
and U16534 (N_16534,N_13912,N_14894);
xnor U16535 (N_16535,N_12823,N_13783);
and U16536 (N_16536,N_13781,N_13382);
and U16537 (N_16537,N_14320,N_13940);
or U16538 (N_16538,N_12224,N_14808);
nor U16539 (N_16539,N_12735,N_13722);
xor U16540 (N_16540,N_14558,N_13530);
and U16541 (N_16541,N_14764,N_13868);
nand U16542 (N_16542,N_12151,N_14021);
nand U16543 (N_16543,N_12729,N_12073);
nand U16544 (N_16544,N_14164,N_12540);
nand U16545 (N_16545,N_14727,N_14549);
nor U16546 (N_16546,N_12950,N_14742);
xor U16547 (N_16547,N_13617,N_13739);
nor U16548 (N_16548,N_12293,N_12716);
or U16549 (N_16549,N_13245,N_14784);
nor U16550 (N_16550,N_12312,N_14905);
nor U16551 (N_16551,N_12161,N_12250);
or U16552 (N_16552,N_14209,N_12776);
and U16553 (N_16553,N_14054,N_12767);
nand U16554 (N_16554,N_12106,N_12844);
nor U16555 (N_16555,N_12376,N_14272);
or U16556 (N_16556,N_12091,N_14278);
nand U16557 (N_16557,N_14788,N_14875);
nand U16558 (N_16558,N_12962,N_13636);
nand U16559 (N_16559,N_14895,N_12361);
xnor U16560 (N_16560,N_14383,N_13640);
and U16561 (N_16561,N_14228,N_14405);
or U16562 (N_16562,N_14792,N_14530);
and U16563 (N_16563,N_13963,N_13141);
or U16564 (N_16564,N_12798,N_14348);
nor U16565 (N_16565,N_14101,N_12836);
and U16566 (N_16566,N_13853,N_14013);
nand U16567 (N_16567,N_12245,N_12897);
or U16568 (N_16568,N_14462,N_12468);
and U16569 (N_16569,N_13628,N_12439);
xnor U16570 (N_16570,N_14303,N_12374);
nor U16571 (N_16571,N_12166,N_12583);
and U16572 (N_16572,N_13656,N_13372);
xnor U16573 (N_16573,N_14380,N_13699);
or U16574 (N_16574,N_13951,N_13036);
xor U16575 (N_16575,N_12879,N_12977);
and U16576 (N_16576,N_14595,N_12611);
or U16577 (N_16577,N_14083,N_14100);
xor U16578 (N_16578,N_14767,N_13866);
xnor U16579 (N_16579,N_12250,N_13601);
and U16580 (N_16580,N_12306,N_12059);
nor U16581 (N_16581,N_13338,N_13172);
nor U16582 (N_16582,N_13424,N_14601);
nand U16583 (N_16583,N_14923,N_14111);
or U16584 (N_16584,N_14225,N_13844);
and U16585 (N_16585,N_14490,N_14354);
nor U16586 (N_16586,N_12214,N_12362);
or U16587 (N_16587,N_13225,N_12363);
nor U16588 (N_16588,N_14756,N_12460);
nand U16589 (N_16589,N_13779,N_12152);
and U16590 (N_16590,N_14569,N_12279);
or U16591 (N_16591,N_12858,N_12285);
xor U16592 (N_16592,N_13914,N_14018);
or U16593 (N_16593,N_13008,N_12921);
or U16594 (N_16594,N_14749,N_12163);
nand U16595 (N_16595,N_13239,N_12275);
xor U16596 (N_16596,N_13250,N_12753);
nand U16597 (N_16597,N_14312,N_13419);
nand U16598 (N_16598,N_13222,N_12662);
and U16599 (N_16599,N_12089,N_13775);
nand U16600 (N_16600,N_12035,N_14759);
or U16601 (N_16601,N_14325,N_12957);
nor U16602 (N_16602,N_13690,N_14380);
nor U16603 (N_16603,N_12359,N_13670);
and U16604 (N_16604,N_14367,N_13066);
nor U16605 (N_16605,N_12445,N_14157);
or U16606 (N_16606,N_12875,N_13768);
or U16607 (N_16607,N_13450,N_13797);
and U16608 (N_16608,N_14137,N_14987);
xnor U16609 (N_16609,N_14500,N_12352);
or U16610 (N_16610,N_13239,N_13594);
xnor U16611 (N_16611,N_14209,N_14704);
or U16612 (N_16612,N_14222,N_12123);
nand U16613 (N_16613,N_12417,N_12592);
and U16614 (N_16614,N_12903,N_14007);
nand U16615 (N_16615,N_12642,N_12693);
or U16616 (N_16616,N_14427,N_14053);
nor U16617 (N_16617,N_12672,N_14210);
and U16618 (N_16618,N_14203,N_14120);
or U16619 (N_16619,N_13024,N_14037);
and U16620 (N_16620,N_13309,N_14290);
and U16621 (N_16621,N_13944,N_14534);
xnor U16622 (N_16622,N_14592,N_13506);
or U16623 (N_16623,N_13442,N_12711);
or U16624 (N_16624,N_12349,N_13780);
and U16625 (N_16625,N_13116,N_12295);
and U16626 (N_16626,N_13207,N_14573);
nor U16627 (N_16627,N_14661,N_14557);
nor U16628 (N_16628,N_12576,N_12697);
nand U16629 (N_16629,N_13726,N_13098);
or U16630 (N_16630,N_13110,N_12626);
nor U16631 (N_16631,N_12883,N_13265);
nor U16632 (N_16632,N_14368,N_13267);
and U16633 (N_16633,N_12680,N_13672);
and U16634 (N_16634,N_14491,N_12625);
nand U16635 (N_16635,N_13053,N_14897);
and U16636 (N_16636,N_12748,N_12498);
xor U16637 (N_16637,N_14021,N_14123);
nand U16638 (N_16638,N_13763,N_13322);
nand U16639 (N_16639,N_13878,N_14929);
and U16640 (N_16640,N_12830,N_13539);
and U16641 (N_16641,N_13643,N_14162);
and U16642 (N_16642,N_13797,N_12303);
xnor U16643 (N_16643,N_12040,N_12465);
nand U16644 (N_16644,N_14994,N_14498);
nand U16645 (N_16645,N_12775,N_13607);
nand U16646 (N_16646,N_13718,N_12806);
nand U16647 (N_16647,N_13144,N_12355);
nand U16648 (N_16648,N_13095,N_14969);
nor U16649 (N_16649,N_12650,N_14101);
xor U16650 (N_16650,N_12556,N_14412);
or U16651 (N_16651,N_14195,N_14444);
nor U16652 (N_16652,N_12857,N_13540);
and U16653 (N_16653,N_14802,N_13533);
nor U16654 (N_16654,N_14130,N_13615);
or U16655 (N_16655,N_13492,N_12902);
xor U16656 (N_16656,N_14969,N_12234);
or U16657 (N_16657,N_14521,N_14110);
xnor U16658 (N_16658,N_14656,N_12673);
nor U16659 (N_16659,N_14586,N_13702);
or U16660 (N_16660,N_12537,N_12531);
or U16661 (N_16661,N_13575,N_14170);
and U16662 (N_16662,N_14059,N_13724);
nor U16663 (N_16663,N_14757,N_13139);
nand U16664 (N_16664,N_14170,N_13287);
nor U16665 (N_16665,N_13619,N_14460);
or U16666 (N_16666,N_12913,N_13415);
nand U16667 (N_16667,N_14895,N_14982);
nand U16668 (N_16668,N_13750,N_14523);
xor U16669 (N_16669,N_12086,N_12939);
and U16670 (N_16670,N_12084,N_14008);
or U16671 (N_16671,N_14552,N_12600);
nor U16672 (N_16672,N_12369,N_12463);
xor U16673 (N_16673,N_13311,N_12910);
nor U16674 (N_16674,N_13502,N_13233);
nand U16675 (N_16675,N_13657,N_12652);
and U16676 (N_16676,N_14869,N_13893);
nand U16677 (N_16677,N_14439,N_13094);
or U16678 (N_16678,N_14556,N_14637);
xnor U16679 (N_16679,N_14363,N_13436);
or U16680 (N_16680,N_14629,N_12583);
and U16681 (N_16681,N_13419,N_14170);
xnor U16682 (N_16682,N_12228,N_14314);
or U16683 (N_16683,N_14155,N_13837);
nand U16684 (N_16684,N_13274,N_13296);
nor U16685 (N_16685,N_14146,N_14773);
nor U16686 (N_16686,N_14805,N_14087);
nor U16687 (N_16687,N_14874,N_13651);
nor U16688 (N_16688,N_12910,N_13161);
and U16689 (N_16689,N_14489,N_14044);
xor U16690 (N_16690,N_12715,N_13000);
nand U16691 (N_16691,N_14247,N_14016);
and U16692 (N_16692,N_13713,N_13931);
nand U16693 (N_16693,N_13103,N_14862);
or U16694 (N_16694,N_12790,N_14554);
nand U16695 (N_16695,N_14868,N_13638);
and U16696 (N_16696,N_14779,N_12443);
xnor U16697 (N_16697,N_12382,N_14525);
nand U16698 (N_16698,N_13462,N_13181);
and U16699 (N_16699,N_13553,N_14384);
xor U16700 (N_16700,N_12545,N_13251);
xor U16701 (N_16701,N_14572,N_13896);
nand U16702 (N_16702,N_14699,N_12946);
or U16703 (N_16703,N_13022,N_12069);
nand U16704 (N_16704,N_14264,N_13542);
or U16705 (N_16705,N_13269,N_13071);
and U16706 (N_16706,N_14937,N_12472);
or U16707 (N_16707,N_13445,N_12947);
and U16708 (N_16708,N_12840,N_12494);
nor U16709 (N_16709,N_14873,N_12838);
xor U16710 (N_16710,N_13696,N_13956);
or U16711 (N_16711,N_13308,N_12179);
xor U16712 (N_16712,N_13983,N_13857);
nor U16713 (N_16713,N_13343,N_14509);
or U16714 (N_16714,N_13137,N_14868);
and U16715 (N_16715,N_14233,N_12520);
or U16716 (N_16716,N_13792,N_12985);
nand U16717 (N_16717,N_14484,N_14423);
or U16718 (N_16718,N_13810,N_14267);
xnor U16719 (N_16719,N_13752,N_13608);
and U16720 (N_16720,N_14649,N_12476);
or U16721 (N_16721,N_12043,N_12939);
nand U16722 (N_16722,N_13793,N_14366);
and U16723 (N_16723,N_14881,N_12965);
and U16724 (N_16724,N_12424,N_12805);
nor U16725 (N_16725,N_14532,N_13542);
and U16726 (N_16726,N_13398,N_12862);
nor U16727 (N_16727,N_12182,N_12418);
nand U16728 (N_16728,N_14955,N_13489);
nand U16729 (N_16729,N_12109,N_13174);
and U16730 (N_16730,N_13293,N_12781);
xor U16731 (N_16731,N_13680,N_13188);
nand U16732 (N_16732,N_14477,N_14100);
and U16733 (N_16733,N_14794,N_12154);
nor U16734 (N_16734,N_13072,N_12725);
nor U16735 (N_16735,N_12241,N_12744);
nand U16736 (N_16736,N_14684,N_14625);
and U16737 (N_16737,N_12057,N_14474);
nand U16738 (N_16738,N_14377,N_14844);
or U16739 (N_16739,N_13025,N_12521);
nor U16740 (N_16740,N_12716,N_12120);
or U16741 (N_16741,N_12822,N_14358);
and U16742 (N_16742,N_13749,N_14353);
xor U16743 (N_16743,N_12755,N_14702);
and U16744 (N_16744,N_14441,N_13542);
and U16745 (N_16745,N_12221,N_12901);
and U16746 (N_16746,N_12956,N_12788);
nor U16747 (N_16747,N_13114,N_12962);
xnor U16748 (N_16748,N_14531,N_14822);
or U16749 (N_16749,N_14468,N_12245);
or U16750 (N_16750,N_14669,N_13215);
and U16751 (N_16751,N_13199,N_14259);
or U16752 (N_16752,N_13750,N_13023);
or U16753 (N_16753,N_13473,N_14948);
or U16754 (N_16754,N_12779,N_12943);
xnor U16755 (N_16755,N_14106,N_13551);
xor U16756 (N_16756,N_12617,N_12379);
nor U16757 (N_16757,N_12054,N_14396);
xnor U16758 (N_16758,N_13899,N_14177);
and U16759 (N_16759,N_13414,N_14962);
xor U16760 (N_16760,N_13299,N_14544);
or U16761 (N_16761,N_12179,N_14256);
nand U16762 (N_16762,N_12473,N_14418);
or U16763 (N_16763,N_13953,N_13778);
xor U16764 (N_16764,N_13750,N_12101);
and U16765 (N_16765,N_13529,N_14112);
nor U16766 (N_16766,N_12563,N_13331);
or U16767 (N_16767,N_13170,N_13204);
nor U16768 (N_16768,N_13995,N_12958);
xor U16769 (N_16769,N_13635,N_12782);
nand U16770 (N_16770,N_12481,N_13212);
or U16771 (N_16771,N_14825,N_14035);
or U16772 (N_16772,N_13876,N_12538);
and U16773 (N_16773,N_14204,N_14111);
and U16774 (N_16774,N_13016,N_12654);
nand U16775 (N_16775,N_13625,N_12098);
or U16776 (N_16776,N_14648,N_12541);
xor U16777 (N_16777,N_12737,N_12161);
and U16778 (N_16778,N_12598,N_14015);
nor U16779 (N_16779,N_12365,N_14133);
or U16780 (N_16780,N_12777,N_13570);
and U16781 (N_16781,N_14443,N_13699);
or U16782 (N_16782,N_14145,N_14585);
nand U16783 (N_16783,N_12030,N_13705);
xor U16784 (N_16784,N_14960,N_13437);
nor U16785 (N_16785,N_13061,N_12029);
xor U16786 (N_16786,N_12891,N_13309);
nand U16787 (N_16787,N_13854,N_14847);
xnor U16788 (N_16788,N_13987,N_13763);
nand U16789 (N_16789,N_12236,N_12441);
xor U16790 (N_16790,N_13042,N_12128);
and U16791 (N_16791,N_12527,N_13248);
nor U16792 (N_16792,N_12728,N_12139);
or U16793 (N_16793,N_13574,N_14152);
and U16794 (N_16794,N_14916,N_12679);
nor U16795 (N_16795,N_12329,N_14653);
and U16796 (N_16796,N_14601,N_14300);
xnor U16797 (N_16797,N_13152,N_14728);
or U16798 (N_16798,N_12837,N_14248);
nand U16799 (N_16799,N_14649,N_13617);
or U16800 (N_16800,N_12580,N_14445);
or U16801 (N_16801,N_14489,N_12054);
or U16802 (N_16802,N_13632,N_14217);
nor U16803 (N_16803,N_12447,N_12756);
nor U16804 (N_16804,N_13961,N_13559);
nor U16805 (N_16805,N_14929,N_12712);
and U16806 (N_16806,N_12878,N_14021);
nand U16807 (N_16807,N_13454,N_13178);
or U16808 (N_16808,N_13634,N_12756);
and U16809 (N_16809,N_14763,N_12564);
nand U16810 (N_16810,N_13504,N_14180);
nand U16811 (N_16811,N_14672,N_14897);
and U16812 (N_16812,N_14029,N_14436);
nor U16813 (N_16813,N_13603,N_12404);
nor U16814 (N_16814,N_14660,N_12458);
and U16815 (N_16815,N_12261,N_14520);
nor U16816 (N_16816,N_12313,N_13885);
nor U16817 (N_16817,N_14533,N_14174);
and U16818 (N_16818,N_12691,N_12591);
nor U16819 (N_16819,N_13807,N_12921);
or U16820 (N_16820,N_12670,N_14467);
nor U16821 (N_16821,N_14884,N_13570);
nor U16822 (N_16822,N_13842,N_12421);
xor U16823 (N_16823,N_14618,N_13805);
and U16824 (N_16824,N_12309,N_14848);
nand U16825 (N_16825,N_12809,N_13632);
xor U16826 (N_16826,N_14253,N_12754);
nand U16827 (N_16827,N_14892,N_14459);
xor U16828 (N_16828,N_12550,N_13708);
or U16829 (N_16829,N_13111,N_12247);
nand U16830 (N_16830,N_12150,N_14127);
nor U16831 (N_16831,N_12498,N_12336);
xor U16832 (N_16832,N_14980,N_13924);
xnor U16833 (N_16833,N_13566,N_12178);
nand U16834 (N_16834,N_14425,N_12834);
or U16835 (N_16835,N_12759,N_12373);
nand U16836 (N_16836,N_13396,N_12069);
and U16837 (N_16837,N_12587,N_14210);
nor U16838 (N_16838,N_14435,N_13604);
and U16839 (N_16839,N_12897,N_13104);
nor U16840 (N_16840,N_12470,N_14873);
nor U16841 (N_16841,N_13876,N_12953);
xor U16842 (N_16842,N_13092,N_14481);
and U16843 (N_16843,N_14767,N_12415);
nand U16844 (N_16844,N_13240,N_13907);
or U16845 (N_16845,N_12401,N_12609);
xnor U16846 (N_16846,N_13477,N_13176);
or U16847 (N_16847,N_14559,N_13606);
or U16848 (N_16848,N_13625,N_12184);
xor U16849 (N_16849,N_12816,N_12082);
and U16850 (N_16850,N_14579,N_14429);
or U16851 (N_16851,N_14921,N_14367);
xor U16852 (N_16852,N_13515,N_13419);
and U16853 (N_16853,N_13061,N_12203);
nor U16854 (N_16854,N_12497,N_12257);
xor U16855 (N_16855,N_13508,N_14950);
nor U16856 (N_16856,N_13344,N_14579);
nand U16857 (N_16857,N_12654,N_14931);
xnor U16858 (N_16858,N_14345,N_14802);
and U16859 (N_16859,N_14960,N_13000);
and U16860 (N_16860,N_13357,N_12830);
nand U16861 (N_16861,N_13004,N_13015);
and U16862 (N_16862,N_14087,N_13854);
nor U16863 (N_16863,N_14209,N_13153);
nand U16864 (N_16864,N_13668,N_13601);
and U16865 (N_16865,N_14356,N_14794);
or U16866 (N_16866,N_13823,N_14371);
and U16867 (N_16867,N_12717,N_14988);
xnor U16868 (N_16868,N_13349,N_14247);
nor U16869 (N_16869,N_12350,N_14481);
or U16870 (N_16870,N_13315,N_14169);
or U16871 (N_16871,N_13230,N_12529);
nor U16872 (N_16872,N_13140,N_12647);
or U16873 (N_16873,N_13167,N_12015);
nor U16874 (N_16874,N_14342,N_13952);
nor U16875 (N_16875,N_13213,N_13734);
nand U16876 (N_16876,N_13197,N_13656);
and U16877 (N_16877,N_13959,N_13322);
and U16878 (N_16878,N_13465,N_14995);
nor U16879 (N_16879,N_13320,N_14552);
xor U16880 (N_16880,N_14644,N_14254);
nand U16881 (N_16881,N_12663,N_13461);
or U16882 (N_16882,N_12527,N_13507);
and U16883 (N_16883,N_14684,N_13125);
nand U16884 (N_16884,N_12892,N_12153);
nor U16885 (N_16885,N_13226,N_12827);
nand U16886 (N_16886,N_14545,N_13926);
nand U16887 (N_16887,N_14955,N_13925);
nand U16888 (N_16888,N_14527,N_12063);
and U16889 (N_16889,N_14902,N_13240);
and U16890 (N_16890,N_14035,N_13243);
nand U16891 (N_16891,N_14574,N_12647);
nand U16892 (N_16892,N_14994,N_14024);
nand U16893 (N_16893,N_13929,N_13800);
or U16894 (N_16894,N_13584,N_14481);
nand U16895 (N_16895,N_14433,N_13027);
or U16896 (N_16896,N_13856,N_12867);
or U16897 (N_16897,N_12621,N_12493);
and U16898 (N_16898,N_13347,N_12129);
and U16899 (N_16899,N_12281,N_12213);
or U16900 (N_16900,N_13371,N_14841);
or U16901 (N_16901,N_13475,N_13570);
nand U16902 (N_16902,N_12824,N_12350);
nor U16903 (N_16903,N_12362,N_14895);
xor U16904 (N_16904,N_13977,N_13551);
nand U16905 (N_16905,N_13176,N_13475);
nor U16906 (N_16906,N_14800,N_13376);
xor U16907 (N_16907,N_14637,N_13036);
xnor U16908 (N_16908,N_14191,N_13476);
or U16909 (N_16909,N_14237,N_14471);
nand U16910 (N_16910,N_13355,N_14676);
and U16911 (N_16911,N_14210,N_13846);
xnor U16912 (N_16912,N_13340,N_12277);
nand U16913 (N_16913,N_14931,N_12613);
nand U16914 (N_16914,N_12485,N_12434);
nor U16915 (N_16915,N_14115,N_12509);
nand U16916 (N_16916,N_12824,N_14856);
and U16917 (N_16917,N_12017,N_13143);
xnor U16918 (N_16918,N_14224,N_13565);
or U16919 (N_16919,N_14593,N_12258);
or U16920 (N_16920,N_12401,N_14473);
nand U16921 (N_16921,N_13857,N_13102);
nor U16922 (N_16922,N_12711,N_14941);
xnor U16923 (N_16923,N_13920,N_14650);
nand U16924 (N_16924,N_14764,N_13181);
and U16925 (N_16925,N_12489,N_12999);
nor U16926 (N_16926,N_12634,N_14633);
xor U16927 (N_16927,N_12232,N_12266);
xor U16928 (N_16928,N_13667,N_12014);
nor U16929 (N_16929,N_13166,N_12802);
or U16930 (N_16930,N_12702,N_13798);
or U16931 (N_16931,N_12817,N_14626);
nand U16932 (N_16932,N_14407,N_14168);
and U16933 (N_16933,N_13060,N_13628);
xnor U16934 (N_16934,N_13382,N_12333);
xnor U16935 (N_16935,N_13883,N_14775);
nor U16936 (N_16936,N_13318,N_12228);
and U16937 (N_16937,N_13745,N_14432);
and U16938 (N_16938,N_14550,N_14742);
and U16939 (N_16939,N_12933,N_14660);
and U16940 (N_16940,N_12116,N_12920);
and U16941 (N_16941,N_13154,N_14268);
and U16942 (N_16942,N_14029,N_12795);
and U16943 (N_16943,N_13980,N_13999);
or U16944 (N_16944,N_14840,N_13084);
and U16945 (N_16945,N_14961,N_14302);
nand U16946 (N_16946,N_14310,N_13073);
or U16947 (N_16947,N_14721,N_12720);
nand U16948 (N_16948,N_12081,N_14008);
or U16949 (N_16949,N_12575,N_14334);
xor U16950 (N_16950,N_13363,N_14245);
or U16951 (N_16951,N_13399,N_14377);
xnor U16952 (N_16952,N_14086,N_13498);
and U16953 (N_16953,N_14149,N_12072);
nand U16954 (N_16954,N_12679,N_13185);
nor U16955 (N_16955,N_14363,N_13999);
and U16956 (N_16956,N_14094,N_14223);
and U16957 (N_16957,N_13288,N_13824);
nand U16958 (N_16958,N_12236,N_12536);
or U16959 (N_16959,N_12337,N_14869);
or U16960 (N_16960,N_13738,N_14386);
nor U16961 (N_16961,N_12059,N_14933);
and U16962 (N_16962,N_14979,N_12718);
and U16963 (N_16963,N_14014,N_13165);
or U16964 (N_16964,N_13277,N_12374);
nand U16965 (N_16965,N_13881,N_14910);
nor U16966 (N_16966,N_14524,N_12915);
and U16967 (N_16967,N_13931,N_14945);
nand U16968 (N_16968,N_14756,N_13868);
or U16969 (N_16969,N_12844,N_12824);
or U16970 (N_16970,N_13360,N_12387);
and U16971 (N_16971,N_13362,N_12822);
nor U16972 (N_16972,N_12962,N_13970);
xor U16973 (N_16973,N_13575,N_13824);
or U16974 (N_16974,N_12644,N_13700);
or U16975 (N_16975,N_13306,N_14010);
nand U16976 (N_16976,N_12416,N_14889);
or U16977 (N_16977,N_14846,N_14967);
xnor U16978 (N_16978,N_12550,N_13819);
xor U16979 (N_16979,N_13135,N_12243);
and U16980 (N_16980,N_13049,N_13989);
and U16981 (N_16981,N_14554,N_14305);
nand U16982 (N_16982,N_12261,N_14640);
or U16983 (N_16983,N_12767,N_12681);
or U16984 (N_16984,N_12778,N_12017);
xor U16985 (N_16985,N_12001,N_13942);
or U16986 (N_16986,N_14019,N_12962);
nand U16987 (N_16987,N_13014,N_14508);
nand U16988 (N_16988,N_14920,N_12213);
and U16989 (N_16989,N_13427,N_14611);
xnor U16990 (N_16990,N_13929,N_14996);
nor U16991 (N_16991,N_12528,N_13906);
nor U16992 (N_16992,N_12910,N_14612);
nand U16993 (N_16993,N_12222,N_12411);
nand U16994 (N_16994,N_13939,N_14662);
nand U16995 (N_16995,N_12960,N_13839);
nor U16996 (N_16996,N_14804,N_12203);
and U16997 (N_16997,N_13581,N_13182);
nor U16998 (N_16998,N_14120,N_13582);
and U16999 (N_16999,N_12705,N_12529);
or U17000 (N_17000,N_13006,N_12012);
or U17001 (N_17001,N_14641,N_12564);
and U17002 (N_17002,N_13747,N_12824);
nand U17003 (N_17003,N_13911,N_13314);
xor U17004 (N_17004,N_12969,N_13701);
nand U17005 (N_17005,N_14702,N_12994);
nand U17006 (N_17006,N_14138,N_13450);
nand U17007 (N_17007,N_13868,N_12961);
xor U17008 (N_17008,N_14497,N_12767);
and U17009 (N_17009,N_14914,N_12549);
or U17010 (N_17010,N_12893,N_12366);
and U17011 (N_17011,N_12495,N_14114);
xor U17012 (N_17012,N_13726,N_12260);
xnor U17013 (N_17013,N_13645,N_12773);
xnor U17014 (N_17014,N_12022,N_14137);
nor U17015 (N_17015,N_14996,N_14903);
or U17016 (N_17016,N_14433,N_13684);
and U17017 (N_17017,N_14317,N_13643);
nand U17018 (N_17018,N_14866,N_13581);
and U17019 (N_17019,N_12403,N_13137);
and U17020 (N_17020,N_13312,N_12277);
xor U17021 (N_17021,N_12184,N_12368);
nor U17022 (N_17022,N_13165,N_12244);
nor U17023 (N_17023,N_12409,N_13604);
xnor U17024 (N_17024,N_12120,N_14908);
nor U17025 (N_17025,N_13286,N_12687);
or U17026 (N_17026,N_12462,N_14412);
or U17027 (N_17027,N_13348,N_12451);
nand U17028 (N_17028,N_13993,N_14224);
or U17029 (N_17029,N_13872,N_12406);
and U17030 (N_17030,N_14308,N_12298);
nor U17031 (N_17031,N_12056,N_12286);
xor U17032 (N_17032,N_13840,N_13744);
or U17033 (N_17033,N_13529,N_13448);
nand U17034 (N_17034,N_12499,N_13002);
nor U17035 (N_17035,N_14664,N_12539);
nor U17036 (N_17036,N_12019,N_14761);
or U17037 (N_17037,N_14526,N_14393);
and U17038 (N_17038,N_12327,N_14899);
xor U17039 (N_17039,N_12415,N_14977);
or U17040 (N_17040,N_14394,N_13267);
and U17041 (N_17041,N_12939,N_14255);
and U17042 (N_17042,N_14786,N_13643);
or U17043 (N_17043,N_14801,N_13187);
or U17044 (N_17044,N_13303,N_12705);
or U17045 (N_17045,N_13708,N_13638);
and U17046 (N_17046,N_14510,N_12301);
xor U17047 (N_17047,N_12288,N_13447);
or U17048 (N_17048,N_13260,N_13411);
xor U17049 (N_17049,N_13993,N_14126);
and U17050 (N_17050,N_12122,N_14435);
nor U17051 (N_17051,N_13692,N_12934);
and U17052 (N_17052,N_14465,N_13548);
nand U17053 (N_17053,N_12969,N_12512);
xor U17054 (N_17054,N_14099,N_12241);
nor U17055 (N_17055,N_13129,N_14922);
xnor U17056 (N_17056,N_12840,N_13310);
or U17057 (N_17057,N_12067,N_12969);
nand U17058 (N_17058,N_13266,N_13476);
or U17059 (N_17059,N_13537,N_12398);
and U17060 (N_17060,N_14290,N_14551);
or U17061 (N_17061,N_14773,N_14015);
or U17062 (N_17062,N_14117,N_13583);
xor U17063 (N_17063,N_14328,N_13799);
and U17064 (N_17064,N_12133,N_12866);
nand U17065 (N_17065,N_13048,N_12970);
xnor U17066 (N_17066,N_12150,N_13914);
nand U17067 (N_17067,N_12504,N_12299);
nand U17068 (N_17068,N_13290,N_14418);
or U17069 (N_17069,N_14078,N_14256);
nor U17070 (N_17070,N_13195,N_12570);
and U17071 (N_17071,N_12815,N_14885);
and U17072 (N_17072,N_14503,N_14251);
nand U17073 (N_17073,N_12152,N_14489);
nor U17074 (N_17074,N_14994,N_14612);
and U17075 (N_17075,N_13672,N_13717);
nand U17076 (N_17076,N_12314,N_14562);
xnor U17077 (N_17077,N_13718,N_14416);
and U17078 (N_17078,N_14950,N_13852);
nand U17079 (N_17079,N_13023,N_12360);
and U17080 (N_17080,N_14303,N_14541);
or U17081 (N_17081,N_13423,N_13750);
nor U17082 (N_17082,N_14338,N_14553);
nand U17083 (N_17083,N_13251,N_13023);
and U17084 (N_17084,N_13508,N_12318);
xor U17085 (N_17085,N_12401,N_12254);
nor U17086 (N_17086,N_12569,N_12186);
xor U17087 (N_17087,N_13954,N_14557);
and U17088 (N_17088,N_14786,N_12473);
nand U17089 (N_17089,N_12936,N_14440);
nand U17090 (N_17090,N_12822,N_12453);
nor U17091 (N_17091,N_12970,N_12265);
nor U17092 (N_17092,N_14080,N_12949);
nand U17093 (N_17093,N_13984,N_14914);
nand U17094 (N_17094,N_13251,N_12853);
and U17095 (N_17095,N_12981,N_12697);
xnor U17096 (N_17096,N_12383,N_13712);
nor U17097 (N_17097,N_14725,N_12807);
and U17098 (N_17098,N_13446,N_12216);
or U17099 (N_17099,N_12876,N_13710);
nand U17100 (N_17100,N_14380,N_13412);
xor U17101 (N_17101,N_13639,N_14504);
or U17102 (N_17102,N_14743,N_14583);
and U17103 (N_17103,N_13637,N_14372);
or U17104 (N_17104,N_13605,N_13567);
nand U17105 (N_17105,N_13372,N_14670);
nand U17106 (N_17106,N_14956,N_14983);
nor U17107 (N_17107,N_14563,N_13353);
nand U17108 (N_17108,N_12854,N_14349);
xor U17109 (N_17109,N_12848,N_12165);
xnor U17110 (N_17110,N_12688,N_14039);
nand U17111 (N_17111,N_12244,N_13410);
nor U17112 (N_17112,N_14686,N_12206);
and U17113 (N_17113,N_13666,N_13347);
and U17114 (N_17114,N_14615,N_14228);
and U17115 (N_17115,N_13393,N_13441);
or U17116 (N_17116,N_12696,N_12432);
nand U17117 (N_17117,N_13046,N_14915);
nand U17118 (N_17118,N_12961,N_12703);
and U17119 (N_17119,N_14769,N_12134);
or U17120 (N_17120,N_12666,N_14064);
and U17121 (N_17121,N_13013,N_14209);
and U17122 (N_17122,N_12391,N_14484);
and U17123 (N_17123,N_12091,N_13181);
and U17124 (N_17124,N_12079,N_14627);
nand U17125 (N_17125,N_12951,N_14661);
and U17126 (N_17126,N_12785,N_12503);
nand U17127 (N_17127,N_12916,N_14055);
and U17128 (N_17128,N_14650,N_14523);
or U17129 (N_17129,N_14788,N_14497);
or U17130 (N_17130,N_12650,N_13179);
nor U17131 (N_17131,N_12802,N_12839);
nor U17132 (N_17132,N_12348,N_13551);
nand U17133 (N_17133,N_12668,N_12159);
nand U17134 (N_17134,N_13721,N_14627);
xnor U17135 (N_17135,N_12198,N_13221);
and U17136 (N_17136,N_14933,N_12535);
and U17137 (N_17137,N_12700,N_13229);
xnor U17138 (N_17138,N_12891,N_12240);
and U17139 (N_17139,N_12814,N_14251);
nor U17140 (N_17140,N_12127,N_14822);
and U17141 (N_17141,N_13240,N_13319);
xnor U17142 (N_17142,N_14670,N_14109);
nand U17143 (N_17143,N_14821,N_12922);
nor U17144 (N_17144,N_13970,N_12233);
and U17145 (N_17145,N_12850,N_13292);
nand U17146 (N_17146,N_14219,N_14777);
nor U17147 (N_17147,N_13438,N_12750);
or U17148 (N_17148,N_14590,N_12757);
and U17149 (N_17149,N_13517,N_14639);
and U17150 (N_17150,N_14843,N_12988);
xor U17151 (N_17151,N_14358,N_12411);
or U17152 (N_17152,N_13947,N_14074);
or U17153 (N_17153,N_13354,N_14243);
and U17154 (N_17154,N_12241,N_13427);
nor U17155 (N_17155,N_12408,N_14951);
nand U17156 (N_17156,N_12546,N_13202);
nand U17157 (N_17157,N_14300,N_12066);
or U17158 (N_17158,N_13347,N_12403);
or U17159 (N_17159,N_13573,N_12704);
nand U17160 (N_17160,N_13967,N_14129);
nor U17161 (N_17161,N_13729,N_14433);
nor U17162 (N_17162,N_14756,N_13968);
and U17163 (N_17163,N_12803,N_14755);
and U17164 (N_17164,N_13286,N_13772);
or U17165 (N_17165,N_13192,N_14593);
xor U17166 (N_17166,N_14982,N_12067);
nand U17167 (N_17167,N_12259,N_14694);
or U17168 (N_17168,N_12942,N_13273);
xor U17169 (N_17169,N_14752,N_12329);
nor U17170 (N_17170,N_14709,N_12878);
and U17171 (N_17171,N_14218,N_14259);
nand U17172 (N_17172,N_12405,N_13618);
nand U17173 (N_17173,N_14065,N_12917);
nand U17174 (N_17174,N_14366,N_14363);
nor U17175 (N_17175,N_14100,N_12687);
and U17176 (N_17176,N_14987,N_14854);
xor U17177 (N_17177,N_14901,N_14851);
and U17178 (N_17178,N_14875,N_12852);
nor U17179 (N_17179,N_13780,N_12616);
or U17180 (N_17180,N_12737,N_13929);
nor U17181 (N_17181,N_12886,N_13975);
and U17182 (N_17182,N_12835,N_13482);
xnor U17183 (N_17183,N_12445,N_14893);
nand U17184 (N_17184,N_14240,N_13354);
nand U17185 (N_17185,N_14745,N_12141);
and U17186 (N_17186,N_13360,N_12767);
or U17187 (N_17187,N_14130,N_13430);
and U17188 (N_17188,N_13005,N_14309);
and U17189 (N_17189,N_13092,N_14463);
nand U17190 (N_17190,N_12911,N_13713);
or U17191 (N_17191,N_12542,N_12214);
xor U17192 (N_17192,N_12652,N_14194);
nand U17193 (N_17193,N_13778,N_14870);
or U17194 (N_17194,N_12846,N_14931);
or U17195 (N_17195,N_13304,N_14333);
and U17196 (N_17196,N_14624,N_12904);
xor U17197 (N_17197,N_12842,N_14231);
xor U17198 (N_17198,N_12150,N_12552);
and U17199 (N_17199,N_13968,N_12319);
nand U17200 (N_17200,N_12854,N_14003);
or U17201 (N_17201,N_13138,N_14030);
nand U17202 (N_17202,N_13704,N_14665);
or U17203 (N_17203,N_12160,N_14346);
nand U17204 (N_17204,N_13513,N_14836);
xnor U17205 (N_17205,N_12800,N_12881);
or U17206 (N_17206,N_14298,N_14512);
nand U17207 (N_17207,N_12712,N_13881);
or U17208 (N_17208,N_13762,N_12279);
or U17209 (N_17209,N_13595,N_13119);
xor U17210 (N_17210,N_13022,N_12057);
or U17211 (N_17211,N_13660,N_14258);
xor U17212 (N_17212,N_12636,N_12966);
xor U17213 (N_17213,N_13280,N_12100);
xor U17214 (N_17214,N_13652,N_13426);
nand U17215 (N_17215,N_14144,N_12442);
nor U17216 (N_17216,N_12244,N_13062);
nand U17217 (N_17217,N_14030,N_12795);
or U17218 (N_17218,N_14596,N_14007);
nand U17219 (N_17219,N_12474,N_13591);
nor U17220 (N_17220,N_13828,N_14221);
and U17221 (N_17221,N_14544,N_12727);
xnor U17222 (N_17222,N_13233,N_13752);
and U17223 (N_17223,N_14016,N_12491);
and U17224 (N_17224,N_13342,N_12604);
nor U17225 (N_17225,N_14913,N_12451);
nor U17226 (N_17226,N_13556,N_12370);
nand U17227 (N_17227,N_14468,N_13207);
xnor U17228 (N_17228,N_13185,N_14085);
and U17229 (N_17229,N_12516,N_14517);
nor U17230 (N_17230,N_13629,N_14792);
or U17231 (N_17231,N_13305,N_14132);
and U17232 (N_17232,N_13331,N_12986);
nor U17233 (N_17233,N_12313,N_13330);
nor U17234 (N_17234,N_14819,N_13531);
nor U17235 (N_17235,N_14233,N_14569);
xnor U17236 (N_17236,N_13947,N_12855);
nand U17237 (N_17237,N_12112,N_12512);
or U17238 (N_17238,N_14299,N_13598);
nor U17239 (N_17239,N_14293,N_13634);
xor U17240 (N_17240,N_12174,N_13896);
nand U17241 (N_17241,N_13579,N_13866);
xor U17242 (N_17242,N_13100,N_14974);
nor U17243 (N_17243,N_12923,N_12164);
nor U17244 (N_17244,N_13229,N_12664);
xor U17245 (N_17245,N_13668,N_14997);
nor U17246 (N_17246,N_13549,N_14952);
and U17247 (N_17247,N_13323,N_14884);
nand U17248 (N_17248,N_14770,N_14983);
and U17249 (N_17249,N_12080,N_12090);
xor U17250 (N_17250,N_14330,N_12302);
and U17251 (N_17251,N_13394,N_12066);
and U17252 (N_17252,N_14150,N_13730);
nor U17253 (N_17253,N_12718,N_12468);
and U17254 (N_17254,N_12836,N_14059);
and U17255 (N_17255,N_13291,N_12249);
nor U17256 (N_17256,N_14557,N_14072);
nor U17257 (N_17257,N_13953,N_12536);
or U17258 (N_17258,N_14741,N_14149);
xnor U17259 (N_17259,N_12147,N_12556);
nand U17260 (N_17260,N_13559,N_13343);
nand U17261 (N_17261,N_13028,N_14343);
xor U17262 (N_17262,N_14673,N_14439);
and U17263 (N_17263,N_14268,N_13759);
and U17264 (N_17264,N_13272,N_13571);
xor U17265 (N_17265,N_12059,N_14678);
nand U17266 (N_17266,N_13413,N_13565);
xor U17267 (N_17267,N_13734,N_14398);
and U17268 (N_17268,N_12037,N_14011);
nor U17269 (N_17269,N_14954,N_13907);
nand U17270 (N_17270,N_14627,N_12985);
and U17271 (N_17271,N_13611,N_14781);
nand U17272 (N_17272,N_13980,N_12781);
and U17273 (N_17273,N_13585,N_13163);
and U17274 (N_17274,N_13118,N_14175);
or U17275 (N_17275,N_14798,N_13380);
nand U17276 (N_17276,N_14549,N_13331);
nor U17277 (N_17277,N_14345,N_13203);
and U17278 (N_17278,N_13609,N_13740);
nand U17279 (N_17279,N_12633,N_13064);
xor U17280 (N_17280,N_13839,N_12534);
nor U17281 (N_17281,N_12998,N_14530);
and U17282 (N_17282,N_13677,N_13603);
and U17283 (N_17283,N_12805,N_14914);
or U17284 (N_17284,N_13216,N_12196);
or U17285 (N_17285,N_13120,N_14804);
nand U17286 (N_17286,N_12548,N_13421);
nor U17287 (N_17287,N_14972,N_13275);
and U17288 (N_17288,N_12877,N_12690);
nand U17289 (N_17289,N_14928,N_14760);
or U17290 (N_17290,N_13320,N_12769);
xor U17291 (N_17291,N_12067,N_13540);
nor U17292 (N_17292,N_14060,N_13391);
or U17293 (N_17293,N_12293,N_14084);
nand U17294 (N_17294,N_13089,N_14452);
nand U17295 (N_17295,N_13229,N_13819);
or U17296 (N_17296,N_13060,N_14097);
nand U17297 (N_17297,N_12261,N_13857);
nor U17298 (N_17298,N_13795,N_13369);
and U17299 (N_17299,N_13417,N_14979);
nor U17300 (N_17300,N_12280,N_13084);
nor U17301 (N_17301,N_13271,N_13292);
and U17302 (N_17302,N_13933,N_13281);
or U17303 (N_17303,N_14949,N_12250);
nand U17304 (N_17304,N_13247,N_14653);
nor U17305 (N_17305,N_12110,N_13550);
xnor U17306 (N_17306,N_12131,N_13270);
or U17307 (N_17307,N_13731,N_12630);
xnor U17308 (N_17308,N_14292,N_13638);
and U17309 (N_17309,N_14667,N_12840);
or U17310 (N_17310,N_12928,N_13528);
nand U17311 (N_17311,N_12780,N_12088);
and U17312 (N_17312,N_12339,N_14081);
nor U17313 (N_17313,N_14789,N_14391);
nand U17314 (N_17314,N_13082,N_14080);
xor U17315 (N_17315,N_13091,N_14602);
xor U17316 (N_17316,N_12142,N_14473);
nor U17317 (N_17317,N_14148,N_14545);
nand U17318 (N_17318,N_13101,N_13420);
nor U17319 (N_17319,N_13917,N_13732);
nor U17320 (N_17320,N_12713,N_14966);
xnor U17321 (N_17321,N_12617,N_12197);
or U17322 (N_17322,N_13076,N_12979);
nor U17323 (N_17323,N_13127,N_12148);
xnor U17324 (N_17324,N_12993,N_13560);
or U17325 (N_17325,N_14318,N_13274);
nor U17326 (N_17326,N_13450,N_13498);
and U17327 (N_17327,N_12064,N_12905);
nand U17328 (N_17328,N_12346,N_13902);
xnor U17329 (N_17329,N_13119,N_13228);
and U17330 (N_17330,N_13356,N_12679);
nor U17331 (N_17331,N_14313,N_14675);
nand U17332 (N_17332,N_12337,N_13610);
nand U17333 (N_17333,N_14364,N_14056);
or U17334 (N_17334,N_13512,N_12266);
nand U17335 (N_17335,N_13613,N_12761);
nand U17336 (N_17336,N_13681,N_12098);
xnor U17337 (N_17337,N_14958,N_13782);
nor U17338 (N_17338,N_12154,N_12305);
and U17339 (N_17339,N_14247,N_12434);
nor U17340 (N_17340,N_14940,N_13095);
xor U17341 (N_17341,N_12125,N_13532);
and U17342 (N_17342,N_14631,N_14355);
nor U17343 (N_17343,N_13013,N_12950);
nand U17344 (N_17344,N_12785,N_12187);
nand U17345 (N_17345,N_13465,N_14593);
nor U17346 (N_17346,N_13312,N_14688);
and U17347 (N_17347,N_14723,N_14594);
xor U17348 (N_17348,N_14207,N_14589);
nand U17349 (N_17349,N_13455,N_14611);
nand U17350 (N_17350,N_14934,N_12088);
xnor U17351 (N_17351,N_13893,N_13679);
or U17352 (N_17352,N_14981,N_13069);
nor U17353 (N_17353,N_13511,N_14437);
and U17354 (N_17354,N_14771,N_13342);
or U17355 (N_17355,N_14487,N_12046);
or U17356 (N_17356,N_13909,N_12930);
nor U17357 (N_17357,N_13660,N_13777);
nand U17358 (N_17358,N_12537,N_13939);
nor U17359 (N_17359,N_14721,N_14852);
and U17360 (N_17360,N_14489,N_14443);
nand U17361 (N_17361,N_12354,N_12941);
xor U17362 (N_17362,N_13529,N_12781);
and U17363 (N_17363,N_12111,N_12951);
nor U17364 (N_17364,N_12909,N_13232);
xnor U17365 (N_17365,N_13836,N_13541);
nor U17366 (N_17366,N_14742,N_12412);
or U17367 (N_17367,N_12543,N_13305);
xnor U17368 (N_17368,N_12199,N_12347);
and U17369 (N_17369,N_13079,N_14714);
nor U17370 (N_17370,N_14162,N_12413);
and U17371 (N_17371,N_14674,N_12492);
or U17372 (N_17372,N_12357,N_13881);
nand U17373 (N_17373,N_14368,N_12889);
or U17374 (N_17374,N_14412,N_14708);
and U17375 (N_17375,N_14818,N_14900);
or U17376 (N_17376,N_13164,N_12742);
and U17377 (N_17377,N_12156,N_13438);
nor U17378 (N_17378,N_13852,N_12045);
xor U17379 (N_17379,N_14572,N_13823);
or U17380 (N_17380,N_14681,N_14170);
nand U17381 (N_17381,N_14882,N_12693);
or U17382 (N_17382,N_14810,N_12145);
and U17383 (N_17383,N_14563,N_13679);
xnor U17384 (N_17384,N_14448,N_14225);
xnor U17385 (N_17385,N_14448,N_14030);
xor U17386 (N_17386,N_14971,N_13779);
or U17387 (N_17387,N_12019,N_14804);
or U17388 (N_17388,N_14436,N_12827);
and U17389 (N_17389,N_14998,N_12136);
xor U17390 (N_17390,N_12164,N_12891);
nand U17391 (N_17391,N_13057,N_13678);
xor U17392 (N_17392,N_13390,N_14691);
xnor U17393 (N_17393,N_13391,N_13664);
or U17394 (N_17394,N_12292,N_12636);
or U17395 (N_17395,N_13920,N_12224);
xor U17396 (N_17396,N_13256,N_14555);
xnor U17397 (N_17397,N_13589,N_13962);
or U17398 (N_17398,N_12160,N_13760);
or U17399 (N_17399,N_12998,N_12951);
or U17400 (N_17400,N_12890,N_14764);
or U17401 (N_17401,N_13832,N_14526);
nor U17402 (N_17402,N_13438,N_13582);
nor U17403 (N_17403,N_13090,N_14663);
xnor U17404 (N_17404,N_14341,N_13062);
xor U17405 (N_17405,N_14888,N_14843);
nand U17406 (N_17406,N_13952,N_13349);
or U17407 (N_17407,N_14611,N_14230);
and U17408 (N_17408,N_12900,N_13246);
xor U17409 (N_17409,N_12024,N_13650);
nand U17410 (N_17410,N_13141,N_14942);
nor U17411 (N_17411,N_12150,N_14330);
or U17412 (N_17412,N_12119,N_13174);
and U17413 (N_17413,N_14332,N_13638);
nor U17414 (N_17414,N_12534,N_12324);
or U17415 (N_17415,N_13054,N_13999);
and U17416 (N_17416,N_13605,N_12262);
xnor U17417 (N_17417,N_14938,N_13977);
nand U17418 (N_17418,N_12168,N_12958);
and U17419 (N_17419,N_12194,N_13951);
xnor U17420 (N_17420,N_12421,N_12736);
and U17421 (N_17421,N_12645,N_14869);
and U17422 (N_17422,N_13768,N_12131);
and U17423 (N_17423,N_13576,N_12607);
or U17424 (N_17424,N_12396,N_13986);
xor U17425 (N_17425,N_13131,N_13063);
nand U17426 (N_17426,N_12698,N_13873);
nand U17427 (N_17427,N_13764,N_14082);
and U17428 (N_17428,N_12434,N_12465);
or U17429 (N_17429,N_13984,N_13367);
xnor U17430 (N_17430,N_13558,N_13668);
nand U17431 (N_17431,N_14578,N_12036);
xnor U17432 (N_17432,N_13822,N_14727);
nor U17433 (N_17433,N_12911,N_13294);
nand U17434 (N_17434,N_14715,N_13625);
nor U17435 (N_17435,N_14371,N_14369);
nand U17436 (N_17436,N_12808,N_12952);
and U17437 (N_17437,N_13566,N_12467);
or U17438 (N_17438,N_14438,N_12845);
nand U17439 (N_17439,N_14560,N_12960);
nand U17440 (N_17440,N_14882,N_13224);
xor U17441 (N_17441,N_14157,N_12702);
and U17442 (N_17442,N_14465,N_12779);
or U17443 (N_17443,N_14163,N_12364);
or U17444 (N_17444,N_13820,N_13414);
and U17445 (N_17445,N_13627,N_14347);
or U17446 (N_17446,N_13992,N_13060);
and U17447 (N_17447,N_14074,N_12172);
xor U17448 (N_17448,N_13631,N_14809);
nand U17449 (N_17449,N_12442,N_12010);
and U17450 (N_17450,N_13815,N_14785);
nor U17451 (N_17451,N_12861,N_12830);
nand U17452 (N_17452,N_13548,N_14928);
nand U17453 (N_17453,N_13092,N_12134);
and U17454 (N_17454,N_12513,N_12105);
or U17455 (N_17455,N_12313,N_14006);
nand U17456 (N_17456,N_13016,N_12773);
and U17457 (N_17457,N_12913,N_13995);
or U17458 (N_17458,N_13252,N_12429);
and U17459 (N_17459,N_14540,N_14720);
and U17460 (N_17460,N_13198,N_14874);
nor U17461 (N_17461,N_14122,N_14761);
and U17462 (N_17462,N_12167,N_12638);
nand U17463 (N_17463,N_13019,N_14714);
and U17464 (N_17464,N_14852,N_13789);
nand U17465 (N_17465,N_12226,N_13269);
xor U17466 (N_17466,N_14759,N_12334);
nand U17467 (N_17467,N_13849,N_14824);
and U17468 (N_17468,N_14070,N_12424);
or U17469 (N_17469,N_12810,N_13939);
or U17470 (N_17470,N_13224,N_13690);
xor U17471 (N_17471,N_13414,N_14778);
or U17472 (N_17472,N_14995,N_12763);
nor U17473 (N_17473,N_14977,N_13102);
xor U17474 (N_17474,N_14269,N_14453);
nor U17475 (N_17475,N_14637,N_13472);
nor U17476 (N_17476,N_12771,N_13209);
xor U17477 (N_17477,N_13319,N_13112);
or U17478 (N_17478,N_12927,N_12750);
or U17479 (N_17479,N_14732,N_12096);
nand U17480 (N_17480,N_12803,N_13026);
xnor U17481 (N_17481,N_13542,N_12425);
nand U17482 (N_17482,N_12728,N_13833);
xnor U17483 (N_17483,N_14676,N_13333);
xor U17484 (N_17484,N_12865,N_12566);
xor U17485 (N_17485,N_12868,N_14249);
nand U17486 (N_17486,N_13800,N_14581);
xnor U17487 (N_17487,N_13923,N_12445);
xor U17488 (N_17488,N_14617,N_12545);
and U17489 (N_17489,N_12422,N_12146);
or U17490 (N_17490,N_14708,N_12785);
or U17491 (N_17491,N_14446,N_13847);
nor U17492 (N_17492,N_13580,N_12966);
or U17493 (N_17493,N_12064,N_13631);
xor U17494 (N_17494,N_13907,N_12556);
xnor U17495 (N_17495,N_14365,N_13181);
and U17496 (N_17496,N_14129,N_12479);
and U17497 (N_17497,N_12842,N_14185);
or U17498 (N_17498,N_12818,N_12752);
nand U17499 (N_17499,N_13924,N_12758);
xnor U17500 (N_17500,N_14104,N_12608);
xnor U17501 (N_17501,N_12918,N_12166);
xor U17502 (N_17502,N_14477,N_13550);
nor U17503 (N_17503,N_14469,N_13459);
and U17504 (N_17504,N_12013,N_12490);
or U17505 (N_17505,N_13464,N_13612);
or U17506 (N_17506,N_14109,N_14700);
nor U17507 (N_17507,N_12010,N_12294);
xor U17508 (N_17508,N_13537,N_13209);
and U17509 (N_17509,N_13834,N_13851);
and U17510 (N_17510,N_12440,N_12706);
nand U17511 (N_17511,N_13298,N_12448);
xor U17512 (N_17512,N_14685,N_14935);
xor U17513 (N_17513,N_14186,N_14265);
nand U17514 (N_17514,N_14737,N_12813);
nor U17515 (N_17515,N_12354,N_14584);
nand U17516 (N_17516,N_12765,N_13705);
and U17517 (N_17517,N_13402,N_13659);
or U17518 (N_17518,N_12970,N_13210);
and U17519 (N_17519,N_12495,N_12712);
nor U17520 (N_17520,N_12707,N_14058);
xor U17521 (N_17521,N_13133,N_12259);
or U17522 (N_17522,N_13823,N_14352);
nand U17523 (N_17523,N_13113,N_13568);
xnor U17524 (N_17524,N_14363,N_13146);
or U17525 (N_17525,N_14377,N_12645);
and U17526 (N_17526,N_14157,N_14568);
or U17527 (N_17527,N_12328,N_12773);
and U17528 (N_17528,N_14349,N_13418);
nand U17529 (N_17529,N_13087,N_12184);
or U17530 (N_17530,N_12456,N_14107);
xnor U17531 (N_17531,N_14756,N_13140);
nand U17532 (N_17532,N_14142,N_13979);
nand U17533 (N_17533,N_12291,N_14535);
and U17534 (N_17534,N_12676,N_13303);
and U17535 (N_17535,N_14302,N_12262);
and U17536 (N_17536,N_12471,N_13708);
nor U17537 (N_17537,N_12480,N_12966);
xnor U17538 (N_17538,N_12960,N_12205);
or U17539 (N_17539,N_12070,N_14600);
nor U17540 (N_17540,N_12830,N_14373);
nand U17541 (N_17541,N_12183,N_14338);
nor U17542 (N_17542,N_14458,N_12201);
nor U17543 (N_17543,N_12373,N_12210);
nand U17544 (N_17544,N_13477,N_12536);
xnor U17545 (N_17545,N_13939,N_14629);
and U17546 (N_17546,N_12597,N_12282);
nor U17547 (N_17547,N_13558,N_12979);
nor U17548 (N_17548,N_12550,N_13945);
nor U17549 (N_17549,N_12736,N_12498);
xor U17550 (N_17550,N_13778,N_13974);
or U17551 (N_17551,N_14659,N_13658);
or U17552 (N_17552,N_13253,N_14365);
nand U17553 (N_17553,N_12296,N_14614);
and U17554 (N_17554,N_12700,N_12918);
xnor U17555 (N_17555,N_13751,N_12058);
or U17556 (N_17556,N_12323,N_14356);
xnor U17557 (N_17557,N_12354,N_14753);
nor U17558 (N_17558,N_14473,N_13090);
or U17559 (N_17559,N_12881,N_12340);
nor U17560 (N_17560,N_13957,N_12908);
nand U17561 (N_17561,N_14231,N_14012);
xor U17562 (N_17562,N_13982,N_12528);
nand U17563 (N_17563,N_14624,N_12898);
or U17564 (N_17564,N_12502,N_12239);
xor U17565 (N_17565,N_14452,N_13587);
nand U17566 (N_17566,N_14728,N_13813);
and U17567 (N_17567,N_12019,N_12863);
nor U17568 (N_17568,N_13421,N_13180);
nand U17569 (N_17569,N_12232,N_14028);
nand U17570 (N_17570,N_13129,N_13246);
xnor U17571 (N_17571,N_12836,N_13717);
and U17572 (N_17572,N_13706,N_12303);
nor U17573 (N_17573,N_14288,N_13643);
or U17574 (N_17574,N_13543,N_14224);
nor U17575 (N_17575,N_14445,N_14285);
and U17576 (N_17576,N_14671,N_14428);
xor U17577 (N_17577,N_12249,N_13204);
nand U17578 (N_17578,N_12637,N_13576);
nor U17579 (N_17579,N_13586,N_13267);
and U17580 (N_17580,N_14796,N_13768);
xnor U17581 (N_17581,N_12903,N_12953);
nand U17582 (N_17582,N_14789,N_12421);
nor U17583 (N_17583,N_12619,N_13986);
and U17584 (N_17584,N_13961,N_12127);
xnor U17585 (N_17585,N_13923,N_14000);
and U17586 (N_17586,N_12087,N_12204);
or U17587 (N_17587,N_13539,N_14033);
nor U17588 (N_17588,N_14130,N_12648);
and U17589 (N_17589,N_14692,N_13385);
or U17590 (N_17590,N_14701,N_12241);
and U17591 (N_17591,N_14051,N_14843);
nor U17592 (N_17592,N_14392,N_12669);
and U17593 (N_17593,N_12784,N_12981);
or U17594 (N_17594,N_12412,N_14606);
nand U17595 (N_17595,N_12309,N_13077);
nor U17596 (N_17596,N_12845,N_13618);
or U17597 (N_17597,N_12527,N_13401);
xnor U17598 (N_17598,N_12865,N_14012);
nand U17599 (N_17599,N_12191,N_13489);
or U17600 (N_17600,N_14973,N_12687);
xor U17601 (N_17601,N_13054,N_14157);
or U17602 (N_17602,N_13467,N_14025);
and U17603 (N_17603,N_13457,N_14910);
and U17604 (N_17604,N_12001,N_12616);
or U17605 (N_17605,N_14548,N_14531);
and U17606 (N_17606,N_14823,N_12123);
or U17607 (N_17607,N_14495,N_14021);
nor U17608 (N_17608,N_13918,N_14192);
xnor U17609 (N_17609,N_13701,N_13668);
nand U17610 (N_17610,N_14604,N_14217);
nand U17611 (N_17611,N_12402,N_14383);
and U17612 (N_17612,N_12767,N_14101);
and U17613 (N_17613,N_13305,N_13632);
nor U17614 (N_17614,N_13598,N_12563);
or U17615 (N_17615,N_12380,N_14280);
nand U17616 (N_17616,N_13077,N_13387);
or U17617 (N_17617,N_14338,N_13563);
and U17618 (N_17618,N_12675,N_12162);
nand U17619 (N_17619,N_13847,N_13432);
nand U17620 (N_17620,N_14408,N_13117);
or U17621 (N_17621,N_14890,N_14689);
and U17622 (N_17622,N_13273,N_13745);
nand U17623 (N_17623,N_12267,N_12665);
xor U17624 (N_17624,N_12608,N_14082);
xnor U17625 (N_17625,N_13307,N_12853);
and U17626 (N_17626,N_14565,N_14423);
nor U17627 (N_17627,N_13612,N_14519);
nand U17628 (N_17628,N_13150,N_14742);
nor U17629 (N_17629,N_13962,N_12015);
nor U17630 (N_17630,N_12084,N_13746);
nor U17631 (N_17631,N_14979,N_12887);
nand U17632 (N_17632,N_13893,N_12931);
nand U17633 (N_17633,N_14897,N_13786);
nor U17634 (N_17634,N_13776,N_13015);
or U17635 (N_17635,N_12724,N_14003);
nor U17636 (N_17636,N_12394,N_14512);
xor U17637 (N_17637,N_13537,N_13255);
xnor U17638 (N_17638,N_12970,N_13221);
nor U17639 (N_17639,N_13605,N_14470);
nand U17640 (N_17640,N_13435,N_14088);
or U17641 (N_17641,N_13168,N_14033);
nor U17642 (N_17642,N_14750,N_14430);
or U17643 (N_17643,N_12205,N_12771);
nor U17644 (N_17644,N_14591,N_13495);
or U17645 (N_17645,N_12268,N_13668);
and U17646 (N_17646,N_12650,N_13322);
or U17647 (N_17647,N_14723,N_14498);
nand U17648 (N_17648,N_12051,N_12235);
nor U17649 (N_17649,N_13303,N_13942);
nand U17650 (N_17650,N_14082,N_13448);
xor U17651 (N_17651,N_14759,N_12520);
xnor U17652 (N_17652,N_12673,N_12929);
nor U17653 (N_17653,N_12790,N_13515);
nor U17654 (N_17654,N_13532,N_13910);
or U17655 (N_17655,N_14441,N_12818);
nor U17656 (N_17656,N_12406,N_12178);
nor U17657 (N_17657,N_13928,N_12662);
and U17658 (N_17658,N_13648,N_14387);
or U17659 (N_17659,N_14940,N_13519);
or U17660 (N_17660,N_14986,N_13534);
or U17661 (N_17661,N_13900,N_12365);
xor U17662 (N_17662,N_12505,N_13482);
and U17663 (N_17663,N_12976,N_12109);
xnor U17664 (N_17664,N_12048,N_12261);
nand U17665 (N_17665,N_14409,N_14812);
and U17666 (N_17666,N_12478,N_14985);
and U17667 (N_17667,N_12998,N_14086);
or U17668 (N_17668,N_12957,N_13896);
or U17669 (N_17669,N_14038,N_14603);
or U17670 (N_17670,N_14697,N_14805);
or U17671 (N_17671,N_13838,N_13800);
nor U17672 (N_17672,N_14186,N_14721);
nand U17673 (N_17673,N_13894,N_12923);
xor U17674 (N_17674,N_12598,N_14513);
nor U17675 (N_17675,N_12936,N_12926);
nor U17676 (N_17676,N_12958,N_13378);
nand U17677 (N_17677,N_13054,N_12052);
nand U17678 (N_17678,N_13525,N_13374);
xor U17679 (N_17679,N_14615,N_12898);
nand U17680 (N_17680,N_12636,N_12475);
or U17681 (N_17681,N_12138,N_14509);
xnor U17682 (N_17682,N_13507,N_13657);
nand U17683 (N_17683,N_12876,N_12412);
nand U17684 (N_17684,N_13684,N_13646);
xor U17685 (N_17685,N_12149,N_14399);
nand U17686 (N_17686,N_12122,N_12944);
xor U17687 (N_17687,N_12225,N_13431);
nor U17688 (N_17688,N_12125,N_13222);
xor U17689 (N_17689,N_13866,N_12145);
or U17690 (N_17690,N_12911,N_12660);
nand U17691 (N_17691,N_14583,N_13264);
and U17692 (N_17692,N_13984,N_14899);
nor U17693 (N_17693,N_12032,N_13142);
nand U17694 (N_17694,N_14130,N_14826);
nand U17695 (N_17695,N_13115,N_14870);
or U17696 (N_17696,N_13013,N_14609);
xnor U17697 (N_17697,N_14167,N_12733);
nor U17698 (N_17698,N_12389,N_12974);
nand U17699 (N_17699,N_13004,N_14404);
nand U17700 (N_17700,N_14385,N_14066);
nand U17701 (N_17701,N_12542,N_13417);
or U17702 (N_17702,N_13456,N_12838);
nand U17703 (N_17703,N_12712,N_13733);
or U17704 (N_17704,N_13012,N_12788);
and U17705 (N_17705,N_12796,N_13082);
and U17706 (N_17706,N_14773,N_14705);
and U17707 (N_17707,N_12832,N_12416);
nand U17708 (N_17708,N_14451,N_13367);
xnor U17709 (N_17709,N_14274,N_12813);
nor U17710 (N_17710,N_13973,N_12261);
xor U17711 (N_17711,N_12418,N_12865);
nor U17712 (N_17712,N_13854,N_14334);
xor U17713 (N_17713,N_13115,N_13876);
nor U17714 (N_17714,N_14116,N_13817);
nand U17715 (N_17715,N_13305,N_12959);
nor U17716 (N_17716,N_14793,N_12266);
and U17717 (N_17717,N_14916,N_12024);
nor U17718 (N_17718,N_12016,N_14272);
nand U17719 (N_17719,N_12649,N_12621);
and U17720 (N_17720,N_14941,N_12424);
nand U17721 (N_17721,N_13585,N_12902);
nor U17722 (N_17722,N_12675,N_13834);
and U17723 (N_17723,N_14506,N_14883);
nor U17724 (N_17724,N_12262,N_13795);
and U17725 (N_17725,N_12757,N_12904);
xnor U17726 (N_17726,N_12503,N_13595);
or U17727 (N_17727,N_14610,N_14352);
nor U17728 (N_17728,N_12794,N_13582);
nand U17729 (N_17729,N_13221,N_13420);
xor U17730 (N_17730,N_12842,N_14413);
and U17731 (N_17731,N_14149,N_12104);
or U17732 (N_17732,N_12371,N_12949);
nor U17733 (N_17733,N_14264,N_14709);
or U17734 (N_17734,N_12451,N_12534);
and U17735 (N_17735,N_12524,N_13058);
xor U17736 (N_17736,N_14374,N_13026);
nor U17737 (N_17737,N_12101,N_12104);
xor U17738 (N_17738,N_14621,N_13510);
xor U17739 (N_17739,N_13934,N_14232);
nor U17740 (N_17740,N_14659,N_12813);
and U17741 (N_17741,N_12567,N_14261);
xnor U17742 (N_17742,N_12982,N_12663);
and U17743 (N_17743,N_12469,N_12967);
xnor U17744 (N_17744,N_12321,N_12108);
and U17745 (N_17745,N_13519,N_14158);
nor U17746 (N_17746,N_14548,N_13806);
and U17747 (N_17747,N_14828,N_14385);
nand U17748 (N_17748,N_12566,N_12879);
xor U17749 (N_17749,N_14922,N_12259);
and U17750 (N_17750,N_13533,N_12692);
and U17751 (N_17751,N_13038,N_14520);
xor U17752 (N_17752,N_13668,N_12006);
xnor U17753 (N_17753,N_13998,N_12416);
or U17754 (N_17754,N_13681,N_12277);
xor U17755 (N_17755,N_12406,N_12708);
or U17756 (N_17756,N_13570,N_12245);
xor U17757 (N_17757,N_14739,N_12633);
and U17758 (N_17758,N_13194,N_13837);
or U17759 (N_17759,N_14653,N_13999);
xor U17760 (N_17760,N_13030,N_12610);
nor U17761 (N_17761,N_13513,N_14660);
xnor U17762 (N_17762,N_12132,N_12974);
and U17763 (N_17763,N_14933,N_14209);
and U17764 (N_17764,N_12219,N_12849);
nand U17765 (N_17765,N_14360,N_14265);
xnor U17766 (N_17766,N_13403,N_13536);
xnor U17767 (N_17767,N_14148,N_12297);
nor U17768 (N_17768,N_12141,N_12111);
xnor U17769 (N_17769,N_13751,N_14390);
nand U17770 (N_17770,N_13751,N_14199);
xnor U17771 (N_17771,N_14753,N_12764);
nand U17772 (N_17772,N_12224,N_13239);
or U17773 (N_17773,N_14779,N_14068);
or U17774 (N_17774,N_12405,N_13379);
nor U17775 (N_17775,N_13060,N_13767);
nor U17776 (N_17776,N_13679,N_13727);
nand U17777 (N_17777,N_13360,N_14149);
or U17778 (N_17778,N_13276,N_14252);
nor U17779 (N_17779,N_13203,N_14778);
nand U17780 (N_17780,N_13708,N_14281);
or U17781 (N_17781,N_12866,N_13745);
nor U17782 (N_17782,N_14261,N_12340);
and U17783 (N_17783,N_14044,N_13125);
nor U17784 (N_17784,N_12372,N_13739);
nor U17785 (N_17785,N_12905,N_14428);
and U17786 (N_17786,N_12265,N_14640);
and U17787 (N_17787,N_13034,N_12251);
or U17788 (N_17788,N_13261,N_13385);
xor U17789 (N_17789,N_14066,N_12797);
nand U17790 (N_17790,N_13683,N_12843);
nor U17791 (N_17791,N_12875,N_13292);
and U17792 (N_17792,N_13005,N_13020);
nor U17793 (N_17793,N_12494,N_14613);
xor U17794 (N_17794,N_14661,N_12903);
or U17795 (N_17795,N_13468,N_12343);
nand U17796 (N_17796,N_13280,N_14788);
and U17797 (N_17797,N_12506,N_12204);
and U17798 (N_17798,N_13613,N_14749);
xnor U17799 (N_17799,N_13825,N_12627);
or U17800 (N_17800,N_14021,N_12301);
nand U17801 (N_17801,N_12783,N_14353);
nand U17802 (N_17802,N_14197,N_14168);
xnor U17803 (N_17803,N_12912,N_12936);
and U17804 (N_17804,N_13911,N_14481);
xor U17805 (N_17805,N_13163,N_13289);
or U17806 (N_17806,N_12403,N_12075);
and U17807 (N_17807,N_13301,N_12869);
and U17808 (N_17808,N_12092,N_13506);
nor U17809 (N_17809,N_12896,N_12037);
and U17810 (N_17810,N_14401,N_13752);
nand U17811 (N_17811,N_13168,N_14872);
xor U17812 (N_17812,N_12728,N_12165);
nand U17813 (N_17813,N_14521,N_13775);
and U17814 (N_17814,N_12228,N_12912);
and U17815 (N_17815,N_12433,N_14802);
xnor U17816 (N_17816,N_12907,N_13217);
or U17817 (N_17817,N_14984,N_12691);
nand U17818 (N_17818,N_12399,N_12989);
nand U17819 (N_17819,N_12118,N_13537);
nor U17820 (N_17820,N_14768,N_13626);
xnor U17821 (N_17821,N_14930,N_12327);
nor U17822 (N_17822,N_12934,N_12819);
nand U17823 (N_17823,N_12546,N_14276);
xnor U17824 (N_17824,N_12738,N_12244);
xnor U17825 (N_17825,N_13922,N_14049);
xor U17826 (N_17826,N_14787,N_14299);
and U17827 (N_17827,N_14956,N_13035);
xor U17828 (N_17828,N_14271,N_14933);
xnor U17829 (N_17829,N_13117,N_12141);
nor U17830 (N_17830,N_14781,N_13030);
or U17831 (N_17831,N_14284,N_12461);
nor U17832 (N_17832,N_13650,N_13872);
or U17833 (N_17833,N_12406,N_14938);
xnor U17834 (N_17834,N_12304,N_13142);
nand U17835 (N_17835,N_12650,N_14783);
nor U17836 (N_17836,N_14077,N_14871);
nor U17837 (N_17837,N_13448,N_14359);
xor U17838 (N_17838,N_14002,N_14151);
nor U17839 (N_17839,N_12036,N_14905);
xor U17840 (N_17840,N_14078,N_14794);
and U17841 (N_17841,N_12233,N_13246);
or U17842 (N_17842,N_12861,N_12279);
and U17843 (N_17843,N_12933,N_12842);
and U17844 (N_17844,N_13082,N_12246);
nor U17845 (N_17845,N_14170,N_12199);
or U17846 (N_17846,N_13581,N_12391);
nor U17847 (N_17847,N_14790,N_14017);
xor U17848 (N_17848,N_13748,N_14249);
and U17849 (N_17849,N_12785,N_14467);
nand U17850 (N_17850,N_12032,N_14540);
and U17851 (N_17851,N_14436,N_13775);
or U17852 (N_17852,N_13823,N_13145);
or U17853 (N_17853,N_12873,N_12447);
xnor U17854 (N_17854,N_12894,N_14972);
nor U17855 (N_17855,N_12165,N_14248);
nand U17856 (N_17856,N_13192,N_14347);
nor U17857 (N_17857,N_14909,N_13747);
xor U17858 (N_17858,N_14578,N_13198);
and U17859 (N_17859,N_14226,N_12021);
nand U17860 (N_17860,N_14818,N_13196);
and U17861 (N_17861,N_14477,N_13515);
and U17862 (N_17862,N_13556,N_14081);
nor U17863 (N_17863,N_13469,N_12114);
or U17864 (N_17864,N_12630,N_12245);
and U17865 (N_17865,N_14001,N_14639);
nand U17866 (N_17866,N_14451,N_13558);
or U17867 (N_17867,N_13411,N_14392);
nor U17868 (N_17868,N_13512,N_13607);
and U17869 (N_17869,N_14921,N_14281);
nor U17870 (N_17870,N_14958,N_14119);
nand U17871 (N_17871,N_14580,N_14178);
or U17872 (N_17872,N_13757,N_12247);
or U17873 (N_17873,N_13041,N_14606);
and U17874 (N_17874,N_12717,N_14082);
nor U17875 (N_17875,N_14645,N_12263);
xor U17876 (N_17876,N_13375,N_13455);
or U17877 (N_17877,N_14744,N_13590);
or U17878 (N_17878,N_12899,N_13976);
nor U17879 (N_17879,N_14316,N_14034);
nor U17880 (N_17880,N_12818,N_13940);
or U17881 (N_17881,N_13567,N_14286);
nand U17882 (N_17882,N_12099,N_12880);
and U17883 (N_17883,N_12986,N_12042);
or U17884 (N_17884,N_13407,N_13261);
nand U17885 (N_17885,N_14882,N_14280);
nand U17886 (N_17886,N_12628,N_13079);
or U17887 (N_17887,N_14253,N_14416);
and U17888 (N_17888,N_14153,N_13947);
and U17889 (N_17889,N_13110,N_14309);
nor U17890 (N_17890,N_14274,N_13148);
nor U17891 (N_17891,N_13472,N_12221);
or U17892 (N_17892,N_14270,N_13947);
or U17893 (N_17893,N_14425,N_13823);
nand U17894 (N_17894,N_14274,N_14561);
and U17895 (N_17895,N_12650,N_14118);
nor U17896 (N_17896,N_14430,N_12526);
and U17897 (N_17897,N_13899,N_14966);
xnor U17898 (N_17898,N_13246,N_12715);
and U17899 (N_17899,N_12221,N_14952);
nand U17900 (N_17900,N_14856,N_13601);
and U17901 (N_17901,N_12038,N_13376);
and U17902 (N_17902,N_12252,N_13600);
and U17903 (N_17903,N_13486,N_14588);
and U17904 (N_17904,N_14385,N_14965);
xnor U17905 (N_17905,N_12991,N_12643);
xnor U17906 (N_17906,N_13365,N_12606);
nand U17907 (N_17907,N_13109,N_13599);
nand U17908 (N_17908,N_12804,N_14973);
or U17909 (N_17909,N_13117,N_13430);
and U17910 (N_17910,N_14747,N_12105);
nor U17911 (N_17911,N_14439,N_12384);
nor U17912 (N_17912,N_13920,N_12836);
nor U17913 (N_17913,N_13784,N_12911);
nor U17914 (N_17914,N_13603,N_13709);
xnor U17915 (N_17915,N_12399,N_13994);
and U17916 (N_17916,N_14042,N_14998);
xnor U17917 (N_17917,N_14886,N_13954);
nor U17918 (N_17918,N_12186,N_12273);
xor U17919 (N_17919,N_12420,N_14408);
xnor U17920 (N_17920,N_13374,N_13370);
and U17921 (N_17921,N_14302,N_12285);
and U17922 (N_17922,N_13911,N_12006);
nand U17923 (N_17923,N_14504,N_14986);
nor U17924 (N_17924,N_13485,N_13677);
and U17925 (N_17925,N_12515,N_12315);
nand U17926 (N_17926,N_13541,N_13811);
nor U17927 (N_17927,N_14689,N_12759);
or U17928 (N_17928,N_14924,N_14435);
nand U17929 (N_17929,N_14283,N_12832);
and U17930 (N_17930,N_14957,N_12986);
nor U17931 (N_17931,N_12208,N_12201);
and U17932 (N_17932,N_14346,N_12211);
nand U17933 (N_17933,N_14331,N_12039);
nand U17934 (N_17934,N_14978,N_13307);
and U17935 (N_17935,N_14389,N_12237);
xnor U17936 (N_17936,N_12090,N_12904);
nand U17937 (N_17937,N_14003,N_14761);
and U17938 (N_17938,N_13294,N_14877);
or U17939 (N_17939,N_12586,N_14019);
xor U17940 (N_17940,N_13402,N_13526);
or U17941 (N_17941,N_12011,N_14641);
and U17942 (N_17942,N_14933,N_14013);
or U17943 (N_17943,N_14985,N_14831);
xnor U17944 (N_17944,N_12735,N_14316);
or U17945 (N_17945,N_13178,N_13595);
or U17946 (N_17946,N_12143,N_12641);
nand U17947 (N_17947,N_13354,N_13345);
or U17948 (N_17948,N_13484,N_13436);
xor U17949 (N_17949,N_14624,N_13301);
or U17950 (N_17950,N_13092,N_14206);
nand U17951 (N_17951,N_14784,N_14626);
nor U17952 (N_17952,N_12544,N_14290);
or U17953 (N_17953,N_13697,N_14908);
or U17954 (N_17954,N_12620,N_13032);
and U17955 (N_17955,N_14328,N_14700);
xnor U17956 (N_17956,N_14714,N_12143);
xor U17957 (N_17957,N_13165,N_14179);
nor U17958 (N_17958,N_13947,N_14574);
or U17959 (N_17959,N_14827,N_14739);
xor U17960 (N_17960,N_12786,N_14788);
nor U17961 (N_17961,N_13151,N_13952);
nor U17962 (N_17962,N_13133,N_13389);
xor U17963 (N_17963,N_12641,N_14558);
nand U17964 (N_17964,N_14646,N_12588);
or U17965 (N_17965,N_13375,N_14022);
nor U17966 (N_17966,N_13795,N_13461);
and U17967 (N_17967,N_12120,N_12901);
xor U17968 (N_17968,N_13867,N_13624);
or U17969 (N_17969,N_14112,N_13459);
nand U17970 (N_17970,N_12007,N_12579);
nor U17971 (N_17971,N_13150,N_13089);
nand U17972 (N_17972,N_12684,N_14364);
nand U17973 (N_17973,N_13191,N_14476);
nand U17974 (N_17974,N_13869,N_12127);
nand U17975 (N_17975,N_14124,N_14103);
xor U17976 (N_17976,N_13924,N_14190);
nand U17977 (N_17977,N_14484,N_12251);
and U17978 (N_17978,N_14657,N_14793);
nor U17979 (N_17979,N_14440,N_14457);
nor U17980 (N_17980,N_12627,N_13694);
xor U17981 (N_17981,N_13112,N_14567);
or U17982 (N_17982,N_12258,N_12101);
xor U17983 (N_17983,N_14356,N_12814);
nor U17984 (N_17984,N_14880,N_13117);
nor U17985 (N_17985,N_14935,N_14828);
and U17986 (N_17986,N_13943,N_13232);
and U17987 (N_17987,N_14844,N_12680);
and U17988 (N_17988,N_14101,N_13102);
xor U17989 (N_17989,N_13130,N_14472);
xor U17990 (N_17990,N_14615,N_12185);
and U17991 (N_17991,N_13876,N_12334);
and U17992 (N_17992,N_13194,N_13372);
and U17993 (N_17993,N_12633,N_12202);
nor U17994 (N_17994,N_13084,N_12166);
or U17995 (N_17995,N_13496,N_13986);
and U17996 (N_17996,N_13235,N_14165);
and U17997 (N_17997,N_12599,N_12512);
xnor U17998 (N_17998,N_13929,N_12146);
and U17999 (N_17999,N_13105,N_12854);
xor U18000 (N_18000,N_16554,N_15963);
nor U18001 (N_18001,N_17970,N_15276);
nor U18002 (N_18002,N_15094,N_17694);
xnor U18003 (N_18003,N_16804,N_17180);
nor U18004 (N_18004,N_17991,N_15071);
nor U18005 (N_18005,N_16197,N_15670);
xor U18006 (N_18006,N_17816,N_16961);
or U18007 (N_18007,N_15910,N_15160);
xnor U18008 (N_18008,N_16512,N_17161);
and U18009 (N_18009,N_15912,N_17939);
nand U18010 (N_18010,N_15344,N_17092);
nand U18011 (N_18011,N_16707,N_17921);
or U18012 (N_18012,N_15602,N_17010);
nor U18013 (N_18013,N_15971,N_17402);
nor U18014 (N_18014,N_16112,N_17914);
nor U18015 (N_18015,N_17143,N_16702);
xor U18016 (N_18016,N_17499,N_16897);
nand U18017 (N_18017,N_16407,N_17496);
or U18018 (N_18018,N_16136,N_16157);
and U18019 (N_18019,N_17788,N_17761);
or U18020 (N_18020,N_17200,N_17481);
or U18021 (N_18021,N_17309,N_17488);
xor U18022 (N_18022,N_15657,N_15023);
xnor U18023 (N_18023,N_16833,N_17288);
nor U18024 (N_18024,N_17450,N_15329);
or U18025 (N_18025,N_17734,N_17426);
xnor U18026 (N_18026,N_16859,N_15612);
nand U18027 (N_18027,N_15949,N_15141);
and U18028 (N_18028,N_15666,N_17222);
xnor U18029 (N_18029,N_16320,N_15114);
or U18030 (N_18030,N_17193,N_16925);
xnor U18031 (N_18031,N_16359,N_15146);
and U18032 (N_18032,N_15957,N_16577);
or U18033 (N_18033,N_16033,N_17836);
xor U18034 (N_18034,N_16392,N_17291);
or U18035 (N_18035,N_16864,N_15998);
nor U18036 (N_18036,N_15645,N_16997);
nand U18037 (N_18037,N_17216,N_15091);
nand U18038 (N_18038,N_15991,N_15954);
nor U18039 (N_18039,N_15376,N_17619);
xnor U18040 (N_18040,N_15567,N_16884);
nand U18041 (N_18041,N_17154,N_16432);
or U18042 (N_18042,N_17243,N_15857);
xnor U18043 (N_18043,N_17775,N_17155);
nand U18044 (N_18044,N_16673,N_15128);
xor U18045 (N_18045,N_15025,N_16663);
xnor U18046 (N_18046,N_16115,N_16789);
nand U18047 (N_18047,N_15327,N_16031);
nor U18048 (N_18048,N_17275,N_16626);
xnor U18049 (N_18049,N_15403,N_16269);
nor U18050 (N_18050,N_17740,N_17937);
xor U18051 (N_18051,N_16694,N_16247);
or U18052 (N_18052,N_16800,N_17702);
xnor U18053 (N_18053,N_15297,N_17475);
nand U18054 (N_18054,N_16920,N_15671);
xnor U18055 (N_18055,N_15153,N_15798);
nor U18056 (N_18056,N_15152,N_15575);
or U18057 (N_18057,N_16250,N_17879);
and U18058 (N_18058,N_15808,N_17037);
and U18059 (N_18059,N_17951,N_17710);
and U18060 (N_18060,N_17729,N_17063);
nand U18061 (N_18061,N_17299,N_17301);
nand U18062 (N_18062,N_16713,N_17576);
nor U18063 (N_18063,N_15404,N_17132);
xnor U18064 (N_18064,N_15188,N_16916);
xor U18065 (N_18065,N_15159,N_16492);
or U18066 (N_18066,N_16449,N_15288);
nand U18067 (N_18067,N_15328,N_17380);
nand U18068 (N_18068,N_15467,N_16922);
or U18069 (N_18069,N_17384,N_17190);
xor U18070 (N_18070,N_17467,N_15417);
xor U18071 (N_18071,N_16621,N_17188);
and U18072 (N_18072,N_17510,N_16443);
xor U18073 (N_18073,N_15945,N_17712);
nor U18074 (N_18074,N_16990,N_16646);
or U18075 (N_18075,N_15975,N_17776);
xnor U18076 (N_18076,N_16245,N_17876);
and U18077 (N_18077,N_15999,N_17428);
or U18078 (N_18078,N_16541,N_16814);
nor U18079 (N_18079,N_16214,N_16519);
xor U18080 (N_18080,N_17144,N_17731);
and U18081 (N_18081,N_15187,N_17007);
xor U18082 (N_18082,N_17432,N_17906);
xor U18083 (N_18083,N_17483,N_16945);
xnor U18084 (N_18084,N_17588,N_17056);
xnor U18085 (N_18085,N_16746,N_15247);
xnor U18086 (N_18086,N_17627,N_16678);
or U18087 (N_18087,N_16855,N_17471);
or U18088 (N_18088,N_17854,N_15885);
nand U18089 (N_18089,N_15075,N_15805);
nor U18090 (N_18090,N_16579,N_16732);
and U18091 (N_18091,N_15295,N_17461);
xnor U18092 (N_18092,N_16275,N_15569);
and U18093 (N_18093,N_17703,N_16476);
and U18094 (N_18094,N_15488,N_17041);
nor U18095 (N_18095,N_16447,N_15844);
nand U18096 (N_18096,N_15773,N_16527);
xor U18097 (N_18097,N_16409,N_16865);
nor U18098 (N_18098,N_15387,N_17016);
nand U18099 (N_18099,N_16711,N_16500);
and U18100 (N_18100,N_16046,N_17520);
xnor U18101 (N_18101,N_16415,N_16977);
or U18102 (N_18102,N_15758,N_15014);
nand U18103 (N_18103,N_17221,N_16330);
and U18104 (N_18104,N_16844,N_15110);
and U18105 (N_18105,N_15699,N_17967);
nand U18106 (N_18106,N_17726,N_17030);
or U18107 (N_18107,N_16040,N_15951);
nand U18108 (N_18108,N_16162,N_17036);
xor U18109 (N_18109,N_17466,N_16216);
nand U18110 (N_18110,N_17374,N_15797);
or U18111 (N_18111,N_16056,N_16687);
xnor U18112 (N_18112,N_16306,N_17187);
or U18113 (N_18113,N_16236,N_16662);
nor U18114 (N_18114,N_16129,N_15219);
and U18115 (N_18115,N_16496,N_15121);
and U18116 (N_18116,N_17548,N_17650);
or U18117 (N_18117,N_15356,N_17283);
nand U18118 (N_18118,N_16367,N_15752);
and U18119 (N_18119,N_17138,N_17070);
or U18120 (N_18120,N_16596,N_15930);
and U18121 (N_18121,N_17868,N_15096);
and U18122 (N_18122,N_16086,N_17071);
xnor U18123 (N_18123,N_16647,N_15068);
and U18124 (N_18124,N_17175,N_17199);
nor U18125 (N_18125,N_15709,N_17617);
or U18126 (N_18126,N_15070,N_15231);
and U18127 (N_18127,N_15464,N_16061);
or U18128 (N_18128,N_15533,N_15063);
nand U18129 (N_18129,N_17434,N_17083);
nor U18130 (N_18130,N_17003,N_17318);
nor U18131 (N_18131,N_17814,N_17556);
nand U18132 (N_18132,N_15543,N_17119);
xnor U18133 (N_18133,N_15561,N_15478);
or U18134 (N_18134,N_17514,N_15795);
nand U18135 (N_18135,N_16140,N_15108);
or U18136 (N_18136,N_16095,N_16340);
nor U18137 (N_18137,N_16907,N_16354);
nor U18138 (N_18138,N_15375,N_15674);
or U18139 (N_18139,N_17074,N_16953);
or U18140 (N_18140,N_16159,N_16516);
nor U18141 (N_18141,N_15350,N_16875);
xnor U18142 (N_18142,N_16421,N_16766);
nor U18143 (N_18143,N_16776,N_16847);
xor U18144 (N_18144,N_15832,N_17172);
and U18145 (N_18145,N_15009,N_15633);
nor U18146 (N_18146,N_15751,N_17508);
and U18147 (N_18147,N_15904,N_17420);
xor U18148 (N_18148,N_17769,N_15320);
nand U18149 (N_18149,N_15200,N_17386);
nand U18150 (N_18150,N_16886,N_17060);
and U18151 (N_18151,N_17176,N_15225);
and U18152 (N_18152,N_17406,N_15580);
or U18153 (N_18153,N_15410,N_17111);
and U18154 (N_18154,N_15800,N_17691);
or U18155 (N_18155,N_15463,N_16104);
and U18156 (N_18156,N_15414,N_15466);
xnor U18157 (N_18157,N_16529,N_17411);
and U18158 (N_18158,N_17821,N_15263);
nand U18159 (N_18159,N_17196,N_17160);
and U18160 (N_18160,N_15066,N_17635);
nand U18161 (N_18161,N_16092,N_15482);
nor U18162 (N_18162,N_16062,N_16866);
nand U18163 (N_18163,N_17944,N_15024);
nand U18164 (N_18164,N_15248,N_16700);
nor U18165 (N_18165,N_16297,N_16989);
xor U18166 (N_18166,N_16353,N_16901);
nor U18167 (N_18167,N_16549,N_17986);
xnor U18168 (N_18168,N_17128,N_16265);
nor U18169 (N_18169,N_16756,N_15815);
or U18170 (N_18170,N_17415,N_15085);
nor U18171 (N_18171,N_17423,N_15245);
nor U18172 (N_18172,N_15677,N_17608);
and U18173 (N_18173,N_17798,N_17053);
or U18174 (N_18174,N_17742,N_16994);
or U18175 (N_18175,N_17271,N_15481);
and U18176 (N_18176,N_15591,N_16173);
nand U18177 (N_18177,N_15166,N_17730);
xnor U18178 (N_18178,N_17898,N_17201);
xnor U18179 (N_18179,N_17760,N_16175);
xor U18180 (N_18180,N_17957,N_17293);
nand U18181 (N_18181,N_15782,N_17335);
nor U18182 (N_18182,N_15544,N_16240);
nand U18183 (N_18183,N_17399,N_17373);
or U18184 (N_18184,N_17048,N_17215);
xor U18185 (N_18185,N_16831,N_17519);
and U18186 (N_18186,N_17897,N_17255);
nand U18187 (N_18187,N_15611,N_15809);
xnor U18188 (N_18188,N_17224,N_16282);
xor U18189 (N_18189,N_15262,N_17503);
nor U18190 (N_18190,N_16422,N_16317);
nor U18191 (N_18191,N_15956,N_17709);
or U18192 (N_18192,N_17085,N_16377);
nor U18193 (N_18193,N_17971,N_16671);
or U18194 (N_18194,N_15652,N_17493);
xnor U18195 (N_18195,N_17727,N_17353);
xor U18196 (N_18196,N_16450,N_17648);
xnor U18197 (N_18197,N_15416,N_17403);
nand U18198 (N_18198,N_17571,N_17717);
and U18199 (N_18199,N_16244,N_16637);
and U18200 (N_18200,N_15541,N_17205);
and U18201 (N_18201,N_16934,N_16771);
and U18202 (N_18202,N_17930,N_17858);
or U18203 (N_18203,N_16352,N_16717);
nand U18204 (N_18204,N_16108,N_15681);
xnor U18205 (N_18205,N_17529,N_16429);
and U18206 (N_18206,N_16283,N_17670);
xnor U18207 (N_18207,N_16440,N_16542);
nor U18208 (N_18208,N_16948,N_15660);
and U18209 (N_18209,N_17330,N_15663);
nand U18210 (N_18210,N_17140,N_17361);
or U18211 (N_18211,N_15624,N_17182);
nand U18212 (N_18212,N_16490,N_17351);
xnor U18213 (N_18213,N_15032,N_16470);
or U18214 (N_18214,N_15801,N_16725);
nand U18215 (N_18215,N_15953,N_17396);
nand U18216 (N_18216,N_17823,N_16648);
nor U18217 (N_18217,N_15545,N_15590);
or U18218 (N_18218,N_17162,N_15233);
nand U18219 (N_18219,N_16345,N_17113);
xor U18220 (N_18220,N_17341,N_16085);
and U18221 (N_18221,N_15948,N_16227);
nor U18222 (N_18222,N_15347,N_17334);
and U18223 (N_18223,N_16419,N_16505);
or U18224 (N_18224,N_15747,N_17297);
nor U18225 (N_18225,N_16551,N_17436);
nand U18226 (N_18226,N_17546,N_16088);
nor U18227 (N_18227,N_17014,N_15040);
nor U18228 (N_18228,N_16399,N_17357);
and U18229 (N_18229,N_16553,N_17312);
nand U18230 (N_18230,N_15315,N_17383);
or U18231 (N_18231,N_16729,N_17072);
or U18232 (N_18232,N_15972,N_16817);
and U18233 (N_18233,N_17468,N_16401);
xor U18234 (N_18234,N_16891,N_17872);
nor U18235 (N_18235,N_16544,N_15348);
nand U18236 (N_18236,N_16444,N_15252);
and U18237 (N_18237,N_15059,N_15104);
and U18238 (N_18238,N_17578,N_16774);
nand U18239 (N_18239,N_17080,N_15651);
or U18240 (N_18240,N_15299,N_16965);
and U18241 (N_18241,N_15579,N_16150);
and U18242 (N_18242,N_15436,N_15157);
or U18243 (N_18243,N_17579,N_16225);
and U18244 (N_18244,N_16737,N_15301);
xnor U18245 (N_18245,N_17961,N_15537);
nor U18246 (N_18246,N_17664,N_17238);
or U18247 (N_18247,N_16810,N_16180);
nand U18248 (N_18248,N_17601,N_15371);
xnor U18249 (N_18249,N_15764,N_16135);
nor U18250 (N_18250,N_16455,N_17629);
and U18251 (N_18251,N_15973,N_17560);
or U18252 (N_18252,N_16777,N_15664);
and U18253 (N_18253,N_16769,N_16193);
nor U18254 (N_18254,N_16581,N_17737);
xor U18255 (N_18255,N_17538,N_17684);
nor U18256 (N_18256,N_15088,N_17225);
nand U18257 (N_18257,N_17981,N_15985);
xnor U18258 (N_18258,N_17804,N_17076);
and U18259 (N_18259,N_17870,N_16107);
nand U18260 (N_18260,N_15163,N_17343);
or U18261 (N_18261,N_16947,N_16261);
and U18262 (N_18262,N_16751,N_16758);
nor U18263 (N_18263,N_15861,N_16940);
xnor U18264 (N_18264,N_17735,N_17460);
nor U18265 (N_18265,N_16044,N_15659);
xnor U18266 (N_18266,N_16828,N_16658);
nor U18267 (N_18267,N_16845,N_15847);
nand U18268 (N_18268,N_15211,N_16363);
or U18269 (N_18269,N_17618,N_15909);
xor U18270 (N_18270,N_15531,N_15803);
nand U18271 (N_18271,N_17218,N_17231);
nor U18272 (N_18272,N_16764,N_17758);
nand U18273 (N_18273,N_15087,N_17485);
nand U18274 (N_18274,N_17605,N_17401);
and U18275 (N_18275,N_15817,N_15846);
and U18276 (N_18276,N_17905,N_17574);
nand U18277 (N_18277,N_17259,N_16651);
nand U18278 (N_18278,N_15309,N_15117);
and U18279 (N_18279,N_16745,N_15287);
and U18280 (N_18280,N_16563,N_17051);
and U18281 (N_18281,N_15272,N_16972);
or U18282 (N_18282,N_15931,N_17536);
xnor U18283 (N_18283,N_16172,N_17120);
nor U18284 (N_18284,N_17077,N_17765);
and U18285 (N_18285,N_16457,N_16358);
or U18286 (N_18286,N_16846,N_15584);
xnor U18287 (N_18287,N_17494,N_17972);
xor U18288 (N_18288,N_15881,N_15177);
nor U18289 (N_18289,N_15449,N_17369);
nand U18290 (N_18290,N_17194,N_16114);
nand U18291 (N_18291,N_15078,N_16942);
nor U18292 (N_18292,N_15065,N_17808);
nor U18293 (N_18293,N_17078,N_15103);
and U18294 (N_18294,N_17491,N_15400);
and U18295 (N_18295,N_17362,N_16735);
nand U18296 (N_18296,N_15422,N_17757);
or U18297 (N_18297,N_17929,N_15813);
xnor U18298 (N_18298,N_17311,N_15997);
nor U18299 (N_18299,N_16686,N_15713);
and U18300 (N_18300,N_17260,N_17178);
or U18301 (N_18301,N_16589,N_17593);
nor U18302 (N_18302,N_17896,N_16278);
nand U18303 (N_18303,N_15194,N_15250);
and U18304 (N_18304,N_17504,N_15044);
or U18305 (N_18305,N_16691,N_16664);
or U18306 (N_18306,N_17746,N_16808);
nand U18307 (N_18307,N_16304,N_17567);
nor U18308 (N_18308,N_16313,N_16073);
or U18309 (N_18309,N_15367,N_16794);
or U18310 (N_18310,N_16856,N_15394);
nor U18311 (N_18311,N_16347,N_15656);
nand U18312 (N_18312,N_16023,N_15908);
xor U18313 (N_18313,N_16127,N_15619);
nor U18314 (N_18314,N_16744,N_15443);
nand U18315 (N_18315,N_15457,N_16234);
xor U18316 (N_18316,N_16154,N_16274);
and U18317 (N_18317,N_17675,N_15538);
xor U18318 (N_18318,N_16991,N_15778);
and U18319 (N_18319,N_15695,N_15921);
and U18320 (N_18320,N_15323,N_17229);
and U18321 (N_18321,N_17697,N_17114);
and U18322 (N_18322,N_17652,N_16381);
nand U18323 (N_18323,N_16030,N_16070);
or U18324 (N_18324,N_15886,N_15691);
nor U18325 (N_18325,N_15831,N_16843);
nand U18326 (N_18326,N_15594,N_15201);
nor U18327 (N_18327,N_16209,N_16398);
nand U18328 (N_18328,N_17705,N_16966);
nand U18329 (N_18329,N_16185,N_17378);
or U18330 (N_18330,N_16018,N_17382);
or U18331 (N_18331,N_16243,N_16933);
nor U18332 (N_18332,N_15130,N_16305);
nand U18333 (N_18333,N_16566,N_15317);
nor U18334 (N_18334,N_15614,N_16893);
nand U18335 (N_18335,N_15833,N_16464);
or U18336 (N_18336,N_15253,N_16229);
xor U18337 (N_18337,N_17342,N_17785);
xnor U18338 (N_18338,N_16680,N_17751);
xnor U18339 (N_18339,N_16650,N_17557);
xor U18340 (N_18340,N_16326,N_17533);
and U18341 (N_18341,N_16821,N_15525);
xor U18342 (N_18342,N_15812,N_16970);
and U18343 (N_18343,N_17098,N_17541);
and U18344 (N_18344,N_16501,N_15551);
or U18345 (N_18345,N_17217,N_17568);
or U18346 (N_18346,N_15702,N_17998);
and U18347 (N_18347,N_16208,N_15916);
xor U18348 (N_18348,N_16649,N_15576);
or U18349 (N_18349,N_16315,N_16284);
nor U18350 (N_18350,N_15868,N_15729);
nor U18351 (N_18351,N_16057,N_17626);
xor U18352 (N_18352,N_15294,N_15362);
or U18353 (N_18353,N_15903,N_15339);
nor U18354 (N_18354,N_16620,N_15938);
xor U18355 (N_18355,N_16726,N_17186);
xor U18356 (N_18356,N_15077,N_16232);
xor U18357 (N_18357,N_15061,N_16543);
and U18358 (N_18358,N_17459,N_17211);
nand U18359 (N_18359,N_17487,N_15598);
nand U18360 (N_18360,N_16477,N_15279);
and U18361 (N_18361,N_16854,N_16985);
xor U18362 (N_18362,N_15462,N_16943);
xnor U18363 (N_18363,N_16210,N_16348);
or U18364 (N_18364,N_16177,N_17204);
nor U18365 (N_18365,N_15895,N_15319);
or U18366 (N_18366,N_15107,N_15582);
xor U18367 (N_18367,N_15136,N_17359);
nand U18368 (N_18368,N_15487,N_15499);
nand U18369 (N_18369,N_16386,N_16653);
or U18370 (N_18370,N_15000,N_16504);
and U18371 (N_18371,N_15051,N_15658);
xor U18372 (N_18372,N_17463,N_17329);
or U18373 (N_18373,N_17988,N_17197);
or U18374 (N_18374,N_16343,N_16684);
and U18375 (N_18375,N_17476,N_15762);
nor U18376 (N_18376,N_17240,N_16390);
or U18377 (N_18377,N_15178,N_17011);
xor U18378 (N_18378,N_15345,N_15304);
nand U18379 (N_18379,N_16849,N_16935);
nand U18380 (N_18380,N_15899,N_17646);
nor U18381 (N_18381,N_15571,N_17319);
xnor U18382 (N_18382,N_17438,N_17871);
or U18383 (N_18383,N_15385,N_17636);
and U18384 (N_18384,N_15980,N_16428);
and U18385 (N_18385,N_17932,N_15140);
and U18386 (N_18386,N_17682,N_17762);
or U18387 (N_18387,N_15202,N_16927);
xnor U18388 (N_18388,N_15244,N_15293);
nand U18389 (N_18389,N_17108,N_15043);
xnor U18390 (N_18390,N_17116,N_16963);
and U18391 (N_18391,N_15306,N_15796);
or U18392 (N_18392,N_17028,N_17805);
xnor U18393 (N_18393,N_16008,N_17976);
or U18394 (N_18394,N_15736,N_15101);
or U18395 (N_18395,N_17999,N_17672);
and U18396 (N_18396,N_16568,N_17867);
nor U18397 (N_18397,N_15568,N_17860);
xor U18398 (N_18398,N_15150,N_15901);
or U18399 (N_18399,N_17997,N_15871);
xor U18400 (N_18400,N_15661,N_15715);
nor U18401 (N_18401,N_15015,N_16017);
nand U18402 (N_18402,N_15447,N_16218);
and U18403 (N_18403,N_17586,N_15669);
nand U18404 (N_18404,N_16618,N_16705);
or U18405 (N_18405,N_17922,N_16546);
xor U18406 (N_18406,N_17572,N_16131);
nor U18407 (N_18407,N_17789,N_16652);
or U18408 (N_18408,N_15316,N_16325);
nand U18409 (N_18409,N_16082,N_17859);
nand U18410 (N_18410,N_15498,N_17370);
or U18411 (N_18411,N_15865,N_17953);
nor U18412 (N_18412,N_17630,N_15278);
xor U18413 (N_18413,N_16871,N_15053);
nor U18414 (N_18414,N_15727,N_15717);
or U18415 (N_18415,N_16411,N_15759);
and U18416 (N_18416,N_16059,N_16176);
or U18417 (N_18417,N_15312,N_16824);
nand U18418 (N_18418,N_17526,N_16502);
xor U18419 (N_18419,N_16335,N_16254);
xnor U18420 (N_18420,N_15923,N_16528);
or U18421 (N_18421,N_16487,N_16486);
or U18422 (N_18422,N_17094,N_17704);
nand U18423 (N_18423,N_17622,N_17797);
xor U18424 (N_18424,N_17449,N_15754);
or U18425 (N_18425,N_17002,N_16242);
or U18426 (N_18426,N_16613,N_16279);
or U18427 (N_18427,N_15753,N_17862);
xor U18428 (N_18428,N_15258,N_15672);
and U18429 (N_18429,N_17550,N_16493);
nand U18430 (N_18430,N_16259,N_17544);
or U18431 (N_18431,N_16143,N_17029);
and U18432 (N_18432,N_16262,N_15355);
and U18433 (N_18433,N_16437,N_15326);
or U18434 (N_18434,N_17109,N_16792);
or U18435 (N_18435,N_15198,N_17430);
nand U18436 (N_18436,N_16644,N_15595);
nand U18437 (N_18437,N_17918,N_15432);
xor U18438 (N_18438,N_16072,N_16010);
and U18439 (N_18439,N_15589,N_16181);
nand U18440 (N_18440,N_16624,N_17666);
or U18441 (N_18441,N_17495,N_16483);
and U18442 (N_18442,N_15185,N_17136);
or U18443 (N_18443,N_16853,N_15036);
nand U18444 (N_18444,N_17549,N_16098);
or U18445 (N_18445,N_17040,N_15450);
and U18446 (N_18446,N_17612,N_15490);
nand U18447 (N_18447,N_17558,N_15418);
xnor U18448 (N_18448,N_17305,N_17017);
or U18449 (N_18449,N_16434,N_16430);
nor U18450 (N_18450,N_15932,N_17958);
and U18451 (N_18451,N_15771,N_15562);
and U18452 (N_18452,N_15678,N_17220);
xor U18453 (N_18453,N_16308,N_16874);
and U18454 (N_18454,N_16454,N_15860);
nand U18455 (N_18455,N_15173,N_16703);
xnor U18456 (N_18456,N_17888,N_17609);
nor U18457 (N_18457,N_15265,N_16427);
nor U18458 (N_18458,N_17582,N_15532);
and U18459 (N_18459,N_15473,N_16075);
nor U18460 (N_18460,N_15118,N_16028);
xor U18461 (N_18461,N_15106,N_16902);
and U18462 (N_18462,N_16382,N_16531);
xnor U18463 (N_18463,N_16582,N_16836);
nor U18464 (N_18464,N_15675,N_17552);
xor U18465 (N_18465,N_17208,N_15520);
or U18466 (N_18466,N_17661,N_16955);
xnor U18467 (N_18467,N_17954,N_15653);
nand U18468 (N_18468,N_17766,N_17728);
nor U18469 (N_18469,N_16042,N_16692);
nand U18470 (N_18470,N_17925,N_15849);
nand U18471 (N_18471,N_15438,N_16721);
xnor U18472 (N_18472,N_16600,N_17207);
and U18473 (N_18473,N_17756,N_16192);
nor U18474 (N_18474,N_16203,N_16882);
or U18475 (N_18475,N_16394,N_15080);
nor U18476 (N_18476,N_16019,N_17893);
xor U18477 (N_18477,N_16069,N_15476);
nor U18478 (N_18478,N_15636,N_16731);
xor U18479 (N_18479,N_17708,N_17393);
nand U18480 (N_18480,N_15465,N_17472);
nor U18481 (N_18481,N_17133,N_17978);
nand U18482 (N_18482,N_15618,N_16158);
nor U18483 (N_18483,N_15994,N_16324);
xnor U18484 (N_18484,N_16050,N_17151);
or U18485 (N_18485,N_17723,N_17427);
nand U18486 (N_18486,N_16812,N_17606);
xnor U18487 (N_18487,N_17409,N_15491);
nor U18488 (N_18488,N_17059,N_17524);
xnor U18489 (N_18489,N_16507,N_15510);
xor U18490 (N_18490,N_15311,N_16573);
nand U18491 (N_18491,N_15891,N_15548);
xor U18492 (N_18492,N_15427,N_15767);
xnor U18493 (N_18493,N_17289,N_17389);
nand U18494 (N_18494,N_15743,N_16199);
nor U18495 (N_18495,N_17469,N_15426);
nor U18496 (N_18496,N_17163,N_16783);
and U18497 (N_18497,N_15934,N_16857);
xor U18498 (N_18498,N_15557,N_17421);
and U18499 (N_18499,N_17148,N_16448);
and U18500 (N_18500,N_15839,N_15226);
xnor U18501 (N_18501,N_16969,N_15468);
xnor U18502 (N_18502,N_15553,N_15804);
and U18503 (N_18503,N_15643,N_15690);
and U18504 (N_18504,N_17096,N_15169);
nand U18505 (N_18505,N_15313,N_16035);
nor U18506 (N_18506,N_15203,N_15003);
nand U18507 (N_18507,N_16083,N_17095);
and U18508 (N_18508,N_16763,N_17101);
nand U18509 (N_18509,N_16149,N_16081);
nor U18510 (N_18510,N_15825,N_17522);
xnor U18511 (N_18511,N_15281,N_15361);
nor U18512 (N_18512,N_15755,N_17165);
nand U18513 (N_18513,N_16190,N_17820);
nor U18514 (N_18514,N_16370,N_15235);
or U18515 (N_18515,N_15256,N_17974);
xor U18516 (N_18516,N_16974,N_17052);
nor U18517 (N_18517,N_16741,N_17512);
and U18518 (N_18518,N_16892,N_17445);
nor U18519 (N_18519,N_17118,N_16978);
nand U18520 (N_18520,N_15719,N_17948);
nand U18521 (N_18521,N_17340,N_17685);
or U18522 (N_18522,N_15848,N_16361);
xor U18523 (N_18523,N_17306,N_15386);
and U18524 (N_18524,N_16263,N_17226);
and U18525 (N_18525,N_16938,N_16205);
or U18526 (N_18526,N_17681,N_16878);
nand U18527 (N_18527,N_17390,N_16230);
nand U18528 (N_18528,N_17157,N_15604);
xor U18529 (N_18529,N_17837,N_15129);
nor U18530 (N_18530,N_15099,N_16887);
and U18531 (N_18531,N_15058,N_15701);
nand U18532 (N_18532,N_15723,N_16580);
xor U18533 (N_18533,N_16597,N_16120);
and U18534 (N_18534,N_17066,N_15193);
or U18535 (N_18535,N_15111,N_15138);
xor U18536 (N_18536,N_17786,N_15283);
xor U18537 (N_18537,N_15277,N_17580);
or U18538 (N_18538,N_16640,N_17625);
and U18539 (N_18539,N_17004,N_17569);
xnor U18540 (N_18540,N_16619,N_17941);
nand U18541 (N_18541,N_17745,N_16813);
and U18542 (N_18542,N_16346,N_16522);
xor U18543 (N_18543,N_17105,N_15119);
or U18544 (N_18544,N_16479,N_16903);
nand U18545 (N_18545,N_17354,N_16740);
nor U18546 (N_18546,N_17425,N_15855);
and U18547 (N_18547,N_16952,N_15894);
and U18548 (N_18548,N_15698,N_16567);
xor U18549 (N_18549,N_16676,N_17674);
nand U18550 (N_18550,N_15401,N_16341);
nand U18551 (N_18551,N_17365,N_17061);
or U18552 (N_18552,N_17802,N_16220);
nand U18553 (N_18553,N_15774,N_15123);
or U18554 (N_18554,N_16445,N_15929);
nand U18555 (N_18555,N_16718,N_15434);
nor U18556 (N_18556,N_16962,N_15732);
or U18557 (N_18557,N_15816,N_15086);
or U18558 (N_18558,N_15013,N_17989);
nor U18559 (N_18559,N_15374,N_15770);
xor U18560 (N_18560,N_17266,N_15834);
xor U18561 (N_18561,N_16089,N_15802);
and U18562 (N_18562,N_16816,N_15946);
nand U18563 (N_18563,N_16144,N_16195);
nand U18564 (N_18564,N_17591,N_16171);
nand U18565 (N_18565,N_17262,N_15654);
nand U18566 (N_18566,N_16539,N_15179);
nand U18567 (N_18567,N_16077,N_15264);
nor U18568 (N_18568,N_16638,N_17435);
or U18569 (N_18569,N_16130,N_16164);
or U18570 (N_18570,N_15703,N_15694);
nor U18571 (N_18571,N_17001,N_15437);
or U18572 (N_18572,N_16369,N_15020);
and U18573 (N_18573,N_15534,N_17046);
xor U18574 (N_18574,N_15708,N_17631);
or U18575 (N_18575,N_16005,N_16782);
xor U18576 (N_18576,N_15859,N_16285);
and U18577 (N_18577,N_15454,N_15693);
nand U18578 (N_18578,N_17082,N_17492);
and U18579 (N_18579,N_16716,N_15982);
and U18580 (N_18580,N_15228,N_16068);
and U18581 (N_18581,N_16986,N_16524);
and U18582 (N_18582,N_17416,N_16622);
nand U18583 (N_18583,N_15500,N_16779);
or U18584 (N_18584,N_15105,N_17811);
or U18585 (N_18585,N_17458,N_15600);
or U18586 (N_18586,N_17454,N_16748);
xor U18587 (N_18587,N_16376,N_17857);
or U18588 (N_18588,N_16908,N_17350);
nand U18589 (N_18589,N_17282,N_15522);
xor U18590 (N_18590,N_16517,N_16043);
xor U18591 (N_18591,N_15034,N_15792);
or U18592 (N_18592,N_17881,N_16045);
or U18593 (N_18593,N_17633,N_15446);
nor U18594 (N_18594,N_16141,N_16099);
and U18595 (N_18595,N_16988,N_15780);
nor U18596 (N_18596,N_17764,N_15814);
and U18597 (N_18597,N_16194,N_15565);
or U18598 (N_18598,N_15866,N_17695);
xor U18599 (N_18599,N_15455,N_15266);
and U18600 (N_18600,N_16174,N_17331);
nand U18601 (N_18601,N_15996,N_16215);
nand U18602 (N_18602,N_16079,N_15113);
nor U18603 (N_18603,N_16281,N_17439);
nand U18604 (N_18604,N_16404,N_16697);
nor U18605 (N_18605,N_17651,N_17024);
or U18606 (N_18606,N_15002,N_16433);
or U18607 (N_18607,N_17812,N_15869);
nand U18608 (N_18608,N_15552,N_15232);
nand U18609 (N_18609,N_17641,N_17690);
xor U18610 (N_18610,N_15234,N_17570);
nor U18611 (N_18611,N_17057,N_17561);
or U18612 (N_18612,N_16395,N_15769);
and U18613 (N_18613,N_16772,N_17081);
nor U18614 (N_18614,N_16511,N_16431);
nor U18615 (N_18615,N_16021,N_17352);
xor U18616 (N_18616,N_15222,N_16316);
nand U18617 (N_18617,N_16788,N_15613);
nand U18618 (N_18618,N_16798,N_15731);
xor U18619 (N_18619,N_17249,N_17559);
or U18620 (N_18620,N_16723,N_16474);
nand U18621 (N_18621,N_17489,N_17594);
xor U18622 (N_18622,N_16163,N_17834);
nand U18623 (N_18623,N_16565,N_17754);
xor U18624 (N_18624,N_16066,N_15342);
nand U18625 (N_18625,N_17358,N_16475);
and U18626 (N_18626,N_15165,N_16182);
nor U18627 (N_18627,N_17296,N_15208);
nand U18628 (N_18628,N_15603,N_16356);
and U18629 (N_18629,N_17725,N_16012);
and U18630 (N_18630,N_16826,N_17599);
or U18631 (N_18631,N_15405,N_15415);
nor U18632 (N_18632,N_17371,N_15213);
and U18633 (N_18633,N_15042,N_17985);
xor U18634 (N_18634,N_16665,N_17112);
and U18635 (N_18635,N_16397,N_16521);
xor U18636 (N_18636,N_15216,N_16037);
and U18637 (N_18637,N_15927,N_16818);
nand U18638 (N_18638,N_17887,N_16572);
and U18639 (N_18639,N_17803,N_17064);
nand U18640 (N_18640,N_15246,N_17772);
nand U18641 (N_18641,N_16586,N_16123);
xnor U18642 (N_18642,N_15484,N_16617);
or U18643 (N_18643,N_15943,N_17553);
and U18644 (N_18644,N_15259,N_16863);
and U18645 (N_18645,N_16538,N_16574);
or U18646 (N_18646,N_15384,N_17049);
and U18647 (N_18647,N_17724,N_16076);
or U18648 (N_18648,N_15243,N_15558);
and U18649 (N_18649,N_16900,N_15480);
xnor U18650 (N_18650,N_16593,N_17295);
xor U18651 (N_18651,N_17457,N_15697);
and U18652 (N_18652,N_16881,N_15388);
nor U18653 (N_18653,N_16168,N_16375);
xnor U18654 (N_18654,N_16630,N_15270);
and U18655 (N_18655,N_17813,N_16736);
nand U18656 (N_18656,N_17833,N_15095);
and U18657 (N_18657,N_16287,N_16312);
xor U18658 (N_18658,N_17210,N_17158);
nor U18659 (N_18659,N_15944,N_16385);
nor U18660 (N_18660,N_15184,N_15721);
xor U18661 (N_18661,N_16576,N_15067);
nand U18662 (N_18662,N_16393,N_16026);
xnor U18663 (N_18663,N_17904,N_15502);
or U18664 (N_18664,N_17145,N_15810);
or U18665 (N_18665,N_16656,N_17307);
nor U18666 (N_18666,N_17250,N_16760);
xor U18667 (N_18667,N_16139,N_16344);
and U18668 (N_18668,N_15696,N_16024);
nor U18669 (N_18669,N_16685,N_17174);
xor U18670 (N_18670,N_16133,N_15424);
nor U18671 (N_18671,N_15517,N_17124);
nand U18672 (N_18672,N_17779,N_17310);
nor U18673 (N_18673,N_17852,N_17509);
or U18674 (N_18674,N_15528,N_17935);
xnor U18675 (N_18675,N_16255,N_15662);
nor U18676 (N_18676,N_17376,N_16889);
and U18677 (N_18677,N_17749,N_16605);
nand U18678 (N_18678,N_15811,N_17799);
and U18679 (N_18679,N_17253,N_15893);
nor U18680 (N_18680,N_17621,N_16489);
and U18681 (N_18681,N_16720,N_17137);
or U18682 (N_18682,N_16829,N_15768);
xor U18683 (N_18683,N_15820,N_16601);
nor U18684 (N_18684,N_17268,N_15599);
xor U18685 (N_18685,N_15154,N_17926);
nor U18686 (N_18686,N_17537,N_16333);
nor U18687 (N_18687,N_17368,N_17321);
nor U18688 (N_18688,N_15738,N_16928);
or U18689 (N_18689,N_15864,N_16213);
nor U18690 (N_18690,N_17106,N_17324);
nor U18691 (N_18691,N_15392,N_16958);
nor U18692 (N_18692,N_16956,N_16587);
and U18693 (N_18693,N_15630,N_16801);
or U18694 (N_18694,N_17794,N_17778);
xnor U18695 (N_18695,N_15615,N_16562);
nor U18696 (N_18696,N_16852,N_17026);
or U18697 (N_18697,N_15383,N_17264);
xnor U18698 (N_18698,N_17298,N_16918);
and U18699 (N_18699,N_15555,N_16585);
nor U18700 (N_18700,N_16767,N_17474);
or U18701 (N_18701,N_16628,N_15433);
and U18702 (N_18702,N_16080,N_17665);
nand U18703 (N_18703,N_16508,N_16053);
xor U18704 (N_18704,N_17515,N_17715);
nand U18705 (N_18705,N_16693,N_17716);
and U18706 (N_18706,N_15607,N_15006);
or U18707 (N_18707,N_15874,N_15214);
or U18708 (N_18708,N_15132,N_17429);
nand U18709 (N_18709,N_16730,N_15835);
and U18710 (N_18710,N_15507,N_15352);
nand U18711 (N_18711,N_16877,N_15207);
and U18712 (N_18712,N_17247,N_16007);
nand U18713 (N_18713,N_16468,N_15254);
xor U18714 (N_18714,N_16862,N_17265);
xnor U18715 (N_18715,N_17949,N_16249);
xor U18716 (N_18716,N_17387,N_16743);
xnor U18717 (N_18717,N_17005,N_17333);
or U18718 (N_18718,N_17027,N_17783);
xnor U18719 (N_18719,N_17156,N_16349);
nand U18720 (N_18720,N_17910,N_15408);
nand U18721 (N_18721,N_17031,N_16768);
nor U18722 (N_18722,N_17920,N_15745);
nand U18723 (N_18723,N_15292,N_17394);
or U18724 (N_18724,N_15076,N_15358);
or U18725 (N_18725,N_16728,N_17008);
nor U18726 (N_18726,N_17655,N_15224);
or U18727 (N_18727,N_17850,N_17841);
or U18728 (N_18728,N_17616,N_16765);
nand U18729 (N_18729,N_16134,N_15227);
nand U18730 (N_18730,N_17130,N_16982);
xnor U18731 (N_18731,N_16441,N_16951);
nor U18732 (N_18732,N_15789,N_15335);
xnor U18733 (N_18733,N_17528,N_16110);
nand U18734 (N_18734,N_16791,N_15756);
or U18735 (N_18735,N_17022,N_15504);
and U18736 (N_18736,N_15242,N_16534);
nand U18737 (N_18737,N_15038,N_17525);
or U18738 (N_18738,N_16301,N_17642);
or U18739 (N_18739,N_16360,N_15883);
xnor U18740 (N_18740,N_16290,N_15937);
nor U18741 (N_18741,N_15593,N_15340);
and U18742 (N_18742,N_15606,N_15714);
xnor U18743 (N_18743,N_17281,N_15882);
or U18744 (N_18744,N_15914,N_16571);
nand U18745 (N_18745,N_16753,N_16913);
nor U18746 (N_18746,N_16712,N_17643);
and U18747 (N_18747,N_15799,N_17824);
and U18748 (N_18748,N_17909,N_15556);
xor U18749 (N_18749,N_17316,N_15289);
and U18750 (N_18750,N_15469,N_15852);
and U18751 (N_18751,N_17448,N_15917);
or U18752 (N_18752,N_16785,N_16446);
and U18753 (N_18753,N_16020,N_17707);
or U18754 (N_18754,N_16458,N_16738);
and U18755 (N_18755,N_17209,N_17901);
nor U18756 (N_18756,N_17099,N_15542);
and U18757 (N_18757,N_15050,N_15486);
nor U18758 (N_18758,N_15546,N_16260);
or U18759 (N_18759,N_17620,N_17656);
nor U18760 (N_18760,N_15257,N_16113);
and U18761 (N_18761,N_17598,N_16293);
xnor U18762 (N_18762,N_15559,N_17624);
and U18763 (N_18763,N_16097,N_17911);
or U18764 (N_18764,N_16412,N_15220);
or U18765 (N_18765,N_16807,N_17069);
nand U18766 (N_18766,N_15638,N_16054);
nor U18767 (N_18767,N_15668,N_16271);
nor U18768 (N_18768,N_16368,N_15915);
nor U18769 (N_18769,N_16184,N_15726);
nand U18770 (N_18770,N_16930,N_17479);
and U18771 (N_18771,N_17796,N_16840);
or U18772 (N_18772,N_15900,N_17032);
xor U18773 (N_18773,N_15445,N_16183);
and U18774 (N_18774,N_17294,N_17623);
or U18775 (N_18775,N_15420,N_16410);
xnor U18776 (N_18776,N_15902,N_17498);
nor U18777 (N_18777,N_15527,N_16924);
nand U18778 (N_18778,N_15563,N_15942);
nor U18779 (N_18779,N_16946,N_17602);
nor U18780 (N_18780,N_16052,N_16701);
or U18781 (N_18781,N_15413,N_17313);
xor U18782 (N_18782,N_16074,N_16207);
and U18783 (N_18783,N_17328,N_17883);
and U18784 (N_18784,N_15019,N_16200);
nand U18785 (N_18785,N_16014,N_16695);
nor U18786 (N_18786,N_15396,N_16709);
xor U18787 (N_18787,N_16118,N_16039);
nor U18788 (N_18788,N_17649,N_17554);
or U18789 (N_18789,N_16964,N_16036);
nand U18790 (N_18790,N_16674,N_17213);
nor U18791 (N_18791,N_17410,N_15016);
and U18792 (N_18792,N_15470,N_15823);
xor U18793 (N_18793,N_16222,N_17565);
or U18794 (N_18794,N_16714,N_17595);
nand U18795 (N_18795,N_17097,N_17966);
xnor U18796 (N_18796,N_17996,N_15397);
nor U18797 (N_18797,N_15640,N_16436);
xor U18798 (N_18798,N_16876,N_17983);
nor U18799 (N_18799,N_17693,N_16983);
nor U18800 (N_18800,N_17270,N_17424);
or U18801 (N_18801,N_15966,N_15627);
or U18802 (N_18802,N_15124,N_17927);
nand U18803 (N_18803,N_15381,N_15592);
and U18804 (N_18804,N_16328,N_15506);
xor U18805 (N_18805,N_17518,N_17667);
and U18806 (N_18806,N_16633,N_17497);
nor U18807 (N_18807,N_16093,N_15564);
or U18808 (N_18808,N_15189,N_17245);
nand U18809 (N_18809,N_15676,N_16602);
xnor U18810 (N_18810,N_15935,N_15237);
and U18811 (N_18811,N_16675,N_17168);
nor U18812 (N_18812,N_15518,N_17600);
nor U18813 (N_18813,N_16481,N_17658);
nor U18814 (N_18814,N_16473,N_15337);
nand U18815 (N_18815,N_15460,N_15617);
xor U18816 (N_18816,N_17395,N_15082);
xor U18817 (N_18817,N_15873,N_16895);
and U18818 (N_18818,N_16478,N_17473);
nor U18819 (N_18819,N_17873,N_16403);
xnor U18820 (N_18820,N_17513,N_15560);
xnor U18821 (N_18821,N_15790,N_17256);
and U18822 (N_18822,N_17683,N_17462);
xnor U18823 (N_18823,N_17973,N_15524);
xor U18824 (N_18824,N_15158,N_16532);
nor U18825 (N_18825,N_16609,N_15161);
nand U18826 (N_18826,N_16762,N_16060);
nand U18827 (N_18827,N_16379,N_16273);
nand U18828 (N_18828,N_17699,N_17615);
xnor U18829 (N_18829,N_17767,N_16503);
and U18830 (N_18830,N_15390,N_17219);
xor U18831 (N_18831,N_15090,N_17654);
nand U18832 (N_18832,N_15239,N_16371);
xor U18833 (N_18833,N_16246,N_17678);
and U18834 (N_18834,N_16048,N_17912);
nand U18835 (N_18835,N_15824,N_15176);
or U18836 (N_18836,N_15635,N_17596);
or U18837 (N_18837,N_16657,N_17451);
nand U18838 (N_18838,N_16256,N_17614);
and U18839 (N_18839,N_16138,N_17317);
and U18840 (N_18840,N_17934,N_16311);
or U18841 (N_18841,N_17257,N_17347);
or U18842 (N_18842,N_15451,N_15494);
nor U18843 (N_18843,N_15147,N_15785);
xnor U18844 (N_18844,N_17869,N_17774);
nand U18845 (N_18845,N_16408,N_16575);
xor U18846 (N_18846,N_17791,N_15144);
or U18847 (N_18847,N_15704,N_17044);
and U18848 (N_18848,N_17828,N_15924);
nor U18849 (N_18849,N_16303,N_17276);
or U18850 (N_18850,N_17968,N_16513);
nand U18851 (N_18851,N_15505,N_15888);
nand U18852 (N_18852,N_16708,N_15887);
nand U18853 (N_18853,N_15489,N_17087);
xnor U18854 (N_18854,N_16944,N_17452);
and U18855 (N_18855,N_17129,N_15321);
or U18856 (N_18856,N_16238,N_15550);
and U18857 (N_18857,N_16219,N_15845);
nand U18858 (N_18858,N_16561,N_15539);
or U18859 (N_18859,N_16309,N_16006);
nor U18860 (N_18860,N_15218,N_17285);
and U18861 (N_18861,N_16839,N_15139);
or U18862 (N_18862,N_17639,N_15425);
nand U18863 (N_18863,N_15970,N_15781);
and U18864 (N_18864,N_15377,N_15969);
or U18865 (N_18865,N_15127,N_17530);
and U18866 (N_18866,N_16608,N_15707);
or U18867 (N_18867,N_15836,N_17198);
and U18868 (N_18868,N_15435,N_15241);
nor U18869 (N_18869,N_16373,N_17277);
nand U18870 (N_18870,N_15341,N_16627);
or U18871 (N_18871,N_15875,N_15905);
nand U18872 (N_18872,N_15906,N_16156);
xor U18873 (N_18873,N_17845,N_16642);
xnor U18874 (N_18874,N_17251,N_17490);
nand U18875 (N_18875,N_17388,N_17743);
xnor U18876 (N_18876,N_15143,N_16905);
nand U18877 (N_18877,N_16105,N_17131);
xnor U18878 (N_18878,N_17248,N_16063);
xnor U18879 (N_18879,N_17752,N_17121);
nand U18880 (N_18880,N_15920,N_15069);
nor U18881 (N_18881,N_16896,N_15821);
nor U18882 (N_18882,N_15974,N_17880);
nand U18883 (N_18883,N_15925,N_15269);
nand U18884 (N_18884,N_15191,N_17523);
xor U18885 (N_18885,N_17237,N_17045);
nor U18886 (N_18886,N_16805,N_16178);
or U18887 (N_18887,N_15419,N_16117);
and U18888 (N_18888,N_16425,N_16936);
nand U18889 (N_18889,N_16032,N_16611);
nand U18890 (N_18890,N_16179,N_17089);
nand U18891 (N_18891,N_15116,N_17900);
or U18892 (N_18892,N_17332,N_17502);
and U18893 (N_18893,N_15503,N_16941);
and U18894 (N_18894,N_16084,N_16338);
xor U18895 (N_18895,N_16276,N_16906);
nand U18896 (N_18896,N_17326,N_15922);
xor U18897 (N_18897,N_17437,N_15761);
or U18898 (N_18898,N_17545,N_17166);
and U18899 (N_18899,N_17777,N_15496);
and U18900 (N_18900,N_16592,N_15428);
nand U18901 (N_18901,N_15411,N_15588);
xnor U18902 (N_18902,N_17982,N_16515);
nor U18903 (N_18903,N_16267,N_16557);
and U18904 (N_18904,N_15162,N_16329);
and U18905 (N_18905,N_16122,N_15223);
xnor U18906 (N_18906,N_15911,N_17680);
nor U18907 (N_18907,N_17647,N_16124);
nand U18908 (N_18908,N_16781,N_15632);
nor U18909 (N_18909,N_15940,N_16595);
or U18910 (N_18910,N_15718,N_16090);
or U18911 (N_18911,N_15330,N_15574);
nand U18912 (N_18912,N_16055,N_17501);
or U18913 (N_18913,N_17258,N_17073);
nor U18914 (N_18914,N_16241,N_15987);
nand U18915 (N_18915,N_16590,N_16472);
and U18916 (N_18916,N_16848,N_17891);
or U18917 (N_18917,N_17815,N_16034);
and U18918 (N_18918,N_17875,N_17962);
or U18919 (N_18919,N_17444,N_15054);
nand U18920 (N_18920,N_15786,N_15913);
xor U18921 (N_18921,N_17668,N_15164);
or U18922 (N_18922,N_16206,N_15679);
or U18923 (N_18923,N_15421,N_17984);
nand U18924 (N_18924,N_16160,N_16950);
nand U18925 (N_18925,N_15398,N_15364);
xor U18926 (N_18926,N_15889,N_17173);
or U18927 (N_18927,N_16939,N_15700);
or U18928 (N_18928,N_16770,N_15181);
and U18929 (N_18929,N_17034,N_16819);
and U18930 (N_18930,N_17753,N_16755);
or U18931 (N_18931,N_16025,N_15060);
or U18932 (N_18932,N_15763,N_16064);
and U18933 (N_18933,N_15807,N_16578);
or U18934 (N_18934,N_16636,N_15260);
and U18935 (N_18935,N_15941,N_15725);
xnor U18936 (N_18936,N_16520,N_17597);
xnor U18937 (N_18937,N_17385,N_17890);
and U18938 (N_18938,N_15622,N_16842);
xor U18939 (N_18939,N_17484,N_15255);
and U18940 (N_18940,N_17955,N_17323);
xor U18941 (N_18941,N_17377,N_16975);
and U18942 (N_18942,N_16835,N_16560);
or U18943 (N_18943,N_17687,N_15064);
xor U18944 (N_18944,N_16423,N_15818);
nor U18945 (N_18945,N_15471,N_15089);
and U18946 (N_18946,N_16911,N_16754);
nor U18947 (N_18947,N_17843,N_16879);
nand U18948 (N_18948,N_15547,N_16253);
xor U18949 (N_18949,N_15325,N_16569);
or U18950 (N_18950,N_15151,N_17290);
nand U18951 (N_18951,N_17562,N_17792);
nor U18952 (N_18952,N_16166,N_16198);
nand U18953 (N_18953,N_16461,N_17659);
or U18954 (N_18954,N_16802,N_17640);
xnor U18955 (N_18955,N_17325,N_16047);
or U18956 (N_18956,N_15382,N_16291);
nor U18957 (N_18957,N_15205,N_17589);
nor U18958 (N_18958,N_17677,N_15540);
nand U18959 (N_18959,N_16722,N_15876);
and U18960 (N_18960,N_17738,N_17058);
or U18961 (N_18961,N_15960,N_17838);
or U18962 (N_18962,N_15448,N_15918);
xor U18963 (N_18963,N_15156,N_15368);
or U18964 (N_18964,N_16332,N_15192);
nand U18965 (N_18965,N_15300,N_16867);
and U18966 (N_18966,N_16632,N_17853);
nand U18967 (N_18967,N_16239,N_15369);
or U18968 (N_18968,N_17913,N_16667);
and U18969 (N_18969,N_17817,N_15155);
nor U18970 (N_18970,N_17135,N_16196);
xnor U18971 (N_18971,N_15298,N_16011);
and U18972 (N_18972,N_15195,N_17945);
nand U18973 (N_18973,N_17142,N_15508);
nor U18974 (N_18974,N_15734,N_17170);
nand U18975 (N_18975,N_16439,N_17477);
nand U18976 (N_18976,N_16683,N_16514);
xor U18977 (N_18977,N_16384,N_17372);
nor U18978 (N_18978,N_15526,N_16161);
nor U18979 (N_18979,N_16299,N_17947);
and U18980 (N_18980,N_15349,N_15354);
nor U18981 (N_18981,N_16467,N_17171);
nor U18982 (N_18982,N_17835,N_17928);
or U18983 (N_18983,N_17093,N_17846);
xnor U18984 (N_18984,N_15989,N_16224);
xor U18985 (N_18985,N_15907,N_17801);
nand U18986 (N_18986,N_15686,N_15513);
or U18987 (N_18987,N_16388,N_16277);
nor U18988 (N_18988,N_15186,N_15685);
or U18989 (N_18989,N_15806,N_15822);
or U18990 (N_18990,N_17771,N_15372);
and U18991 (N_18991,N_17679,N_15536);
nor U18992 (N_18992,N_17923,N_17013);
and U18993 (N_18993,N_16629,N_16607);
xor U18994 (N_18994,N_15240,N_15007);
nor U18995 (N_18995,N_17239,N_17686);
and U18996 (N_18996,N_17338,N_17272);
nand U18997 (N_18997,N_17539,N_16830);
or U18998 (N_18998,N_16823,N_17701);
or U18999 (N_18999,N_16594,N_16300);
xnor U19000 (N_19000,N_16327,N_16223);
or U19001 (N_19001,N_16067,N_15477);
nand U19002 (N_19002,N_15047,N_16993);
nand U19003 (N_19003,N_16706,N_15794);
nand U19004 (N_19004,N_16235,N_16237);
nor U19005 (N_19005,N_15628,N_16336);
or U19006 (N_19006,N_17110,N_15856);
xor U19007 (N_19007,N_15290,N_16832);
nand U19008 (N_19008,N_16899,N_16825);
or U19009 (N_19009,N_15629,N_16506);
nand U19010 (N_19010,N_17671,N_17090);
nand U19011 (N_19011,N_15098,N_15965);
nor U19012 (N_19012,N_17840,N_17360);
nand U19013 (N_19013,N_16971,N_16491);
and U19014 (N_19014,N_15609,N_15453);
and U19015 (N_19015,N_17000,N_16931);
nor U19016 (N_19016,N_16533,N_17644);
xnor U19017 (N_19017,N_17965,N_15784);
xnor U19018 (N_19018,N_15441,N_16000);
nor U19019 (N_19019,N_17744,N_16898);
and U19020 (N_19020,N_17607,N_17246);
xor U19021 (N_19021,N_16153,N_16495);
xor U19022 (N_19022,N_16257,N_16167);
nand U19023 (N_19023,N_15452,N_17575);
or U19024 (N_19024,N_16272,N_15961);
nand U19025 (N_19025,N_15456,N_15461);
xnor U19026 (N_19026,N_17719,N_17706);
xnor U19027 (N_19027,N_16704,N_17581);
and U19028 (N_19028,N_15744,N_17874);
nor U19029 (N_19029,N_15049,N_16202);
or U19030 (N_19030,N_16350,N_15440);
and U19031 (N_19031,N_17829,N_15322);
nand U19032 (N_19032,N_16919,N_17592);
and U19033 (N_19033,N_15365,N_16957);
or U19034 (N_19034,N_16322,N_17848);
xor U19035 (N_19035,N_16319,N_15017);
xor U19036 (N_19036,N_16041,N_15271);
nor U19037 (N_19037,N_17741,N_17995);
nor U19038 (N_19038,N_16121,N_16137);
and U19039 (N_19039,N_17851,N_16288);
nand U19040 (N_19040,N_16465,N_15872);
xnor U19041 (N_19041,N_15585,N_15079);
xor U19042 (N_19042,N_15608,N_17025);
nand U19043 (N_19043,N_15175,N_15854);
and U19044 (N_19044,N_17414,N_15648);
nand U19045 (N_19045,N_16610,N_16351);
xnor U19046 (N_19046,N_17584,N_17748);
and U19047 (N_19047,N_17638,N_15431);
and U19048 (N_19048,N_16451,N_17940);
nand U19049 (N_19049,N_16413,N_16909);
xor U19050 (N_19050,N_17894,N_17628);
xor U19051 (N_19051,N_15072,N_15229);
xnor U19052 (N_19052,N_15018,N_15081);
xor U19053 (N_19053,N_16682,N_15133);
xnor U19054 (N_19054,N_16482,N_16155);
xnor U19055 (N_19055,N_16820,N_15212);
or U19056 (N_19056,N_16424,N_15765);
xnor U19057 (N_19057,N_17714,N_17907);
or U19058 (N_19058,N_17747,N_16666);
nand U19059 (N_19059,N_16126,N_15642);
and U19060 (N_19060,N_16251,N_15055);
and U19061 (N_19061,N_17146,N_16525);
nor U19062 (N_19062,N_17603,N_17711);
and U19063 (N_19063,N_16639,N_17800);
nor U19064 (N_19064,N_17039,N_16880);
and U19065 (N_19065,N_17500,N_15581);
xnor U19066 (N_19066,N_15261,N_16058);
or U19067 (N_19067,N_16310,N_16298);
nand U19068 (N_19068,N_15314,N_17938);
xnor U19069 (N_19069,N_17364,N_16414);
xor U19070 (N_19070,N_15183,N_15634);
nor U19071 (N_19071,N_15172,N_16302);
and U19072 (N_19072,N_17339,N_17287);
xnor U19073 (N_19073,N_15221,N_15760);
or U19074 (N_19074,N_15877,N_15373);
or U19075 (N_19075,N_15977,N_17203);
and U19076 (N_19076,N_17189,N_15509);
xnor U19077 (N_19077,N_16634,N_15967);
xor U19078 (N_19078,N_16530,N_15174);
xor U19079 (N_19079,N_17886,N_15750);
or U19080 (N_19080,N_16987,N_17849);
nor U19081 (N_19081,N_16459,N_17422);
nor U19082 (N_19082,N_17657,N_16102);
xor U19083 (N_19083,N_15647,N_17228);
or U19084 (N_19084,N_17583,N_16917);
nor U19085 (N_19085,N_16438,N_16606);
and U19086 (N_19086,N_16545,N_15168);
or U19087 (N_19087,N_15549,N_17696);
nor U19088 (N_19088,N_16612,N_16796);
nor U19089 (N_19089,N_16148,N_15870);
nand U19090 (N_19090,N_15366,N_17336);
or U19091 (N_19091,N_16497,N_15010);
nor U19092 (N_19092,N_15649,N_15958);
nor U19093 (N_19093,N_15981,N_17844);
xnor U19094 (N_19094,N_15273,N_15409);
xor U19095 (N_19095,N_17736,N_16850);
and U19096 (N_19096,N_15093,N_16655);
xor U19097 (N_19097,N_16689,N_17542);
nor U19098 (N_19098,N_15879,N_16391);
and U19099 (N_19099,N_15444,N_17866);
or U19100 (N_19100,N_15120,N_16616);
and U19101 (N_19101,N_15074,N_15748);
nand U19102 (N_19102,N_17585,N_16374);
and U19103 (N_19103,N_15206,N_17993);
nand U19104 (N_19104,N_16949,N_15712);
nand U19105 (N_19105,N_15863,N_15783);
or U19106 (N_19106,N_16416,N_15880);
xor U19107 (N_19107,N_16078,N_15134);
or U19108 (N_19108,N_17431,N_16873);
nor U19109 (N_19109,N_16087,N_17346);
or U19110 (N_19110,N_15495,N_15919);
xnor U19111 (N_19111,N_17304,N_17123);
or U19112 (N_19112,N_16654,N_17899);
nor U19113 (N_19113,N_17232,N_17267);
and U19114 (N_19114,N_17020,N_17810);
and U19115 (N_19115,N_15302,N_17300);
nand U19116 (N_19116,N_17826,N_15275);
nor U19117 (N_19117,N_15073,N_15037);
xnor U19118 (N_19118,N_15370,N_16699);
xnor U19119 (N_19119,N_15787,N_15631);
xor U19120 (N_19120,N_16838,N_17086);
or U19121 (N_19121,N_15291,N_15171);
nand U19122 (N_19122,N_16231,N_16270);
xnor U19123 (N_19123,N_17956,N_16331);
nand U19124 (N_19124,N_17280,N_17104);
and U19125 (N_19125,N_17915,N_17054);
xnor U19126 (N_19126,N_16923,N_17632);
nand U19127 (N_19127,N_16294,N_17269);
xnor U19128 (N_19128,N_17464,N_16002);
and U19129 (N_19129,N_15993,N_17885);
and U19130 (N_19130,N_16536,N_15724);
xnor U19131 (N_19131,N_15182,N_16890);
xor U19132 (N_19132,N_17946,N_16426);
or U19133 (N_19133,N_15583,N_15475);
or U19134 (N_19134,N_15483,N_16258);
nor U19135 (N_19135,N_15928,N_15022);
and U19136 (N_19136,N_16915,N_16834);
xor U19137 (N_19137,N_17322,N_15199);
nor U19138 (N_19138,N_15351,N_17807);
nor U19139 (N_19139,N_17669,N_17442);
and U19140 (N_19140,N_15236,N_17573);
nand U19141 (N_19141,N_17292,N_17102);
nand U19142 (N_19142,N_15625,N_15720);
or U19143 (N_19143,N_16100,N_16803);
nand U19144 (N_19144,N_16286,N_17540);
nand U19145 (N_19145,N_16526,N_16547);
or U19146 (N_19146,N_17413,N_15268);
xor U19147 (N_19147,N_17692,N_17405);
or U19148 (N_19148,N_15610,N_17770);
nand U19149 (N_19149,N_17963,N_16396);
and U19150 (N_19150,N_17349,N_17990);
nand U19151 (N_19151,N_16998,N_17547);
nand U19152 (N_19152,N_17278,N_17610);
or U19153 (N_19153,N_15554,N_16968);
nand U19154 (N_19154,N_16378,N_17551);
xor U19155 (N_19155,N_15170,N_17230);
or U19156 (N_19156,N_15705,N_15238);
and U19157 (N_19157,N_16463,N_15439);
or U19158 (N_19158,N_16217,N_17534);
nand U19159 (N_19159,N_16119,N_15492);
nand U19160 (N_19160,N_15102,N_16670);
nand U19161 (N_19161,N_15282,N_16860);
xor U19162 (N_19162,N_16366,N_15230);
xor U19163 (N_19163,N_17831,N_15308);
nand U19164 (N_19164,N_16471,N_15947);
nor U19165 (N_19165,N_15655,N_17212);
nor U19166 (N_19166,N_16435,N_17367);
or U19167 (N_19167,N_17952,N_15497);
nor U19168 (N_19168,N_17700,N_17830);
nor U19169 (N_19169,N_15684,N_15057);
xnor U19170 (N_19170,N_16631,N_15267);
and U19171 (N_19171,N_16984,N_16509);
or U19172 (N_19172,N_17455,N_17235);
or U19173 (N_19173,N_16757,N_15285);
xnor U19174 (N_19174,N_16960,N_15722);
and U19175 (N_19175,N_17252,N_17863);
nor U19176 (N_19176,N_15334,N_17392);
nor U19177 (N_19177,N_17223,N_16065);
or U19178 (N_19178,N_17877,N_17698);
xnor U19179 (N_19179,N_16926,N_17864);
nand U19180 (N_19180,N_15035,N_17447);
nor U19181 (N_19181,N_15843,N_16761);
nor U19182 (N_19182,N_16837,N_17975);
or U19183 (N_19183,N_15115,N_17977);
and U19184 (N_19184,N_15601,N_15737);
xnor U19185 (N_19185,N_16841,N_16742);
or U19186 (N_19186,N_16498,N_17379);
and U19187 (N_19187,N_15092,N_17100);
nand U19188 (N_19188,N_16795,N_16793);
nand U19189 (N_19189,N_17169,N_17126);
nand U19190 (N_19190,N_16559,N_16727);
nand U19191 (N_19191,N_17465,N_15682);
nand U19192 (N_19192,N_17532,N_17147);
nor U19193 (N_19193,N_16266,N_17412);
xor U19194 (N_19194,N_17564,N_16022);
or U19195 (N_19195,N_15125,N_15976);
or U19196 (N_19196,N_15274,N_15850);
or U19197 (N_19197,N_17739,N_15990);
nor U19198 (N_19198,N_17183,N_16672);
nand U19199 (N_19199,N_16466,N_16318);
and U19200 (N_19200,N_16420,N_15515);
and U19201 (N_19201,N_17441,N_15992);
xor U19202 (N_19202,N_16357,N_15097);
xor U19203 (N_19203,N_15573,N_15280);
or U19204 (N_19204,N_17507,N_16188);
nor U19205 (N_19205,N_16264,N_16125);
nor U19206 (N_19206,N_15665,N_17167);
and U19207 (N_19207,N_17832,N_15741);
or U19208 (N_19208,N_17689,N_16488);
or U19209 (N_19209,N_15983,N_15641);
nor U19210 (N_19210,N_16661,N_15251);
xnor U19211 (N_19211,N_15380,N_15867);
and U19212 (N_19212,N_15210,N_15305);
and U19213 (N_19213,N_16749,N_16339);
nand U19214 (N_19214,N_16211,N_15474);
nand U19215 (N_19215,N_17750,N_15359);
nand U19216 (N_19216,N_17019,N_17134);
or U19217 (N_19217,N_16790,N_17878);
xnor U19218 (N_19218,N_17012,N_15135);
nand U19219 (N_19219,N_16759,N_16456);
nand U19220 (N_19220,N_17486,N_17273);
xnor U19221 (N_19221,N_15793,N_16013);
nand U19222 (N_19222,N_17721,N_17214);
xnor U19223 (N_19223,N_17787,N_17865);
and U19224 (N_19224,N_17676,N_16101);
and U19225 (N_19225,N_15939,N_15711);
or U19226 (N_19226,N_17375,N_17637);
xor U19227 (N_19227,N_17244,N_16815);
nand U19228 (N_19228,N_17337,N_17535);
or U19229 (N_19229,N_17839,N_17908);
xor U19230 (N_19230,N_17302,N_16872);
and U19231 (N_19231,N_17782,N_16452);
nor U19232 (N_19232,N_15149,N_15616);
or U19233 (N_19233,N_16453,N_16681);
and U19234 (N_19234,N_17924,N_15008);
and U19235 (N_19235,N_17065,N_16615);
nor U19236 (N_19236,N_16201,N_17440);
and U19237 (N_19237,N_15819,N_16584);
nand U19238 (N_19238,N_17933,N_16550);
xnor U19239 (N_19239,N_16715,N_15514);
and U19240 (N_19240,N_17994,N_17236);
and U19241 (N_19241,N_16787,N_17308);
and U19242 (N_19242,N_15578,N_17773);
nor U19243 (N_19243,N_15791,N_17006);
xnor U19244 (N_19244,N_17950,N_17780);
and U19245 (N_19245,N_17453,N_15209);
or U19246 (N_19246,N_17042,N_17284);
xor U19247 (N_19247,N_15479,N_16780);
xor U19248 (N_19248,N_17759,N_15984);
and U19249 (N_19249,N_16603,N_15858);
or U19250 (N_19250,N_17327,N_15892);
and U19251 (N_19251,N_15827,N_16116);
and U19252 (N_19252,N_15898,N_17720);
nand U19253 (N_19253,N_17784,N_17960);
xor U19254 (N_19254,N_17068,N_17919);
nor U19255 (N_19255,N_17164,N_17917);
nand U19256 (N_19256,N_15523,N_17400);
nor U19257 (N_19257,N_17856,N_16499);
xnor U19258 (N_19258,N_16510,N_17662);
or U19259 (N_19259,N_16786,N_16811);
or U19260 (N_19260,N_17663,N_17480);
nand U19261 (N_19261,N_15357,N_17234);
and U19262 (N_19262,N_17505,N_15988);
or U19263 (N_19263,N_17673,N_17809);
and U19264 (N_19264,N_15395,N_17023);
xor U19265 (N_19265,N_16518,N_15062);
nand U19266 (N_19266,N_16564,N_15180);
nor U19267 (N_19267,N_15363,N_15742);
or U19268 (N_19268,N_17261,N_15529);
and U19269 (N_19269,N_15485,N_15122);
and U19270 (N_19270,N_16967,N_15955);
or U19271 (N_19271,N_17763,N_16128);
nor U19272 (N_19272,N_16992,N_17191);
or U19273 (N_19273,N_16937,N_15572);
and U19274 (N_19274,N_15391,N_16418);
and U19275 (N_19275,N_17511,N_16170);
and U19276 (N_19276,N_17822,N_16252);
xnor U19277 (N_19277,N_17795,N_17344);
and U19278 (N_19278,N_17407,N_15423);
nor U19279 (N_19279,N_16635,N_16696);
and U19280 (N_19280,N_15639,N_17009);
nand U19281 (N_19281,N_17320,N_16645);
nor U19282 (N_19282,N_15145,N_16187);
nand U19283 (N_19283,N_16604,N_16494);
nand U19284 (N_19284,N_16280,N_16996);
nor U19285 (N_19285,N_17055,N_15733);
or U19286 (N_19286,N_16822,N_16910);
xor U19287 (N_19287,N_16296,N_15683);
and U19288 (N_19288,N_15429,N_16535);
nand U19289 (N_19289,N_15570,N_17241);
nor U19290 (N_19290,N_16979,N_17531);
and U19291 (N_19291,N_16710,N_16827);
nand U19292 (N_19292,N_16204,N_16660);
and U19293 (N_19293,N_17263,N_17521);
or U19294 (N_19294,N_16954,N_15710);
xnor U19295 (N_19295,N_16337,N_17075);
nor U19296 (N_19296,N_16734,N_16558);
nand U19297 (N_19297,N_16885,N_17125);
and U19298 (N_19298,N_17818,N_16583);
nor U19299 (N_19299,N_16921,N_15324);
nor U19300 (N_19300,N_15012,N_16355);
nand U19301 (N_19301,N_17062,N_15688);
and U19302 (N_19302,N_15215,N_16191);
nand U19303 (N_19303,N_16049,N_16484);
or U19304 (N_19304,N_17847,N_16001);
nand U19305 (N_19305,N_17122,N_16851);
nand U19306 (N_19306,N_15333,N_16480);
nor U19307 (N_19307,N_16537,N_17021);
or U19308 (N_19308,N_15535,N_16146);
and U19309 (N_19309,N_16221,N_16894);
and U19310 (N_19310,N_15851,N_15379);
and U19311 (N_19311,N_15338,N_17018);
nor U19312 (N_19312,N_17855,N_15706);
xnor U19313 (N_19313,N_17793,N_15730);
nand U19314 (N_19314,N_16799,N_16186);
xnor U19315 (N_19315,N_15056,N_17903);
nor U19316 (N_19316,N_16307,N_15148);
nor U19317 (N_19317,N_17084,N_15493);
and U19318 (N_19318,N_16292,N_16548);
nand U19319 (N_19319,N_15964,N_17768);
nor U19320 (N_19320,N_16321,N_17889);
nor U19321 (N_19321,N_16690,N_17517);
or U19322 (N_19322,N_16071,N_16556);
or U19323 (N_19323,N_16462,N_17356);
and U19324 (N_19324,N_15353,N_15650);
xnor U19325 (N_19325,N_15412,N_15776);
nor U19326 (N_19326,N_15962,N_15620);
and U19327 (N_19327,N_15936,N_16679);
and U19328 (N_19328,N_15689,N_16669);
nand U19329 (N_19329,N_17315,N_16096);
and U19330 (N_19330,N_16362,N_15897);
nor U19331 (N_19331,N_15196,N_16623);
or U19332 (N_19332,N_17722,N_16334);
and U19333 (N_19333,N_15878,N_16598);
nand U19334 (N_19334,N_16151,N_16233);
or U19335 (N_19335,N_17604,N_15644);
nor U19336 (N_19336,N_16009,N_15137);
and U19337 (N_19337,N_15399,N_17381);
and U19338 (N_19338,N_17506,N_17861);
nor U19339 (N_19339,N_15190,N_15605);
nand U19340 (N_19340,N_16103,N_15472);
xnor U19341 (N_19341,N_15501,N_15687);
and U19342 (N_19342,N_16389,N_15986);
and U19343 (N_19343,N_16289,N_15621);
nand U19344 (N_19344,N_16555,N_17688);
xnor U19345 (N_19345,N_16323,N_17348);
nand U19346 (N_19346,N_17419,N_15332);
and U19347 (N_19347,N_15027,N_17404);
and U19348 (N_19348,N_16976,N_16169);
and U19349 (N_19349,N_17577,N_15766);
and U19350 (N_19350,N_17563,N_17653);
nand U19351 (N_19351,N_15566,N_17149);
nand U19352 (N_19352,N_16038,N_16228);
xor U19353 (N_19353,N_15838,N_17366);
nand U19354 (N_19354,N_15284,N_15788);
xnor U19355 (N_19355,N_16485,N_16912);
nand U19356 (N_19356,N_17274,N_15100);
xor U19357 (N_19357,N_16523,N_15511);
or U19358 (N_19358,N_15749,N_15896);
or U19359 (N_19359,N_16027,N_15519);
nand U19360 (N_19360,N_16406,N_16132);
or U19361 (N_19361,N_16775,N_16724);
and U19362 (N_19362,N_15430,N_16870);
or U19363 (N_19363,N_15826,N_17050);
xor U19364 (N_19364,N_16268,N_16599);
or U19365 (N_19365,N_16417,N_15828);
or U19366 (N_19366,N_17482,N_15521);
and U19367 (N_19367,N_17397,N_17363);
nor U19368 (N_19368,N_17882,N_16004);
nand U19369 (N_19369,N_15052,N_15167);
and U19370 (N_19370,N_15626,N_17033);
and U19371 (N_19371,N_15307,N_15623);
nor U19372 (N_19372,N_15360,N_17177);
or U19373 (N_19373,N_17611,N_16469);
nand U19374 (N_19374,N_16973,N_17139);
nor U19375 (N_19375,N_16145,N_17942);
and U19376 (N_19376,N_15197,N_17153);
xnor U19377 (N_19377,N_17790,N_16932);
and U19378 (N_19378,N_15978,N_15597);
and U19379 (N_19379,N_17227,N_17179);
and U19380 (N_19380,N_16460,N_16784);
or U19381 (N_19381,N_17150,N_15045);
xor U19382 (N_19382,N_16189,N_16698);
or U19383 (N_19383,N_17433,N_15303);
or U19384 (N_19384,N_17279,N_16861);
xor U19385 (N_19385,N_16806,N_16212);
nor U19386 (N_19386,N_16733,N_15728);
or U19387 (N_19387,N_15378,N_17107);
nand U19388 (N_19388,N_16614,N_17733);
xor U19389 (N_19389,N_17566,N_15829);
nand U19390 (N_19390,N_16091,N_15249);
and U19391 (N_19391,N_16442,N_16797);
nand U19392 (N_19392,N_17242,N_17979);
nand U19393 (N_19393,N_15926,N_15204);
and U19394 (N_19394,N_17038,N_17067);
xnor U19395 (N_19395,N_15890,N_16752);
and U19396 (N_19396,N_16995,N_16552);
and U19397 (N_19397,N_17206,N_15131);
and U19398 (N_19398,N_16314,N_15021);
nand U19399 (N_19399,N_16015,N_15853);
and U19400 (N_19400,N_15577,N_16641);
nor U19401 (N_19401,N_17964,N_15772);
nor U19402 (N_19402,N_16625,N_17902);
or U19403 (N_19403,N_17345,N_15033);
or U19404 (N_19404,N_15692,N_17969);
nand U19405 (N_19405,N_15039,N_15011);
or U19406 (N_19406,N_15005,N_15673);
nand U19407 (N_19407,N_17713,N_16999);
and U19408 (N_19408,N_17088,N_16109);
xnor U19409 (N_19409,N_15979,N_15933);
and U19410 (N_19410,N_16868,N_17355);
and U19411 (N_19411,N_16380,N_16372);
xnor U19412 (N_19412,N_15126,N_15884);
nand U19413 (N_19413,N_15830,N_15775);
xnor U19414 (N_19414,N_15735,N_15779);
nand U19415 (N_19415,N_16248,N_15777);
nor U19416 (N_19416,N_15318,N_17035);
and U19417 (N_19417,N_15046,N_15646);
and U19418 (N_19418,N_17470,N_15837);
or U19419 (N_19419,N_17936,N_15587);
nor U19420 (N_19420,N_16981,N_17079);
xor U19421 (N_19421,N_17115,N_16773);
or U19422 (N_19422,N_16111,N_15030);
nor U19423 (N_19423,N_17286,N_17408);
or U19424 (N_19424,N_17043,N_16914);
xor U19425 (N_19425,N_16959,N_17827);
or U19426 (N_19426,N_17516,N_16226);
and U19427 (N_19427,N_17825,N_16588);
nor U19428 (N_19428,N_15842,N_15840);
nand U19429 (N_19429,N_17117,N_17943);
nor U19430 (N_19430,N_17233,N_15407);
nand U19431 (N_19431,N_17645,N_16888);
and U19432 (N_19432,N_17417,N_17959);
nand U19433 (N_19433,N_15343,N_17718);
and U19434 (N_19434,N_16106,N_15512);
and U19435 (N_19435,N_16739,N_15995);
nand U19436 (N_19436,N_15740,N_15026);
or U19437 (N_19437,N_15286,N_15389);
nor U19438 (N_19438,N_17732,N_15336);
or U19439 (N_19439,N_15028,N_17443);
nand U19440 (N_19440,N_17590,N_15516);
xor U19441 (N_19441,N_17980,N_16402);
nor U19442 (N_19442,N_17819,N_17555);
and U19443 (N_19443,N_15959,N_16869);
nor U19444 (N_19444,N_17103,N_17587);
nand U19445 (N_19445,N_16904,N_17202);
xor U19446 (N_19446,N_17892,N_17254);
xnor U19447 (N_19447,N_15112,N_15459);
and U19448 (N_19448,N_17527,N_15757);
or U19449 (N_19449,N_17047,N_17634);
xnor U19450 (N_19450,N_17181,N_15841);
nand U19451 (N_19451,N_16677,N_15346);
nor U19452 (N_19452,N_15586,N_16668);
xnor U19453 (N_19453,N_17931,N_15716);
or U19454 (N_19454,N_15739,N_16570);
nor U19455 (N_19455,N_16387,N_15402);
nor U19456 (N_19456,N_15393,N_17987);
or U19457 (N_19457,N_15142,N_15331);
xor U19458 (N_19458,N_16747,N_17613);
or U19459 (N_19459,N_16929,N_17141);
or U19460 (N_19460,N_15310,N_16591);
nor U19461 (N_19461,N_16750,N_16540);
or U19462 (N_19462,N_16152,N_16016);
xnor U19463 (N_19463,N_15217,N_17806);
and U19464 (N_19464,N_16383,N_16094);
and U19465 (N_19465,N_17152,N_17314);
nor U19466 (N_19466,N_15680,N_15950);
nand U19467 (N_19467,N_15029,N_15004);
nand U19468 (N_19468,N_17916,N_16147);
and U19469 (N_19469,N_17755,N_17895);
and U19470 (N_19470,N_17456,N_16165);
or U19471 (N_19471,N_16980,N_17195);
and U19472 (N_19472,N_16643,N_15048);
nor U19473 (N_19473,N_17391,N_16003);
nor U19474 (N_19474,N_17184,N_17127);
or U19475 (N_19475,N_17398,N_17185);
or U19476 (N_19476,N_15968,N_16342);
nand U19477 (N_19477,N_17159,N_15952);
nor U19478 (N_19478,N_15001,N_16400);
nand U19479 (N_19479,N_17543,N_16778);
nand U19480 (N_19480,N_15109,N_17091);
and U19481 (N_19481,N_15637,N_15596);
and U19482 (N_19482,N_16364,N_17418);
or U19483 (N_19483,N_15083,N_16295);
xnor U19484 (N_19484,N_15862,N_16883);
nor U19485 (N_19485,N_15458,N_15031);
or U19486 (N_19486,N_16405,N_15041);
xor U19487 (N_19487,N_15667,N_16365);
xnor U19488 (N_19488,N_17781,N_16029);
nor U19489 (N_19489,N_17303,N_15746);
and U19490 (N_19490,N_17192,N_16809);
or U19491 (N_19491,N_16688,N_16858);
nor U19492 (N_19492,N_15442,N_15296);
xnor U19493 (N_19493,N_17015,N_17660);
or U19494 (N_19494,N_17478,N_15406);
nor U19495 (N_19495,N_17992,N_15530);
nand U19496 (N_19496,N_17842,N_15084);
nand U19497 (N_19497,N_17446,N_17884);
nor U19498 (N_19498,N_16659,N_16719);
or U19499 (N_19499,N_16051,N_16142);
xor U19500 (N_19500,N_16728,N_15184);
and U19501 (N_19501,N_15043,N_15589);
nand U19502 (N_19502,N_17416,N_17348);
and U19503 (N_19503,N_15221,N_17939);
or U19504 (N_19504,N_17054,N_16079);
and U19505 (N_19505,N_15198,N_16512);
xnor U19506 (N_19506,N_16289,N_16953);
and U19507 (N_19507,N_15363,N_17058);
or U19508 (N_19508,N_16874,N_17797);
and U19509 (N_19509,N_16251,N_15450);
or U19510 (N_19510,N_17080,N_17803);
nor U19511 (N_19511,N_15610,N_17215);
xnor U19512 (N_19512,N_17903,N_16719);
nor U19513 (N_19513,N_16358,N_15306);
nor U19514 (N_19514,N_16642,N_17182);
nand U19515 (N_19515,N_17341,N_16832);
and U19516 (N_19516,N_15534,N_16039);
nand U19517 (N_19517,N_17088,N_16269);
or U19518 (N_19518,N_15382,N_16030);
xnor U19519 (N_19519,N_16820,N_16695);
nand U19520 (N_19520,N_16290,N_15500);
and U19521 (N_19521,N_16952,N_15938);
or U19522 (N_19522,N_16543,N_17913);
and U19523 (N_19523,N_17439,N_17409);
xnor U19524 (N_19524,N_15646,N_16112);
xor U19525 (N_19525,N_16868,N_16473);
nand U19526 (N_19526,N_16514,N_16443);
or U19527 (N_19527,N_15928,N_15951);
nor U19528 (N_19528,N_17212,N_17921);
or U19529 (N_19529,N_17504,N_15277);
or U19530 (N_19530,N_16266,N_17188);
and U19531 (N_19531,N_15332,N_15330);
nand U19532 (N_19532,N_16364,N_15178);
and U19533 (N_19533,N_16539,N_16266);
xor U19534 (N_19534,N_17833,N_16365);
xor U19535 (N_19535,N_17476,N_17363);
nand U19536 (N_19536,N_17557,N_17220);
nand U19537 (N_19537,N_16207,N_15077);
or U19538 (N_19538,N_15964,N_17693);
nand U19539 (N_19539,N_16466,N_16349);
or U19540 (N_19540,N_15884,N_15151);
and U19541 (N_19541,N_15231,N_16706);
and U19542 (N_19542,N_15888,N_15853);
and U19543 (N_19543,N_16010,N_17989);
nor U19544 (N_19544,N_16809,N_17861);
and U19545 (N_19545,N_17941,N_15662);
and U19546 (N_19546,N_16193,N_17817);
nand U19547 (N_19547,N_16334,N_16413);
or U19548 (N_19548,N_15113,N_15618);
and U19549 (N_19549,N_17476,N_17875);
or U19550 (N_19550,N_16209,N_17207);
and U19551 (N_19551,N_17645,N_17218);
xor U19552 (N_19552,N_15308,N_15526);
nand U19553 (N_19553,N_17061,N_16021);
xor U19554 (N_19554,N_16973,N_15164);
nand U19555 (N_19555,N_15642,N_16706);
nor U19556 (N_19556,N_16267,N_16382);
nand U19557 (N_19557,N_17464,N_17727);
or U19558 (N_19558,N_16184,N_16332);
and U19559 (N_19559,N_17136,N_17899);
xor U19560 (N_19560,N_17447,N_17558);
xnor U19561 (N_19561,N_16859,N_17966);
and U19562 (N_19562,N_16890,N_15933);
nand U19563 (N_19563,N_16464,N_17556);
nand U19564 (N_19564,N_17488,N_16665);
xor U19565 (N_19565,N_16542,N_16201);
nor U19566 (N_19566,N_15681,N_17005);
nor U19567 (N_19567,N_16018,N_15208);
and U19568 (N_19568,N_15554,N_15750);
or U19569 (N_19569,N_16154,N_16466);
xnor U19570 (N_19570,N_17853,N_16354);
nand U19571 (N_19571,N_17632,N_17971);
and U19572 (N_19572,N_15823,N_16663);
and U19573 (N_19573,N_17093,N_15194);
and U19574 (N_19574,N_17655,N_17563);
or U19575 (N_19575,N_15786,N_15748);
nand U19576 (N_19576,N_15662,N_17434);
nand U19577 (N_19577,N_16015,N_17433);
xor U19578 (N_19578,N_15307,N_16096);
nor U19579 (N_19579,N_17160,N_15291);
xnor U19580 (N_19580,N_16703,N_17949);
xnor U19581 (N_19581,N_17830,N_16425);
nand U19582 (N_19582,N_15994,N_17811);
or U19583 (N_19583,N_16870,N_15999);
nand U19584 (N_19584,N_15690,N_16602);
xnor U19585 (N_19585,N_16213,N_17167);
xor U19586 (N_19586,N_17499,N_17172);
and U19587 (N_19587,N_17012,N_15863);
xnor U19588 (N_19588,N_15167,N_15361);
and U19589 (N_19589,N_17227,N_15709);
and U19590 (N_19590,N_15433,N_15360);
and U19591 (N_19591,N_15337,N_17259);
or U19592 (N_19592,N_16435,N_17922);
and U19593 (N_19593,N_15373,N_16167);
nand U19594 (N_19594,N_17133,N_17818);
or U19595 (N_19595,N_16872,N_17635);
or U19596 (N_19596,N_15943,N_17929);
xor U19597 (N_19597,N_17221,N_16194);
or U19598 (N_19598,N_15583,N_16354);
nor U19599 (N_19599,N_17000,N_17915);
or U19600 (N_19600,N_17876,N_15929);
nand U19601 (N_19601,N_16591,N_15842);
xnor U19602 (N_19602,N_16157,N_16441);
xor U19603 (N_19603,N_15681,N_16728);
nand U19604 (N_19604,N_16125,N_15381);
and U19605 (N_19605,N_15734,N_16345);
and U19606 (N_19606,N_17164,N_17966);
or U19607 (N_19607,N_17101,N_15116);
and U19608 (N_19608,N_16922,N_15924);
and U19609 (N_19609,N_15455,N_16067);
and U19610 (N_19610,N_15411,N_17115);
nand U19611 (N_19611,N_15634,N_17548);
xnor U19612 (N_19612,N_17724,N_17626);
nor U19613 (N_19613,N_16150,N_16774);
nor U19614 (N_19614,N_16276,N_16788);
and U19615 (N_19615,N_16203,N_17796);
and U19616 (N_19616,N_16720,N_16863);
xor U19617 (N_19617,N_15942,N_15690);
xor U19618 (N_19618,N_15742,N_15139);
and U19619 (N_19619,N_17001,N_15819);
or U19620 (N_19620,N_15803,N_17533);
and U19621 (N_19621,N_15903,N_17275);
nand U19622 (N_19622,N_17135,N_15644);
nand U19623 (N_19623,N_16760,N_15772);
nand U19624 (N_19624,N_17763,N_15813);
and U19625 (N_19625,N_16907,N_17507);
nor U19626 (N_19626,N_16567,N_17266);
or U19627 (N_19627,N_17777,N_15725);
xnor U19628 (N_19628,N_16545,N_15930);
nor U19629 (N_19629,N_16242,N_17153);
nand U19630 (N_19630,N_16306,N_16558);
xor U19631 (N_19631,N_17277,N_15616);
xnor U19632 (N_19632,N_16634,N_15275);
and U19633 (N_19633,N_16193,N_15276);
nor U19634 (N_19634,N_16310,N_15436);
xor U19635 (N_19635,N_17508,N_15542);
or U19636 (N_19636,N_15148,N_16999);
and U19637 (N_19637,N_15461,N_16384);
or U19638 (N_19638,N_17375,N_17236);
nor U19639 (N_19639,N_15543,N_16498);
nor U19640 (N_19640,N_16165,N_15031);
and U19641 (N_19641,N_16788,N_15472);
nor U19642 (N_19642,N_16924,N_16931);
nand U19643 (N_19643,N_17717,N_16456);
nor U19644 (N_19644,N_15294,N_16918);
or U19645 (N_19645,N_16111,N_17104);
xor U19646 (N_19646,N_15304,N_15609);
or U19647 (N_19647,N_16723,N_15711);
nor U19648 (N_19648,N_16383,N_15224);
or U19649 (N_19649,N_16818,N_16000);
or U19650 (N_19650,N_16543,N_16353);
or U19651 (N_19651,N_17105,N_17711);
nand U19652 (N_19652,N_16222,N_16664);
or U19653 (N_19653,N_16071,N_16938);
and U19654 (N_19654,N_15178,N_16683);
or U19655 (N_19655,N_16735,N_17388);
and U19656 (N_19656,N_16265,N_17488);
xnor U19657 (N_19657,N_15890,N_16599);
and U19658 (N_19658,N_17024,N_17573);
nor U19659 (N_19659,N_16022,N_17431);
xor U19660 (N_19660,N_17637,N_17883);
or U19661 (N_19661,N_16662,N_17804);
and U19662 (N_19662,N_17347,N_17890);
nor U19663 (N_19663,N_17905,N_16992);
nand U19664 (N_19664,N_15071,N_15091);
nand U19665 (N_19665,N_17948,N_16818);
nor U19666 (N_19666,N_15196,N_15205);
xor U19667 (N_19667,N_16291,N_17687);
nand U19668 (N_19668,N_17822,N_15508);
xor U19669 (N_19669,N_15986,N_17124);
xor U19670 (N_19670,N_16613,N_17453);
and U19671 (N_19671,N_17733,N_15654);
xnor U19672 (N_19672,N_17823,N_15914);
and U19673 (N_19673,N_15870,N_15738);
and U19674 (N_19674,N_17548,N_15733);
nand U19675 (N_19675,N_16732,N_16549);
nand U19676 (N_19676,N_16078,N_17662);
or U19677 (N_19677,N_15798,N_16312);
xnor U19678 (N_19678,N_17124,N_15821);
and U19679 (N_19679,N_15544,N_17244);
and U19680 (N_19680,N_16360,N_16915);
xor U19681 (N_19681,N_15494,N_16634);
and U19682 (N_19682,N_16280,N_17972);
or U19683 (N_19683,N_17116,N_17646);
xor U19684 (N_19684,N_17824,N_15688);
or U19685 (N_19685,N_17147,N_15557);
nand U19686 (N_19686,N_17157,N_17447);
and U19687 (N_19687,N_16690,N_17292);
nor U19688 (N_19688,N_15759,N_15807);
and U19689 (N_19689,N_15176,N_15921);
nor U19690 (N_19690,N_17010,N_15928);
nand U19691 (N_19691,N_16973,N_16742);
nand U19692 (N_19692,N_17714,N_17969);
and U19693 (N_19693,N_17539,N_16614);
nor U19694 (N_19694,N_16855,N_16150);
and U19695 (N_19695,N_17439,N_15830);
and U19696 (N_19696,N_15437,N_16879);
or U19697 (N_19697,N_15995,N_17154);
nor U19698 (N_19698,N_15405,N_16838);
nor U19699 (N_19699,N_15039,N_17030);
nand U19700 (N_19700,N_17269,N_17231);
nor U19701 (N_19701,N_16614,N_15650);
nand U19702 (N_19702,N_16122,N_16887);
or U19703 (N_19703,N_15570,N_16191);
nor U19704 (N_19704,N_17541,N_15798);
or U19705 (N_19705,N_16060,N_16990);
or U19706 (N_19706,N_15746,N_17729);
nor U19707 (N_19707,N_17464,N_15275);
and U19708 (N_19708,N_17885,N_15013);
or U19709 (N_19709,N_16124,N_17561);
xor U19710 (N_19710,N_15690,N_15812);
or U19711 (N_19711,N_17391,N_17050);
nand U19712 (N_19712,N_17911,N_16354);
xnor U19713 (N_19713,N_16608,N_16190);
xnor U19714 (N_19714,N_16103,N_16154);
nor U19715 (N_19715,N_17785,N_17427);
nand U19716 (N_19716,N_17330,N_15343);
or U19717 (N_19717,N_16307,N_15564);
xnor U19718 (N_19718,N_16797,N_15978);
nor U19719 (N_19719,N_15161,N_16719);
nand U19720 (N_19720,N_17837,N_17503);
nor U19721 (N_19721,N_15794,N_16085);
and U19722 (N_19722,N_16491,N_17076);
xnor U19723 (N_19723,N_17735,N_17019);
nand U19724 (N_19724,N_16188,N_16795);
nand U19725 (N_19725,N_15311,N_15857);
and U19726 (N_19726,N_15773,N_17832);
nor U19727 (N_19727,N_17960,N_16424);
nand U19728 (N_19728,N_15813,N_16767);
nand U19729 (N_19729,N_17663,N_17893);
and U19730 (N_19730,N_15224,N_15275);
and U19731 (N_19731,N_17905,N_15722);
or U19732 (N_19732,N_16924,N_17868);
nor U19733 (N_19733,N_17636,N_16523);
and U19734 (N_19734,N_16439,N_16377);
nor U19735 (N_19735,N_15423,N_16142);
xnor U19736 (N_19736,N_17170,N_16305);
nor U19737 (N_19737,N_16112,N_15655);
or U19738 (N_19738,N_15127,N_16426);
or U19739 (N_19739,N_16806,N_16171);
xor U19740 (N_19740,N_17827,N_15445);
xnor U19741 (N_19741,N_15653,N_17736);
nand U19742 (N_19742,N_15256,N_17137);
nand U19743 (N_19743,N_16440,N_15994);
or U19744 (N_19744,N_16575,N_17772);
nor U19745 (N_19745,N_17144,N_16756);
and U19746 (N_19746,N_15696,N_16738);
nand U19747 (N_19747,N_17943,N_17373);
and U19748 (N_19748,N_15754,N_15520);
xnor U19749 (N_19749,N_17173,N_15163);
and U19750 (N_19750,N_15045,N_15782);
or U19751 (N_19751,N_15298,N_16581);
and U19752 (N_19752,N_15763,N_17295);
xor U19753 (N_19753,N_17014,N_17495);
or U19754 (N_19754,N_16699,N_16031);
and U19755 (N_19755,N_15827,N_15669);
xor U19756 (N_19756,N_17403,N_16574);
xnor U19757 (N_19757,N_17977,N_16979);
xnor U19758 (N_19758,N_17063,N_16524);
nand U19759 (N_19759,N_15382,N_17534);
or U19760 (N_19760,N_15818,N_17669);
or U19761 (N_19761,N_16502,N_17849);
and U19762 (N_19762,N_15298,N_17923);
and U19763 (N_19763,N_17479,N_15793);
or U19764 (N_19764,N_17876,N_15921);
nand U19765 (N_19765,N_16627,N_16770);
nand U19766 (N_19766,N_17881,N_16727);
and U19767 (N_19767,N_17203,N_16533);
xnor U19768 (N_19768,N_16853,N_16781);
xor U19769 (N_19769,N_17875,N_17666);
xnor U19770 (N_19770,N_16966,N_15793);
nor U19771 (N_19771,N_15933,N_16586);
and U19772 (N_19772,N_16438,N_15404);
and U19773 (N_19773,N_15809,N_15221);
xor U19774 (N_19774,N_17571,N_15257);
and U19775 (N_19775,N_17862,N_17950);
or U19776 (N_19776,N_17808,N_16991);
nand U19777 (N_19777,N_15120,N_15459);
xor U19778 (N_19778,N_15723,N_16558);
nor U19779 (N_19779,N_17535,N_15649);
xnor U19780 (N_19780,N_17222,N_15392);
xor U19781 (N_19781,N_16289,N_16531);
xor U19782 (N_19782,N_16228,N_16124);
and U19783 (N_19783,N_17719,N_17174);
nand U19784 (N_19784,N_17922,N_17933);
nor U19785 (N_19785,N_17203,N_17214);
nand U19786 (N_19786,N_15805,N_16530);
xnor U19787 (N_19787,N_15069,N_15180);
or U19788 (N_19788,N_15351,N_17226);
nand U19789 (N_19789,N_15491,N_16220);
or U19790 (N_19790,N_15662,N_17405);
and U19791 (N_19791,N_15145,N_15964);
nand U19792 (N_19792,N_17690,N_17036);
or U19793 (N_19793,N_16762,N_15841);
or U19794 (N_19794,N_16392,N_17152);
xor U19795 (N_19795,N_17233,N_17591);
nand U19796 (N_19796,N_15564,N_17535);
and U19797 (N_19797,N_17503,N_15357);
or U19798 (N_19798,N_15905,N_17390);
nor U19799 (N_19799,N_16323,N_17031);
nand U19800 (N_19800,N_16096,N_16429);
nor U19801 (N_19801,N_17344,N_17085);
nor U19802 (N_19802,N_17505,N_15335);
or U19803 (N_19803,N_15098,N_15695);
or U19804 (N_19804,N_16557,N_17234);
or U19805 (N_19805,N_16458,N_15247);
xor U19806 (N_19806,N_16654,N_15655);
nand U19807 (N_19807,N_16730,N_15589);
xnor U19808 (N_19808,N_17930,N_16262);
nor U19809 (N_19809,N_15910,N_16415);
or U19810 (N_19810,N_16368,N_17909);
and U19811 (N_19811,N_16023,N_16217);
and U19812 (N_19812,N_17646,N_16529);
nand U19813 (N_19813,N_16423,N_16087);
nor U19814 (N_19814,N_15952,N_15576);
nor U19815 (N_19815,N_15545,N_17454);
nand U19816 (N_19816,N_16129,N_15947);
nor U19817 (N_19817,N_15438,N_15129);
nor U19818 (N_19818,N_15623,N_16903);
and U19819 (N_19819,N_16790,N_16809);
or U19820 (N_19820,N_17750,N_15097);
nor U19821 (N_19821,N_17170,N_17706);
and U19822 (N_19822,N_16584,N_17546);
nand U19823 (N_19823,N_17556,N_17240);
nor U19824 (N_19824,N_17165,N_16323);
xnor U19825 (N_19825,N_15957,N_15746);
and U19826 (N_19826,N_17422,N_15536);
and U19827 (N_19827,N_17090,N_17546);
nand U19828 (N_19828,N_17619,N_16620);
xor U19829 (N_19829,N_16125,N_17025);
and U19830 (N_19830,N_17354,N_17995);
nor U19831 (N_19831,N_15050,N_15850);
nand U19832 (N_19832,N_17976,N_17900);
xnor U19833 (N_19833,N_16398,N_17599);
or U19834 (N_19834,N_16519,N_17009);
or U19835 (N_19835,N_15531,N_15250);
xnor U19836 (N_19836,N_16794,N_16793);
and U19837 (N_19837,N_17827,N_16788);
nor U19838 (N_19838,N_15934,N_15519);
and U19839 (N_19839,N_17268,N_16762);
nand U19840 (N_19840,N_17531,N_16897);
xnor U19841 (N_19841,N_17619,N_17264);
xor U19842 (N_19842,N_17229,N_15187);
or U19843 (N_19843,N_15295,N_16776);
or U19844 (N_19844,N_17689,N_16394);
and U19845 (N_19845,N_15274,N_17920);
xnor U19846 (N_19846,N_17581,N_15944);
and U19847 (N_19847,N_16829,N_17134);
and U19848 (N_19848,N_15681,N_17937);
or U19849 (N_19849,N_17783,N_15251);
nor U19850 (N_19850,N_15983,N_17411);
or U19851 (N_19851,N_15591,N_16296);
nand U19852 (N_19852,N_17326,N_17342);
xnor U19853 (N_19853,N_15330,N_17481);
nor U19854 (N_19854,N_17395,N_17747);
or U19855 (N_19855,N_15619,N_16979);
and U19856 (N_19856,N_17727,N_17840);
nand U19857 (N_19857,N_17320,N_17900);
or U19858 (N_19858,N_15905,N_17470);
xnor U19859 (N_19859,N_17554,N_17092);
or U19860 (N_19860,N_17843,N_16861);
nor U19861 (N_19861,N_17623,N_16391);
and U19862 (N_19862,N_17138,N_15726);
and U19863 (N_19863,N_16194,N_15403);
or U19864 (N_19864,N_17697,N_16966);
or U19865 (N_19865,N_15177,N_17808);
and U19866 (N_19866,N_17944,N_15569);
and U19867 (N_19867,N_15465,N_17630);
and U19868 (N_19868,N_15236,N_16804);
nor U19869 (N_19869,N_17532,N_17393);
xnor U19870 (N_19870,N_15876,N_15886);
nor U19871 (N_19871,N_16003,N_15725);
nor U19872 (N_19872,N_17650,N_16003);
nor U19873 (N_19873,N_16634,N_16778);
nand U19874 (N_19874,N_15523,N_15652);
nor U19875 (N_19875,N_16458,N_17345);
xor U19876 (N_19876,N_17907,N_16599);
or U19877 (N_19877,N_16967,N_17134);
nand U19878 (N_19878,N_17339,N_17583);
or U19879 (N_19879,N_16568,N_15268);
and U19880 (N_19880,N_17826,N_17050);
xor U19881 (N_19881,N_16864,N_16547);
xor U19882 (N_19882,N_16782,N_17492);
or U19883 (N_19883,N_16870,N_17790);
or U19884 (N_19884,N_15922,N_17367);
nand U19885 (N_19885,N_15655,N_15431);
and U19886 (N_19886,N_15245,N_16571);
and U19887 (N_19887,N_15906,N_17640);
nor U19888 (N_19888,N_15256,N_16399);
nor U19889 (N_19889,N_17788,N_15920);
nor U19890 (N_19890,N_16029,N_15501);
xnor U19891 (N_19891,N_17288,N_16556);
or U19892 (N_19892,N_15752,N_15889);
xnor U19893 (N_19893,N_17233,N_16309);
nor U19894 (N_19894,N_17438,N_16051);
or U19895 (N_19895,N_16444,N_17717);
xnor U19896 (N_19896,N_16420,N_17000);
and U19897 (N_19897,N_17369,N_15440);
nor U19898 (N_19898,N_15933,N_17246);
nand U19899 (N_19899,N_16374,N_17079);
and U19900 (N_19900,N_17126,N_16092);
and U19901 (N_19901,N_16113,N_15948);
nand U19902 (N_19902,N_17936,N_16040);
xnor U19903 (N_19903,N_16282,N_17541);
or U19904 (N_19904,N_15643,N_16828);
xor U19905 (N_19905,N_15746,N_16654);
nand U19906 (N_19906,N_15740,N_17542);
or U19907 (N_19907,N_17662,N_15808);
nor U19908 (N_19908,N_17782,N_17439);
or U19909 (N_19909,N_16893,N_17871);
or U19910 (N_19910,N_17008,N_16373);
or U19911 (N_19911,N_17190,N_15821);
nor U19912 (N_19912,N_15000,N_17110);
nor U19913 (N_19913,N_16070,N_15939);
xor U19914 (N_19914,N_16537,N_15560);
nand U19915 (N_19915,N_16355,N_15286);
nand U19916 (N_19916,N_15259,N_15208);
xnor U19917 (N_19917,N_15938,N_16290);
nand U19918 (N_19918,N_17779,N_16554);
xnor U19919 (N_19919,N_16644,N_17392);
or U19920 (N_19920,N_16490,N_17759);
and U19921 (N_19921,N_17515,N_16100);
and U19922 (N_19922,N_16169,N_17100);
nor U19923 (N_19923,N_15872,N_15860);
nor U19924 (N_19924,N_15165,N_15816);
xor U19925 (N_19925,N_16584,N_16496);
or U19926 (N_19926,N_15869,N_17943);
nand U19927 (N_19927,N_17204,N_16852);
nor U19928 (N_19928,N_16517,N_15928);
nor U19929 (N_19929,N_16934,N_16227);
nand U19930 (N_19930,N_15959,N_17857);
and U19931 (N_19931,N_16368,N_15068);
nor U19932 (N_19932,N_17922,N_17683);
nand U19933 (N_19933,N_16706,N_15579);
nand U19934 (N_19934,N_16657,N_15207);
nand U19935 (N_19935,N_15446,N_17070);
nor U19936 (N_19936,N_16857,N_16727);
and U19937 (N_19937,N_15392,N_17669);
nand U19938 (N_19938,N_16631,N_16275);
and U19939 (N_19939,N_15417,N_17314);
nor U19940 (N_19940,N_16255,N_17079);
and U19941 (N_19941,N_17103,N_17019);
nand U19942 (N_19942,N_17032,N_16426);
nor U19943 (N_19943,N_15424,N_17447);
or U19944 (N_19944,N_16091,N_15407);
nand U19945 (N_19945,N_15775,N_17421);
and U19946 (N_19946,N_15431,N_16986);
nand U19947 (N_19947,N_16186,N_15942);
or U19948 (N_19948,N_16948,N_16748);
nand U19949 (N_19949,N_15420,N_16101);
nor U19950 (N_19950,N_15013,N_16416);
xor U19951 (N_19951,N_15825,N_17970);
nor U19952 (N_19952,N_17929,N_15227);
nand U19953 (N_19953,N_16069,N_15056);
nand U19954 (N_19954,N_16905,N_16547);
nor U19955 (N_19955,N_17400,N_15371);
or U19956 (N_19956,N_15088,N_16217);
xor U19957 (N_19957,N_17812,N_16348);
xnor U19958 (N_19958,N_16039,N_17951);
nand U19959 (N_19959,N_17963,N_15720);
or U19960 (N_19960,N_16014,N_17122);
nor U19961 (N_19961,N_15432,N_15453);
and U19962 (N_19962,N_15854,N_16168);
nand U19963 (N_19963,N_17751,N_17463);
nand U19964 (N_19964,N_15101,N_17816);
and U19965 (N_19965,N_15255,N_17971);
nand U19966 (N_19966,N_16364,N_17502);
and U19967 (N_19967,N_17500,N_17030);
or U19968 (N_19968,N_15480,N_16699);
nand U19969 (N_19969,N_16084,N_17259);
nor U19970 (N_19970,N_17700,N_17000);
or U19971 (N_19971,N_15013,N_16187);
nor U19972 (N_19972,N_15989,N_15959);
nor U19973 (N_19973,N_17838,N_15164);
or U19974 (N_19974,N_17570,N_15147);
xor U19975 (N_19975,N_17192,N_16298);
and U19976 (N_19976,N_15998,N_16146);
nor U19977 (N_19977,N_15383,N_17280);
and U19978 (N_19978,N_17594,N_15765);
or U19979 (N_19979,N_17462,N_17351);
nand U19980 (N_19980,N_16169,N_16306);
nand U19981 (N_19981,N_15962,N_17190);
or U19982 (N_19982,N_15211,N_16114);
and U19983 (N_19983,N_16599,N_16346);
or U19984 (N_19984,N_15978,N_17925);
nand U19985 (N_19985,N_15520,N_16098);
nor U19986 (N_19986,N_15360,N_16612);
xor U19987 (N_19987,N_16475,N_16555);
xor U19988 (N_19988,N_15779,N_16289);
xor U19989 (N_19989,N_16078,N_16419);
nor U19990 (N_19990,N_15568,N_15401);
xor U19991 (N_19991,N_16927,N_16135);
nand U19992 (N_19992,N_17632,N_17317);
and U19993 (N_19993,N_15696,N_17621);
or U19994 (N_19994,N_15007,N_17301);
and U19995 (N_19995,N_16365,N_16537);
or U19996 (N_19996,N_15138,N_15481);
and U19997 (N_19997,N_15109,N_15439);
nand U19998 (N_19998,N_17386,N_16050);
xor U19999 (N_19999,N_15793,N_16544);
nand U20000 (N_20000,N_16013,N_15885);
or U20001 (N_20001,N_15085,N_17947);
nor U20002 (N_20002,N_15616,N_17770);
nor U20003 (N_20003,N_17594,N_17338);
xnor U20004 (N_20004,N_17426,N_17966);
nand U20005 (N_20005,N_16305,N_15419);
or U20006 (N_20006,N_16504,N_15130);
or U20007 (N_20007,N_15140,N_15121);
or U20008 (N_20008,N_17267,N_17910);
and U20009 (N_20009,N_17474,N_17795);
and U20010 (N_20010,N_17090,N_16640);
nor U20011 (N_20011,N_17217,N_15518);
nand U20012 (N_20012,N_16366,N_15272);
and U20013 (N_20013,N_17181,N_15223);
and U20014 (N_20014,N_16723,N_17737);
nor U20015 (N_20015,N_17259,N_15062);
nand U20016 (N_20016,N_17243,N_15542);
and U20017 (N_20017,N_17598,N_17765);
and U20018 (N_20018,N_15889,N_16498);
xor U20019 (N_20019,N_17752,N_17847);
or U20020 (N_20020,N_16751,N_17174);
nand U20021 (N_20021,N_17666,N_17514);
or U20022 (N_20022,N_15718,N_17461);
nor U20023 (N_20023,N_15377,N_17059);
and U20024 (N_20024,N_16953,N_15865);
xor U20025 (N_20025,N_17289,N_16032);
or U20026 (N_20026,N_15626,N_15238);
and U20027 (N_20027,N_17242,N_15693);
xnor U20028 (N_20028,N_16834,N_15170);
nand U20029 (N_20029,N_16216,N_15811);
nor U20030 (N_20030,N_17664,N_15490);
or U20031 (N_20031,N_16637,N_16693);
xor U20032 (N_20032,N_16491,N_15813);
nand U20033 (N_20033,N_17175,N_16641);
nor U20034 (N_20034,N_15283,N_17994);
xor U20035 (N_20035,N_16894,N_15375);
and U20036 (N_20036,N_17280,N_16479);
or U20037 (N_20037,N_17497,N_16130);
or U20038 (N_20038,N_17913,N_17947);
nand U20039 (N_20039,N_17780,N_16522);
xnor U20040 (N_20040,N_15375,N_16892);
nand U20041 (N_20041,N_15682,N_15755);
and U20042 (N_20042,N_15884,N_15840);
and U20043 (N_20043,N_16234,N_17437);
nor U20044 (N_20044,N_15292,N_15254);
and U20045 (N_20045,N_16503,N_17135);
nor U20046 (N_20046,N_17701,N_16337);
xor U20047 (N_20047,N_15853,N_15090);
and U20048 (N_20048,N_15245,N_15158);
and U20049 (N_20049,N_15799,N_16817);
nor U20050 (N_20050,N_17193,N_17929);
nand U20051 (N_20051,N_16704,N_17815);
nand U20052 (N_20052,N_16548,N_17854);
or U20053 (N_20053,N_16371,N_17253);
xnor U20054 (N_20054,N_16600,N_16075);
xor U20055 (N_20055,N_16657,N_16185);
nor U20056 (N_20056,N_15530,N_16334);
or U20057 (N_20057,N_15637,N_17189);
nor U20058 (N_20058,N_15593,N_16043);
and U20059 (N_20059,N_16563,N_15674);
and U20060 (N_20060,N_16568,N_17914);
or U20061 (N_20061,N_15428,N_16071);
nand U20062 (N_20062,N_16888,N_15487);
xnor U20063 (N_20063,N_17909,N_16403);
nand U20064 (N_20064,N_17425,N_15019);
nand U20065 (N_20065,N_16630,N_15816);
nand U20066 (N_20066,N_16233,N_16098);
xnor U20067 (N_20067,N_15057,N_16362);
or U20068 (N_20068,N_16443,N_15041);
nand U20069 (N_20069,N_16793,N_17898);
xor U20070 (N_20070,N_15410,N_15337);
or U20071 (N_20071,N_16224,N_15059);
xor U20072 (N_20072,N_17569,N_17756);
or U20073 (N_20073,N_15690,N_15564);
xor U20074 (N_20074,N_16432,N_16982);
xor U20075 (N_20075,N_15893,N_15773);
or U20076 (N_20076,N_16136,N_15624);
nand U20077 (N_20077,N_17834,N_17745);
xnor U20078 (N_20078,N_15901,N_16969);
or U20079 (N_20079,N_17335,N_15239);
xor U20080 (N_20080,N_17839,N_15161);
or U20081 (N_20081,N_15262,N_17588);
xor U20082 (N_20082,N_16715,N_15178);
or U20083 (N_20083,N_15298,N_17144);
nand U20084 (N_20084,N_16500,N_15545);
nor U20085 (N_20085,N_15784,N_17464);
xor U20086 (N_20086,N_16028,N_15366);
xnor U20087 (N_20087,N_17352,N_15205);
and U20088 (N_20088,N_17890,N_15835);
and U20089 (N_20089,N_16463,N_15647);
nand U20090 (N_20090,N_16903,N_17157);
nor U20091 (N_20091,N_17456,N_16542);
and U20092 (N_20092,N_16459,N_17120);
and U20093 (N_20093,N_17617,N_17944);
or U20094 (N_20094,N_17593,N_17133);
nand U20095 (N_20095,N_15041,N_17426);
nor U20096 (N_20096,N_17080,N_16090);
nor U20097 (N_20097,N_15296,N_16538);
nand U20098 (N_20098,N_17648,N_15990);
nor U20099 (N_20099,N_17091,N_15864);
xnor U20100 (N_20100,N_16959,N_15166);
nand U20101 (N_20101,N_16016,N_17840);
nor U20102 (N_20102,N_15296,N_15655);
xor U20103 (N_20103,N_16201,N_15185);
nand U20104 (N_20104,N_16312,N_15234);
and U20105 (N_20105,N_17953,N_15254);
and U20106 (N_20106,N_17597,N_15791);
nand U20107 (N_20107,N_16673,N_16034);
xnor U20108 (N_20108,N_16060,N_16028);
nor U20109 (N_20109,N_16546,N_15652);
xor U20110 (N_20110,N_15770,N_15152);
or U20111 (N_20111,N_16355,N_15169);
nor U20112 (N_20112,N_15766,N_16593);
or U20113 (N_20113,N_16075,N_15133);
nand U20114 (N_20114,N_15560,N_17130);
xor U20115 (N_20115,N_16784,N_15952);
or U20116 (N_20116,N_17477,N_17901);
nand U20117 (N_20117,N_16083,N_16135);
or U20118 (N_20118,N_17683,N_15079);
xnor U20119 (N_20119,N_15600,N_17668);
and U20120 (N_20120,N_16050,N_16979);
nor U20121 (N_20121,N_17001,N_16768);
xnor U20122 (N_20122,N_17122,N_16843);
nor U20123 (N_20123,N_17635,N_16434);
nor U20124 (N_20124,N_17289,N_15601);
xor U20125 (N_20125,N_15661,N_15008);
xor U20126 (N_20126,N_15409,N_16305);
nand U20127 (N_20127,N_17588,N_15238);
nor U20128 (N_20128,N_15010,N_17903);
xor U20129 (N_20129,N_16816,N_17870);
nor U20130 (N_20130,N_15257,N_17229);
or U20131 (N_20131,N_17393,N_17337);
xnor U20132 (N_20132,N_15695,N_16293);
nor U20133 (N_20133,N_17775,N_17329);
nor U20134 (N_20134,N_16428,N_17793);
or U20135 (N_20135,N_15580,N_17620);
or U20136 (N_20136,N_16745,N_17147);
nand U20137 (N_20137,N_16898,N_15231);
nand U20138 (N_20138,N_17557,N_17718);
or U20139 (N_20139,N_15756,N_15764);
nand U20140 (N_20140,N_15748,N_17089);
nor U20141 (N_20141,N_16565,N_17431);
nand U20142 (N_20142,N_17619,N_17415);
or U20143 (N_20143,N_15631,N_16691);
nand U20144 (N_20144,N_15984,N_15401);
or U20145 (N_20145,N_17512,N_15939);
nor U20146 (N_20146,N_15149,N_17452);
or U20147 (N_20147,N_17991,N_17286);
nor U20148 (N_20148,N_16853,N_17512);
and U20149 (N_20149,N_16713,N_17609);
or U20150 (N_20150,N_15160,N_15752);
xor U20151 (N_20151,N_16822,N_16866);
or U20152 (N_20152,N_17854,N_15032);
nand U20153 (N_20153,N_16376,N_16968);
nand U20154 (N_20154,N_15530,N_15784);
and U20155 (N_20155,N_17062,N_17388);
nand U20156 (N_20156,N_17159,N_17090);
nand U20157 (N_20157,N_16941,N_15923);
xor U20158 (N_20158,N_16018,N_16566);
xor U20159 (N_20159,N_17503,N_17312);
nand U20160 (N_20160,N_17966,N_16180);
or U20161 (N_20161,N_17938,N_15240);
nand U20162 (N_20162,N_16356,N_15659);
nand U20163 (N_20163,N_17236,N_15968);
and U20164 (N_20164,N_16466,N_17886);
or U20165 (N_20165,N_15024,N_16066);
xnor U20166 (N_20166,N_15770,N_15222);
and U20167 (N_20167,N_16085,N_17344);
nand U20168 (N_20168,N_16041,N_16424);
and U20169 (N_20169,N_15166,N_16140);
or U20170 (N_20170,N_16580,N_15135);
xnor U20171 (N_20171,N_15221,N_16110);
or U20172 (N_20172,N_17174,N_17715);
and U20173 (N_20173,N_15295,N_17923);
or U20174 (N_20174,N_15353,N_17770);
xor U20175 (N_20175,N_16323,N_15544);
nor U20176 (N_20176,N_17639,N_17036);
or U20177 (N_20177,N_17813,N_15715);
and U20178 (N_20178,N_15833,N_17186);
xnor U20179 (N_20179,N_15758,N_16481);
nand U20180 (N_20180,N_17717,N_17040);
nand U20181 (N_20181,N_17501,N_15811);
nor U20182 (N_20182,N_17462,N_16886);
or U20183 (N_20183,N_17132,N_16271);
or U20184 (N_20184,N_16229,N_17190);
or U20185 (N_20185,N_16615,N_16095);
xor U20186 (N_20186,N_15720,N_15719);
and U20187 (N_20187,N_17821,N_15467);
and U20188 (N_20188,N_16333,N_17067);
or U20189 (N_20189,N_15818,N_16401);
or U20190 (N_20190,N_15562,N_17596);
and U20191 (N_20191,N_16880,N_15551);
nor U20192 (N_20192,N_15803,N_15159);
nor U20193 (N_20193,N_17259,N_15152);
or U20194 (N_20194,N_17002,N_15375);
and U20195 (N_20195,N_16577,N_17499);
and U20196 (N_20196,N_16092,N_17936);
xnor U20197 (N_20197,N_16732,N_17926);
xnor U20198 (N_20198,N_15121,N_16528);
nand U20199 (N_20199,N_15310,N_16354);
and U20200 (N_20200,N_15294,N_17465);
nor U20201 (N_20201,N_16130,N_15228);
nand U20202 (N_20202,N_15230,N_17290);
nor U20203 (N_20203,N_17865,N_16221);
or U20204 (N_20204,N_15678,N_15583);
and U20205 (N_20205,N_15944,N_16643);
nor U20206 (N_20206,N_16661,N_17985);
nand U20207 (N_20207,N_17086,N_17795);
nor U20208 (N_20208,N_16768,N_17535);
nand U20209 (N_20209,N_16621,N_16422);
or U20210 (N_20210,N_16350,N_16011);
and U20211 (N_20211,N_17176,N_15922);
or U20212 (N_20212,N_16179,N_16431);
nor U20213 (N_20213,N_15870,N_16287);
or U20214 (N_20214,N_15769,N_16126);
nand U20215 (N_20215,N_15614,N_16460);
nor U20216 (N_20216,N_16205,N_16625);
and U20217 (N_20217,N_16845,N_15073);
or U20218 (N_20218,N_15084,N_17959);
and U20219 (N_20219,N_17717,N_17884);
and U20220 (N_20220,N_15039,N_17606);
xnor U20221 (N_20221,N_15409,N_17357);
and U20222 (N_20222,N_17225,N_15429);
nor U20223 (N_20223,N_17300,N_15830);
nor U20224 (N_20224,N_17071,N_16241);
nand U20225 (N_20225,N_15238,N_16265);
nor U20226 (N_20226,N_15473,N_15067);
and U20227 (N_20227,N_17842,N_17212);
and U20228 (N_20228,N_17928,N_17559);
nor U20229 (N_20229,N_17665,N_16217);
nor U20230 (N_20230,N_16135,N_17054);
nor U20231 (N_20231,N_16500,N_15302);
or U20232 (N_20232,N_17589,N_16341);
and U20233 (N_20233,N_15311,N_16688);
or U20234 (N_20234,N_15184,N_17386);
xnor U20235 (N_20235,N_17553,N_15986);
nor U20236 (N_20236,N_17290,N_17042);
nor U20237 (N_20237,N_17481,N_16584);
xnor U20238 (N_20238,N_15449,N_16351);
or U20239 (N_20239,N_16341,N_17724);
xnor U20240 (N_20240,N_16538,N_17952);
xnor U20241 (N_20241,N_17750,N_17357);
nand U20242 (N_20242,N_17322,N_16699);
nand U20243 (N_20243,N_16775,N_15305);
and U20244 (N_20244,N_16275,N_17522);
and U20245 (N_20245,N_15993,N_15300);
nor U20246 (N_20246,N_17578,N_16636);
xor U20247 (N_20247,N_17478,N_15956);
nor U20248 (N_20248,N_15210,N_17213);
or U20249 (N_20249,N_15477,N_15940);
or U20250 (N_20250,N_17845,N_15051);
or U20251 (N_20251,N_15052,N_17815);
or U20252 (N_20252,N_15092,N_15303);
xnor U20253 (N_20253,N_15166,N_15950);
xnor U20254 (N_20254,N_17080,N_16914);
xor U20255 (N_20255,N_15885,N_16937);
nor U20256 (N_20256,N_16637,N_16750);
nor U20257 (N_20257,N_17832,N_16995);
xor U20258 (N_20258,N_15541,N_16858);
nand U20259 (N_20259,N_16175,N_17458);
nand U20260 (N_20260,N_16199,N_17460);
nand U20261 (N_20261,N_16077,N_17631);
and U20262 (N_20262,N_16581,N_15205);
nor U20263 (N_20263,N_15086,N_17775);
xnor U20264 (N_20264,N_16075,N_17547);
and U20265 (N_20265,N_17165,N_17295);
nor U20266 (N_20266,N_15865,N_16464);
or U20267 (N_20267,N_15725,N_17188);
or U20268 (N_20268,N_17773,N_16108);
nand U20269 (N_20269,N_15059,N_17762);
and U20270 (N_20270,N_15551,N_15922);
or U20271 (N_20271,N_16648,N_17355);
and U20272 (N_20272,N_16002,N_15106);
nor U20273 (N_20273,N_17012,N_16409);
xnor U20274 (N_20274,N_17512,N_16117);
nand U20275 (N_20275,N_16260,N_15564);
and U20276 (N_20276,N_16314,N_16294);
nor U20277 (N_20277,N_15382,N_16166);
or U20278 (N_20278,N_17297,N_17599);
nor U20279 (N_20279,N_15696,N_15123);
nand U20280 (N_20280,N_16966,N_16037);
nand U20281 (N_20281,N_17426,N_15741);
nor U20282 (N_20282,N_15337,N_17157);
and U20283 (N_20283,N_15448,N_15308);
nor U20284 (N_20284,N_16643,N_15015);
nand U20285 (N_20285,N_17640,N_16323);
nor U20286 (N_20286,N_15366,N_17763);
or U20287 (N_20287,N_16025,N_16663);
nor U20288 (N_20288,N_16187,N_16575);
and U20289 (N_20289,N_17380,N_16386);
or U20290 (N_20290,N_17763,N_16239);
and U20291 (N_20291,N_16245,N_16368);
nor U20292 (N_20292,N_17157,N_15664);
xnor U20293 (N_20293,N_15981,N_17477);
and U20294 (N_20294,N_17575,N_15390);
and U20295 (N_20295,N_16287,N_16520);
or U20296 (N_20296,N_17497,N_16134);
or U20297 (N_20297,N_15706,N_15398);
nor U20298 (N_20298,N_16978,N_17100);
and U20299 (N_20299,N_15064,N_15343);
nor U20300 (N_20300,N_16600,N_15496);
nand U20301 (N_20301,N_17440,N_15956);
nor U20302 (N_20302,N_15804,N_15853);
nor U20303 (N_20303,N_16131,N_17398);
and U20304 (N_20304,N_16785,N_15138);
nand U20305 (N_20305,N_16033,N_16933);
nor U20306 (N_20306,N_16560,N_16115);
or U20307 (N_20307,N_16531,N_15807);
nor U20308 (N_20308,N_15450,N_15204);
and U20309 (N_20309,N_17434,N_16182);
and U20310 (N_20310,N_17472,N_16250);
and U20311 (N_20311,N_15593,N_16816);
nor U20312 (N_20312,N_16999,N_16460);
and U20313 (N_20313,N_16502,N_16049);
xnor U20314 (N_20314,N_17622,N_15281);
nand U20315 (N_20315,N_16783,N_16337);
or U20316 (N_20316,N_15419,N_16785);
nand U20317 (N_20317,N_16252,N_17839);
and U20318 (N_20318,N_17043,N_16270);
xnor U20319 (N_20319,N_16816,N_16843);
xnor U20320 (N_20320,N_15446,N_16073);
nand U20321 (N_20321,N_16334,N_17950);
or U20322 (N_20322,N_17490,N_16914);
nor U20323 (N_20323,N_17138,N_16518);
nor U20324 (N_20324,N_15461,N_16485);
or U20325 (N_20325,N_17098,N_16358);
nor U20326 (N_20326,N_16113,N_16520);
or U20327 (N_20327,N_16009,N_15739);
and U20328 (N_20328,N_17904,N_17199);
nor U20329 (N_20329,N_15348,N_17480);
and U20330 (N_20330,N_17750,N_16013);
nor U20331 (N_20331,N_16319,N_17356);
xnor U20332 (N_20332,N_17478,N_16038);
nor U20333 (N_20333,N_17409,N_16405);
xor U20334 (N_20334,N_16634,N_16999);
nand U20335 (N_20335,N_17885,N_15265);
nand U20336 (N_20336,N_16096,N_15611);
nor U20337 (N_20337,N_17809,N_15854);
nand U20338 (N_20338,N_15917,N_16934);
xor U20339 (N_20339,N_15645,N_16784);
nand U20340 (N_20340,N_16161,N_17622);
or U20341 (N_20341,N_15389,N_17537);
or U20342 (N_20342,N_17687,N_15128);
or U20343 (N_20343,N_16920,N_15424);
nand U20344 (N_20344,N_15620,N_16854);
or U20345 (N_20345,N_16594,N_16304);
nor U20346 (N_20346,N_16756,N_17821);
nand U20347 (N_20347,N_17907,N_16361);
nor U20348 (N_20348,N_15382,N_16161);
xnor U20349 (N_20349,N_17645,N_15852);
or U20350 (N_20350,N_17874,N_16769);
nor U20351 (N_20351,N_17377,N_17934);
nor U20352 (N_20352,N_16551,N_16862);
nand U20353 (N_20353,N_16195,N_17241);
nor U20354 (N_20354,N_17848,N_16915);
or U20355 (N_20355,N_15183,N_17185);
nor U20356 (N_20356,N_17335,N_17209);
or U20357 (N_20357,N_15314,N_15523);
or U20358 (N_20358,N_17163,N_17686);
nor U20359 (N_20359,N_17940,N_17889);
or U20360 (N_20360,N_17046,N_17709);
xnor U20361 (N_20361,N_17907,N_16450);
nand U20362 (N_20362,N_17834,N_16386);
nand U20363 (N_20363,N_16360,N_17736);
nand U20364 (N_20364,N_16607,N_17326);
nor U20365 (N_20365,N_16727,N_17753);
nand U20366 (N_20366,N_15042,N_15693);
xnor U20367 (N_20367,N_15102,N_15097);
or U20368 (N_20368,N_15055,N_15034);
nor U20369 (N_20369,N_16943,N_16525);
and U20370 (N_20370,N_16760,N_16088);
xnor U20371 (N_20371,N_16118,N_15341);
or U20372 (N_20372,N_15970,N_15570);
nor U20373 (N_20373,N_15746,N_15809);
nor U20374 (N_20374,N_16343,N_17247);
nand U20375 (N_20375,N_17644,N_16404);
xnor U20376 (N_20376,N_16882,N_16558);
or U20377 (N_20377,N_16159,N_17110);
and U20378 (N_20378,N_15682,N_16769);
and U20379 (N_20379,N_16844,N_15112);
nand U20380 (N_20380,N_16888,N_16701);
and U20381 (N_20381,N_15214,N_17152);
xor U20382 (N_20382,N_16242,N_16858);
nand U20383 (N_20383,N_16198,N_17241);
xor U20384 (N_20384,N_17255,N_15973);
or U20385 (N_20385,N_17550,N_15941);
nor U20386 (N_20386,N_16333,N_17926);
and U20387 (N_20387,N_15648,N_16149);
or U20388 (N_20388,N_17520,N_16980);
and U20389 (N_20389,N_16766,N_15748);
and U20390 (N_20390,N_15140,N_15568);
nand U20391 (N_20391,N_16937,N_15773);
xnor U20392 (N_20392,N_16932,N_16455);
and U20393 (N_20393,N_16942,N_15853);
xnor U20394 (N_20394,N_17787,N_17758);
nor U20395 (N_20395,N_16841,N_17836);
nor U20396 (N_20396,N_17472,N_17598);
nand U20397 (N_20397,N_17318,N_17076);
and U20398 (N_20398,N_16453,N_16550);
and U20399 (N_20399,N_16582,N_16378);
nand U20400 (N_20400,N_17465,N_16822);
and U20401 (N_20401,N_15102,N_16680);
and U20402 (N_20402,N_17766,N_16040);
and U20403 (N_20403,N_16161,N_17524);
nor U20404 (N_20404,N_15804,N_15349);
nand U20405 (N_20405,N_17594,N_15376);
nor U20406 (N_20406,N_17841,N_15994);
nor U20407 (N_20407,N_17930,N_16517);
nor U20408 (N_20408,N_17976,N_16181);
and U20409 (N_20409,N_15244,N_16434);
nor U20410 (N_20410,N_16628,N_15578);
nor U20411 (N_20411,N_15312,N_16088);
and U20412 (N_20412,N_17991,N_17390);
nor U20413 (N_20413,N_17608,N_16146);
xnor U20414 (N_20414,N_17259,N_15109);
nor U20415 (N_20415,N_16081,N_15422);
nor U20416 (N_20416,N_15897,N_16973);
or U20417 (N_20417,N_15591,N_15361);
xor U20418 (N_20418,N_17826,N_15081);
and U20419 (N_20419,N_17154,N_17355);
nand U20420 (N_20420,N_16891,N_15273);
nor U20421 (N_20421,N_15453,N_15862);
nand U20422 (N_20422,N_17050,N_17741);
xor U20423 (N_20423,N_15888,N_17172);
xor U20424 (N_20424,N_16414,N_15376);
and U20425 (N_20425,N_15640,N_17237);
and U20426 (N_20426,N_15855,N_15125);
nand U20427 (N_20427,N_17290,N_17159);
or U20428 (N_20428,N_17354,N_16677);
nand U20429 (N_20429,N_15158,N_17826);
and U20430 (N_20430,N_15699,N_15126);
nand U20431 (N_20431,N_15072,N_16024);
and U20432 (N_20432,N_16114,N_16112);
or U20433 (N_20433,N_17934,N_15559);
and U20434 (N_20434,N_17842,N_16292);
nand U20435 (N_20435,N_16970,N_16045);
xor U20436 (N_20436,N_15357,N_16577);
nor U20437 (N_20437,N_17598,N_16417);
or U20438 (N_20438,N_17817,N_17962);
xor U20439 (N_20439,N_15875,N_17755);
nand U20440 (N_20440,N_16263,N_16266);
or U20441 (N_20441,N_15258,N_15564);
and U20442 (N_20442,N_17196,N_15922);
xor U20443 (N_20443,N_15297,N_16577);
nor U20444 (N_20444,N_16428,N_16860);
nor U20445 (N_20445,N_16411,N_16780);
xnor U20446 (N_20446,N_17361,N_17578);
nand U20447 (N_20447,N_15089,N_15470);
nand U20448 (N_20448,N_16542,N_16609);
nor U20449 (N_20449,N_16249,N_15879);
nand U20450 (N_20450,N_16933,N_15050);
nor U20451 (N_20451,N_17514,N_17312);
nand U20452 (N_20452,N_16957,N_16826);
and U20453 (N_20453,N_15806,N_16525);
xor U20454 (N_20454,N_16756,N_16882);
nor U20455 (N_20455,N_17902,N_16990);
xnor U20456 (N_20456,N_15546,N_16796);
or U20457 (N_20457,N_15365,N_16714);
and U20458 (N_20458,N_17273,N_17484);
nor U20459 (N_20459,N_17082,N_15898);
or U20460 (N_20460,N_15610,N_17498);
nor U20461 (N_20461,N_17196,N_17675);
xor U20462 (N_20462,N_16409,N_17734);
or U20463 (N_20463,N_15938,N_17659);
nand U20464 (N_20464,N_15136,N_15320);
xnor U20465 (N_20465,N_17194,N_16896);
nand U20466 (N_20466,N_16425,N_17703);
nor U20467 (N_20467,N_17322,N_17795);
nand U20468 (N_20468,N_17674,N_16655);
and U20469 (N_20469,N_16972,N_17747);
or U20470 (N_20470,N_16748,N_15913);
nand U20471 (N_20471,N_17191,N_15582);
nor U20472 (N_20472,N_16322,N_17811);
and U20473 (N_20473,N_16742,N_17806);
nor U20474 (N_20474,N_15785,N_16096);
and U20475 (N_20475,N_16831,N_15406);
or U20476 (N_20476,N_15200,N_15180);
and U20477 (N_20477,N_17857,N_15004);
xnor U20478 (N_20478,N_17874,N_17586);
nand U20479 (N_20479,N_17657,N_16277);
nand U20480 (N_20480,N_15757,N_17490);
nor U20481 (N_20481,N_15268,N_15145);
nand U20482 (N_20482,N_17120,N_15670);
nand U20483 (N_20483,N_17847,N_15348);
and U20484 (N_20484,N_15036,N_17931);
xor U20485 (N_20485,N_16138,N_15186);
or U20486 (N_20486,N_17532,N_16088);
xnor U20487 (N_20487,N_16058,N_16630);
and U20488 (N_20488,N_15602,N_15567);
nand U20489 (N_20489,N_16851,N_15106);
nand U20490 (N_20490,N_15584,N_15626);
nor U20491 (N_20491,N_16721,N_15152);
and U20492 (N_20492,N_17418,N_16223);
xnor U20493 (N_20493,N_17197,N_17541);
or U20494 (N_20494,N_15374,N_16467);
or U20495 (N_20495,N_16712,N_16612);
and U20496 (N_20496,N_17767,N_16322);
or U20497 (N_20497,N_16752,N_17341);
nor U20498 (N_20498,N_16476,N_17614);
or U20499 (N_20499,N_15165,N_16697);
nor U20500 (N_20500,N_15972,N_15712);
nor U20501 (N_20501,N_17920,N_17628);
nand U20502 (N_20502,N_17377,N_16165);
and U20503 (N_20503,N_17601,N_17013);
xnor U20504 (N_20504,N_15449,N_17417);
xor U20505 (N_20505,N_17819,N_16439);
nand U20506 (N_20506,N_17646,N_15363);
and U20507 (N_20507,N_15151,N_15184);
xor U20508 (N_20508,N_15264,N_17115);
and U20509 (N_20509,N_17892,N_15157);
and U20510 (N_20510,N_16216,N_16121);
nand U20511 (N_20511,N_15407,N_17835);
xor U20512 (N_20512,N_16748,N_16970);
or U20513 (N_20513,N_16421,N_17793);
and U20514 (N_20514,N_16065,N_17757);
and U20515 (N_20515,N_15798,N_15933);
nor U20516 (N_20516,N_16182,N_16408);
and U20517 (N_20517,N_15484,N_17557);
xnor U20518 (N_20518,N_15018,N_16225);
nand U20519 (N_20519,N_15173,N_16866);
nand U20520 (N_20520,N_16653,N_15456);
or U20521 (N_20521,N_15391,N_15491);
nor U20522 (N_20522,N_17602,N_15564);
nand U20523 (N_20523,N_16370,N_16472);
nand U20524 (N_20524,N_17471,N_16419);
nor U20525 (N_20525,N_16265,N_17411);
nand U20526 (N_20526,N_17943,N_17502);
xnor U20527 (N_20527,N_15130,N_16806);
or U20528 (N_20528,N_15085,N_17827);
nor U20529 (N_20529,N_16031,N_16638);
nand U20530 (N_20530,N_16323,N_16991);
or U20531 (N_20531,N_15074,N_16704);
nor U20532 (N_20532,N_16080,N_16167);
or U20533 (N_20533,N_17554,N_17036);
xor U20534 (N_20534,N_16733,N_16912);
xnor U20535 (N_20535,N_17719,N_16783);
xor U20536 (N_20536,N_16748,N_15980);
or U20537 (N_20537,N_17190,N_16534);
xnor U20538 (N_20538,N_17977,N_17560);
nor U20539 (N_20539,N_17982,N_16214);
or U20540 (N_20540,N_17874,N_15514);
and U20541 (N_20541,N_17306,N_16629);
nand U20542 (N_20542,N_16516,N_17517);
xor U20543 (N_20543,N_16719,N_17713);
or U20544 (N_20544,N_17666,N_16637);
or U20545 (N_20545,N_17353,N_17812);
xnor U20546 (N_20546,N_16244,N_16293);
or U20547 (N_20547,N_17720,N_16771);
xnor U20548 (N_20548,N_17426,N_16668);
nor U20549 (N_20549,N_15682,N_16206);
nand U20550 (N_20550,N_17261,N_17050);
nand U20551 (N_20551,N_17321,N_16549);
xor U20552 (N_20552,N_15679,N_15341);
nand U20553 (N_20553,N_17696,N_17450);
or U20554 (N_20554,N_16473,N_16652);
xnor U20555 (N_20555,N_15702,N_15212);
or U20556 (N_20556,N_16615,N_17550);
xnor U20557 (N_20557,N_17655,N_17244);
xor U20558 (N_20558,N_15540,N_16270);
xnor U20559 (N_20559,N_16629,N_16899);
and U20560 (N_20560,N_15657,N_15239);
xnor U20561 (N_20561,N_15472,N_17611);
or U20562 (N_20562,N_16238,N_15619);
or U20563 (N_20563,N_15486,N_15052);
nand U20564 (N_20564,N_15924,N_17299);
nand U20565 (N_20565,N_17435,N_16193);
nor U20566 (N_20566,N_15854,N_15668);
nor U20567 (N_20567,N_16362,N_17522);
and U20568 (N_20568,N_17400,N_17235);
nand U20569 (N_20569,N_16408,N_17687);
xnor U20570 (N_20570,N_17304,N_16503);
xnor U20571 (N_20571,N_15033,N_15373);
nor U20572 (N_20572,N_16006,N_15697);
nor U20573 (N_20573,N_16876,N_15269);
and U20574 (N_20574,N_16261,N_16373);
or U20575 (N_20575,N_16450,N_15818);
nor U20576 (N_20576,N_16424,N_15925);
nor U20577 (N_20577,N_16256,N_16819);
and U20578 (N_20578,N_17858,N_15289);
and U20579 (N_20579,N_15683,N_16683);
nand U20580 (N_20580,N_16448,N_16744);
or U20581 (N_20581,N_17410,N_17734);
nor U20582 (N_20582,N_16026,N_15445);
nand U20583 (N_20583,N_15758,N_16878);
nand U20584 (N_20584,N_17492,N_15728);
xnor U20585 (N_20585,N_17806,N_17715);
or U20586 (N_20586,N_16554,N_15103);
nor U20587 (N_20587,N_16970,N_15703);
nor U20588 (N_20588,N_15116,N_17064);
xnor U20589 (N_20589,N_16055,N_17700);
xor U20590 (N_20590,N_15357,N_16114);
and U20591 (N_20591,N_16953,N_15495);
xnor U20592 (N_20592,N_17524,N_15990);
nor U20593 (N_20593,N_17666,N_15351);
nand U20594 (N_20594,N_17593,N_15440);
nand U20595 (N_20595,N_16079,N_15727);
or U20596 (N_20596,N_15275,N_16473);
nor U20597 (N_20597,N_17306,N_15435);
xnor U20598 (N_20598,N_17882,N_17394);
xor U20599 (N_20599,N_16257,N_17449);
nor U20600 (N_20600,N_17308,N_15919);
nor U20601 (N_20601,N_17294,N_15087);
and U20602 (N_20602,N_15800,N_15034);
and U20603 (N_20603,N_16170,N_15476);
nor U20604 (N_20604,N_15008,N_15302);
nor U20605 (N_20605,N_15076,N_17201);
and U20606 (N_20606,N_15664,N_15057);
and U20607 (N_20607,N_17128,N_15303);
xor U20608 (N_20608,N_15145,N_16091);
and U20609 (N_20609,N_16320,N_17137);
nor U20610 (N_20610,N_16735,N_15372);
xor U20611 (N_20611,N_15481,N_16768);
nor U20612 (N_20612,N_17638,N_15819);
or U20613 (N_20613,N_16351,N_16037);
and U20614 (N_20614,N_16894,N_17454);
nand U20615 (N_20615,N_17307,N_17247);
or U20616 (N_20616,N_16805,N_17515);
xor U20617 (N_20617,N_15648,N_15430);
nor U20618 (N_20618,N_17335,N_15012);
or U20619 (N_20619,N_17511,N_17566);
xor U20620 (N_20620,N_16530,N_15944);
and U20621 (N_20621,N_17621,N_16767);
or U20622 (N_20622,N_16605,N_17276);
nand U20623 (N_20623,N_16824,N_17876);
nand U20624 (N_20624,N_17627,N_15685);
nand U20625 (N_20625,N_15377,N_17551);
and U20626 (N_20626,N_16814,N_16050);
and U20627 (N_20627,N_16914,N_16894);
nor U20628 (N_20628,N_17298,N_16870);
or U20629 (N_20629,N_16400,N_16100);
and U20630 (N_20630,N_17787,N_16563);
or U20631 (N_20631,N_17943,N_17494);
nand U20632 (N_20632,N_17778,N_15400);
and U20633 (N_20633,N_17468,N_16115);
and U20634 (N_20634,N_15071,N_17693);
and U20635 (N_20635,N_16635,N_15018);
nor U20636 (N_20636,N_17920,N_17396);
or U20637 (N_20637,N_16659,N_17306);
nand U20638 (N_20638,N_16647,N_15260);
and U20639 (N_20639,N_16108,N_16255);
or U20640 (N_20640,N_15799,N_15668);
or U20641 (N_20641,N_17289,N_17228);
nand U20642 (N_20642,N_15250,N_15187);
or U20643 (N_20643,N_16699,N_16736);
or U20644 (N_20644,N_16070,N_17187);
xnor U20645 (N_20645,N_17562,N_16387);
or U20646 (N_20646,N_15684,N_16361);
or U20647 (N_20647,N_15126,N_15410);
and U20648 (N_20648,N_16479,N_15334);
and U20649 (N_20649,N_16140,N_15056);
xor U20650 (N_20650,N_17720,N_16933);
nand U20651 (N_20651,N_16932,N_16136);
and U20652 (N_20652,N_15121,N_17161);
nor U20653 (N_20653,N_15454,N_16563);
xnor U20654 (N_20654,N_17693,N_15204);
and U20655 (N_20655,N_17759,N_15761);
nand U20656 (N_20656,N_15934,N_16513);
and U20657 (N_20657,N_15164,N_17952);
nor U20658 (N_20658,N_17404,N_15826);
or U20659 (N_20659,N_15047,N_16826);
nor U20660 (N_20660,N_16301,N_17166);
or U20661 (N_20661,N_15237,N_17658);
nor U20662 (N_20662,N_16615,N_17208);
and U20663 (N_20663,N_16877,N_15702);
nor U20664 (N_20664,N_16268,N_15171);
nand U20665 (N_20665,N_15446,N_16872);
nand U20666 (N_20666,N_16558,N_15651);
nand U20667 (N_20667,N_16562,N_16176);
nor U20668 (N_20668,N_15961,N_17387);
or U20669 (N_20669,N_16443,N_15211);
xor U20670 (N_20670,N_16707,N_15499);
nor U20671 (N_20671,N_15820,N_16380);
nand U20672 (N_20672,N_17703,N_16487);
nor U20673 (N_20673,N_17083,N_17245);
nor U20674 (N_20674,N_17109,N_15655);
xnor U20675 (N_20675,N_15100,N_15297);
or U20676 (N_20676,N_16974,N_16740);
nand U20677 (N_20677,N_15800,N_16792);
nand U20678 (N_20678,N_17136,N_15996);
nor U20679 (N_20679,N_16042,N_15471);
nor U20680 (N_20680,N_15289,N_16081);
nand U20681 (N_20681,N_15800,N_16150);
or U20682 (N_20682,N_16989,N_17844);
or U20683 (N_20683,N_15084,N_16750);
and U20684 (N_20684,N_15356,N_15153);
nor U20685 (N_20685,N_17267,N_16978);
nor U20686 (N_20686,N_17554,N_16675);
or U20687 (N_20687,N_15627,N_15038);
and U20688 (N_20688,N_15656,N_15837);
nand U20689 (N_20689,N_16374,N_15054);
nor U20690 (N_20690,N_16188,N_16593);
nand U20691 (N_20691,N_15703,N_17269);
xor U20692 (N_20692,N_15617,N_15414);
or U20693 (N_20693,N_15375,N_16461);
nand U20694 (N_20694,N_17655,N_16359);
nand U20695 (N_20695,N_16987,N_15864);
or U20696 (N_20696,N_16940,N_15416);
nor U20697 (N_20697,N_17208,N_16654);
or U20698 (N_20698,N_15640,N_15169);
or U20699 (N_20699,N_17588,N_16907);
xnor U20700 (N_20700,N_17088,N_15637);
or U20701 (N_20701,N_16387,N_15422);
nand U20702 (N_20702,N_17972,N_15243);
and U20703 (N_20703,N_15640,N_17818);
nand U20704 (N_20704,N_16100,N_15469);
and U20705 (N_20705,N_17180,N_15587);
or U20706 (N_20706,N_15934,N_15518);
or U20707 (N_20707,N_16797,N_16147);
nand U20708 (N_20708,N_15008,N_15575);
or U20709 (N_20709,N_16888,N_17223);
nand U20710 (N_20710,N_15322,N_17173);
xnor U20711 (N_20711,N_15790,N_17078);
nor U20712 (N_20712,N_16509,N_15255);
nor U20713 (N_20713,N_15317,N_15984);
or U20714 (N_20714,N_15315,N_17559);
or U20715 (N_20715,N_15899,N_15503);
nand U20716 (N_20716,N_16485,N_15432);
nor U20717 (N_20717,N_16411,N_15059);
xnor U20718 (N_20718,N_15372,N_16510);
xor U20719 (N_20719,N_15383,N_15079);
xor U20720 (N_20720,N_16309,N_17069);
xor U20721 (N_20721,N_16147,N_15515);
or U20722 (N_20722,N_16317,N_17486);
and U20723 (N_20723,N_16804,N_17736);
or U20724 (N_20724,N_17058,N_17602);
and U20725 (N_20725,N_16550,N_15989);
xnor U20726 (N_20726,N_16570,N_15716);
nand U20727 (N_20727,N_15224,N_16854);
or U20728 (N_20728,N_15713,N_17735);
and U20729 (N_20729,N_16102,N_15356);
nand U20730 (N_20730,N_15982,N_16934);
or U20731 (N_20731,N_16912,N_17627);
and U20732 (N_20732,N_17727,N_15343);
and U20733 (N_20733,N_16763,N_16583);
or U20734 (N_20734,N_16467,N_15877);
and U20735 (N_20735,N_16117,N_16756);
nand U20736 (N_20736,N_17159,N_15470);
and U20737 (N_20737,N_16641,N_15607);
or U20738 (N_20738,N_16126,N_17562);
nor U20739 (N_20739,N_17058,N_16435);
xor U20740 (N_20740,N_15097,N_15926);
and U20741 (N_20741,N_16248,N_15541);
xor U20742 (N_20742,N_16207,N_16451);
and U20743 (N_20743,N_15285,N_16566);
nor U20744 (N_20744,N_16662,N_15334);
xnor U20745 (N_20745,N_15925,N_15411);
and U20746 (N_20746,N_16924,N_16431);
or U20747 (N_20747,N_17301,N_15651);
xnor U20748 (N_20748,N_17149,N_17408);
or U20749 (N_20749,N_16614,N_17366);
nand U20750 (N_20750,N_15008,N_17997);
or U20751 (N_20751,N_15133,N_15719);
nand U20752 (N_20752,N_16424,N_16179);
or U20753 (N_20753,N_15961,N_17401);
nor U20754 (N_20754,N_17108,N_17598);
and U20755 (N_20755,N_15203,N_17667);
nand U20756 (N_20756,N_17871,N_15409);
nand U20757 (N_20757,N_15817,N_17304);
nor U20758 (N_20758,N_16100,N_16844);
and U20759 (N_20759,N_17045,N_16565);
and U20760 (N_20760,N_16926,N_15547);
or U20761 (N_20761,N_17952,N_15951);
xnor U20762 (N_20762,N_17965,N_16478);
xnor U20763 (N_20763,N_16624,N_17275);
nor U20764 (N_20764,N_15057,N_17879);
and U20765 (N_20765,N_17480,N_16829);
nand U20766 (N_20766,N_16589,N_15091);
or U20767 (N_20767,N_16043,N_15047);
and U20768 (N_20768,N_17018,N_17549);
nand U20769 (N_20769,N_15414,N_17598);
or U20770 (N_20770,N_17085,N_16070);
or U20771 (N_20771,N_17355,N_16583);
nor U20772 (N_20772,N_16118,N_16865);
xnor U20773 (N_20773,N_15526,N_17699);
xnor U20774 (N_20774,N_16501,N_15041);
nand U20775 (N_20775,N_16271,N_17512);
nor U20776 (N_20776,N_15323,N_17934);
nor U20777 (N_20777,N_15079,N_16349);
xor U20778 (N_20778,N_17606,N_15752);
nand U20779 (N_20779,N_15715,N_17538);
or U20780 (N_20780,N_15443,N_17425);
xnor U20781 (N_20781,N_17721,N_17745);
and U20782 (N_20782,N_17009,N_15302);
nand U20783 (N_20783,N_16107,N_15695);
and U20784 (N_20784,N_15821,N_15328);
nor U20785 (N_20785,N_17547,N_17595);
xor U20786 (N_20786,N_16601,N_16684);
nand U20787 (N_20787,N_17266,N_16367);
or U20788 (N_20788,N_15231,N_15156);
nor U20789 (N_20789,N_17899,N_16305);
and U20790 (N_20790,N_17959,N_15143);
nand U20791 (N_20791,N_15172,N_16011);
nor U20792 (N_20792,N_16436,N_15174);
nor U20793 (N_20793,N_17011,N_17393);
xnor U20794 (N_20794,N_16314,N_16522);
xor U20795 (N_20795,N_16842,N_15093);
or U20796 (N_20796,N_15364,N_15665);
xnor U20797 (N_20797,N_15723,N_15570);
or U20798 (N_20798,N_15615,N_16886);
xor U20799 (N_20799,N_15358,N_17800);
or U20800 (N_20800,N_16907,N_15410);
nor U20801 (N_20801,N_15762,N_16936);
or U20802 (N_20802,N_17348,N_17294);
and U20803 (N_20803,N_15066,N_16525);
xnor U20804 (N_20804,N_16906,N_17754);
or U20805 (N_20805,N_15080,N_15167);
nor U20806 (N_20806,N_17638,N_16894);
and U20807 (N_20807,N_16433,N_17012);
or U20808 (N_20808,N_16811,N_15909);
xor U20809 (N_20809,N_15603,N_15204);
and U20810 (N_20810,N_16812,N_16678);
and U20811 (N_20811,N_16143,N_17785);
nor U20812 (N_20812,N_17457,N_15768);
xnor U20813 (N_20813,N_17615,N_17095);
nand U20814 (N_20814,N_15512,N_16765);
xor U20815 (N_20815,N_17993,N_15487);
nor U20816 (N_20816,N_16783,N_16243);
nor U20817 (N_20817,N_15088,N_17191);
and U20818 (N_20818,N_16081,N_17023);
xnor U20819 (N_20819,N_17516,N_17566);
nor U20820 (N_20820,N_17689,N_16795);
and U20821 (N_20821,N_16241,N_15810);
xnor U20822 (N_20822,N_17270,N_17267);
or U20823 (N_20823,N_16851,N_16127);
nor U20824 (N_20824,N_15486,N_17672);
or U20825 (N_20825,N_16471,N_16052);
and U20826 (N_20826,N_15785,N_16237);
nor U20827 (N_20827,N_17635,N_17193);
nor U20828 (N_20828,N_17601,N_16835);
xnor U20829 (N_20829,N_17068,N_16803);
or U20830 (N_20830,N_15822,N_17618);
nand U20831 (N_20831,N_16506,N_16463);
nand U20832 (N_20832,N_17729,N_15389);
nand U20833 (N_20833,N_16101,N_17936);
xnor U20834 (N_20834,N_17378,N_17770);
xor U20835 (N_20835,N_16639,N_16725);
xnor U20836 (N_20836,N_17891,N_17926);
xor U20837 (N_20837,N_15639,N_15755);
nor U20838 (N_20838,N_15069,N_17427);
or U20839 (N_20839,N_16401,N_15721);
or U20840 (N_20840,N_15975,N_16171);
and U20841 (N_20841,N_15964,N_17466);
nand U20842 (N_20842,N_16730,N_17847);
nand U20843 (N_20843,N_16974,N_17343);
nor U20844 (N_20844,N_16761,N_17441);
and U20845 (N_20845,N_17119,N_16176);
xnor U20846 (N_20846,N_15029,N_16774);
or U20847 (N_20847,N_17807,N_17988);
and U20848 (N_20848,N_15647,N_16185);
nor U20849 (N_20849,N_16510,N_16982);
nand U20850 (N_20850,N_16647,N_15228);
nor U20851 (N_20851,N_17402,N_16849);
nor U20852 (N_20852,N_17145,N_15624);
xnor U20853 (N_20853,N_15478,N_16273);
nand U20854 (N_20854,N_17001,N_15363);
and U20855 (N_20855,N_16386,N_15720);
or U20856 (N_20856,N_15391,N_16437);
or U20857 (N_20857,N_17999,N_16566);
or U20858 (N_20858,N_17285,N_16472);
nand U20859 (N_20859,N_16233,N_17730);
or U20860 (N_20860,N_16792,N_15863);
or U20861 (N_20861,N_15262,N_16248);
or U20862 (N_20862,N_17833,N_17748);
or U20863 (N_20863,N_16813,N_17972);
nand U20864 (N_20864,N_15889,N_16315);
or U20865 (N_20865,N_15280,N_17204);
or U20866 (N_20866,N_16922,N_16694);
xor U20867 (N_20867,N_15012,N_15104);
xnor U20868 (N_20868,N_16273,N_17694);
and U20869 (N_20869,N_16685,N_16597);
nand U20870 (N_20870,N_15027,N_15159);
xor U20871 (N_20871,N_16017,N_15315);
nand U20872 (N_20872,N_16487,N_17070);
and U20873 (N_20873,N_17367,N_15918);
nand U20874 (N_20874,N_17338,N_17047);
and U20875 (N_20875,N_16319,N_17292);
xnor U20876 (N_20876,N_16063,N_15429);
or U20877 (N_20877,N_17791,N_15831);
xor U20878 (N_20878,N_16041,N_15121);
or U20879 (N_20879,N_17287,N_16333);
or U20880 (N_20880,N_17024,N_16630);
or U20881 (N_20881,N_16170,N_15335);
or U20882 (N_20882,N_15092,N_16840);
xor U20883 (N_20883,N_16029,N_15970);
nor U20884 (N_20884,N_17580,N_15133);
xnor U20885 (N_20885,N_15298,N_15158);
nand U20886 (N_20886,N_16170,N_16490);
and U20887 (N_20887,N_15770,N_15923);
and U20888 (N_20888,N_17337,N_17779);
and U20889 (N_20889,N_16511,N_15398);
nand U20890 (N_20890,N_16827,N_15609);
xor U20891 (N_20891,N_17553,N_16793);
and U20892 (N_20892,N_17626,N_16710);
or U20893 (N_20893,N_16527,N_15984);
nor U20894 (N_20894,N_15445,N_17813);
and U20895 (N_20895,N_15496,N_16700);
xor U20896 (N_20896,N_16906,N_16738);
xor U20897 (N_20897,N_15532,N_15497);
or U20898 (N_20898,N_17116,N_15216);
nor U20899 (N_20899,N_17014,N_16939);
and U20900 (N_20900,N_17898,N_17493);
and U20901 (N_20901,N_15572,N_17249);
xnor U20902 (N_20902,N_16493,N_15933);
xnor U20903 (N_20903,N_17828,N_16586);
nand U20904 (N_20904,N_17579,N_15376);
or U20905 (N_20905,N_17614,N_16827);
or U20906 (N_20906,N_16605,N_17521);
nand U20907 (N_20907,N_15342,N_15794);
xnor U20908 (N_20908,N_16594,N_16485);
nand U20909 (N_20909,N_17273,N_15313);
nor U20910 (N_20910,N_16989,N_17228);
xnor U20911 (N_20911,N_17749,N_16910);
and U20912 (N_20912,N_15630,N_16831);
xor U20913 (N_20913,N_16496,N_16049);
and U20914 (N_20914,N_17249,N_15006);
or U20915 (N_20915,N_15544,N_17985);
and U20916 (N_20916,N_16790,N_16440);
nand U20917 (N_20917,N_17083,N_15081);
nor U20918 (N_20918,N_15997,N_16599);
nor U20919 (N_20919,N_17799,N_16313);
nand U20920 (N_20920,N_15247,N_15451);
nand U20921 (N_20921,N_16671,N_17879);
nand U20922 (N_20922,N_16294,N_17266);
nand U20923 (N_20923,N_16818,N_16585);
nor U20924 (N_20924,N_17333,N_15725);
nor U20925 (N_20925,N_17294,N_15506);
nand U20926 (N_20926,N_15212,N_15926);
nand U20927 (N_20927,N_17147,N_17357);
xor U20928 (N_20928,N_15173,N_17651);
xnor U20929 (N_20929,N_16641,N_15554);
or U20930 (N_20930,N_15715,N_16464);
xor U20931 (N_20931,N_15500,N_16626);
nand U20932 (N_20932,N_17293,N_16231);
nand U20933 (N_20933,N_15583,N_15184);
xor U20934 (N_20934,N_15710,N_17777);
xnor U20935 (N_20935,N_16741,N_16189);
and U20936 (N_20936,N_16945,N_15550);
nor U20937 (N_20937,N_17787,N_15299);
nand U20938 (N_20938,N_17396,N_15413);
xor U20939 (N_20939,N_16003,N_17419);
nor U20940 (N_20940,N_16661,N_15523);
nand U20941 (N_20941,N_17052,N_16630);
or U20942 (N_20942,N_16313,N_16130);
nand U20943 (N_20943,N_17934,N_17768);
or U20944 (N_20944,N_16640,N_16051);
xor U20945 (N_20945,N_16042,N_16592);
nand U20946 (N_20946,N_17443,N_16044);
and U20947 (N_20947,N_16087,N_16638);
and U20948 (N_20948,N_15185,N_16611);
nor U20949 (N_20949,N_17819,N_15113);
nand U20950 (N_20950,N_17423,N_16582);
and U20951 (N_20951,N_16484,N_15143);
nand U20952 (N_20952,N_15908,N_17956);
nand U20953 (N_20953,N_16897,N_15123);
xor U20954 (N_20954,N_15606,N_17001);
nor U20955 (N_20955,N_16455,N_16354);
nor U20956 (N_20956,N_15493,N_15732);
nand U20957 (N_20957,N_17437,N_15394);
nor U20958 (N_20958,N_15528,N_15059);
or U20959 (N_20959,N_16781,N_16787);
nor U20960 (N_20960,N_16365,N_16616);
nand U20961 (N_20961,N_15688,N_15624);
nand U20962 (N_20962,N_15691,N_15772);
nand U20963 (N_20963,N_17489,N_17870);
nand U20964 (N_20964,N_16550,N_17555);
and U20965 (N_20965,N_15096,N_16913);
or U20966 (N_20966,N_16009,N_17078);
xnor U20967 (N_20967,N_15505,N_15218);
nor U20968 (N_20968,N_16196,N_15135);
or U20969 (N_20969,N_16349,N_17277);
and U20970 (N_20970,N_16049,N_16105);
or U20971 (N_20971,N_16346,N_17058);
nand U20972 (N_20972,N_16705,N_15363);
and U20973 (N_20973,N_15990,N_15666);
nand U20974 (N_20974,N_17191,N_15234);
and U20975 (N_20975,N_16692,N_17779);
nand U20976 (N_20976,N_16848,N_16408);
nor U20977 (N_20977,N_16912,N_16162);
or U20978 (N_20978,N_15425,N_16951);
or U20979 (N_20979,N_15649,N_17386);
nor U20980 (N_20980,N_17272,N_16625);
nand U20981 (N_20981,N_15617,N_15628);
and U20982 (N_20982,N_15212,N_17996);
nor U20983 (N_20983,N_17262,N_15946);
xor U20984 (N_20984,N_16334,N_15487);
nor U20985 (N_20985,N_16651,N_15504);
or U20986 (N_20986,N_17858,N_17259);
nand U20987 (N_20987,N_15081,N_17015);
nor U20988 (N_20988,N_17860,N_17145);
nand U20989 (N_20989,N_16714,N_16920);
nand U20990 (N_20990,N_16458,N_16536);
and U20991 (N_20991,N_16480,N_17856);
nand U20992 (N_20992,N_16250,N_17977);
nor U20993 (N_20993,N_17106,N_17361);
xor U20994 (N_20994,N_15080,N_15676);
nand U20995 (N_20995,N_16428,N_16239);
xor U20996 (N_20996,N_15292,N_15091);
nand U20997 (N_20997,N_17356,N_17841);
and U20998 (N_20998,N_15189,N_16883);
nand U20999 (N_20999,N_15953,N_17766);
nor U21000 (N_21000,N_20149,N_18209);
or U21001 (N_21001,N_19087,N_20059);
nor U21002 (N_21002,N_20005,N_18363);
xnor U21003 (N_21003,N_19484,N_18996);
or U21004 (N_21004,N_18952,N_19657);
nor U21005 (N_21005,N_18116,N_19521);
xor U21006 (N_21006,N_20802,N_18678);
xor U21007 (N_21007,N_20848,N_18989);
or U21008 (N_21008,N_20258,N_18111);
nand U21009 (N_21009,N_18080,N_18014);
or U21010 (N_21010,N_18763,N_19110);
or U21011 (N_21011,N_19019,N_20702);
nor U21012 (N_21012,N_19530,N_18561);
nand U21013 (N_21013,N_20766,N_19612);
nor U21014 (N_21014,N_20656,N_19046);
or U21015 (N_21015,N_18956,N_18479);
xnor U21016 (N_21016,N_18125,N_20754);
nand U21017 (N_21017,N_19355,N_19440);
nand U21018 (N_21018,N_20081,N_18666);
nand U21019 (N_21019,N_20763,N_18445);
nand U21020 (N_21020,N_18260,N_20071);
nand U21021 (N_21021,N_18647,N_18810);
nand U21022 (N_21022,N_19899,N_18423);
xnor U21023 (N_21023,N_20843,N_18041);
and U21024 (N_21024,N_18685,N_19061);
or U21025 (N_21025,N_20202,N_19838);
and U21026 (N_21026,N_20811,N_19850);
xnor U21027 (N_21027,N_18292,N_18094);
and U21028 (N_21028,N_20490,N_20627);
or U21029 (N_21029,N_18305,N_20900);
xnor U21030 (N_21030,N_20143,N_20680);
and U21031 (N_21031,N_20929,N_20123);
nand U21032 (N_21032,N_19175,N_19207);
and U21033 (N_21033,N_19450,N_20536);
and U21034 (N_21034,N_19621,N_19870);
nand U21035 (N_21035,N_19787,N_18715);
nand U21036 (N_21036,N_19893,N_18807);
nor U21037 (N_21037,N_20065,N_19684);
xor U21038 (N_21038,N_18833,N_19430);
or U21039 (N_21039,N_19610,N_20860);
or U21040 (N_21040,N_18386,N_19401);
and U21041 (N_21041,N_19834,N_19723);
xnor U21042 (N_21042,N_18006,N_18454);
nor U21043 (N_21043,N_18039,N_19068);
and U21044 (N_21044,N_19164,N_19976);
xor U21045 (N_21045,N_20155,N_18540);
nor U21046 (N_21046,N_19362,N_20245);
nor U21047 (N_21047,N_20611,N_19736);
nor U21048 (N_21048,N_19074,N_18299);
nor U21049 (N_21049,N_18916,N_20338);
nand U21050 (N_21050,N_19921,N_19309);
or U21051 (N_21051,N_18408,N_20376);
nor U21052 (N_21052,N_19597,N_19528);
and U21053 (N_21053,N_20320,N_18905);
or U21054 (N_21054,N_18102,N_18017);
and U21055 (N_21055,N_19819,N_18681);
nand U21056 (N_21056,N_20000,N_18696);
and U21057 (N_21057,N_20344,N_20184);
and U21058 (N_21058,N_18473,N_18107);
nand U21059 (N_21059,N_18573,N_20664);
or U21060 (N_21060,N_19457,N_19849);
nor U21061 (N_21061,N_18712,N_18320);
nor U21062 (N_21062,N_20021,N_19713);
or U21063 (N_21063,N_18166,N_19628);
or U21064 (N_21064,N_19885,N_20046);
and U21065 (N_21065,N_19718,N_18227);
nand U21066 (N_21066,N_20424,N_18021);
or U21067 (N_21067,N_20354,N_20359);
nand U21068 (N_21068,N_20989,N_19947);
and U21069 (N_21069,N_18372,N_19459);
or U21070 (N_21070,N_18362,N_19318);
xnor U21071 (N_21071,N_20417,N_20820);
and U21072 (N_21072,N_18951,N_20215);
nor U21073 (N_21073,N_19384,N_18512);
or U21074 (N_21074,N_19030,N_18811);
nand U21075 (N_21075,N_20581,N_19800);
and U21076 (N_21076,N_19872,N_18237);
nand U21077 (N_21077,N_18564,N_19648);
nand U21078 (N_21078,N_18592,N_20412);
nor U21079 (N_21079,N_18649,N_20111);
xor U21080 (N_21080,N_19058,N_19571);
or U21081 (N_21081,N_18694,N_18535);
xnor U21082 (N_21082,N_18353,N_20995);
xor U21083 (N_21083,N_20119,N_19176);
xnor U21084 (N_21084,N_18067,N_18603);
nor U21085 (N_21085,N_20661,N_19351);
xor U21086 (N_21086,N_20686,N_20604);
nor U21087 (N_21087,N_19620,N_19290);
or U21088 (N_21088,N_19428,N_19051);
and U21089 (N_21089,N_18528,N_20413);
xnor U21090 (N_21090,N_18416,N_19367);
nand U21091 (N_21091,N_20431,N_19514);
and U21092 (N_21092,N_20363,N_20899);
nor U21093 (N_21093,N_18691,N_18848);
nor U21094 (N_21094,N_20148,N_19063);
xor U21095 (N_21095,N_20284,N_20409);
and U21096 (N_21096,N_19577,N_18218);
xor U21097 (N_21097,N_20550,N_19879);
nand U21098 (N_21098,N_18663,N_20405);
xnor U21099 (N_21099,N_18293,N_20554);
xor U21100 (N_21100,N_18387,N_18341);
and U21101 (N_21101,N_18967,N_19468);
nand U21102 (N_21102,N_19288,N_19234);
nand U21103 (N_21103,N_19582,N_18314);
or U21104 (N_21104,N_18415,N_19762);
nor U21105 (N_21105,N_20573,N_20404);
and U21106 (N_21106,N_18627,N_20523);
and U21107 (N_21107,N_19091,N_18259);
xnor U21108 (N_21108,N_19790,N_18802);
and U21109 (N_21109,N_18994,N_19499);
nand U21110 (N_21110,N_18165,N_20542);
and U21111 (N_21111,N_18104,N_20653);
or U21112 (N_21112,N_20788,N_20122);
nor U21113 (N_21113,N_19596,N_20855);
nand U21114 (N_21114,N_20785,N_20677);
nand U21115 (N_21115,N_19174,N_18239);
or U21116 (N_21116,N_19845,N_18539);
and U21117 (N_21117,N_18901,N_18674);
and U21118 (N_21118,N_20027,N_20538);
or U21119 (N_21119,N_19279,N_19554);
nand U21120 (N_21120,N_20817,N_20952);
xor U21121 (N_21121,N_18171,N_18906);
or U21122 (N_21122,N_20243,N_20017);
xor U21123 (N_21123,N_20458,N_18448);
and U21124 (N_21124,N_18738,N_18949);
and U21125 (N_21125,N_20968,N_20369);
xor U21126 (N_21126,N_18709,N_19121);
and U21127 (N_21127,N_19922,N_20316);
xor U21128 (N_21128,N_18378,N_19996);
nor U21129 (N_21129,N_20084,N_19746);
nand U21130 (N_21130,N_19203,N_18370);
and U21131 (N_21131,N_18861,N_18894);
nand U21132 (N_21132,N_20662,N_19296);
xnor U21133 (N_21133,N_20882,N_18354);
nand U21134 (N_21134,N_19465,N_19536);
and U21135 (N_21135,N_20399,N_20827);
nand U21136 (N_21136,N_19667,N_20228);
nor U21137 (N_21137,N_19520,N_20553);
and U21138 (N_21138,N_18523,N_20673);
or U21139 (N_21139,N_20225,N_19890);
or U21140 (N_21140,N_20714,N_20566);
nand U21141 (N_21141,N_18971,N_19054);
and U21142 (N_21142,N_20274,N_19044);
or U21143 (N_21143,N_20290,N_18244);
nor U21144 (N_21144,N_18915,N_20312);
and U21145 (N_21145,N_19122,N_20837);
xor U21146 (N_21146,N_19389,N_20423);
or U21147 (N_21147,N_18112,N_19316);
nand U21148 (N_21148,N_20339,N_18163);
nand U21149 (N_21149,N_19274,N_20346);
nor U21150 (N_21150,N_19242,N_19509);
xor U21151 (N_21151,N_20500,N_20620);
and U21152 (N_21152,N_20983,N_18789);
nor U21153 (N_21153,N_18824,N_19353);
and U21154 (N_21154,N_20194,N_20772);
and U21155 (N_21155,N_19263,N_18505);
or U21156 (N_21156,N_19594,N_20138);
xor U21157 (N_21157,N_19154,N_18957);
xor U21158 (N_21158,N_18657,N_18942);
xor U21159 (N_21159,N_18057,N_19625);
or U21160 (N_21160,N_19972,N_20237);
and U21161 (N_21161,N_19480,N_19140);
or U21162 (N_21162,N_19780,N_20925);
and U21163 (N_21163,N_20305,N_20188);
and U21164 (N_21164,N_19150,N_20422);
or U21165 (N_21165,N_19265,N_20307);
nor U21166 (N_21166,N_19130,N_18889);
nor U21167 (N_21167,N_20246,N_20161);
and U21168 (N_21168,N_18913,N_18404);
nor U21169 (N_21169,N_20966,N_18725);
nor U21170 (N_21170,N_18149,N_18365);
and U21171 (N_21171,N_20867,N_20883);
xnor U21172 (N_21172,N_18297,N_20833);
xnor U21173 (N_21173,N_20878,N_19075);
or U21174 (N_21174,N_20561,N_20019);
or U21175 (N_21175,N_19337,N_20715);
nand U21176 (N_21176,N_20321,N_19682);
nand U21177 (N_21177,N_20574,N_20247);
xor U21178 (N_21178,N_19171,N_19519);
xor U21179 (N_21179,N_18975,N_20341);
nand U21180 (N_21180,N_19772,N_20951);
xnor U21181 (N_21181,N_19705,N_18780);
or U21182 (N_21182,N_19675,N_20251);
or U21183 (N_21183,N_20986,N_20777);
nand U21184 (N_21184,N_18252,N_20740);
nor U21185 (N_21185,N_20541,N_18938);
xor U21186 (N_21186,N_18834,N_20803);
nor U21187 (N_21187,N_19936,N_18823);
xnor U21188 (N_21188,N_19141,N_18108);
xor U21189 (N_21189,N_18818,N_18472);
nor U21190 (N_21190,N_18839,N_19711);
xor U21191 (N_21191,N_19848,N_18958);
or U21192 (N_21192,N_18702,N_20804);
and U21193 (N_21193,N_18250,N_20999);
xor U21194 (N_21194,N_19617,N_19832);
or U21195 (N_21195,N_20436,N_18753);
or U21196 (N_21196,N_19956,N_18424);
or U21197 (N_21197,N_19760,N_18869);
xnor U21198 (N_21198,N_19844,N_18455);
xor U21199 (N_21199,N_20825,N_19346);
nor U21200 (N_21200,N_20203,N_18434);
nand U21201 (N_21201,N_20594,N_18483);
xor U21202 (N_21202,N_20061,N_20041);
and U21203 (N_21203,N_19204,N_20637);
nand U21204 (N_21204,N_19822,N_19402);
or U21205 (N_21205,N_18706,N_19634);
nand U21206 (N_21206,N_20643,N_19754);
nand U21207 (N_21207,N_18837,N_18574);
or U21208 (N_21208,N_20013,N_20921);
and U21209 (N_21209,N_19877,N_20231);
and U21210 (N_21210,N_18337,N_19314);
or U21211 (N_21211,N_18055,N_19418);
nand U21212 (N_21212,N_20419,N_19456);
and U21213 (N_21213,N_19205,N_19359);
xnor U21214 (N_21214,N_18462,N_18632);
and U21215 (N_21215,N_20014,N_20414);
nand U21216 (N_21216,N_18150,N_19120);
xor U21217 (N_21217,N_19920,N_20216);
nor U21218 (N_21218,N_18376,N_19502);
or U21219 (N_21219,N_18982,N_20392);
xor U21220 (N_21220,N_19538,N_18233);
xor U21221 (N_21221,N_18096,N_19158);
xor U21222 (N_21222,N_20403,N_19285);
nor U21223 (N_21223,N_20515,N_18842);
nor U21224 (N_21224,N_18158,N_20390);
or U21225 (N_21225,N_18282,N_18182);
nand U21226 (N_21226,N_19949,N_20557);
nand U21227 (N_21227,N_20205,N_18127);
and U21228 (N_21228,N_19233,N_19769);
nand U21229 (N_21229,N_18984,N_20087);
or U21230 (N_21230,N_20963,N_18832);
or U21231 (N_21231,N_20514,N_18684);
or U21232 (N_21232,N_18911,N_19335);
and U21233 (N_21233,N_18413,N_18075);
nor U21234 (N_21234,N_19250,N_20336);
nand U21235 (N_21235,N_20908,N_19108);
nor U21236 (N_21236,N_19858,N_19761);
nand U21237 (N_21237,N_19157,N_18133);
and U21238 (N_21238,N_18480,N_19077);
and U21239 (N_21239,N_20654,N_18430);
and U21240 (N_21240,N_18411,N_18170);
nand U21241 (N_21241,N_18855,N_18746);
nor U21242 (N_21242,N_19574,N_18863);
or U21243 (N_21243,N_20296,N_20893);
or U21244 (N_21244,N_19312,N_20823);
and U21245 (N_21245,N_18486,N_19493);
xnor U21246 (N_21246,N_20310,N_20281);
nor U21247 (N_21247,N_20889,N_18331);
nand U21248 (N_21248,N_19276,N_20191);
or U21249 (N_21249,N_20475,N_20055);
nand U21250 (N_21250,N_18397,N_20004);
xnor U21251 (N_21251,N_20181,N_18587);
or U21252 (N_21252,N_20787,N_18526);
nand U21253 (N_21253,N_18966,N_18000);
nand U21254 (N_21254,N_18860,N_20576);
xor U21255 (N_21255,N_18608,N_20668);
and U21256 (N_21256,N_19286,N_20744);
xnor U21257 (N_21257,N_20020,N_19050);
or U21258 (N_21258,N_18446,N_18868);
and U21259 (N_21259,N_18936,N_20672);
xor U21260 (N_21260,N_20375,N_20998);
and U21261 (N_21261,N_19467,N_19038);
xor U21262 (N_21262,N_20992,N_19368);
xnor U21263 (N_21263,N_20374,N_18497);
nand U21264 (N_21264,N_20110,N_20224);
or U21265 (N_21265,N_20851,N_18114);
nor U21266 (N_21266,N_19891,N_18840);
nand U21267 (N_21267,N_20764,N_19706);
or U21268 (N_21268,N_18164,N_18676);
and U21269 (N_21269,N_18302,N_20497);
nor U21270 (N_21270,N_20208,N_18640);
nand U21271 (N_21271,N_20568,N_19636);
nand U21272 (N_21272,N_18760,N_18216);
or U21273 (N_21273,N_18719,N_18558);
nand U21274 (N_21274,N_18440,N_20189);
nand U21275 (N_21275,N_18503,N_20901);
or U21276 (N_21276,N_20845,N_19466);
nand U21277 (N_21277,N_19445,N_19100);
xor U21278 (N_21278,N_18826,N_19930);
nand U21279 (N_21279,N_19095,N_19869);
xor U21280 (N_21280,N_18447,N_19151);
nand U21281 (N_21281,N_18669,N_19585);
nor U21282 (N_21282,N_19173,N_20147);
xnor U21283 (N_21283,N_20166,N_18687);
or U21284 (N_21284,N_18582,N_19002);
nand U21285 (N_21285,N_19975,N_20979);
and U21286 (N_21286,N_19562,N_18658);
xor U21287 (N_21287,N_18286,N_18585);
nor U21288 (N_21288,N_20325,N_18972);
nand U21289 (N_21289,N_19918,N_18744);
or U21290 (N_21290,N_18531,N_18814);
xor U21291 (N_21291,N_20815,N_20552);
nand U21292 (N_21292,N_18101,N_18267);
nor U21293 (N_21293,N_19887,N_18374);
xnor U21294 (N_21294,N_20349,N_18619);
nor U21295 (N_21295,N_18279,N_19251);
and U21296 (N_21296,N_20578,N_20335);
xor U21297 (N_21297,N_19471,N_19994);
and U21298 (N_21298,N_18532,N_20612);
and U21299 (N_21299,N_20904,N_18110);
xnor U21300 (N_21300,N_18550,N_20253);
and U21301 (N_21301,N_19550,N_19488);
nand U21302 (N_21302,N_18697,N_19565);
nand U21303 (N_21303,N_20941,N_18510);
xnor U21304 (N_21304,N_18891,N_20731);
nand U21305 (N_21305,N_19511,N_18403);
nor U21306 (N_21306,N_18740,N_20076);
xor U21307 (N_21307,N_19661,N_20558);
or U21308 (N_21308,N_20563,N_20050);
nand U21309 (N_21309,N_19958,N_20355);
nor U21310 (N_21310,N_18401,N_19155);
xnor U21311 (N_21311,N_20660,N_19474);
or U21312 (N_21312,N_19375,N_19651);
xnor U21313 (N_21313,N_18226,N_18596);
xor U21314 (N_21314,N_20283,N_18867);
nor U21315 (N_21315,N_18143,N_19070);
nand U21316 (N_21316,N_19733,N_18886);
xnor U21317 (N_21317,N_19900,N_20476);
nand U21318 (N_21318,N_18169,N_18620);
nor U21319 (N_21319,N_20493,N_19454);
nor U21320 (N_21320,N_18529,N_18487);
and U21321 (N_21321,N_19576,N_20555);
and U21322 (N_21322,N_20547,N_20711);
and U21323 (N_21323,N_19386,N_18993);
and U21324 (N_21324,N_19256,N_19541);
nor U21325 (N_21325,N_20725,N_20728);
nor U21326 (N_21326,N_18935,N_20010);
or U21327 (N_21327,N_20154,N_20141);
nor U21328 (N_21328,N_18283,N_18659);
nor U21329 (N_21329,N_20306,N_19461);
and U21330 (N_21330,N_18008,N_19813);
nor U21331 (N_21331,N_20751,N_20749);
xor U21332 (N_21332,N_18634,N_19045);
or U21333 (N_21333,N_19567,N_20774);
and U21334 (N_21334,N_19939,N_19280);
xor U21335 (N_21335,N_20093,N_19348);
xor U21336 (N_21336,N_19794,N_19593);
or U21337 (N_21337,N_19752,N_18928);
and U21338 (N_21338,N_20796,N_20935);
nor U21339 (N_21339,N_18843,N_18326);
nor U21340 (N_21340,N_18074,N_19810);
nor U21341 (N_21341,N_18918,N_20142);
and U21342 (N_21342,N_20511,N_18323);
xor U21343 (N_21343,N_20330,N_20930);
and U21344 (N_21344,N_18650,N_19107);
nor U21345 (N_21345,N_20276,N_18546);
or U21346 (N_21346,N_19246,N_18545);
or U21347 (N_21347,N_19799,N_20539);
nor U21348 (N_21348,N_19017,N_19604);
nand U21349 (N_21349,N_18167,N_19808);
and U21350 (N_21350,N_20077,N_18764);
and U21351 (N_21351,N_18792,N_18191);
xnor U21352 (N_21352,N_18775,N_18513);
nand U21353 (N_21353,N_18849,N_18900);
nor U21354 (N_21354,N_20880,N_19609);
or U21355 (N_21355,N_20967,N_18741);
xnor U21356 (N_21356,N_20810,N_20256);
and U21357 (N_21357,N_20640,N_18670);
nand U21358 (N_21358,N_18138,N_20881);
or U21359 (N_21359,N_20844,N_18005);
and U21360 (N_21360,N_18072,N_18999);
and U21361 (N_21361,N_18973,N_20757);
and U21362 (N_21362,N_18425,N_18025);
nand U21363 (N_21363,N_18668,N_19886);
nand U21364 (N_21364,N_19543,N_19724);
nor U21365 (N_21365,N_19915,N_18334);
or U21366 (N_21366,N_18667,N_18082);
nor U21367 (N_21367,N_18895,N_18866);
nor U21368 (N_21368,N_19805,N_20759);
nand U21369 (N_21369,N_20875,N_20377);
and U21370 (N_21370,N_19267,N_20502);
nor U21371 (N_21371,N_19653,N_20970);
and U21372 (N_21372,N_18258,N_19340);
and U21373 (N_21373,N_20190,N_20795);
and U21374 (N_21374,N_19605,N_19964);
and U21375 (N_21375,N_19113,N_18607);
xnor U21376 (N_21376,N_20927,N_19277);
nand U21377 (N_21377,N_18452,N_20097);
and U21378 (N_21378,N_20758,N_20070);
xor U21379 (N_21379,N_20408,N_19708);
xor U21380 (N_21380,N_19134,N_18172);
or U21381 (N_21381,N_18909,N_19901);
nor U21382 (N_21382,N_18470,N_18004);
and U21383 (N_21383,N_19144,N_20703);
nor U21384 (N_21384,N_19181,N_19961);
nor U21385 (N_21385,N_20100,N_18943);
xor U21386 (N_21386,N_20674,N_19487);
nand U21387 (N_21387,N_20048,N_18042);
nand U21388 (N_21388,N_20863,N_18145);
nor U21389 (N_21389,N_19252,N_20736);
nor U21390 (N_21390,N_19298,N_18019);
and U21391 (N_21391,N_18405,N_18736);
nand U21392 (N_21392,N_18872,N_20364);
and U21393 (N_21393,N_18808,N_18638);
nand U21394 (N_21394,N_19435,N_18517);
nor U21395 (N_21395,N_18593,N_18793);
or U21396 (N_21396,N_19142,N_18393);
nor U21397 (N_21397,N_19331,N_20192);
xnor U21398 (N_21398,N_20615,N_18555);
nor U21399 (N_21399,N_18536,N_19236);
nor U21400 (N_21400,N_18129,N_18914);
or U21401 (N_21401,N_20508,N_19463);
xnor U21402 (N_21402,N_18466,N_18050);
xnor U21403 (N_21403,N_19944,N_20849);
nand U21404 (N_21404,N_19734,N_20426);
nand U21405 (N_21405,N_19965,N_19545);
and U21406 (N_21406,N_20721,N_18348);
and U21407 (N_21407,N_20486,N_20962);
nor U21408 (N_21408,N_18449,N_20261);
nor U21409 (N_21409,N_20768,N_18484);
nor U21410 (N_21410,N_18257,N_20314);
xnor U21411 (N_21411,N_20152,N_18247);
or U21412 (N_21412,N_18859,N_20445);
nor U21413 (N_21413,N_20478,N_19637);
xor U21414 (N_21414,N_18242,N_20540);
or U21415 (N_21415,N_18622,N_18502);
nand U21416 (N_21416,N_20869,N_19300);
nor U21417 (N_21417,N_20443,N_18439);
nand U21418 (N_21418,N_20808,N_18134);
xor U21419 (N_21419,N_18987,N_20971);
and U21420 (N_21420,N_19553,N_20226);
xnor U21421 (N_21421,N_18677,N_18930);
or U21422 (N_21422,N_19764,N_18752);
nor U21423 (N_21423,N_19307,N_20584);
xnor U21424 (N_21424,N_18174,N_19105);
or U21425 (N_21425,N_20895,N_20145);
xor U21426 (N_21426,N_19911,N_20183);
nor U21427 (N_21427,N_18369,N_18825);
nor U21428 (N_21428,N_20397,N_20572);
or U21429 (N_21429,N_19513,N_20974);
xor U21430 (N_21430,N_18481,N_20577);
nor U21431 (N_21431,N_18488,N_20201);
nor U21432 (N_21432,N_18965,N_20695);
nor U21433 (N_21433,N_20760,N_20864);
and U21434 (N_21434,N_18407,N_19037);
xnor U21435 (N_21435,N_20285,N_19152);
nor U21436 (N_21436,N_18309,N_18850);
nor U21437 (N_21437,N_18395,N_19627);
nor U21438 (N_21438,N_18318,N_19273);
nand U21439 (N_21439,N_18568,N_19365);
nand U21440 (N_21440,N_20433,N_18287);
and U21441 (N_21441,N_19913,N_20460);
nor U21442 (N_21442,N_18804,N_18076);
nor U21443 (N_21443,N_19327,N_18092);
and U21444 (N_21444,N_18519,N_19129);
xor U21445 (N_21445,N_19117,N_19618);
and U21446 (N_21446,N_20273,N_20300);
or U21447 (N_21447,N_18576,N_19977);
nor U21448 (N_21448,N_19725,N_18713);
nand U21449 (N_21449,N_20272,N_19052);
or U21450 (N_21450,N_18051,N_19629);
nand U21451 (N_21451,N_20856,N_18921);
or U21452 (N_21452,N_20726,N_19559);
and U21453 (N_21453,N_19674,N_19592);
nor U21454 (N_21454,N_18128,N_20832);
nor U21455 (N_21455,N_20733,N_18155);
xnor U21456 (N_21456,N_19426,N_18782);
and U21457 (N_21457,N_19504,N_20678);
nand U21458 (N_21458,N_18360,N_18224);
xnor U21459 (N_21459,N_18817,N_19506);
and U21460 (N_21460,N_20126,N_18594);
xor U21461 (N_21461,N_20260,N_19540);
and U21462 (N_21462,N_20168,N_19161);
or U21463 (N_21463,N_20133,N_20692);
or U21464 (N_21464,N_20955,N_19168);
and U21465 (N_21465,N_19243,N_19906);
xor U21466 (N_21466,N_20386,N_20708);
and U21467 (N_21467,N_19012,N_20473);
or U21468 (N_21468,N_18489,N_18419);
and U21469 (N_21469,N_19115,N_19059);
and U21470 (N_21470,N_18181,N_20988);
nor U21471 (N_21471,N_18241,N_18986);
or U21472 (N_21472,N_18053,N_20337);
and U21473 (N_21473,N_19929,N_19581);
and U21474 (N_21474,N_19926,N_19735);
or U21475 (N_21475,N_18500,N_20079);
xor U21476 (N_21476,N_20469,N_18245);
or U21477 (N_21477,N_19833,N_18195);
or U21478 (N_21478,N_20689,N_18788);
nand U21479 (N_21479,N_18106,N_19908);
nor U21480 (N_21480,N_18893,N_19195);
nand U21481 (N_21481,N_18152,N_18321);
xor U21482 (N_21482,N_19579,N_20452);
and U21483 (N_21483,N_19614,N_20297);
nor U21484 (N_21484,N_20470,N_19392);
nand U21485 (N_21485,N_19694,N_19013);
nor U21486 (N_21486,N_20602,N_18277);
or U21487 (N_21487,N_20829,N_18841);
and U21488 (N_21488,N_19334,N_18530);
nand U21489 (N_21489,N_19730,N_20938);
nand U21490 (N_21490,N_18431,N_18049);
nor U21491 (N_21491,N_18566,N_20984);
nor U21492 (N_21492,N_18621,N_20852);
and U21493 (N_21493,N_20214,N_19721);
and U21494 (N_21494,N_19957,N_20915);
xor U21495 (N_21495,N_19678,N_18997);
and U21496 (N_21496,N_18838,N_19497);
nor U21497 (N_21497,N_20537,N_18361);
xor U21498 (N_21498,N_19971,N_20366);
nand U21499 (N_21499,N_20543,N_19967);
nand U21500 (N_21500,N_20533,N_19919);
and U21501 (N_21501,N_18240,N_19272);
nand U21502 (N_21502,N_18007,N_18828);
nor U21503 (N_21503,N_18235,N_20813);
xnor U21504 (N_21504,N_20448,N_18246);
or U21505 (N_21505,N_19518,N_18924);
xor U21506 (N_21506,N_19624,N_19998);
nand U21507 (N_21507,N_18506,N_20230);
nand U21508 (N_21508,N_20780,N_20472);
nor U21509 (N_21509,N_19479,N_19112);
and U21510 (N_21510,N_18148,N_19015);
nor U21511 (N_21511,N_20569,N_19162);
and U21512 (N_21512,N_19874,N_20373);
and U21513 (N_21513,N_19685,N_19671);
or U21514 (N_21514,N_19807,N_20911);
nor U21515 (N_21515,N_19222,N_20741);
or U21516 (N_21516,N_19160,N_18325);
or U21517 (N_21517,N_20451,N_19380);
nor U21518 (N_21518,N_18024,N_19925);
xor U21519 (N_21519,N_20965,N_19768);
and U21520 (N_21520,N_19910,N_20350);
nand U21521 (N_21521,N_18047,N_20663);
nor U21522 (N_21522,N_18016,N_20480);
xnor U21523 (N_21523,N_19186,N_19404);
xnor U21524 (N_21524,N_19599,N_20199);
xnor U21525 (N_21525,N_19003,N_20564);
nor U21526 (N_21526,N_19086,N_18606);
xnor U21527 (N_21527,N_20635,N_20873);
xor U21528 (N_21528,N_18873,N_20607);
or U21529 (N_21529,N_19345,N_20106);
or U21530 (N_21530,N_19793,N_19644);
and U21531 (N_21531,N_20464,N_20343);
nand U21532 (N_21532,N_18995,N_20991);
xor U21533 (N_21533,N_19544,N_18645);
nand U21534 (N_21534,N_20716,N_20806);
and U21535 (N_21535,N_20614,N_20610);
nand U21536 (N_21536,N_19744,N_20091);
nand U21537 (N_21537,N_18482,N_18743);
and U21538 (N_21538,N_20854,N_18623);
or U21539 (N_21539,N_20858,N_20068);
nor U21540 (N_21540,N_18056,N_19235);
or U21541 (N_21541,N_20114,N_18180);
nor U21542 (N_21542,N_19098,N_18979);
nand U21543 (N_21543,N_20380,N_19639);
xnor U21544 (N_21544,N_19294,N_20108);
or U21545 (N_21545,N_20559,N_20370);
nand U21546 (N_21546,N_19374,N_19570);
or U21547 (N_21547,N_19261,N_18346);
and U21548 (N_21548,N_18926,N_20116);
nand U21549 (N_21549,N_19601,N_20358);
nor U21550 (N_21550,N_18198,N_19219);
or U21551 (N_21551,N_18980,N_18761);
and U21552 (N_21552,N_18060,N_20322);
nor U21553 (N_21553,N_19000,N_18123);
xnor U21554 (N_21554,N_18686,N_20029);
xor U21555 (N_21555,N_20179,N_18813);
xnor U21556 (N_21556,N_20720,N_20738);
nor U21557 (N_21557,N_19770,N_20289);
and U21558 (N_21558,N_20709,N_20428);
nor U21559 (N_21559,N_19783,N_19909);
and U21560 (N_21560,N_18160,N_20159);
or U21561 (N_21561,N_20688,N_18070);
nor U21562 (N_21562,N_18421,N_19476);
nor U21563 (N_21563,N_19410,N_18990);
or U21564 (N_21564,N_18144,N_18192);
nand U21565 (N_21565,N_20799,N_19189);
or U21566 (N_21566,N_20007,N_18892);
nand U21567 (N_21567,N_20682,N_20069);
nor U21568 (N_21568,N_18272,N_20579);
nor U21569 (N_21569,N_20313,N_19271);
or U21570 (N_21570,N_20888,N_20826);
xnor U21571 (N_21571,N_20924,N_19361);
nand U21572 (N_21572,N_19253,N_18562);
xnor U21573 (N_21573,N_20195,N_19992);
nor U21574 (N_21574,N_18551,N_20121);
nor U21575 (N_21575,N_18249,N_18151);
and U21576 (N_21576,N_19875,N_18600);
and U21577 (N_21577,N_20990,N_20582);
or U21578 (N_21578,N_18700,N_18727);
or U21579 (N_21579,N_20649,N_20421);
nor U21580 (N_21580,N_18208,N_20269);
xor U21581 (N_21581,N_20128,N_19633);
and U21582 (N_21582,N_18950,N_20870);
and U21583 (N_21583,N_19704,N_18307);
and U21584 (N_21584,N_18812,N_20402);
or U21585 (N_21585,N_19319,N_19281);
nor U21586 (N_21586,N_18091,N_19275);
nand U21587 (N_21587,N_19710,N_20964);
or U21588 (N_21588,N_20850,N_20646);
nor U21589 (N_21589,N_19914,N_19873);
nand U21590 (N_21590,N_18858,N_18460);
xor U21591 (N_21591,N_19011,N_20934);
xnor U21592 (N_21592,N_19446,N_18953);
nor U21593 (N_21593,N_18547,N_18754);
and U21594 (N_21594,N_18864,N_18073);
and U21595 (N_21595,N_20887,N_19356);
xnor U21596 (N_21596,N_20909,N_18710);
nand U21597 (N_21597,N_18265,N_18013);
and U21598 (N_21598,N_19515,N_20427);
nand U21599 (N_21599,N_20588,N_18580);
or U21600 (N_21600,N_20494,N_20903);
nor U21601 (N_21601,N_20248,N_20236);
and U21602 (N_21602,N_19933,N_20471);
and U21603 (N_21603,N_18992,N_18219);
and U21604 (N_21604,N_19215,N_19424);
nand U21605 (N_21605,N_19194,N_19691);
and U21606 (N_21606,N_20619,N_20288);
xnor U21607 (N_21607,N_20894,N_19049);
and U21608 (N_21608,N_20841,N_18437);
and U21609 (N_21609,N_19485,N_18306);
nor U21610 (N_21610,N_19608,N_19436);
and U21611 (N_21611,N_18961,N_18022);
nand U21612 (N_21612,N_18015,N_19131);
and U21613 (N_21613,N_19983,N_18147);
xor U21614 (N_21614,N_19935,N_20645);
nand U21615 (N_21615,N_20266,N_18162);
nand U21616 (N_21616,N_19212,N_20389);
xor U21617 (N_21617,N_19820,N_18698);
nand U21618 (N_21618,N_18998,N_20042);
nand U21619 (N_21619,N_19007,N_19741);
nor U21620 (N_21620,N_19434,N_18368);
xnor U21621 (N_21621,N_20210,N_19237);
nor U21622 (N_21622,N_20522,N_19473);
and U21623 (N_21623,N_19496,N_19963);
nand U21624 (N_21624,N_18830,N_19357);
nor U21625 (N_21625,N_19383,N_19857);
nand U21626 (N_21626,N_20585,N_20846);
nor U21627 (N_21627,N_18829,N_20118);
nor U21628 (N_21628,N_20771,N_20008);
or U21629 (N_21629,N_19630,N_20838);
or U21630 (N_21630,N_18578,N_18945);
nand U21631 (N_21631,N_18090,N_18052);
xor U21632 (N_21632,N_18498,N_18255);
xor U21633 (N_21633,N_20509,N_18173);
nand U21634 (N_21634,N_20223,N_19756);
and U21635 (N_21635,N_20498,N_20099);
and U21636 (N_21636,N_19864,N_19505);
xor U21637 (N_21637,N_18494,N_19381);
or U21638 (N_21638,N_19643,N_19638);
and U21639 (N_21639,N_20626,N_20016);
or U21640 (N_21640,N_20734,N_18471);
nand U21641 (N_21641,N_19092,N_19245);
nor U21642 (N_21642,N_18068,N_18071);
and U21643 (N_21643,N_20876,N_19689);
xnor U21644 (N_21644,N_18396,N_20271);
nor U21645 (N_21645,N_20270,N_19247);
and U21646 (N_21646,N_19923,N_20078);
xnor U21647 (N_21647,N_19025,N_20756);
or U21648 (N_21648,N_20442,N_20605);
nand U21649 (N_21649,N_18294,N_19449);
nand U21650 (N_21650,N_20367,N_20931);
nand U21651 (N_21651,N_20006,N_20765);
nand U21652 (N_21652,N_18786,N_20437);
xor U21653 (N_21653,N_18029,N_19697);
or U21654 (N_21654,N_18981,N_18137);
xnor U21655 (N_21655,N_19895,N_20124);
and U21656 (N_21656,N_19884,N_18878);
xnor U21657 (N_21657,N_18313,N_19672);
nor U21658 (N_21658,N_20528,N_18617);
or U21659 (N_21659,N_18364,N_18771);
nand U21660 (N_21660,N_18382,N_19184);
or U21661 (N_21661,N_20311,N_18153);
or U21662 (N_21662,N_18748,N_18827);
nand U21663 (N_21663,N_18204,N_19740);
xnor U21664 (N_21664,N_18874,N_19987);
xnor U21665 (N_21665,N_19517,N_20063);
xnor U21666 (N_21666,N_20836,N_20054);
nor U21667 (N_21667,N_20356,N_18085);
xor U21668 (N_21668,N_18507,N_18714);
or U21669 (N_21669,N_19358,N_20907);
and U21670 (N_21670,N_20665,N_18845);
or U21671 (N_21671,N_19322,N_20510);
xor U21672 (N_21672,N_19221,N_20357);
nand U21673 (N_21673,N_19525,N_18871);
or U21674 (N_21674,N_20022,N_18962);
and U21675 (N_21675,N_18777,N_18345);
nand U21676 (N_21676,N_18630,N_19460);
nor U21677 (N_21677,N_18876,N_18350);
nor U21678 (N_21678,N_19425,N_19178);
nand U21679 (N_21679,N_20801,N_19081);
or U21680 (N_21680,N_20629,N_19111);
and U21681 (N_21681,N_19677,N_18046);
nand U21682 (N_21682,N_20919,N_20707);
and U21683 (N_21683,N_20752,N_19417);
nand U21684 (N_21684,N_18554,N_19403);
xor U21685 (N_21685,N_19293,N_18816);
or U21686 (N_21686,N_19508,N_19244);
nand U21687 (N_21687,N_20861,N_19227);
xor U21688 (N_21688,N_18624,N_20696);
or U21689 (N_21689,N_19606,N_18210);
nor U21690 (N_21690,N_18009,N_20450);
and U21691 (N_21691,N_18538,N_19680);
nor U21692 (N_21692,N_18038,N_19719);
nor U21693 (N_21693,N_20229,N_20135);
nor U21694 (N_21694,N_19882,N_20853);
xor U21695 (N_21695,N_19336,N_20565);
nor U21696 (N_21696,N_18176,N_20685);
nand U21697 (N_21697,N_20302,N_19622);
xnor U21698 (N_21698,N_20267,N_19116);
or U21699 (N_21699,N_18351,N_20291);
xnor U21700 (N_21700,N_19934,N_18194);
or U21701 (N_21701,N_18774,N_18983);
and U21702 (N_21702,N_20683,N_20748);
xor U21703 (N_21703,N_20221,N_19344);
xnor U21704 (N_21704,N_19489,N_20319);
nor U21705 (N_21705,N_18642,N_18904);
or U21706 (N_21706,N_20279,N_19148);
or U21707 (N_21707,N_20342,N_19777);
and U21708 (N_21708,N_18444,N_20747);
or U21709 (N_21709,N_18140,N_19470);
xnor U21710 (N_21710,N_20792,N_18105);
nor U21711 (N_21711,N_20015,N_20507);
xor U21712 (N_21712,N_19343,N_19586);
and U21713 (N_21713,N_19533,N_19670);
xnor U21714 (N_21714,N_18520,N_20975);
and U21715 (N_21715,N_18319,N_19532);
nor U21716 (N_21716,N_20567,N_20529);
or U21717 (N_21717,N_18214,N_18790);
xnor U21718 (N_21718,N_20468,N_19647);
or U21719 (N_21719,N_19867,N_18394);
and U21720 (N_21720,N_19619,N_19224);
or U21721 (N_21721,N_19206,N_19902);
and U21722 (N_21722,N_19220,N_18335);
xnor U21723 (N_21723,N_18784,N_19478);
and U21724 (N_21724,N_18063,N_20781);
xor U21725 (N_21725,N_19812,N_20939);
or U21726 (N_21726,N_20044,N_18040);
nor U21727 (N_21727,N_19325,N_18625);
nand U21728 (N_21728,N_20890,N_19659);
nand U21729 (N_21729,N_19945,N_19196);
and U21730 (N_21730,N_20681,N_18504);
xor U21731 (N_21731,N_20718,N_18679);
nor U21732 (N_21732,N_18660,N_18602);
nand U21733 (N_21733,N_20517,N_18095);
and U21734 (N_21734,N_20217,N_20286);
and U21735 (N_21735,N_20308,N_18932);
nand U21736 (N_21736,N_19654,N_19163);
or U21737 (N_21737,N_20329,N_19492);
xor U21738 (N_21738,N_18135,N_20254);
nor U21739 (N_21739,N_18117,N_20655);
and U21740 (N_21740,N_20457,N_18010);
or U21741 (N_21741,N_18796,N_19385);
xor U21742 (N_21742,N_19500,N_18084);
nor U21743 (N_21743,N_18877,N_18549);
or U21744 (N_21744,N_20842,N_19803);
nand U21745 (N_21745,N_19198,N_20847);
nand U21746 (N_21746,N_19749,N_19228);
or U21747 (N_21747,N_19818,N_19066);
nand U21748 (N_21748,N_20884,N_20137);
or U21749 (N_21749,N_19193,N_18200);
nor U21750 (N_21750,N_20105,N_20621);
xor U21751 (N_21751,N_18835,N_18762);
nand U21752 (N_21752,N_19714,N_19603);
nand U21753 (N_21753,N_19557,N_19974);
nand U21754 (N_21754,N_20043,N_18963);
nand U21755 (N_21755,N_18815,N_19048);
nand U21756 (N_21756,N_19165,N_19103);
or U21757 (N_21757,N_20011,N_19982);
or U21758 (N_21758,N_18389,N_19715);
or U21759 (N_21759,N_19871,N_20130);
xor U21760 (N_21760,N_19916,N_19208);
xor U21761 (N_21761,N_18723,N_20659);
xor U21762 (N_21762,N_18937,N_20031);
and U21763 (N_21763,N_19156,N_18159);
nand U21764 (N_21764,N_19414,N_19774);
or U21765 (N_21765,N_18119,N_18342);
nor U21766 (N_21766,N_19411,N_18616);
or U21767 (N_21767,N_18189,N_18367);
nand U21768 (N_21768,N_18717,N_19510);
xor U21769 (N_21769,N_19709,N_18595);
and U21770 (N_21770,N_18977,N_18865);
xor U21771 (N_21771,N_19067,N_20255);
xor U21772 (N_21772,N_20400,N_20944);
nor U21773 (N_21773,N_20171,N_20315);
nand U21774 (N_21774,N_19124,N_18605);
nand U21775 (N_21775,N_20178,N_19836);
or U21776 (N_21776,N_18328,N_20047);
or U21777 (N_21777,N_20560,N_19408);
nand U21778 (N_21778,N_20292,N_18034);
or U21779 (N_21779,N_19123,N_18718);
and U21780 (N_21780,N_18079,N_19432);
or U21781 (N_21781,N_19778,N_19213);
nor U21782 (N_21782,N_18799,N_19753);
and U21783 (N_21783,N_18922,N_19767);
nor U21784 (N_21784,N_18797,N_20958);
nand U21785 (N_21785,N_18311,N_19094);
and U21786 (N_21786,N_18896,N_20282);
or U21787 (N_21787,N_20455,N_20461);
xor U21788 (N_21788,N_20499,N_19082);
or U21789 (N_21789,N_19865,N_20036);
and U21790 (N_21790,N_18575,N_19824);
nor U21791 (N_21791,N_18854,N_18944);
and U21792 (N_21792,N_20694,N_20033);
nand U21793 (N_21793,N_18641,N_20805);
nand U21794 (N_21794,N_20474,N_19306);
nor U21795 (N_21795,N_20198,N_18254);
and U21796 (N_21796,N_20092,N_18541);
nand U21797 (N_21797,N_18183,N_19370);
xnor U21798 (N_21798,N_20932,N_20519);
nor U21799 (N_21799,N_20395,N_19016);
or U21800 (N_21800,N_20429,N_19024);
and U21801 (N_21801,N_18820,N_19702);
nand U21802 (N_21802,N_18238,N_18384);
nor U21803 (N_21803,N_18043,N_20082);
nand U21804 (N_21804,N_19283,N_19185);
nand U21805 (N_21805,N_20710,N_18707);
and U21806 (N_21806,N_18589,N_18457);
or U21807 (N_21807,N_18653,N_20959);
and U21808 (N_21808,N_19377,N_19372);
or U21809 (N_21809,N_18186,N_20551);
and U21810 (N_21810,N_19785,N_18491);
nor U21811 (N_21811,N_18635,N_18801);
xor U21812 (N_21812,N_20318,N_19595);
or U21813 (N_21813,N_19257,N_20024);
and U21814 (N_21814,N_19026,N_20323);
and U21815 (N_21815,N_18045,N_18441);
or U21816 (N_21816,N_18373,N_20616);
and U21817 (N_21817,N_19262,N_18093);
or U21818 (N_21818,N_19060,N_19311);
or U21819 (N_21819,N_20613,N_19759);
nor U21820 (N_21820,N_20704,N_20298);
and U21821 (N_21821,N_18450,N_18232);
nand U21822 (N_21822,N_20238,N_20441);
xor U21823 (N_21823,N_20232,N_19249);
nand U21824 (N_21824,N_20956,N_18730);
and U21825 (N_21825,N_18190,N_20327);
nor U21826 (N_21826,N_18948,N_19655);
or U21827 (N_21827,N_19631,N_18610);
or U21828 (N_21828,N_20489,N_19320);
or U21829 (N_21829,N_19031,N_20032);
nor U21830 (N_21830,N_18103,N_19940);
and U21831 (N_21831,N_20712,N_18857);
or U21832 (N_21832,N_18643,N_19959);
nand U21833 (N_21833,N_19814,N_18509);
xnor U21834 (N_21834,N_19692,N_20362);
and U21835 (N_21835,N_18661,N_19575);
and U21836 (N_21836,N_19782,N_19966);
xor U21837 (N_21837,N_19429,N_18584);
nor U21838 (N_21838,N_18356,N_19376);
xor U21839 (N_21839,N_19989,N_19907);
or U21840 (N_21840,N_19928,N_19223);
nand U21841 (N_21841,N_20617,N_20920);
and U21842 (N_21842,N_20053,N_18298);
and U21843 (N_21843,N_18193,N_19695);
xor U21844 (N_21844,N_19090,N_20698);
xnor U21845 (N_21845,N_18349,N_20730);
nand U21846 (N_21846,N_20520,N_18212);
and U21847 (N_21847,N_18202,N_20454);
xor U21848 (N_21848,N_20516,N_20165);
nor U21849 (N_21849,N_19611,N_20371);
nor U21850 (N_21850,N_20746,N_20058);
nand U21851 (N_21851,N_18385,N_20012);
nand U21852 (N_21852,N_20885,N_20512);
nor U21853 (N_21853,N_18003,N_19438);
nor U21854 (N_21854,N_19342,N_18631);
or U21855 (N_21855,N_19743,N_19969);
xnor U21856 (N_21856,N_19991,N_19153);
nand U21857 (N_21857,N_19555,N_20671);
nand U21858 (N_21858,N_19531,N_18338);
or U21859 (N_21859,N_18317,N_18968);
and U21860 (N_21860,N_20222,N_19645);
xnor U21861 (N_21861,N_19119,N_20586);
xnor U21862 (N_21862,N_20057,N_18571);
or U21863 (N_21863,N_19482,N_19781);
xnor U21864 (N_21864,N_19079,N_20086);
xnor U21865 (N_21865,N_19954,N_20822);
xor U21866 (N_21866,N_18388,N_20295);
or U21867 (N_21867,N_20278,N_20177);
or U21868 (N_21868,N_20868,N_19825);
or U21869 (N_21869,N_19569,N_20090);
or U21870 (N_21870,N_19469,N_20948);
or U21871 (N_21871,N_19897,N_19354);
and U21872 (N_21872,N_20351,N_18941);
nor U21873 (N_21873,N_19363,N_20173);
or U21874 (N_21874,N_18139,N_18923);
or U21875 (N_21875,N_20484,N_20632);
or U21876 (N_21876,N_19065,N_19441);
or U21877 (N_21877,N_18069,N_19029);
nand U21878 (N_21878,N_19656,N_18228);
xor U21879 (N_21879,N_19868,N_18693);
or U21880 (N_21880,N_18991,N_20831);
and U21881 (N_21881,N_18295,N_20928);
nor U21882 (N_21882,N_18701,N_18451);
nand U21883 (N_21883,N_18175,N_19950);
nand U21884 (N_21884,N_19475,N_19248);
nor U21885 (N_21885,N_18436,N_20104);
or U21886 (N_21886,N_20548,N_19854);
and U21887 (N_21887,N_20782,N_19995);
and U21888 (N_21888,N_20684,N_18636);
and U21889 (N_21889,N_19102,N_18130);
nor U21890 (N_21890,N_18567,N_18708);
nand U21891 (N_21891,N_18002,N_20793);
or U21892 (N_21892,N_18414,N_18682);
nand U21893 (N_21893,N_19360,N_20667);
nand U21894 (N_21894,N_19828,N_19779);
nand U21895 (N_21895,N_19416,N_18201);
or U21896 (N_21896,N_18275,N_18795);
nor U21897 (N_21897,N_18203,N_19537);
and U21898 (N_21898,N_19955,N_20623);
xnor U21899 (N_21899,N_20809,N_20789);
and U21900 (N_21900,N_20722,N_18168);
xor U21901 (N_21901,N_20372,N_20218);
nor U21902 (N_21902,N_18565,N_20485);
nand U21903 (N_21903,N_20742,N_19732);
nor U21904 (N_21904,N_18604,N_20980);
nand U21905 (N_21905,N_19758,N_18412);
nor U21906 (N_21906,N_18467,N_19413);
nor U21907 (N_21907,N_18031,N_19529);
and U21908 (N_21908,N_18492,N_18648);
or U21909 (N_21909,N_18819,N_20002);
or U21910 (N_21910,N_19823,N_19742);
and U21911 (N_21911,N_18124,N_18734);
xor U21912 (N_21912,N_20293,N_20797);
and U21913 (N_21913,N_19200,N_18501);
or U21914 (N_21914,N_18300,N_18065);
nor U21915 (N_21915,N_18081,N_18033);
nand U21916 (N_21916,N_19167,N_20735);
xor U21917 (N_21917,N_18315,N_18927);
nor U21918 (N_21918,N_19861,N_20294);
nand U21919 (N_21919,N_18525,N_19388);
and U21920 (N_21920,N_20657,N_18508);
or U21921 (N_21921,N_18077,N_19613);
xnor U21922 (N_21922,N_19953,N_19566);
and U21923 (N_21923,N_20252,N_20648);
nor U21924 (N_21924,N_19101,N_19106);
nor U21925 (N_21925,N_20098,N_19001);
or U21926 (N_21926,N_18703,N_19341);
nand U21927 (N_21927,N_20546,N_18933);
nor U21928 (N_21928,N_18377,N_19590);
and U21929 (N_21929,N_19917,N_18156);
nor U21930 (N_21930,N_19412,N_18671);
and U21931 (N_21931,N_20977,N_19811);
nand U21932 (N_21932,N_18432,N_19789);
nand U21933 (N_21933,N_18347,N_18846);
xor U21934 (N_21934,N_19548,N_19126);
xor U21935 (N_21935,N_19040,N_18120);
nor U21936 (N_21936,N_20589,N_18557);
or U21937 (N_21937,N_18733,N_20127);
or U21938 (N_21938,N_20562,N_20724);
xnor U21939 (N_21939,N_20886,N_20545);
nor U21940 (N_21940,N_18456,N_19587);
and U21941 (N_21941,N_19329,N_18464);
or U21942 (N_21942,N_19169,N_20241);
nor U21943 (N_21943,N_18898,N_20150);
and U21944 (N_21944,N_20946,N_20361);
and U21945 (N_21945,N_20828,N_20088);
and U21946 (N_21946,N_19491,N_20786);
nand U21947 (N_21947,N_19795,N_18355);
xor U21948 (N_21948,N_20467,N_18281);
xor U21949 (N_21949,N_18429,N_18409);
nand U21950 (N_21950,N_20690,N_20587);
or U21951 (N_21951,N_19942,N_18785);
nor U21952 (N_21952,N_20600,N_20233);
or U21953 (N_21953,N_20679,N_18803);
xor U21954 (N_21954,N_20717,N_20544);
nor U21955 (N_21955,N_18711,N_18929);
and U21956 (N_21956,N_18474,N_20669);
or U21957 (N_21957,N_19788,N_18086);
nand U21958 (N_21958,N_19211,N_18310);
nor U21959 (N_21959,N_19801,N_20034);
or U21960 (N_21960,N_18264,N_18322);
or U21961 (N_21961,N_20556,N_18947);
xnor U21962 (N_21962,N_19616,N_19563);
xnor U21963 (N_21963,N_19352,N_20487);
xor U21964 (N_21964,N_18225,N_18485);
nand U21965 (N_21965,N_18885,N_20769);
or U21966 (N_21966,N_19669,N_18902);
nor U21967 (N_21967,N_20085,N_20891);
or U21968 (N_21968,N_19339,N_18662);
and U21969 (N_21969,N_19366,N_19534);
nor U21970 (N_21970,N_19802,N_19635);
and U21971 (N_21971,N_19722,N_19841);
nand U21972 (N_21972,N_18583,N_19948);
and U21973 (N_21973,N_20134,N_20365);
nor U21974 (N_21974,N_18559,N_20658);
xnor U21975 (N_21975,N_18939,N_20456);
or U21976 (N_21976,N_20933,N_19830);
or U21977 (N_21977,N_20197,N_18054);
xor U21978 (N_21978,N_19707,N_20038);
nor U21979 (N_21979,N_18495,N_19839);
nand U21980 (N_21980,N_20040,N_20153);
xor U21981 (N_21981,N_20030,N_19973);
and U21982 (N_21982,N_20705,N_18609);
nor U21983 (N_21983,N_20993,N_20723);
and U21984 (N_21984,N_18142,N_20244);
or U21985 (N_21985,N_19135,N_19023);
and U21986 (N_21986,N_18268,N_20750);
nand U21987 (N_21987,N_18735,N_18121);
xor U21988 (N_21988,N_20333,N_19898);
nor U21989 (N_21989,N_20593,N_20549);
nor U21990 (N_21990,N_20592,N_18327);
xnor U21991 (N_21991,N_18988,N_19988);
or U21992 (N_21992,N_20755,N_19036);
or U21993 (N_21993,N_19127,N_18664);
nor U21994 (N_21994,N_20591,N_19217);
and U21995 (N_21995,N_20524,N_19260);
and U21996 (N_21996,N_19665,N_19188);
xor U21997 (N_21997,N_18522,N_18903);
nor U21998 (N_21998,N_20530,N_19646);
nand U21999 (N_21999,N_18652,N_19210);
xnor U22000 (N_22000,N_18721,N_18136);
nand U22001 (N_22001,N_19085,N_19985);
and U22002 (N_22002,N_19846,N_19326);
nor U22003 (N_22003,N_18028,N_20101);
nand U22004 (N_22004,N_19516,N_20503);
and U22005 (N_22005,N_20693,N_20892);
or U22006 (N_22006,N_20240,N_20234);
xor U22007 (N_22007,N_20700,N_20132);
xnor U22008 (N_22008,N_20348,N_20976);
and U22009 (N_22009,N_19927,N_20383);
or U22010 (N_22010,N_20947,N_18969);
nor U22011 (N_22011,N_19230,N_20025);
or U22012 (N_22012,N_19750,N_20347);
nand U22013 (N_22013,N_19727,N_19423);
nor U22014 (N_22014,N_18438,N_19159);
nor U22015 (N_22015,N_20212,N_18908);
and U22016 (N_22016,N_19904,N_18882);
and U22017 (N_22017,N_20872,N_18059);
nor U22018 (N_22018,N_18847,N_19398);
xnor U22019 (N_22019,N_20739,N_19986);
and U22020 (N_22020,N_19006,N_18126);
xnor U22021 (N_22021,N_19535,N_19888);
nand U22022 (N_22022,N_20912,N_20407);
and U22023 (N_22023,N_19128,N_19549);
nor U22024 (N_22024,N_20056,N_19962);
nor U22025 (N_22025,N_19080,N_18934);
nand U22026 (N_22026,N_19748,N_20834);
and U22027 (N_22027,N_19981,N_18852);
and U22028 (N_22028,N_20953,N_18330);
nor U22029 (N_22029,N_19350,N_19658);
and U22030 (N_22030,N_20776,N_20518);
xnor U22031 (N_22031,N_20622,N_18581);
nor U22032 (N_22032,N_19993,N_18757);
nand U22033 (N_22033,N_19668,N_18806);
xnor U22034 (N_22034,N_20994,N_18427);
xor U22035 (N_22035,N_20916,N_18461);
xor U22036 (N_22036,N_20917,N_19269);
nor U22037 (N_22037,N_18490,N_19878);
xor U22038 (N_22038,N_18463,N_20304);
or U22039 (N_22039,N_18030,N_20465);
or U22040 (N_22040,N_20652,N_20599);
or U22041 (N_22041,N_20905,N_19241);
nor U22042 (N_22042,N_20035,N_19420);
or U22043 (N_22043,N_20115,N_19932);
xor U22044 (N_22044,N_18672,N_20727);
or U22045 (N_22045,N_20463,N_18087);
and U22046 (N_22046,N_19472,N_18262);
xor U22047 (N_22047,N_20113,N_19332);
or U22048 (N_22048,N_18766,N_18115);
xnor U22049 (N_22049,N_19093,N_18146);
nand U22050 (N_22050,N_19179,N_18560);
nand U22051 (N_22051,N_18726,N_19542);
or U22052 (N_22052,N_19757,N_18358);
and U22053 (N_22053,N_20438,N_20580);
or U22054 (N_22054,N_20625,N_19097);
nor U22055 (N_22055,N_18954,N_20534);
or U22056 (N_22056,N_20368,N_18976);
xnor U22057 (N_22057,N_20830,N_19951);
nor U22058 (N_22058,N_18511,N_18230);
xor U22059 (N_22059,N_19145,N_20360);
nand U22060 (N_22060,N_19323,N_18270);
nand U22061 (N_22061,N_20960,N_19010);
xor U22062 (N_22062,N_18339,N_19512);
nor U22063 (N_22063,N_20571,N_20973);
and U22064 (N_22064,N_19136,N_18088);
and U22065 (N_22065,N_18750,N_18537);
and U22066 (N_22066,N_18552,N_19308);
nand U22067 (N_22067,N_20303,N_18831);
or U22068 (N_22068,N_20083,N_20151);
or U22069 (N_22069,N_20125,N_19304);
or U22070 (N_22070,N_20603,N_18058);
xor U22071 (N_22071,N_18316,N_19632);
nor U22072 (N_22072,N_19662,N_20073);
nand U22073 (N_22073,N_19731,N_20488);
and U22074 (N_22074,N_20479,N_19806);
xor U22075 (N_22075,N_19047,N_18359);
xor U22076 (N_22076,N_18044,N_19523);
nand U22077 (N_22077,N_20324,N_18768);
or U22078 (N_22078,N_18304,N_20525);
xor U22079 (N_22079,N_18261,N_20481);
xor U22080 (N_22080,N_19062,N_18122);
xnor U22081 (N_22081,N_18765,N_19197);
xnor U22082 (N_22082,N_19043,N_18626);
nand U22083 (N_22083,N_18745,N_19607);
xor U22084 (N_22084,N_18426,N_20263);
and U22085 (N_22085,N_20352,N_19866);
xor U22086 (N_22086,N_20169,N_19199);
and U22087 (N_22087,N_18266,N_19990);
and U22088 (N_22088,N_18689,N_20331);
nor U22089 (N_22089,N_20264,N_20819);
or U22090 (N_22090,N_19690,N_20913);
xor U22091 (N_22091,N_18274,N_19328);
xor U22092 (N_22092,N_20982,N_18269);
xor U22093 (N_22093,N_18215,N_18794);
or U22094 (N_22094,N_19580,N_19664);
nand U22095 (N_22095,N_18118,N_20862);
or U22096 (N_22096,N_19546,N_19399);
and U22097 (N_22097,N_20985,N_18514);
nor U22098 (N_22098,N_19084,N_18375);
nand U22099 (N_22099,N_18196,N_19301);
nand U22100 (N_22100,N_19903,N_20387);
nand U22101 (N_22101,N_18184,N_19860);
xnor U22102 (N_22102,N_19591,N_19310);
nand U22103 (N_22103,N_19187,N_18380);
nand U22104 (N_22104,N_20160,N_20940);
and U22105 (N_22105,N_20379,N_19856);
nor U22106 (N_22106,N_19192,N_19568);
or U22107 (N_22107,N_18556,N_18724);
nand U22108 (N_22108,N_18290,N_19666);
and U22109 (N_22109,N_20446,N_19486);
and U22110 (N_22110,N_20317,N_18611);
and U22111 (N_22111,N_20388,N_18366);
nor U22112 (N_22112,N_18553,N_18758);
xnor U22113 (N_22113,N_20491,N_18772);
or U22114 (N_22114,N_20644,N_19458);
xnor U22115 (N_22115,N_18946,N_19855);
nand U22116 (N_22116,N_20987,N_20638);
nor U22117 (N_22117,N_20926,N_20328);
and U22118 (N_22118,N_19232,N_19712);
nand U22119 (N_22119,N_18291,N_19552);
or U22120 (N_22120,N_20206,N_18716);
nor U22121 (N_22121,N_18066,N_20595);
nor U22122 (N_22122,N_20675,N_20418);
or U22123 (N_22123,N_18618,N_20140);
and U22124 (N_22124,N_20275,N_19447);
nor U22125 (N_22125,N_20066,N_18881);
xnor U22126 (N_22126,N_18179,N_18207);
nand U22127 (N_22127,N_19798,N_20120);
xor U22128 (N_22128,N_18654,N_20495);
xor U22129 (N_22129,N_18418,N_19524);
nand U22130 (N_22130,N_20447,N_19738);
nor U22131 (N_22131,N_19558,N_19809);
xor U22132 (N_22132,N_19745,N_19028);
nand U22133 (N_22133,N_18332,N_20023);
xnor U22134 (N_22134,N_18805,N_20570);
nor U22135 (N_22135,N_19766,N_18579);
nor U22136 (N_22136,N_19970,N_19946);
nand U22137 (N_22137,N_19686,N_20062);
xor U22138 (N_22138,N_19289,N_18442);
nand U22139 (N_22139,N_20879,N_20596);
or U22140 (N_22140,N_19477,N_20639);
or U22141 (N_22141,N_18205,N_19673);
nand U22142 (N_22142,N_18435,N_20770);
xor U22143 (N_22143,N_20094,N_18154);
or U22144 (N_22144,N_18178,N_18747);
or U22145 (N_22145,N_19464,N_19847);
or U22146 (N_22146,N_19172,N_19391);
xor U22147 (N_22147,N_18769,N_19315);
nor U22148 (N_22148,N_20706,N_19397);
and U22149 (N_22149,N_20691,N_18211);
nor U22150 (N_22150,N_19573,N_18516);
nand U22151 (N_22151,N_18767,N_20326);
or U22152 (N_22152,N_18544,N_19560);
nand U22153 (N_22153,N_18699,N_19373);
or U22154 (N_22154,N_18614,N_19313);
nand U22155 (N_22155,N_19364,N_18974);
and U22156 (N_22156,N_20186,N_19451);
nand U22157 (N_22157,N_19892,N_20631);
nor U22158 (N_22158,N_18739,N_19831);
and U22159 (N_22159,N_18221,N_19804);
and U22160 (N_22160,N_20257,N_20112);
nor U22161 (N_22161,N_19952,N_19292);
nand U22162 (N_22162,N_18271,N_18459);
xnor U22163 (N_22163,N_20003,N_20211);
nor U22164 (N_22164,N_18692,N_20072);
or U22165 (N_22165,N_19863,N_20954);
and U22166 (N_22166,N_20902,N_18188);
nand U22167 (N_22167,N_20937,N_18887);
and U22168 (N_22168,N_18276,N_19378);
xor U22169 (N_22169,N_18020,N_18064);
nand U22170 (N_22170,N_20923,N_19626);
and U22171 (N_22171,N_19835,N_19937);
xor U22172 (N_22172,N_18157,N_20401);
xor U22173 (N_22173,N_18428,N_18875);
nand U22174 (N_22174,N_20535,N_19688);
or U22175 (N_22175,N_20411,N_19076);
nor U22176 (N_22176,N_20840,N_19791);
xnor U22177 (N_22177,N_19180,N_18851);
xor U22178 (N_22178,N_20779,N_18773);
nand U22179 (N_22179,N_18113,N_18985);
and U22180 (N_22180,N_18675,N_19005);
or U22181 (N_22181,N_20773,N_19717);
xor U22182 (N_22182,N_18217,N_18940);
and U22183 (N_22183,N_19679,N_20957);
and U22184 (N_22184,N_19291,N_19146);
nand U22185 (N_22185,N_18964,N_19507);
or U22186 (N_22186,N_19201,N_18779);
or U22187 (N_22187,N_19027,N_20532);
xnor U22188 (N_22188,N_20176,N_19268);
xnor U22189 (N_22189,N_19501,N_20753);
xnor U22190 (N_22190,N_19883,N_18199);
or U22191 (N_22191,N_18231,N_19905);
xor U22192 (N_22192,N_19455,N_20103);
nand U22193 (N_22193,N_19797,N_20897);
nor U22194 (N_22194,N_18599,N_19078);
xor U22195 (N_22195,N_19409,N_19218);
or U22196 (N_22196,N_18821,N_20978);
or U22197 (N_22197,N_19739,N_19371);
and U22198 (N_22198,N_19042,N_19615);
nand U22199 (N_22199,N_18731,N_20394);
nand U22200 (N_22200,N_19776,N_18312);
or U22201 (N_22201,N_20466,N_18836);
nor U22202 (N_22202,N_19726,N_19104);
or U22203 (N_22203,N_18586,N_19650);
or U22204 (N_22204,N_19266,N_20001);
nor U22205 (N_22205,N_20334,N_19912);
nand U22206 (N_22206,N_20575,N_19572);
and U22207 (N_22207,N_19170,N_18570);
nor U22208 (N_22208,N_20670,N_20743);
and U22209 (N_22209,N_20634,N_19980);
nand U22210 (N_22210,N_18433,N_19395);
and U22211 (N_22211,N_18344,N_20262);
xnor U22212 (N_22212,N_18285,N_20641);
or U22213 (N_22213,N_20521,N_19602);
xnor U22214 (N_22214,N_19109,N_18612);
nor U22215 (N_22215,N_19317,N_20609);
nor U22216 (N_22216,N_20432,N_19960);
nand U22217 (N_22217,N_20729,N_19771);
xor U22218 (N_22218,N_20874,N_20200);
nor U22219 (N_22219,N_19598,N_20037);
or U22220 (N_22220,N_18011,N_18234);
nor U22221 (N_22221,N_18499,N_19270);
or U22222 (N_22222,N_18062,N_18220);
nand U22223 (N_22223,N_19009,N_20865);
or U22224 (N_22224,N_19837,N_20790);
nor U22225 (N_22225,N_20193,N_20918);
nor U22226 (N_22226,N_19114,N_18680);
and U22227 (N_22227,N_19442,N_19258);
nand U22228 (N_22228,N_19676,N_18109);
xor U22229 (N_22229,N_18301,N_18910);
and U22230 (N_22230,N_20406,N_18542);
xor U22231 (N_22231,N_19649,N_19393);
nor U22232 (N_22232,N_20095,N_20170);
or U22233 (N_22233,N_19687,N_20227);
xnor U22234 (N_22234,N_18477,N_19008);
nand U22235 (N_22235,N_20896,N_20167);
or U22236 (N_22236,N_18185,N_19941);
nand U22237 (N_22237,N_19997,N_19439);
nor U22238 (N_22238,N_18883,N_20910);
xor U22239 (N_22239,N_19018,N_18704);
and U22240 (N_22240,N_18749,N_20943);
or U22241 (N_22241,N_18897,N_18078);
nor U22242 (N_22242,N_18644,N_20332);
or U22243 (N_22243,N_20162,N_19394);
nand U22244 (N_22244,N_19069,N_19584);
nand U22245 (N_22245,N_20814,N_20219);
nand U22246 (N_22246,N_20798,N_18381);
and U22247 (N_22247,N_20052,N_18303);
and U22248 (N_22248,N_19979,N_18141);
nand U22249 (N_22249,N_20039,N_18809);
nand U22250 (N_22250,N_18187,N_19231);
nand U22251 (N_22251,N_18959,N_20415);
nor U22252 (N_22252,N_18781,N_18931);
or U22253 (N_22253,N_19984,N_20701);
or U22254 (N_22254,N_20174,N_19138);
nor U22255 (N_22255,N_20385,N_20816);
or U22256 (N_22256,N_18336,N_18637);
and U22257 (N_22257,N_19133,N_20067);
or U22258 (N_22258,N_20026,N_18791);
nor U22259 (N_22259,N_19238,N_20398);
nand U22260 (N_22260,N_19881,N_20969);
nor U22261 (N_22261,N_19287,N_19083);
nor U22262 (N_22262,N_20666,N_18880);
nor U22263 (N_22263,N_18289,N_20018);
nor U22264 (N_22264,N_18656,N_19183);
or U22265 (N_22265,N_20453,N_19427);
and U22266 (N_22266,N_18907,N_19551);
nor U22267 (N_22267,N_20839,N_20462);
nor U22268 (N_22268,N_18329,N_19522);
xor U22269 (N_22269,N_20396,N_19014);
or U22270 (N_22270,N_19747,N_20651);
nor U22271 (N_22271,N_20107,N_20309);
or U22272 (N_22272,N_18263,N_19240);
or U22273 (N_22273,N_20871,N_18099);
xor U22274 (N_22274,N_19703,N_19938);
xor U22275 (N_22275,N_18673,N_18284);
nand U22276 (N_22276,N_19004,N_19448);
or U22277 (N_22277,N_18925,N_19035);
xnor U22278 (N_22278,N_20997,N_18655);
and U22279 (N_22279,N_18688,N_19729);
nor U22280 (N_22280,N_18890,N_19387);
nor U22281 (N_22281,N_20187,N_19589);
xnor U22282 (N_22282,N_20249,N_20906);
nand U22283 (N_22283,N_20606,N_18639);
xor U22284 (N_22284,N_18633,N_20821);
and U22285 (N_22285,N_19073,N_18524);
or U22286 (N_22286,N_19765,N_19400);
xnor U22287 (N_22287,N_18787,N_18770);
or U22288 (N_22288,N_19020,N_19321);
or U22289 (N_22289,N_20185,N_20049);
or U22290 (N_22290,N_19481,N_19347);
xnor U22291 (N_22291,N_19924,N_19330);
nor U22292 (N_22292,N_19816,N_19896);
and U22293 (N_22293,N_20060,N_19297);
and U22294 (N_22294,N_20239,N_18800);
and U22295 (N_22295,N_20410,N_20857);
nor U22296 (N_22296,N_19349,N_19642);
or U22297 (N_22297,N_19032,N_18534);
nand U22298 (N_22298,N_20761,N_20209);
and U22299 (N_22299,N_19225,N_18651);
and U22300 (N_22300,N_19763,N_20378);
and U22301 (N_22301,N_20713,N_18422);
nand U22302 (N_22302,N_18515,N_20382);
and U22303 (N_22303,N_20859,N_20642);
xnor U22304 (N_22304,N_20972,N_20449);
nor U22305 (N_22305,N_18197,N_19021);
nand U22306 (N_22306,N_18027,N_19071);
or U22307 (N_22307,N_18399,N_20597);
or U22308 (N_22308,N_18572,N_19255);
nand U22309 (N_22309,N_20163,N_20157);
xor U22310 (N_22310,N_18251,N_19829);
nand U22311 (N_22311,N_18340,N_20583);
and U22312 (N_22312,N_19299,N_20425);
nor U22313 (N_22313,N_19437,N_18888);
and U22314 (N_22314,N_18862,N_20791);
nor U22315 (N_22315,N_18683,N_18798);
xnor U22316 (N_22316,N_19406,N_18280);
and U22317 (N_22317,N_18273,N_20096);
or U22318 (N_22318,N_19333,N_19415);
xor U22319 (N_22319,N_18759,N_18256);
xnor U22320 (N_22320,N_18468,N_20136);
or U22321 (N_22321,N_20265,N_18083);
and U22322 (N_22322,N_20778,N_18391);
or U22323 (N_22323,N_19039,N_18569);
nor U22324 (N_22324,N_18756,N_20483);
xnor U22325 (N_22325,N_19641,N_18577);
nor U22326 (N_22326,N_19495,N_19784);
xor U22327 (N_22327,N_18601,N_20505);
xor U22328 (N_22328,N_20172,N_19452);
xnor U22329 (N_22329,N_19089,N_19494);
nor U22330 (N_22330,N_19503,N_18778);
nor U22331 (N_22331,N_20416,N_18597);
or U22332 (N_22332,N_19660,N_18018);
and U22333 (N_22333,N_18023,N_19407);
and U22334 (N_22334,N_20647,N_19578);
nor U22335 (N_22335,N_18458,N_19862);
nor U22336 (N_22336,N_20391,N_18518);
and U22337 (N_22337,N_20381,N_19698);
or U22338 (N_22338,N_18392,N_20080);
nand U22339 (N_22339,N_18856,N_18177);
nand U22340 (N_22340,N_19498,N_18493);
nor U22341 (N_22341,N_18161,N_20922);
and U22342 (N_22342,N_19139,N_20459);
nor U22343 (N_22343,N_19876,N_19390);
nand U22344 (N_22344,N_20235,N_18417);
nor U22345 (N_22345,N_20117,N_19462);
and U22346 (N_22346,N_19264,N_19033);
and U22347 (N_22347,N_19239,N_20762);
xor U22348 (N_22348,N_20045,N_19055);
nor U22349 (N_22349,N_18970,N_19278);
nand U22350 (N_22350,N_19623,N_18278);
or U22351 (N_22351,N_19840,N_20818);
nor U22352 (N_22352,N_19999,N_18012);
nand U22353 (N_22353,N_20444,N_20434);
nor U22354 (N_22354,N_19143,N_20526);
and U22355 (N_22355,N_18097,N_19405);
or U22356 (N_22356,N_20676,N_20767);
nor U22357 (N_22357,N_20089,N_19041);
or U22358 (N_22358,N_20299,N_20259);
nand U22359 (N_22359,N_18400,N_19851);
nor U22360 (N_22360,N_19728,N_19259);
and U22361 (N_22361,N_18722,N_20835);
and U22362 (N_22362,N_20699,N_19701);
xnor U22363 (N_22363,N_19056,N_19053);
xnor U22364 (N_22364,N_19931,N_18035);
and U22365 (N_22365,N_19096,N_20936);
and U22366 (N_22366,N_19226,N_19853);
or U22367 (N_22367,N_19490,N_19786);
xor U22368 (N_22368,N_20353,N_20687);
nor U22369 (N_22369,N_18590,N_19132);
and U22370 (N_22370,N_18343,N_18037);
xnor U22371 (N_22371,N_18695,N_19826);
xnor U22372 (N_22372,N_19216,N_20345);
or U22373 (N_22373,N_19064,N_19792);
xor U22374 (N_22374,N_20624,N_20775);
nor U22375 (N_22375,N_20393,N_18223);
and U22376 (N_22376,N_19034,N_19483);
xor U22377 (N_22377,N_19382,N_18646);
nand U22378 (N_22378,N_19817,N_18476);
xnor U22379 (N_22379,N_18131,N_20182);
xor U22380 (N_22380,N_19880,N_20129);
xnor U22381 (N_22381,N_18543,N_19640);
and U22382 (N_22382,N_20628,N_18465);
nor U22383 (N_22383,N_18563,N_18100);
or U22384 (N_22384,N_20131,N_20618);
nand U22385 (N_22385,N_20950,N_20719);
and U22386 (N_22386,N_19166,N_18729);
and U22387 (N_22387,N_18253,N_19303);
nor U22388 (N_22388,N_20384,N_19088);
or U22389 (N_22389,N_18061,N_20220);
xnor U22390 (N_22390,N_18615,N_18705);
or U22391 (N_22391,N_19137,N_19229);
nand U22392 (N_22392,N_19539,N_20598);
nor U22393 (N_22393,N_20800,N_20156);
and U22394 (N_22394,N_19182,N_20590);
and U22395 (N_22395,N_20439,N_20280);
and U22396 (N_22396,N_19209,N_18955);
and U22397 (N_22397,N_18919,N_18478);
nand U22398 (N_22398,N_20277,N_20981);
nand U22399 (N_22399,N_20196,N_19453);
xnor U22400 (N_22400,N_19099,N_19681);
xnor U22401 (N_22401,N_18308,N_18236);
nand U22402 (N_22402,N_18521,N_18737);
and U22403 (N_22403,N_20075,N_20268);
or U22404 (N_22404,N_18036,N_18089);
nand U22405 (N_22405,N_20807,N_19827);
xor U22406 (N_22406,N_20028,N_20945);
nand U22407 (N_22407,N_18665,N_19147);
or U22408 (N_22408,N_20435,N_19842);
nor U22409 (N_22409,N_18098,N_18978);
or U22410 (N_22410,N_19125,N_19284);
or U22411 (N_22411,N_20630,N_19443);
and U22412 (N_22412,N_19177,N_18048);
xor U22413 (N_22413,N_18206,N_18629);
nand U22414 (N_22414,N_20914,N_19396);
and U22415 (N_22415,N_18870,N_19588);
or U22416 (N_22416,N_20942,N_18783);
nand U22417 (N_22417,N_20783,N_19796);
nor U22418 (N_22418,N_20207,N_20496);
and U22419 (N_22419,N_19421,N_18899);
xnor U22420 (N_22420,N_18371,N_20636);
xnor U22421 (N_22421,N_20477,N_20501);
xor U22422 (N_22422,N_19696,N_19699);
or U22423 (N_22423,N_18920,N_20074);
and U22424 (N_22424,N_18690,N_19700);
or U22425 (N_22425,N_20697,N_19894);
nor U22426 (N_22426,N_18406,N_19214);
xor U22427 (N_22427,N_18296,N_19843);
nor U22428 (N_22428,N_20180,N_19968);
and U22429 (N_22429,N_18379,N_19852);
xor U22430 (N_22430,N_20287,N_19149);
and U22431 (N_22431,N_18960,N_18001);
and U22432 (N_22432,N_19072,N_20420);
xnor U22433 (N_22433,N_18243,N_19561);
nor U22434 (N_22434,N_18879,N_18751);
nor U22435 (N_22435,N_18732,N_18402);
xor U22436 (N_22436,N_18742,N_20139);
nand U22437 (N_22437,N_19022,N_18248);
or U22438 (N_22438,N_18390,N_20745);
nor U22439 (N_22439,N_18443,N_20482);
xor U22440 (N_22440,N_19422,N_18496);
nand U22441 (N_22441,N_19821,N_19716);
xor U22442 (N_22442,N_20430,N_18588);
xnor U22443 (N_22443,N_19720,N_18628);
xnor U22444 (N_22444,N_19859,N_18613);
and U22445 (N_22445,N_19583,N_20996);
nor U22446 (N_22446,N_19737,N_18598);
xnor U22447 (N_22447,N_18324,N_20737);
nor U22448 (N_22448,N_18352,N_19526);
nand U22449 (N_22449,N_20213,N_19191);
nand U22450 (N_22450,N_19433,N_20784);
nand U22451 (N_22451,N_20009,N_19663);
xnor U22452 (N_22452,N_18728,N_18591);
xnor U22453 (N_22453,N_18776,N_20506);
or U22454 (N_22454,N_18853,N_19773);
nand U22455 (N_22455,N_19683,N_18229);
or U22456 (N_22456,N_20513,N_20144);
xnor U22457 (N_22457,N_20824,N_20250);
and U22458 (N_22458,N_19431,N_18333);
xor U22459 (N_22459,N_20527,N_19305);
nand U22460 (N_22460,N_19556,N_18844);
nand U22461 (N_22461,N_19600,N_20812);
nor U22462 (N_22462,N_19282,N_18912);
or U22463 (N_22463,N_20051,N_19444);
or U22464 (N_22464,N_20794,N_20531);
xor U22465 (N_22465,N_18469,N_18213);
and U22466 (N_22466,N_19379,N_18533);
and U22467 (N_22467,N_20158,N_18548);
or U22468 (N_22468,N_20650,N_18527);
or U22469 (N_22469,N_18032,N_19202);
nor U22470 (N_22470,N_18026,N_19118);
nor U22471 (N_22471,N_20102,N_18475);
xor U22472 (N_22472,N_20633,N_20242);
and U22473 (N_22473,N_18822,N_20732);
and U22474 (N_22474,N_19775,N_20877);
or U22475 (N_22475,N_20898,N_20492);
nor U22476 (N_22476,N_18884,N_19815);
and U22477 (N_22477,N_19755,N_20109);
xnor U22478 (N_22478,N_20949,N_19751);
or U22479 (N_22479,N_18410,N_20301);
or U22480 (N_22480,N_19369,N_19564);
nor U22481 (N_22481,N_20961,N_18453);
and U22482 (N_22482,N_19652,N_18398);
xor U22483 (N_22483,N_18917,N_18420);
or U22484 (N_22484,N_19419,N_20164);
nor U22485 (N_22485,N_19254,N_19978);
nor U22486 (N_22486,N_19295,N_18755);
xnor U22487 (N_22487,N_18288,N_20601);
xor U22488 (N_22488,N_19302,N_19693);
nand U22489 (N_22489,N_19943,N_18132);
nand U22490 (N_22490,N_18720,N_19527);
or U22491 (N_22491,N_20504,N_18222);
or U22492 (N_22492,N_20064,N_19547);
nor U22493 (N_22493,N_19324,N_20608);
or U22494 (N_22494,N_19190,N_20440);
and U22495 (N_22495,N_18357,N_20866);
xnor U22496 (N_22496,N_20340,N_18383);
and U22497 (N_22497,N_19057,N_20146);
nor U22498 (N_22498,N_19338,N_19889);
and U22499 (N_22499,N_20204,N_20175);
nor U22500 (N_22500,N_18379,N_19549);
nor U22501 (N_22501,N_20072,N_18451);
nor U22502 (N_22502,N_20574,N_18966);
nor U22503 (N_22503,N_19841,N_19201);
xor U22504 (N_22504,N_19293,N_19373);
or U22505 (N_22505,N_20253,N_18145);
xor U22506 (N_22506,N_19334,N_18423);
nor U22507 (N_22507,N_19479,N_19884);
xor U22508 (N_22508,N_20504,N_20745);
nor U22509 (N_22509,N_19163,N_18447);
or U22510 (N_22510,N_20690,N_19711);
or U22511 (N_22511,N_20208,N_18713);
or U22512 (N_22512,N_19640,N_19432);
xor U22513 (N_22513,N_19532,N_18508);
nand U22514 (N_22514,N_19923,N_19406);
nor U22515 (N_22515,N_20172,N_20654);
nand U22516 (N_22516,N_18909,N_18543);
nor U22517 (N_22517,N_20428,N_18984);
or U22518 (N_22518,N_20240,N_18488);
nand U22519 (N_22519,N_20113,N_18309);
xor U22520 (N_22520,N_20295,N_20587);
nand U22521 (N_22521,N_20260,N_18378);
nor U22522 (N_22522,N_19113,N_18902);
and U22523 (N_22523,N_19490,N_19979);
nor U22524 (N_22524,N_19958,N_18719);
nand U22525 (N_22525,N_19106,N_18243);
or U22526 (N_22526,N_18951,N_20152);
xor U22527 (N_22527,N_20989,N_20445);
or U22528 (N_22528,N_19698,N_19056);
nand U22529 (N_22529,N_20468,N_18052);
nand U22530 (N_22530,N_20748,N_18222);
or U22531 (N_22531,N_19359,N_19327);
xor U22532 (N_22532,N_19268,N_18387);
nand U22533 (N_22533,N_18270,N_18567);
xor U22534 (N_22534,N_18338,N_18923);
or U22535 (N_22535,N_19839,N_20617);
xor U22536 (N_22536,N_19527,N_19470);
or U22537 (N_22537,N_18962,N_19176);
nor U22538 (N_22538,N_18627,N_18390);
nor U22539 (N_22539,N_19173,N_20529);
and U22540 (N_22540,N_19365,N_19627);
nand U22541 (N_22541,N_20173,N_18031);
nand U22542 (N_22542,N_20526,N_18213);
and U22543 (N_22543,N_19942,N_20895);
nor U22544 (N_22544,N_20296,N_18552);
nor U22545 (N_22545,N_18999,N_19608);
xnor U22546 (N_22546,N_19257,N_20382);
xnor U22547 (N_22547,N_19579,N_19544);
nor U22548 (N_22548,N_19709,N_18373);
xor U22549 (N_22549,N_19267,N_20056);
xor U22550 (N_22550,N_20615,N_18271);
or U22551 (N_22551,N_19090,N_18105);
xnor U22552 (N_22552,N_18267,N_19582);
nor U22553 (N_22553,N_18803,N_19583);
or U22554 (N_22554,N_19128,N_18674);
nand U22555 (N_22555,N_18436,N_20196);
nor U22556 (N_22556,N_19062,N_18501);
nand U22557 (N_22557,N_19829,N_19100);
nor U22558 (N_22558,N_20635,N_19348);
nor U22559 (N_22559,N_18958,N_20001);
or U22560 (N_22560,N_18632,N_20213);
nor U22561 (N_22561,N_18708,N_20527);
nor U22562 (N_22562,N_20968,N_19668);
or U22563 (N_22563,N_19473,N_18177);
and U22564 (N_22564,N_19284,N_19605);
xor U22565 (N_22565,N_20932,N_18818);
nand U22566 (N_22566,N_18362,N_20959);
nor U22567 (N_22567,N_20755,N_19707);
nand U22568 (N_22568,N_20026,N_20916);
and U22569 (N_22569,N_18827,N_20468);
or U22570 (N_22570,N_18986,N_18818);
nand U22571 (N_22571,N_19920,N_19832);
and U22572 (N_22572,N_18806,N_18319);
nor U22573 (N_22573,N_20206,N_19524);
xor U22574 (N_22574,N_18678,N_18770);
nand U22575 (N_22575,N_20359,N_18466);
xor U22576 (N_22576,N_20887,N_20690);
nor U22577 (N_22577,N_18284,N_20871);
and U22578 (N_22578,N_20715,N_19331);
nand U22579 (N_22579,N_20239,N_19735);
nand U22580 (N_22580,N_18438,N_20006);
or U22581 (N_22581,N_19576,N_20106);
and U22582 (N_22582,N_19548,N_20159);
nor U22583 (N_22583,N_20020,N_18894);
xor U22584 (N_22584,N_18528,N_19539);
or U22585 (N_22585,N_19268,N_18110);
nor U22586 (N_22586,N_18269,N_20148);
and U22587 (N_22587,N_19624,N_18962);
nor U22588 (N_22588,N_20504,N_18665);
or U22589 (N_22589,N_20431,N_20428);
nand U22590 (N_22590,N_20787,N_20276);
xnor U22591 (N_22591,N_19321,N_19161);
xor U22592 (N_22592,N_18038,N_20678);
or U22593 (N_22593,N_20456,N_18910);
and U22594 (N_22594,N_20820,N_18130);
or U22595 (N_22595,N_19648,N_18807);
and U22596 (N_22596,N_20287,N_20892);
nand U22597 (N_22597,N_20376,N_19224);
or U22598 (N_22598,N_18209,N_20815);
and U22599 (N_22599,N_19537,N_20214);
nor U22600 (N_22600,N_18143,N_19682);
nand U22601 (N_22601,N_18823,N_19463);
xor U22602 (N_22602,N_19460,N_19378);
nand U22603 (N_22603,N_19135,N_19899);
and U22604 (N_22604,N_19802,N_18846);
xnor U22605 (N_22605,N_18045,N_18663);
or U22606 (N_22606,N_18611,N_18314);
and U22607 (N_22607,N_20362,N_20224);
xor U22608 (N_22608,N_19531,N_19462);
and U22609 (N_22609,N_20739,N_19901);
or U22610 (N_22610,N_18085,N_20699);
xnor U22611 (N_22611,N_18428,N_20078);
or U22612 (N_22612,N_18655,N_20184);
nand U22613 (N_22613,N_19322,N_18508);
or U22614 (N_22614,N_19510,N_18281);
nor U22615 (N_22615,N_20076,N_20916);
and U22616 (N_22616,N_18935,N_20050);
nor U22617 (N_22617,N_19245,N_18220);
and U22618 (N_22618,N_19165,N_18006);
nand U22619 (N_22619,N_19791,N_20950);
or U22620 (N_22620,N_20999,N_19678);
xor U22621 (N_22621,N_20290,N_18732);
nand U22622 (N_22622,N_20116,N_19711);
nor U22623 (N_22623,N_18345,N_18622);
or U22624 (N_22624,N_19886,N_19878);
xor U22625 (N_22625,N_20233,N_19182);
nor U22626 (N_22626,N_19664,N_18421);
or U22627 (N_22627,N_18104,N_18106);
or U22628 (N_22628,N_18546,N_20486);
and U22629 (N_22629,N_20044,N_20735);
xnor U22630 (N_22630,N_18324,N_19132);
xnor U22631 (N_22631,N_18921,N_19746);
nor U22632 (N_22632,N_18787,N_19900);
xnor U22633 (N_22633,N_19148,N_19966);
xor U22634 (N_22634,N_18012,N_18538);
xor U22635 (N_22635,N_18839,N_20194);
and U22636 (N_22636,N_19179,N_20482);
nand U22637 (N_22637,N_20988,N_20432);
nor U22638 (N_22638,N_18295,N_20868);
nor U22639 (N_22639,N_18233,N_19845);
xor U22640 (N_22640,N_18473,N_18831);
nand U22641 (N_22641,N_20823,N_19677);
and U22642 (N_22642,N_19684,N_18220);
xor U22643 (N_22643,N_20527,N_20156);
or U22644 (N_22644,N_20636,N_20791);
nand U22645 (N_22645,N_20705,N_18367);
and U22646 (N_22646,N_18699,N_18737);
xor U22647 (N_22647,N_19769,N_19370);
and U22648 (N_22648,N_20908,N_18992);
nor U22649 (N_22649,N_20989,N_20439);
or U22650 (N_22650,N_20799,N_18394);
and U22651 (N_22651,N_18121,N_20605);
nor U22652 (N_22652,N_19916,N_20478);
or U22653 (N_22653,N_20368,N_20598);
nand U22654 (N_22654,N_18408,N_19761);
xor U22655 (N_22655,N_18819,N_19234);
or U22656 (N_22656,N_18108,N_19872);
xor U22657 (N_22657,N_20737,N_19701);
nor U22658 (N_22658,N_20045,N_20407);
nor U22659 (N_22659,N_19067,N_20584);
nand U22660 (N_22660,N_20155,N_19305);
nand U22661 (N_22661,N_19022,N_18867);
nand U22662 (N_22662,N_20637,N_19999);
nand U22663 (N_22663,N_20324,N_18571);
and U22664 (N_22664,N_18174,N_18673);
and U22665 (N_22665,N_20749,N_18484);
nand U22666 (N_22666,N_19048,N_19778);
or U22667 (N_22667,N_19068,N_20911);
or U22668 (N_22668,N_20298,N_18355);
or U22669 (N_22669,N_20920,N_18108);
or U22670 (N_22670,N_19548,N_20284);
nor U22671 (N_22671,N_19699,N_20429);
or U22672 (N_22672,N_20278,N_20919);
xnor U22673 (N_22673,N_19397,N_18007);
and U22674 (N_22674,N_19833,N_20942);
and U22675 (N_22675,N_19050,N_18092);
nor U22676 (N_22676,N_18283,N_18089);
or U22677 (N_22677,N_18518,N_19418);
nor U22678 (N_22678,N_18825,N_19886);
xnor U22679 (N_22679,N_18819,N_18965);
xnor U22680 (N_22680,N_20480,N_19117);
xnor U22681 (N_22681,N_19073,N_18851);
xor U22682 (N_22682,N_19390,N_18139);
nor U22683 (N_22683,N_18007,N_19991);
nand U22684 (N_22684,N_20103,N_18142);
nor U22685 (N_22685,N_19492,N_18142);
nor U22686 (N_22686,N_19697,N_20504);
nand U22687 (N_22687,N_18385,N_19147);
nand U22688 (N_22688,N_18955,N_20289);
and U22689 (N_22689,N_18866,N_18551);
and U22690 (N_22690,N_18205,N_19337);
xor U22691 (N_22691,N_18209,N_20612);
or U22692 (N_22692,N_19331,N_19601);
nor U22693 (N_22693,N_20180,N_18861);
or U22694 (N_22694,N_20413,N_20955);
nor U22695 (N_22695,N_19619,N_20056);
and U22696 (N_22696,N_18554,N_19430);
and U22697 (N_22697,N_20680,N_20060);
xnor U22698 (N_22698,N_18288,N_20118);
nand U22699 (N_22699,N_19016,N_20812);
and U22700 (N_22700,N_18003,N_18171);
nand U22701 (N_22701,N_20577,N_20251);
and U22702 (N_22702,N_18572,N_19120);
nand U22703 (N_22703,N_19035,N_20841);
or U22704 (N_22704,N_19569,N_19214);
nand U22705 (N_22705,N_19260,N_19252);
xnor U22706 (N_22706,N_18293,N_20475);
nand U22707 (N_22707,N_20478,N_19582);
and U22708 (N_22708,N_19905,N_20965);
and U22709 (N_22709,N_20810,N_18472);
xnor U22710 (N_22710,N_20159,N_19612);
or U22711 (N_22711,N_18451,N_19557);
nand U22712 (N_22712,N_18503,N_20424);
or U22713 (N_22713,N_19337,N_20345);
or U22714 (N_22714,N_19396,N_20868);
nor U22715 (N_22715,N_19290,N_20759);
xnor U22716 (N_22716,N_18522,N_18266);
nand U22717 (N_22717,N_19638,N_19079);
nor U22718 (N_22718,N_19677,N_20995);
xnor U22719 (N_22719,N_20671,N_20412);
xnor U22720 (N_22720,N_18976,N_20822);
nand U22721 (N_22721,N_18620,N_18714);
or U22722 (N_22722,N_18115,N_18253);
nor U22723 (N_22723,N_19829,N_18179);
nor U22724 (N_22724,N_20642,N_19409);
nor U22725 (N_22725,N_18661,N_20071);
xnor U22726 (N_22726,N_19096,N_18000);
nor U22727 (N_22727,N_20270,N_18245);
nor U22728 (N_22728,N_20687,N_18865);
and U22729 (N_22729,N_20675,N_18308);
and U22730 (N_22730,N_20829,N_19893);
nand U22731 (N_22731,N_18223,N_19790);
nand U22732 (N_22732,N_18921,N_19856);
or U22733 (N_22733,N_19256,N_19199);
xnor U22734 (N_22734,N_20391,N_19453);
nand U22735 (N_22735,N_20451,N_18680);
and U22736 (N_22736,N_19446,N_20557);
and U22737 (N_22737,N_20081,N_20990);
xor U22738 (N_22738,N_19746,N_18989);
xnor U22739 (N_22739,N_19414,N_20002);
or U22740 (N_22740,N_19629,N_18820);
xor U22741 (N_22741,N_20907,N_18002);
or U22742 (N_22742,N_20700,N_18877);
nand U22743 (N_22743,N_18239,N_19656);
nor U22744 (N_22744,N_20029,N_18894);
xnor U22745 (N_22745,N_20701,N_18822);
nand U22746 (N_22746,N_18629,N_19676);
and U22747 (N_22747,N_20337,N_19218);
and U22748 (N_22748,N_18557,N_19098);
or U22749 (N_22749,N_18216,N_20093);
xnor U22750 (N_22750,N_18517,N_20515);
and U22751 (N_22751,N_19297,N_19994);
nor U22752 (N_22752,N_18226,N_18307);
xnor U22753 (N_22753,N_19316,N_20974);
or U22754 (N_22754,N_18220,N_20860);
xor U22755 (N_22755,N_18069,N_18068);
xnor U22756 (N_22756,N_19934,N_20735);
nand U22757 (N_22757,N_20103,N_19135);
and U22758 (N_22758,N_20266,N_18085);
and U22759 (N_22759,N_20573,N_18640);
xnor U22760 (N_22760,N_19223,N_20509);
xnor U22761 (N_22761,N_19491,N_20328);
nand U22762 (N_22762,N_18937,N_20057);
nand U22763 (N_22763,N_20017,N_19548);
nand U22764 (N_22764,N_18507,N_19394);
or U22765 (N_22765,N_20013,N_19964);
and U22766 (N_22766,N_18634,N_20947);
xnor U22767 (N_22767,N_18311,N_19195);
and U22768 (N_22768,N_20631,N_20522);
xor U22769 (N_22769,N_18766,N_19678);
and U22770 (N_22770,N_19135,N_19686);
or U22771 (N_22771,N_18228,N_18621);
and U22772 (N_22772,N_19371,N_18263);
and U22773 (N_22773,N_19627,N_19775);
nand U22774 (N_22774,N_18500,N_18690);
xnor U22775 (N_22775,N_18326,N_18974);
nand U22776 (N_22776,N_20530,N_18341);
nor U22777 (N_22777,N_18979,N_18191);
nand U22778 (N_22778,N_19461,N_19538);
or U22779 (N_22779,N_18444,N_18691);
or U22780 (N_22780,N_19963,N_18847);
or U22781 (N_22781,N_19112,N_20030);
or U22782 (N_22782,N_19951,N_20384);
xnor U22783 (N_22783,N_20777,N_19719);
or U22784 (N_22784,N_20493,N_18000);
or U22785 (N_22785,N_18863,N_19503);
nand U22786 (N_22786,N_19787,N_18909);
and U22787 (N_22787,N_20144,N_20721);
nand U22788 (N_22788,N_18525,N_18712);
or U22789 (N_22789,N_18686,N_18696);
or U22790 (N_22790,N_19804,N_19414);
xor U22791 (N_22791,N_18223,N_18800);
xor U22792 (N_22792,N_20793,N_20011);
xor U22793 (N_22793,N_19253,N_20626);
nor U22794 (N_22794,N_19263,N_18110);
and U22795 (N_22795,N_20846,N_19033);
and U22796 (N_22796,N_19282,N_19951);
or U22797 (N_22797,N_19643,N_18355);
nor U22798 (N_22798,N_19769,N_19952);
nand U22799 (N_22799,N_20903,N_19056);
and U22800 (N_22800,N_19416,N_19507);
nand U22801 (N_22801,N_18016,N_20933);
nand U22802 (N_22802,N_19765,N_18053);
or U22803 (N_22803,N_20869,N_20193);
nand U22804 (N_22804,N_18309,N_20804);
xor U22805 (N_22805,N_20369,N_19973);
xnor U22806 (N_22806,N_18119,N_20339);
and U22807 (N_22807,N_20110,N_18877);
or U22808 (N_22808,N_18981,N_19420);
nand U22809 (N_22809,N_18815,N_20344);
nor U22810 (N_22810,N_19957,N_18686);
xnor U22811 (N_22811,N_20937,N_18711);
xnor U22812 (N_22812,N_19255,N_20578);
nand U22813 (N_22813,N_19524,N_19658);
and U22814 (N_22814,N_20037,N_20067);
nand U22815 (N_22815,N_18004,N_20626);
xor U22816 (N_22816,N_20728,N_18121);
xor U22817 (N_22817,N_18773,N_19864);
nand U22818 (N_22818,N_18275,N_19897);
nor U22819 (N_22819,N_18561,N_18653);
nor U22820 (N_22820,N_19617,N_19301);
xor U22821 (N_22821,N_18266,N_20927);
or U22822 (N_22822,N_19456,N_18721);
nand U22823 (N_22823,N_18500,N_18806);
xor U22824 (N_22824,N_18665,N_19281);
xor U22825 (N_22825,N_19212,N_19326);
and U22826 (N_22826,N_20431,N_18904);
or U22827 (N_22827,N_20284,N_19871);
nand U22828 (N_22828,N_20265,N_19773);
and U22829 (N_22829,N_19723,N_18081);
and U22830 (N_22830,N_19268,N_18707);
xnor U22831 (N_22831,N_19537,N_20584);
xor U22832 (N_22832,N_18554,N_18051);
nor U22833 (N_22833,N_20544,N_19933);
and U22834 (N_22834,N_18704,N_19755);
nand U22835 (N_22835,N_19680,N_19970);
nor U22836 (N_22836,N_18463,N_20549);
xor U22837 (N_22837,N_19384,N_19004);
and U22838 (N_22838,N_18400,N_18403);
nand U22839 (N_22839,N_20827,N_19690);
and U22840 (N_22840,N_18054,N_19948);
nor U22841 (N_22841,N_18759,N_18509);
nor U22842 (N_22842,N_19216,N_19151);
xnor U22843 (N_22843,N_18135,N_19528);
or U22844 (N_22844,N_19514,N_18996);
nor U22845 (N_22845,N_19615,N_18048);
or U22846 (N_22846,N_18479,N_20899);
xnor U22847 (N_22847,N_20536,N_18805);
nor U22848 (N_22848,N_18009,N_18745);
xnor U22849 (N_22849,N_19197,N_18752);
nand U22850 (N_22850,N_20107,N_20819);
and U22851 (N_22851,N_20404,N_20421);
or U22852 (N_22852,N_18450,N_20761);
nor U22853 (N_22853,N_19665,N_20673);
nor U22854 (N_22854,N_20521,N_20798);
and U22855 (N_22855,N_19757,N_20925);
xnor U22856 (N_22856,N_19929,N_18409);
nand U22857 (N_22857,N_19742,N_18104);
nand U22858 (N_22858,N_18764,N_19750);
or U22859 (N_22859,N_20697,N_20039);
nand U22860 (N_22860,N_20728,N_19660);
nand U22861 (N_22861,N_19247,N_18645);
or U22862 (N_22862,N_18639,N_19009);
or U22863 (N_22863,N_20573,N_20610);
xor U22864 (N_22864,N_20494,N_20072);
nor U22865 (N_22865,N_19338,N_19513);
or U22866 (N_22866,N_19968,N_18846);
nand U22867 (N_22867,N_20092,N_20051);
nor U22868 (N_22868,N_20776,N_20980);
nor U22869 (N_22869,N_19247,N_18232);
nor U22870 (N_22870,N_19406,N_18612);
nand U22871 (N_22871,N_20750,N_20437);
xor U22872 (N_22872,N_19791,N_18609);
xor U22873 (N_22873,N_20016,N_18118);
or U22874 (N_22874,N_18944,N_19028);
nor U22875 (N_22875,N_19277,N_18450);
xnor U22876 (N_22876,N_18791,N_18707);
nand U22877 (N_22877,N_20205,N_18303);
and U22878 (N_22878,N_19924,N_18903);
or U22879 (N_22879,N_18137,N_19835);
and U22880 (N_22880,N_18166,N_18357);
nor U22881 (N_22881,N_18821,N_19720);
xor U22882 (N_22882,N_18395,N_20735);
or U22883 (N_22883,N_19783,N_19545);
nor U22884 (N_22884,N_18054,N_20682);
and U22885 (N_22885,N_20027,N_18078);
xor U22886 (N_22886,N_19401,N_19241);
nor U22887 (N_22887,N_20890,N_20591);
xor U22888 (N_22888,N_20428,N_18018);
nand U22889 (N_22889,N_19360,N_19291);
nor U22890 (N_22890,N_20563,N_19332);
nand U22891 (N_22891,N_20206,N_18627);
and U22892 (N_22892,N_20291,N_18829);
and U22893 (N_22893,N_20882,N_18734);
xor U22894 (N_22894,N_18128,N_20729);
or U22895 (N_22895,N_19487,N_18677);
nor U22896 (N_22896,N_19492,N_19334);
xnor U22897 (N_22897,N_19158,N_20102);
xnor U22898 (N_22898,N_20764,N_18579);
xor U22899 (N_22899,N_19795,N_20553);
nand U22900 (N_22900,N_18931,N_19010);
xor U22901 (N_22901,N_18076,N_20343);
or U22902 (N_22902,N_20366,N_18013);
xnor U22903 (N_22903,N_19085,N_19700);
and U22904 (N_22904,N_19571,N_20815);
xor U22905 (N_22905,N_20783,N_19142);
nand U22906 (N_22906,N_18331,N_19494);
nand U22907 (N_22907,N_19346,N_20747);
and U22908 (N_22908,N_20047,N_19871);
xor U22909 (N_22909,N_18525,N_18191);
xnor U22910 (N_22910,N_18563,N_18078);
xor U22911 (N_22911,N_18164,N_18729);
nand U22912 (N_22912,N_20110,N_19931);
nand U22913 (N_22913,N_18934,N_18705);
nor U22914 (N_22914,N_20284,N_20075);
or U22915 (N_22915,N_20001,N_19597);
or U22916 (N_22916,N_19632,N_18883);
nor U22917 (N_22917,N_19749,N_18607);
xor U22918 (N_22918,N_19601,N_18272);
xnor U22919 (N_22919,N_20023,N_19685);
xnor U22920 (N_22920,N_19468,N_19393);
or U22921 (N_22921,N_18960,N_20220);
nand U22922 (N_22922,N_18726,N_19074);
nor U22923 (N_22923,N_20227,N_19078);
nor U22924 (N_22924,N_18707,N_20051);
xor U22925 (N_22925,N_19190,N_20468);
or U22926 (N_22926,N_19543,N_20400);
nor U22927 (N_22927,N_19057,N_18825);
xnor U22928 (N_22928,N_18005,N_20312);
or U22929 (N_22929,N_20601,N_19701);
nand U22930 (N_22930,N_19157,N_20116);
nor U22931 (N_22931,N_19506,N_20945);
and U22932 (N_22932,N_20677,N_18195);
xor U22933 (N_22933,N_20444,N_18281);
and U22934 (N_22934,N_19808,N_19116);
nand U22935 (N_22935,N_19160,N_18199);
xnor U22936 (N_22936,N_20715,N_18912);
and U22937 (N_22937,N_19849,N_19281);
and U22938 (N_22938,N_20802,N_20373);
xor U22939 (N_22939,N_20519,N_18296);
xnor U22940 (N_22940,N_18004,N_20488);
or U22941 (N_22941,N_20862,N_20366);
and U22942 (N_22942,N_18813,N_19903);
xor U22943 (N_22943,N_18307,N_20085);
xor U22944 (N_22944,N_20818,N_19684);
and U22945 (N_22945,N_19723,N_19099);
and U22946 (N_22946,N_18705,N_18108);
nand U22947 (N_22947,N_19097,N_19162);
nor U22948 (N_22948,N_19566,N_20407);
nor U22949 (N_22949,N_20427,N_20498);
nor U22950 (N_22950,N_18120,N_19377);
nand U22951 (N_22951,N_20982,N_18225);
nor U22952 (N_22952,N_18169,N_19187);
and U22953 (N_22953,N_20587,N_18301);
and U22954 (N_22954,N_20808,N_19156);
and U22955 (N_22955,N_19925,N_19320);
nor U22956 (N_22956,N_20798,N_18714);
nor U22957 (N_22957,N_20355,N_19838);
nand U22958 (N_22958,N_18276,N_20725);
nor U22959 (N_22959,N_20552,N_20303);
or U22960 (N_22960,N_20496,N_18431);
xnor U22961 (N_22961,N_20119,N_20826);
and U22962 (N_22962,N_19688,N_20958);
nand U22963 (N_22963,N_18539,N_18193);
nor U22964 (N_22964,N_18979,N_20244);
or U22965 (N_22965,N_18139,N_19101);
xnor U22966 (N_22966,N_20244,N_20305);
nor U22967 (N_22967,N_19822,N_20790);
nand U22968 (N_22968,N_20370,N_19361);
xnor U22969 (N_22969,N_20308,N_19715);
and U22970 (N_22970,N_19186,N_19078);
or U22971 (N_22971,N_20418,N_18886);
and U22972 (N_22972,N_19019,N_18220);
nand U22973 (N_22973,N_19197,N_18140);
and U22974 (N_22974,N_18424,N_20047);
xor U22975 (N_22975,N_18757,N_18886);
nand U22976 (N_22976,N_19733,N_20198);
or U22977 (N_22977,N_19801,N_20239);
and U22978 (N_22978,N_19827,N_20299);
xor U22979 (N_22979,N_20544,N_18732);
xor U22980 (N_22980,N_19426,N_20846);
nor U22981 (N_22981,N_20877,N_19236);
nand U22982 (N_22982,N_19565,N_18399);
and U22983 (N_22983,N_19631,N_19091);
or U22984 (N_22984,N_20440,N_19848);
or U22985 (N_22985,N_19689,N_18671);
xnor U22986 (N_22986,N_20176,N_19625);
or U22987 (N_22987,N_18866,N_20094);
nand U22988 (N_22988,N_18085,N_20403);
and U22989 (N_22989,N_20007,N_18633);
nor U22990 (N_22990,N_19071,N_18844);
or U22991 (N_22991,N_18684,N_18895);
or U22992 (N_22992,N_20371,N_20950);
and U22993 (N_22993,N_20523,N_18171);
nand U22994 (N_22994,N_19674,N_18841);
nor U22995 (N_22995,N_19893,N_18843);
xor U22996 (N_22996,N_20639,N_19735);
or U22997 (N_22997,N_18302,N_20114);
nor U22998 (N_22998,N_18937,N_19270);
xor U22999 (N_22999,N_19257,N_19049);
nand U23000 (N_23000,N_20555,N_19932);
xor U23001 (N_23001,N_20545,N_18061);
xor U23002 (N_23002,N_19780,N_20020);
or U23003 (N_23003,N_18294,N_18239);
or U23004 (N_23004,N_18652,N_20567);
and U23005 (N_23005,N_20529,N_18480);
xnor U23006 (N_23006,N_20025,N_19261);
nor U23007 (N_23007,N_18841,N_20071);
nand U23008 (N_23008,N_20109,N_20137);
nor U23009 (N_23009,N_20532,N_18478);
nor U23010 (N_23010,N_20618,N_18775);
nor U23011 (N_23011,N_18311,N_18838);
nor U23012 (N_23012,N_20445,N_20828);
nor U23013 (N_23013,N_19566,N_20215);
xnor U23014 (N_23014,N_18878,N_20931);
nor U23015 (N_23015,N_18876,N_18371);
and U23016 (N_23016,N_18627,N_18527);
xor U23017 (N_23017,N_20408,N_18287);
nand U23018 (N_23018,N_20981,N_19010);
xnor U23019 (N_23019,N_19731,N_19049);
nand U23020 (N_23020,N_19294,N_19355);
xor U23021 (N_23021,N_20414,N_20921);
nand U23022 (N_23022,N_18584,N_19498);
and U23023 (N_23023,N_19098,N_20912);
and U23024 (N_23024,N_20508,N_18185);
or U23025 (N_23025,N_19811,N_20554);
xnor U23026 (N_23026,N_20458,N_20099);
and U23027 (N_23027,N_20561,N_18624);
xor U23028 (N_23028,N_18306,N_18424);
or U23029 (N_23029,N_18921,N_19328);
nand U23030 (N_23030,N_20669,N_19805);
and U23031 (N_23031,N_19109,N_20217);
nand U23032 (N_23032,N_20087,N_19373);
nand U23033 (N_23033,N_20994,N_18701);
and U23034 (N_23034,N_18920,N_18689);
nand U23035 (N_23035,N_19011,N_20915);
xor U23036 (N_23036,N_20414,N_20590);
nor U23037 (N_23037,N_18286,N_19003);
or U23038 (N_23038,N_19759,N_19502);
nand U23039 (N_23039,N_18939,N_19633);
nand U23040 (N_23040,N_20563,N_18497);
xnor U23041 (N_23041,N_19949,N_18207);
xor U23042 (N_23042,N_18832,N_19291);
nor U23043 (N_23043,N_18404,N_20272);
and U23044 (N_23044,N_18668,N_20977);
nor U23045 (N_23045,N_18680,N_19888);
or U23046 (N_23046,N_18890,N_19954);
and U23047 (N_23047,N_19866,N_19790);
xnor U23048 (N_23048,N_18192,N_20768);
or U23049 (N_23049,N_18093,N_19883);
nand U23050 (N_23050,N_20735,N_19527);
nand U23051 (N_23051,N_19480,N_19388);
nor U23052 (N_23052,N_19134,N_18294);
nand U23053 (N_23053,N_20333,N_18753);
nand U23054 (N_23054,N_19134,N_20417);
or U23055 (N_23055,N_20452,N_19316);
nand U23056 (N_23056,N_18605,N_20016);
nand U23057 (N_23057,N_18848,N_18689);
nor U23058 (N_23058,N_20398,N_20564);
nor U23059 (N_23059,N_20280,N_18177);
xnor U23060 (N_23060,N_18569,N_19701);
xor U23061 (N_23061,N_20701,N_20646);
and U23062 (N_23062,N_19716,N_20755);
and U23063 (N_23063,N_19025,N_19995);
nand U23064 (N_23064,N_19826,N_20607);
and U23065 (N_23065,N_18072,N_20034);
or U23066 (N_23066,N_20487,N_18788);
and U23067 (N_23067,N_20871,N_18025);
and U23068 (N_23068,N_18251,N_20712);
or U23069 (N_23069,N_19044,N_18462);
nor U23070 (N_23070,N_20247,N_19560);
xnor U23071 (N_23071,N_19271,N_18864);
or U23072 (N_23072,N_18567,N_19841);
and U23073 (N_23073,N_18334,N_20092);
nor U23074 (N_23074,N_20240,N_18875);
nor U23075 (N_23075,N_18644,N_18862);
or U23076 (N_23076,N_19311,N_20891);
xnor U23077 (N_23077,N_20610,N_18743);
and U23078 (N_23078,N_20167,N_20450);
xor U23079 (N_23079,N_20787,N_18246);
and U23080 (N_23080,N_20559,N_18528);
nand U23081 (N_23081,N_19286,N_20311);
nor U23082 (N_23082,N_19300,N_20653);
xnor U23083 (N_23083,N_19376,N_20180);
nor U23084 (N_23084,N_18306,N_19892);
and U23085 (N_23085,N_18293,N_19502);
or U23086 (N_23086,N_20409,N_19664);
and U23087 (N_23087,N_18219,N_19917);
nor U23088 (N_23088,N_20131,N_19468);
nor U23089 (N_23089,N_18291,N_18358);
or U23090 (N_23090,N_18300,N_20102);
and U23091 (N_23091,N_20683,N_20010);
nand U23092 (N_23092,N_20943,N_18671);
nor U23093 (N_23093,N_19658,N_20690);
xnor U23094 (N_23094,N_20328,N_19481);
nand U23095 (N_23095,N_19631,N_18711);
and U23096 (N_23096,N_19157,N_20104);
xor U23097 (N_23097,N_18790,N_20120);
nor U23098 (N_23098,N_20058,N_18301);
xor U23099 (N_23099,N_19670,N_20747);
nand U23100 (N_23100,N_20276,N_19776);
xnor U23101 (N_23101,N_18016,N_19391);
nor U23102 (N_23102,N_18379,N_20227);
nand U23103 (N_23103,N_19970,N_19868);
xnor U23104 (N_23104,N_20049,N_20346);
and U23105 (N_23105,N_19151,N_20205);
or U23106 (N_23106,N_18869,N_19021);
and U23107 (N_23107,N_18617,N_20037);
nor U23108 (N_23108,N_18249,N_19516);
and U23109 (N_23109,N_19112,N_18046);
nand U23110 (N_23110,N_19852,N_20603);
and U23111 (N_23111,N_18596,N_20749);
and U23112 (N_23112,N_20785,N_20014);
or U23113 (N_23113,N_20734,N_20091);
nor U23114 (N_23114,N_19298,N_20191);
and U23115 (N_23115,N_18233,N_18781);
xor U23116 (N_23116,N_19574,N_19249);
xor U23117 (N_23117,N_18449,N_19733);
nand U23118 (N_23118,N_19349,N_19472);
nand U23119 (N_23119,N_20827,N_18359);
or U23120 (N_23120,N_20372,N_20753);
nand U23121 (N_23121,N_18825,N_20718);
or U23122 (N_23122,N_18944,N_20723);
nand U23123 (N_23123,N_18672,N_18664);
and U23124 (N_23124,N_19504,N_20174);
and U23125 (N_23125,N_19094,N_20444);
xor U23126 (N_23126,N_19892,N_20333);
nor U23127 (N_23127,N_20368,N_18842);
nand U23128 (N_23128,N_19175,N_20239);
or U23129 (N_23129,N_19808,N_18653);
nor U23130 (N_23130,N_20855,N_19002);
and U23131 (N_23131,N_19111,N_18275);
nor U23132 (N_23132,N_20773,N_19065);
and U23133 (N_23133,N_19180,N_19722);
xnor U23134 (N_23134,N_19391,N_20615);
and U23135 (N_23135,N_20966,N_18482);
nand U23136 (N_23136,N_18583,N_18783);
nand U23137 (N_23137,N_20531,N_20054);
nand U23138 (N_23138,N_19671,N_20173);
nand U23139 (N_23139,N_20572,N_20169);
and U23140 (N_23140,N_20747,N_19659);
and U23141 (N_23141,N_20589,N_20378);
nor U23142 (N_23142,N_18841,N_20241);
xnor U23143 (N_23143,N_18237,N_20836);
or U23144 (N_23144,N_19989,N_18504);
and U23145 (N_23145,N_19195,N_20438);
nand U23146 (N_23146,N_20872,N_18440);
xor U23147 (N_23147,N_20093,N_19168);
nor U23148 (N_23148,N_19562,N_19926);
nand U23149 (N_23149,N_18513,N_20443);
xor U23150 (N_23150,N_18735,N_18345);
or U23151 (N_23151,N_20947,N_19845);
nand U23152 (N_23152,N_19309,N_18214);
or U23153 (N_23153,N_18722,N_18439);
xnor U23154 (N_23154,N_20743,N_20573);
nor U23155 (N_23155,N_19960,N_20253);
xnor U23156 (N_23156,N_18637,N_20499);
nand U23157 (N_23157,N_19855,N_20842);
xnor U23158 (N_23158,N_18593,N_18845);
nand U23159 (N_23159,N_20161,N_19166);
or U23160 (N_23160,N_18097,N_20287);
xnor U23161 (N_23161,N_18542,N_19147);
or U23162 (N_23162,N_18982,N_18223);
xnor U23163 (N_23163,N_20700,N_18810);
or U23164 (N_23164,N_20887,N_18236);
and U23165 (N_23165,N_18507,N_18165);
nand U23166 (N_23166,N_20984,N_19602);
or U23167 (N_23167,N_18625,N_19999);
or U23168 (N_23168,N_19761,N_19187);
xor U23169 (N_23169,N_20361,N_20068);
nor U23170 (N_23170,N_20264,N_18967);
xor U23171 (N_23171,N_18774,N_20254);
and U23172 (N_23172,N_20817,N_19628);
or U23173 (N_23173,N_19435,N_19254);
nor U23174 (N_23174,N_19696,N_18663);
xor U23175 (N_23175,N_20150,N_18633);
and U23176 (N_23176,N_19261,N_20903);
and U23177 (N_23177,N_19842,N_19784);
nand U23178 (N_23178,N_18993,N_19992);
xor U23179 (N_23179,N_19226,N_20692);
and U23180 (N_23180,N_20547,N_19325);
nor U23181 (N_23181,N_18831,N_18347);
nor U23182 (N_23182,N_20829,N_18149);
and U23183 (N_23183,N_20069,N_18351);
nor U23184 (N_23184,N_20946,N_18297);
or U23185 (N_23185,N_18221,N_19081);
and U23186 (N_23186,N_20819,N_20078);
or U23187 (N_23187,N_20328,N_20987);
or U23188 (N_23188,N_18273,N_18105);
nand U23189 (N_23189,N_19244,N_18937);
nor U23190 (N_23190,N_19167,N_18516);
nor U23191 (N_23191,N_20154,N_18700);
and U23192 (N_23192,N_20905,N_18983);
nor U23193 (N_23193,N_20756,N_18560);
xor U23194 (N_23194,N_18988,N_19633);
xor U23195 (N_23195,N_18032,N_19870);
nand U23196 (N_23196,N_20895,N_18792);
nand U23197 (N_23197,N_18961,N_18451);
nand U23198 (N_23198,N_20000,N_19522);
and U23199 (N_23199,N_20047,N_20668);
xor U23200 (N_23200,N_20432,N_20124);
nand U23201 (N_23201,N_18769,N_18475);
nor U23202 (N_23202,N_20057,N_19327);
nand U23203 (N_23203,N_20641,N_20887);
or U23204 (N_23204,N_18283,N_18864);
and U23205 (N_23205,N_20614,N_19153);
nor U23206 (N_23206,N_20502,N_19521);
and U23207 (N_23207,N_18596,N_20967);
nor U23208 (N_23208,N_18722,N_20213);
and U23209 (N_23209,N_18376,N_19433);
and U23210 (N_23210,N_20893,N_20602);
xor U23211 (N_23211,N_20296,N_19978);
xnor U23212 (N_23212,N_19183,N_18337);
nor U23213 (N_23213,N_18907,N_18710);
xnor U23214 (N_23214,N_20553,N_18743);
and U23215 (N_23215,N_19362,N_18928);
nor U23216 (N_23216,N_18167,N_18265);
xnor U23217 (N_23217,N_18747,N_19649);
nor U23218 (N_23218,N_19233,N_20643);
and U23219 (N_23219,N_18449,N_19338);
and U23220 (N_23220,N_19324,N_18945);
nand U23221 (N_23221,N_18412,N_19549);
or U23222 (N_23222,N_19261,N_19648);
and U23223 (N_23223,N_20656,N_19428);
and U23224 (N_23224,N_18240,N_20571);
nor U23225 (N_23225,N_18410,N_20712);
and U23226 (N_23226,N_19529,N_19376);
and U23227 (N_23227,N_18540,N_20000);
and U23228 (N_23228,N_18345,N_19407);
nand U23229 (N_23229,N_19487,N_19272);
nor U23230 (N_23230,N_20215,N_20923);
xor U23231 (N_23231,N_19087,N_19322);
or U23232 (N_23232,N_19347,N_19674);
or U23233 (N_23233,N_18003,N_18864);
nand U23234 (N_23234,N_18308,N_18058);
xor U23235 (N_23235,N_20123,N_18811);
nand U23236 (N_23236,N_18693,N_20412);
and U23237 (N_23237,N_18792,N_20365);
and U23238 (N_23238,N_19234,N_18179);
and U23239 (N_23239,N_19789,N_20770);
nor U23240 (N_23240,N_18834,N_20127);
nor U23241 (N_23241,N_18797,N_18241);
and U23242 (N_23242,N_20453,N_20259);
or U23243 (N_23243,N_18966,N_18423);
xnor U23244 (N_23244,N_19942,N_20328);
xor U23245 (N_23245,N_18241,N_19889);
nor U23246 (N_23246,N_20575,N_20186);
xor U23247 (N_23247,N_18547,N_19035);
or U23248 (N_23248,N_18770,N_19877);
and U23249 (N_23249,N_18438,N_19142);
and U23250 (N_23250,N_18945,N_20041);
or U23251 (N_23251,N_19607,N_19336);
and U23252 (N_23252,N_20951,N_19689);
nor U23253 (N_23253,N_18500,N_20939);
xnor U23254 (N_23254,N_19588,N_19950);
or U23255 (N_23255,N_19669,N_19249);
xnor U23256 (N_23256,N_18700,N_18216);
xor U23257 (N_23257,N_18761,N_20354);
or U23258 (N_23258,N_18548,N_18851);
xnor U23259 (N_23259,N_20752,N_19444);
or U23260 (N_23260,N_18773,N_18808);
nor U23261 (N_23261,N_19790,N_20576);
and U23262 (N_23262,N_20254,N_20927);
nor U23263 (N_23263,N_19722,N_20969);
xor U23264 (N_23264,N_19814,N_20300);
xor U23265 (N_23265,N_18312,N_20589);
nand U23266 (N_23266,N_19296,N_19656);
or U23267 (N_23267,N_19347,N_20535);
or U23268 (N_23268,N_19700,N_18481);
or U23269 (N_23269,N_18343,N_19318);
or U23270 (N_23270,N_20689,N_20017);
nand U23271 (N_23271,N_20771,N_20158);
and U23272 (N_23272,N_20845,N_19235);
or U23273 (N_23273,N_18101,N_18069);
xnor U23274 (N_23274,N_19882,N_19554);
or U23275 (N_23275,N_20119,N_19554);
nand U23276 (N_23276,N_18092,N_19706);
and U23277 (N_23277,N_19990,N_19120);
nor U23278 (N_23278,N_20782,N_18928);
and U23279 (N_23279,N_20794,N_18141);
and U23280 (N_23280,N_20816,N_18508);
xor U23281 (N_23281,N_20679,N_20865);
and U23282 (N_23282,N_19989,N_20065);
xor U23283 (N_23283,N_18690,N_20370);
and U23284 (N_23284,N_19875,N_20356);
and U23285 (N_23285,N_18779,N_19059);
nand U23286 (N_23286,N_20769,N_19853);
nor U23287 (N_23287,N_19197,N_18469);
nor U23288 (N_23288,N_18815,N_20972);
xor U23289 (N_23289,N_19352,N_18817);
or U23290 (N_23290,N_18295,N_20293);
nor U23291 (N_23291,N_18611,N_20893);
xor U23292 (N_23292,N_19697,N_18660);
nand U23293 (N_23293,N_19864,N_20532);
nand U23294 (N_23294,N_19594,N_20987);
xor U23295 (N_23295,N_19985,N_19181);
xor U23296 (N_23296,N_18132,N_18938);
and U23297 (N_23297,N_20114,N_20349);
nand U23298 (N_23298,N_20956,N_20364);
nor U23299 (N_23299,N_20711,N_18645);
and U23300 (N_23300,N_20455,N_20671);
nand U23301 (N_23301,N_19279,N_20468);
xnor U23302 (N_23302,N_20621,N_20773);
nand U23303 (N_23303,N_19129,N_18742);
nand U23304 (N_23304,N_18057,N_18699);
or U23305 (N_23305,N_20800,N_19078);
nand U23306 (N_23306,N_19168,N_19547);
nand U23307 (N_23307,N_19251,N_20718);
or U23308 (N_23308,N_18645,N_20068);
or U23309 (N_23309,N_18693,N_20669);
nand U23310 (N_23310,N_20324,N_18473);
and U23311 (N_23311,N_19531,N_20729);
or U23312 (N_23312,N_20380,N_18112);
xor U23313 (N_23313,N_20106,N_20121);
or U23314 (N_23314,N_18764,N_20459);
or U23315 (N_23315,N_20905,N_19202);
xnor U23316 (N_23316,N_20369,N_20705);
or U23317 (N_23317,N_18916,N_18725);
xnor U23318 (N_23318,N_20450,N_19682);
or U23319 (N_23319,N_18496,N_18220);
and U23320 (N_23320,N_18710,N_19654);
nor U23321 (N_23321,N_20157,N_18398);
nand U23322 (N_23322,N_18979,N_19741);
and U23323 (N_23323,N_19379,N_20435);
or U23324 (N_23324,N_20193,N_18135);
or U23325 (N_23325,N_18633,N_19305);
or U23326 (N_23326,N_19550,N_18347);
or U23327 (N_23327,N_18522,N_20555);
and U23328 (N_23328,N_20618,N_20412);
and U23329 (N_23329,N_20311,N_18499);
nor U23330 (N_23330,N_20035,N_19973);
nor U23331 (N_23331,N_19131,N_18864);
or U23332 (N_23332,N_19809,N_19959);
nor U23333 (N_23333,N_18605,N_20578);
and U23334 (N_23334,N_18377,N_19351);
xor U23335 (N_23335,N_20288,N_19049);
or U23336 (N_23336,N_18552,N_19564);
or U23337 (N_23337,N_18778,N_20305);
nor U23338 (N_23338,N_19796,N_20342);
xnor U23339 (N_23339,N_20114,N_18989);
xnor U23340 (N_23340,N_20515,N_18391);
nor U23341 (N_23341,N_20020,N_20133);
nor U23342 (N_23342,N_20798,N_19182);
xor U23343 (N_23343,N_19544,N_20447);
xnor U23344 (N_23344,N_20473,N_19909);
nor U23345 (N_23345,N_18557,N_20845);
nand U23346 (N_23346,N_18625,N_20176);
nor U23347 (N_23347,N_18928,N_18948);
and U23348 (N_23348,N_20138,N_18988);
or U23349 (N_23349,N_18189,N_20171);
nand U23350 (N_23350,N_19811,N_18201);
nand U23351 (N_23351,N_20208,N_20161);
and U23352 (N_23352,N_20648,N_18987);
or U23353 (N_23353,N_18864,N_19495);
xor U23354 (N_23354,N_18336,N_18875);
and U23355 (N_23355,N_19468,N_19136);
nand U23356 (N_23356,N_18057,N_19321);
or U23357 (N_23357,N_18122,N_20326);
and U23358 (N_23358,N_19601,N_19302);
or U23359 (N_23359,N_18457,N_19219);
or U23360 (N_23360,N_18013,N_19395);
or U23361 (N_23361,N_20878,N_18074);
nor U23362 (N_23362,N_20835,N_19673);
or U23363 (N_23363,N_20122,N_19513);
xor U23364 (N_23364,N_19980,N_18922);
xnor U23365 (N_23365,N_18876,N_20536);
or U23366 (N_23366,N_20885,N_18892);
xnor U23367 (N_23367,N_20658,N_19925);
nand U23368 (N_23368,N_18853,N_19774);
or U23369 (N_23369,N_18830,N_19954);
nand U23370 (N_23370,N_18605,N_18842);
xor U23371 (N_23371,N_20511,N_20933);
nor U23372 (N_23372,N_20418,N_20054);
and U23373 (N_23373,N_18817,N_18876);
and U23374 (N_23374,N_19554,N_18911);
and U23375 (N_23375,N_18911,N_19085);
nand U23376 (N_23376,N_20799,N_19969);
nor U23377 (N_23377,N_20536,N_18997);
nor U23378 (N_23378,N_19462,N_19527);
and U23379 (N_23379,N_18501,N_19863);
xnor U23380 (N_23380,N_19411,N_19472);
xnor U23381 (N_23381,N_18959,N_19997);
nand U23382 (N_23382,N_19944,N_20003);
or U23383 (N_23383,N_20052,N_18890);
or U23384 (N_23384,N_19354,N_18362);
and U23385 (N_23385,N_19116,N_20869);
and U23386 (N_23386,N_19985,N_19770);
nand U23387 (N_23387,N_20891,N_19871);
xor U23388 (N_23388,N_18159,N_19856);
nor U23389 (N_23389,N_19077,N_20169);
and U23390 (N_23390,N_19533,N_18929);
nor U23391 (N_23391,N_20573,N_19150);
xor U23392 (N_23392,N_18307,N_18713);
nand U23393 (N_23393,N_20977,N_18532);
xnor U23394 (N_23394,N_18612,N_18841);
xnor U23395 (N_23395,N_20403,N_20570);
or U23396 (N_23396,N_19241,N_20252);
xor U23397 (N_23397,N_19193,N_18547);
xor U23398 (N_23398,N_19531,N_18812);
xor U23399 (N_23399,N_18643,N_20062);
xor U23400 (N_23400,N_19253,N_20423);
nor U23401 (N_23401,N_20452,N_20482);
nor U23402 (N_23402,N_20808,N_18644);
xor U23403 (N_23403,N_19971,N_18581);
and U23404 (N_23404,N_18714,N_20096);
xnor U23405 (N_23405,N_19623,N_20214);
and U23406 (N_23406,N_18007,N_19970);
or U23407 (N_23407,N_18715,N_18328);
nor U23408 (N_23408,N_20316,N_18225);
nor U23409 (N_23409,N_20057,N_18961);
nor U23410 (N_23410,N_19034,N_18800);
and U23411 (N_23411,N_19829,N_18333);
xor U23412 (N_23412,N_19880,N_19484);
or U23413 (N_23413,N_19017,N_19793);
and U23414 (N_23414,N_18245,N_20418);
and U23415 (N_23415,N_19412,N_19020);
and U23416 (N_23416,N_19884,N_19276);
nor U23417 (N_23417,N_18750,N_20321);
or U23418 (N_23418,N_18160,N_19590);
xor U23419 (N_23419,N_19953,N_19802);
and U23420 (N_23420,N_20463,N_18980);
and U23421 (N_23421,N_20609,N_19187);
nand U23422 (N_23422,N_20321,N_20819);
xnor U23423 (N_23423,N_18614,N_18599);
nor U23424 (N_23424,N_19281,N_20803);
xnor U23425 (N_23425,N_18059,N_20107);
and U23426 (N_23426,N_19842,N_20116);
nand U23427 (N_23427,N_20216,N_19162);
nor U23428 (N_23428,N_19452,N_18502);
and U23429 (N_23429,N_18635,N_20153);
xor U23430 (N_23430,N_18389,N_18661);
nand U23431 (N_23431,N_19326,N_19584);
nand U23432 (N_23432,N_20332,N_19191);
and U23433 (N_23433,N_18807,N_19989);
xor U23434 (N_23434,N_20327,N_18288);
nand U23435 (N_23435,N_19770,N_18322);
or U23436 (N_23436,N_18214,N_18383);
nor U23437 (N_23437,N_20321,N_19745);
nand U23438 (N_23438,N_20438,N_20086);
nor U23439 (N_23439,N_20942,N_18663);
and U23440 (N_23440,N_20798,N_18475);
nand U23441 (N_23441,N_19619,N_20049);
or U23442 (N_23442,N_20430,N_18015);
xnor U23443 (N_23443,N_18297,N_18400);
xor U23444 (N_23444,N_20957,N_20655);
or U23445 (N_23445,N_18001,N_19511);
or U23446 (N_23446,N_20478,N_19394);
nand U23447 (N_23447,N_18746,N_18798);
and U23448 (N_23448,N_20065,N_19171);
and U23449 (N_23449,N_18661,N_19940);
nor U23450 (N_23450,N_18859,N_18239);
and U23451 (N_23451,N_18310,N_19191);
and U23452 (N_23452,N_18294,N_19455);
xor U23453 (N_23453,N_18086,N_19149);
nor U23454 (N_23454,N_18224,N_18043);
and U23455 (N_23455,N_20632,N_18385);
xnor U23456 (N_23456,N_19016,N_18881);
and U23457 (N_23457,N_18004,N_18554);
or U23458 (N_23458,N_19261,N_18060);
nand U23459 (N_23459,N_18218,N_18753);
or U23460 (N_23460,N_18088,N_19269);
nor U23461 (N_23461,N_20440,N_19316);
nor U23462 (N_23462,N_18407,N_19600);
and U23463 (N_23463,N_18590,N_18493);
xnor U23464 (N_23464,N_20257,N_19658);
and U23465 (N_23465,N_18127,N_20022);
xor U23466 (N_23466,N_19751,N_18256);
xnor U23467 (N_23467,N_19106,N_20183);
xor U23468 (N_23468,N_18382,N_18650);
and U23469 (N_23469,N_19492,N_18311);
xor U23470 (N_23470,N_19491,N_18211);
and U23471 (N_23471,N_19885,N_18061);
xnor U23472 (N_23472,N_18860,N_19319);
or U23473 (N_23473,N_18269,N_18763);
and U23474 (N_23474,N_20516,N_18474);
and U23475 (N_23475,N_19057,N_18189);
nor U23476 (N_23476,N_18449,N_18730);
nand U23477 (N_23477,N_18692,N_18989);
and U23478 (N_23478,N_18282,N_18902);
nor U23479 (N_23479,N_18703,N_19187);
and U23480 (N_23480,N_19718,N_20079);
and U23481 (N_23481,N_19458,N_20080);
nand U23482 (N_23482,N_18031,N_18756);
xnor U23483 (N_23483,N_19858,N_18373);
or U23484 (N_23484,N_20099,N_19340);
and U23485 (N_23485,N_19584,N_19687);
nand U23486 (N_23486,N_20650,N_19071);
or U23487 (N_23487,N_19525,N_18853);
nor U23488 (N_23488,N_18641,N_20360);
and U23489 (N_23489,N_18351,N_20781);
nand U23490 (N_23490,N_18896,N_19280);
nor U23491 (N_23491,N_20467,N_19491);
xnor U23492 (N_23492,N_18505,N_19572);
and U23493 (N_23493,N_19405,N_20430);
nand U23494 (N_23494,N_19900,N_20231);
xor U23495 (N_23495,N_19941,N_20575);
and U23496 (N_23496,N_18278,N_19208);
and U23497 (N_23497,N_18357,N_19150);
and U23498 (N_23498,N_20935,N_20918);
and U23499 (N_23499,N_18653,N_19112);
and U23500 (N_23500,N_20470,N_19493);
nor U23501 (N_23501,N_19635,N_20677);
or U23502 (N_23502,N_20776,N_20800);
nor U23503 (N_23503,N_18807,N_20604);
xor U23504 (N_23504,N_18059,N_19197);
nand U23505 (N_23505,N_18080,N_18399);
and U23506 (N_23506,N_20763,N_20725);
xnor U23507 (N_23507,N_20186,N_18452);
or U23508 (N_23508,N_19660,N_20667);
or U23509 (N_23509,N_18301,N_18881);
or U23510 (N_23510,N_18998,N_19140);
nand U23511 (N_23511,N_18448,N_19594);
nand U23512 (N_23512,N_19494,N_19628);
nand U23513 (N_23513,N_18594,N_20869);
nor U23514 (N_23514,N_20075,N_20125);
or U23515 (N_23515,N_19403,N_20210);
nor U23516 (N_23516,N_18008,N_19063);
and U23517 (N_23517,N_18811,N_19439);
or U23518 (N_23518,N_19632,N_18156);
and U23519 (N_23519,N_19589,N_20803);
nand U23520 (N_23520,N_18467,N_19364);
xnor U23521 (N_23521,N_19591,N_19076);
or U23522 (N_23522,N_18696,N_18419);
or U23523 (N_23523,N_20448,N_20767);
nor U23524 (N_23524,N_20418,N_18993);
nor U23525 (N_23525,N_20591,N_18157);
nand U23526 (N_23526,N_18690,N_19323);
or U23527 (N_23527,N_18876,N_20759);
xnor U23528 (N_23528,N_20071,N_18018);
and U23529 (N_23529,N_20186,N_18527);
nand U23530 (N_23530,N_20924,N_20222);
xor U23531 (N_23531,N_19888,N_18143);
and U23532 (N_23532,N_18406,N_19663);
or U23533 (N_23533,N_19060,N_20743);
xor U23534 (N_23534,N_20382,N_20791);
nor U23535 (N_23535,N_18054,N_19119);
nand U23536 (N_23536,N_20970,N_20680);
and U23537 (N_23537,N_20366,N_20643);
or U23538 (N_23538,N_20795,N_18381);
nand U23539 (N_23539,N_18712,N_20571);
or U23540 (N_23540,N_19538,N_18054);
nand U23541 (N_23541,N_18148,N_18788);
xor U23542 (N_23542,N_20274,N_19807);
or U23543 (N_23543,N_20504,N_20876);
or U23544 (N_23544,N_19841,N_18002);
nor U23545 (N_23545,N_19038,N_20722);
and U23546 (N_23546,N_20626,N_19220);
and U23547 (N_23547,N_18545,N_19620);
nand U23548 (N_23548,N_19490,N_20628);
and U23549 (N_23549,N_19397,N_19039);
nor U23550 (N_23550,N_19717,N_18353);
and U23551 (N_23551,N_19199,N_19887);
nor U23552 (N_23552,N_20422,N_19713);
nor U23553 (N_23553,N_18148,N_18898);
nand U23554 (N_23554,N_20292,N_20865);
nor U23555 (N_23555,N_19575,N_19484);
nand U23556 (N_23556,N_20971,N_18262);
xnor U23557 (N_23557,N_18848,N_20729);
nand U23558 (N_23558,N_19442,N_20049);
and U23559 (N_23559,N_18661,N_18433);
or U23560 (N_23560,N_19286,N_20391);
and U23561 (N_23561,N_19776,N_20026);
or U23562 (N_23562,N_18021,N_20932);
nand U23563 (N_23563,N_18348,N_18980);
and U23564 (N_23564,N_19930,N_20542);
or U23565 (N_23565,N_20733,N_18255);
and U23566 (N_23566,N_18711,N_18977);
and U23567 (N_23567,N_18526,N_19734);
and U23568 (N_23568,N_18392,N_18561);
xnor U23569 (N_23569,N_19376,N_20172);
nor U23570 (N_23570,N_19841,N_18133);
nor U23571 (N_23571,N_20466,N_20440);
xor U23572 (N_23572,N_18228,N_20963);
or U23573 (N_23573,N_19403,N_20158);
nand U23574 (N_23574,N_19655,N_19613);
nand U23575 (N_23575,N_18143,N_20086);
nand U23576 (N_23576,N_18241,N_18158);
xor U23577 (N_23577,N_19849,N_20374);
nor U23578 (N_23578,N_19530,N_18501);
nand U23579 (N_23579,N_18008,N_18880);
nand U23580 (N_23580,N_18499,N_18008);
or U23581 (N_23581,N_20610,N_19297);
nor U23582 (N_23582,N_18951,N_18402);
or U23583 (N_23583,N_19171,N_20478);
or U23584 (N_23584,N_19569,N_18751);
and U23585 (N_23585,N_19252,N_18767);
and U23586 (N_23586,N_19086,N_19340);
or U23587 (N_23587,N_19481,N_18064);
and U23588 (N_23588,N_19755,N_20450);
and U23589 (N_23589,N_19395,N_20897);
nand U23590 (N_23590,N_18694,N_20004);
nand U23591 (N_23591,N_18040,N_20853);
nand U23592 (N_23592,N_20319,N_20381);
and U23593 (N_23593,N_20326,N_19617);
nand U23594 (N_23594,N_19905,N_20024);
nand U23595 (N_23595,N_18079,N_19268);
or U23596 (N_23596,N_18982,N_18995);
nand U23597 (N_23597,N_20158,N_19404);
nor U23598 (N_23598,N_20559,N_20573);
or U23599 (N_23599,N_20090,N_19941);
and U23600 (N_23600,N_19950,N_20276);
and U23601 (N_23601,N_19021,N_18354);
nand U23602 (N_23602,N_18658,N_20352);
nand U23603 (N_23603,N_19335,N_19090);
nand U23604 (N_23604,N_20786,N_20291);
nor U23605 (N_23605,N_18541,N_18172);
xor U23606 (N_23606,N_19025,N_20500);
nor U23607 (N_23607,N_19019,N_20533);
nor U23608 (N_23608,N_20903,N_20228);
nand U23609 (N_23609,N_20011,N_20424);
nor U23610 (N_23610,N_20844,N_20412);
and U23611 (N_23611,N_19426,N_20003);
nor U23612 (N_23612,N_20793,N_20096);
xor U23613 (N_23613,N_20278,N_20570);
and U23614 (N_23614,N_20318,N_19770);
or U23615 (N_23615,N_20954,N_19679);
nor U23616 (N_23616,N_18330,N_18508);
nor U23617 (N_23617,N_20558,N_18688);
nor U23618 (N_23618,N_18971,N_20081);
and U23619 (N_23619,N_18646,N_18595);
and U23620 (N_23620,N_20682,N_19856);
nand U23621 (N_23621,N_20280,N_20633);
nor U23622 (N_23622,N_19394,N_18510);
or U23623 (N_23623,N_20866,N_19941);
or U23624 (N_23624,N_20601,N_19155);
nor U23625 (N_23625,N_19900,N_20853);
nor U23626 (N_23626,N_19781,N_18696);
and U23627 (N_23627,N_19384,N_18874);
nand U23628 (N_23628,N_18483,N_19195);
nor U23629 (N_23629,N_20845,N_19434);
nand U23630 (N_23630,N_19611,N_18541);
nand U23631 (N_23631,N_19510,N_19191);
xnor U23632 (N_23632,N_20717,N_20038);
nor U23633 (N_23633,N_20169,N_18499);
nor U23634 (N_23634,N_18809,N_18900);
xnor U23635 (N_23635,N_20964,N_18766);
nand U23636 (N_23636,N_20299,N_18780);
xnor U23637 (N_23637,N_19443,N_18188);
nor U23638 (N_23638,N_18076,N_18341);
nor U23639 (N_23639,N_19491,N_18844);
and U23640 (N_23640,N_20341,N_20490);
xnor U23641 (N_23641,N_20861,N_18033);
or U23642 (N_23642,N_20757,N_19080);
xnor U23643 (N_23643,N_18108,N_20618);
and U23644 (N_23644,N_19190,N_19599);
or U23645 (N_23645,N_19343,N_18455);
nand U23646 (N_23646,N_20157,N_18044);
or U23647 (N_23647,N_19257,N_19639);
xnor U23648 (N_23648,N_19024,N_20352);
nand U23649 (N_23649,N_20059,N_18916);
or U23650 (N_23650,N_20839,N_18195);
and U23651 (N_23651,N_19819,N_20590);
xor U23652 (N_23652,N_20392,N_18647);
nand U23653 (N_23653,N_20797,N_18017);
nor U23654 (N_23654,N_19061,N_18168);
and U23655 (N_23655,N_20610,N_18128);
or U23656 (N_23656,N_18219,N_20871);
or U23657 (N_23657,N_18124,N_19699);
nor U23658 (N_23658,N_20964,N_20412);
nor U23659 (N_23659,N_20712,N_19105);
nor U23660 (N_23660,N_20051,N_19977);
xnor U23661 (N_23661,N_20235,N_19074);
xnor U23662 (N_23662,N_20250,N_18584);
xor U23663 (N_23663,N_18948,N_20544);
nor U23664 (N_23664,N_20445,N_19680);
and U23665 (N_23665,N_19042,N_20533);
xor U23666 (N_23666,N_19553,N_19704);
and U23667 (N_23667,N_18010,N_20904);
nand U23668 (N_23668,N_18716,N_20776);
xnor U23669 (N_23669,N_20211,N_18299);
and U23670 (N_23670,N_19464,N_19102);
and U23671 (N_23671,N_19926,N_20012);
nand U23672 (N_23672,N_20803,N_18242);
and U23673 (N_23673,N_19541,N_18478);
xor U23674 (N_23674,N_19457,N_20769);
xor U23675 (N_23675,N_20347,N_19276);
or U23676 (N_23676,N_20462,N_20216);
nand U23677 (N_23677,N_19485,N_20634);
xnor U23678 (N_23678,N_19969,N_19429);
nand U23679 (N_23679,N_19819,N_18723);
xnor U23680 (N_23680,N_18635,N_18845);
or U23681 (N_23681,N_18723,N_20415);
or U23682 (N_23682,N_20572,N_18212);
or U23683 (N_23683,N_18808,N_18126);
xor U23684 (N_23684,N_19869,N_18884);
nor U23685 (N_23685,N_20807,N_20114);
or U23686 (N_23686,N_18920,N_20161);
xor U23687 (N_23687,N_20729,N_20884);
or U23688 (N_23688,N_18134,N_20816);
nor U23689 (N_23689,N_18144,N_20279);
nand U23690 (N_23690,N_20633,N_19387);
nor U23691 (N_23691,N_18489,N_19128);
or U23692 (N_23692,N_20042,N_20070);
nand U23693 (N_23693,N_20726,N_19489);
xor U23694 (N_23694,N_18888,N_18129);
or U23695 (N_23695,N_19307,N_19564);
or U23696 (N_23696,N_19755,N_19316);
nor U23697 (N_23697,N_19720,N_20778);
and U23698 (N_23698,N_19646,N_19699);
nor U23699 (N_23699,N_20702,N_20771);
or U23700 (N_23700,N_18034,N_20603);
and U23701 (N_23701,N_19057,N_20964);
xnor U23702 (N_23702,N_19795,N_19141);
or U23703 (N_23703,N_18306,N_20965);
nor U23704 (N_23704,N_18637,N_19487);
nand U23705 (N_23705,N_18122,N_20150);
or U23706 (N_23706,N_19911,N_20089);
nor U23707 (N_23707,N_18729,N_18181);
nand U23708 (N_23708,N_19948,N_18780);
or U23709 (N_23709,N_19053,N_20333);
and U23710 (N_23710,N_19750,N_18961);
and U23711 (N_23711,N_20216,N_18427);
nand U23712 (N_23712,N_19660,N_18775);
nand U23713 (N_23713,N_19218,N_18078);
nand U23714 (N_23714,N_20552,N_20715);
nand U23715 (N_23715,N_18857,N_19287);
or U23716 (N_23716,N_18996,N_18219);
nand U23717 (N_23717,N_19916,N_20642);
xnor U23718 (N_23718,N_19353,N_20694);
and U23719 (N_23719,N_18746,N_19184);
nand U23720 (N_23720,N_18942,N_18425);
and U23721 (N_23721,N_18994,N_20705);
or U23722 (N_23722,N_18013,N_19203);
xnor U23723 (N_23723,N_19341,N_18709);
or U23724 (N_23724,N_18156,N_18092);
and U23725 (N_23725,N_18477,N_18389);
nor U23726 (N_23726,N_19680,N_20992);
xnor U23727 (N_23727,N_18258,N_19459);
nand U23728 (N_23728,N_20778,N_20352);
xnor U23729 (N_23729,N_18028,N_18439);
or U23730 (N_23730,N_19396,N_18677);
nor U23731 (N_23731,N_20150,N_19298);
xnor U23732 (N_23732,N_18057,N_19559);
nor U23733 (N_23733,N_19429,N_20673);
and U23734 (N_23734,N_18806,N_20078);
xor U23735 (N_23735,N_18221,N_19509);
nand U23736 (N_23736,N_18927,N_19138);
nor U23737 (N_23737,N_19136,N_18291);
and U23738 (N_23738,N_18789,N_18170);
nand U23739 (N_23739,N_20006,N_20285);
nor U23740 (N_23740,N_20198,N_20391);
or U23741 (N_23741,N_20758,N_20245);
nand U23742 (N_23742,N_20825,N_20681);
nor U23743 (N_23743,N_19422,N_19455);
and U23744 (N_23744,N_20635,N_19191);
nand U23745 (N_23745,N_19376,N_20808);
and U23746 (N_23746,N_18085,N_18096);
nor U23747 (N_23747,N_19354,N_20636);
nor U23748 (N_23748,N_18802,N_20810);
nand U23749 (N_23749,N_18031,N_20473);
nor U23750 (N_23750,N_18510,N_20429);
xnor U23751 (N_23751,N_20221,N_20200);
xnor U23752 (N_23752,N_20696,N_18978);
or U23753 (N_23753,N_19690,N_20445);
xor U23754 (N_23754,N_20933,N_20224);
nand U23755 (N_23755,N_19072,N_20583);
nand U23756 (N_23756,N_19977,N_19410);
xnor U23757 (N_23757,N_18217,N_18299);
nand U23758 (N_23758,N_20359,N_20463);
or U23759 (N_23759,N_20241,N_18415);
or U23760 (N_23760,N_18452,N_19043);
xnor U23761 (N_23761,N_20787,N_20236);
xor U23762 (N_23762,N_18192,N_20551);
xnor U23763 (N_23763,N_19760,N_20174);
and U23764 (N_23764,N_19408,N_19416);
nand U23765 (N_23765,N_19213,N_20951);
nor U23766 (N_23766,N_19418,N_19531);
nand U23767 (N_23767,N_18149,N_19448);
or U23768 (N_23768,N_20230,N_20462);
nor U23769 (N_23769,N_20105,N_18032);
nand U23770 (N_23770,N_18073,N_18299);
or U23771 (N_23771,N_20460,N_20156);
nand U23772 (N_23772,N_20661,N_20236);
or U23773 (N_23773,N_20807,N_19621);
and U23774 (N_23774,N_18635,N_20085);
xnor U23775 (N_23775,N_19582,N_20277);
xor U23776 (N_23776,N_20636,N_19697);
and U23777 (N_23777,N_19621,N_18450);
nand U23778 (N_23778,N_19167,N_20349);
and U23779 (N_23779,N_20129,N_20591);
nor U23780 (N_23780,N_18670,N_18408);
and U23781 (N_23781,N_20007,N_20705);
nor U23782 (N_23782,N_18146,N_20468);
or U23783 (N_23783,N_18817,N_19792);
nor U23784 (N_23784,N_19368,N_20651);
xor U23785 (N_23785,N_20414,N_19773);
xnor U23786 (N_23786,N_19828,N_18366);
xnor U23787 (N_23787,N_18826,N_18063);
and U23788 (N_23788,N_19902,N_20910);
and U23789 (N_23789,N_19229,N_20249);
or U23790 (N_23790,N_20546,N_20534);
nor U23791 (N_23791,N_19072,N_20209);
or U23792 (N_23792,N_20417,N_19801);
xor U23793 (N_23793,N_20093,N_18613);
nand U23794 (N_23794,N_18738,N_18097);
nor U23795 (N_23795,N_20578,N_20673);
or U23796 (N_23796,N_18671,N_19880);
and U23797 (N_23797,N_18257,N_19595);
and U23798 (N_23798,N_18433,N_19532);
and U23799 (N_23799,N_20574,N_18923);
xnor U23800 (N_23800,N_18046,N_20942);
xor U23801 (N_23801,N_18378,N_18319);
nand U23802 (N_23802,N_18705,N_20570);
xor U23803 (N_23803,N_18377,N_20354);
and U23804 (N_23804,N_18753,N_20503);
xor U23805 (N_23805,N_20012,N_20773);
nor U23806 (N_23806,N_18378,N_18023);
and U23807 (N_23807,N_19480,N_18916);
xnor U23808 (N_23808,N_20445,N_20553);
or U23809 (N_23809,N_19124,N_19672);
xor U23810 (N_23810,N_18193,N_20252);
or U23811 (N_23811,N_19287,N_18957);
nand U23812 (N_23812,N_18269,N_20856);
or U23813 (N_23813,N_19888,N_18440);
nand U23814 (N_23814,N_19892,N_20891);
and U23815 (N_23815,N_18663,N_19079);
and U23816 (N_23816,N_19288,N_18992);
nand U23817 (N_23817,N_20575,N_18635);
nand U23818 (N_23818,N_18233,N_18656);
and U23819 (N_23819,N_20803,N_18742);
xor U23820 (N_23820,N_19587,N_19076);
and U23821 (N_23821,N_18377,N_20823);
or U23822 (N_23822,N_18936,N_19708);
nand U23823 (N_23823,N_18628,N_18368);
nor U23824 (N_23824,N_18027,N_19390);
nand U23825 (N_23825,N_19114,N_20207);
nor U23826 (N_23826,N_18426,N_19699);
or U23827 (N_23827,N_18448,N_19347);
nand U23828 (N_23828,N_20485,N_19425);
nor U23829 (N_23829,N_18615,N_19910);
and U23830 (N_23830,N_19119,N_20167);
nand U23831 (N_23831,N_19210,N_19098);
and U23832 (N_23832,N_20900,N_20877);
or U23833 (N_23833,N_19019,N_19422);
and U23834 (N_23834,N_19536,N_18908);
xor U23835 (N_23835,N_20315,N_18387);
xnor U23836 (N_23836,N_18023,N_20866);
and U23837 (N_23837,N_19612,N_18776);
or U23838 (N_23838,N_18687,N_20742);
nand U23839 (N_23839,N_18693,N_19781);
or U23840 (N_23840,N_19573,N_18796);
or U23841 (N_23841,N_18468,N_19381);
and U23842 (N_23842,N_20547,N_18045);
nor U23843 (N_23843,N_20509,N_20057);
xnor U23844 (N_23844,N_18561,N_19894);
nor U23845 (N_23845,N_19314,N_19862);
nor U23846 (N_23846,N_19354,N_19580);
nor U23847 (N_23847,N_19363,N_18859);
or U23848 (N_23848,N_18626,N_19028);
xor U23849 (N_23849,N_19543,N_18510);
xor U23850 (N_23850,N_20469,N_20381);
or U23851 (N_23851,N_20659,N_20991);
nand U23852 (N_23852,N_20571,N_18258);
and U23853 (N_23853,N_18003,N_18120);
xnor U23854 (N_23854,N_19200,N_20020);
xor U23855 (N_23855,N_18942,N_18656);
nand U23856 (N_23856,N_20735,N_19418);
xnor U23857 (N_23857,N_19502,N_18786);
xor U23858 (N_23858,N_19123,N_18639);
nand U23859 (N_23859,N_20773,N_18472);
nand U23860 (N_23860,N_20005,N_19346);
or U23861 (N_23861,N_20497,N_18619);
nand U23862 (N_23862,N_20176,N_19729);
or U23863 (N_23863,N_19427,N_18876);
and U23864 (N_23864,N_20314,N_19615);
xnor U23865 (N_23865,N_19825,N_20856);
and U23866 (N_23866,N_18701,N_18402);
nand U23867 (N_23867,N_19834,N_20148);
nor U23868 (N_23868,N_20593,N_20676);
nand U23869 (N_23869,N_19287,N_20088);
nand U23870 (N_23870,N_19573,N_19822);
xor U23871 (N_23871,N_20737,N_19301);
and U23872 (N_23872,N_18951,N_18837);
or U23873 (N_23873,N_19503,N_19358);
xnor U23874 (N_23874,N_19308,N_20300);
xnor U23875 (N_23875,N_18713,N_20978);
xor U23876 (N_23876,N_18596,N_19333);
or U23877 (N_23877,N_20802,N_18134);
or U23878 (N_23878,N_19753,N_18717);
nor U23879 (N_23879,N_20155,N_20725);
nand U23880 (N_23880,N_20214,N_18387);
nand U23881 (N_23881,N_18531,N_20250);
and U23882 (N_23882,N_20374,N_19867);
nor U23883 (N_23883,N_18130,N_20187);
nand U23884 (N_23884,N_20356,N_19265);
xnor U23885 (N_23885,N_18098,N_19872);
nand U23886 (N_23886,N_19698,N_19689);
xor U23887 (N_23887,N_19796,N_20131);
and U23888 (N_23888,N_19533,N_19753);
nand U23889 (N_23889,N_18519,N_18062);
nand U23890 (N_23890,N_20766,N_18818);
nor U23891 (N_23891,N_20843,N_18184);
nor U23892 (N_23892,N_18595,N_18005);
nand U23893 (N_23893,N_18485,N_19127);
nor U23894 (N_23894,N_18768,N_18166);
or U23895 (N_23895,N_19636,N_20578);
xor U23896 (N_23896,N_19952,N_20065);
nor U23897 (N_23897,N_19071,N_18952);
xor U23898 (N_23898,N_18322,N_19396);
nor U23899 (N_23899,N_19972,N_20764);
xor U23900 (N_23900,N_20485,N_18806);
nor U23901 (N_23901,N_18669,N_19986);
and U23902 (N_23902,N_19456,N_20574);
and U23903 (N_23903,N_19673,N_18212);
nor U23904 (N_23904,N_18947,N_18952);
or U23905 (N_23905,N_20274,N_20740);
or U23906 (N_23906,N_19308,N_20188);
nand U23907 (N_23907,N_20999,N_18655);
or U23908 (N_23908,N_18502,N_18626);
xnor U23909 (N_23909,N_18101,N_19536);
xnor U23910 (N_23910,N_20266,N_19744);
nand U23911 (N_23911,N_19518,N_19955);
or U23912 (N_23912,N_19518,N_19464);
and U23913 (N_23913,N_19531,N_19305);
and U23914 (N_23914,N_19717,N_19062);
xor U23915 (N_23915,N_20173,N_20865);
or U23916 (N_23916,N_20044,N_19520);
nand U23917 (N_23917,N_19827,N_20339);
and U23918 (N_23918,N_20765,N_20928);
xnor U23919 (N_23919,N_20162,N_20566);
nor U23920 (N_23920,N_18333,N_19613);
or U23921 (N_23921,N_19189,N_18297);
or U23922 (N_23922,N_19076,N_18759);
nor U23923 (N_23923,N_20598,N_19941);
xnor U23924 (N_23924,N_20779,N_18448);
nand U23925 (N_23925,N_20645,N_19663);
and U23926 (N_23926,N_20881,N_20232);
and U23927 (N_23927,N_18012,N_20427);
and U23928 (N_23928,N_20110,N_19030);
nor U23929 (N_23929,N_19880,N_18766);
nand U23930 (N_23930,N_19415,N_18017);
or U23931 (N_23931,N_20727,N_19530);
or U23932 (N_23932,N_19959,N_19788);
nor U23933 (N_23933,N_20703,N_19330);
nand U23934 (N_23934,N_20937,N_18840);
xor U23935 (N_23935,N_19997,N_19184);
nand U23936 (N_23936,N_20127,N_20616);
and U23937 (N_23937,N_19057,N_19712);
xor U23938 (N_23938,N_19159,N_18635);
nand U23939 (N_23939,N_20282,N_20469);
and U23940 (N_23940,N_18243,N_19695);
nand U23941 (N_23941,N_20136,N_18090);
xnor U23942 (N_23942,N_20751,N_18651);
xnor U23943 (N_23943,N_18534,N_20576);
and U23944 (N_23944,N_19845,N_20815);
nor U23945 (N_23945,N_20811,N_18624);
xor U23946 (N_23946,N_20597,N_18242);
xnor U23947 (N_23947,N_20100,N_18458);
nor U23948 (N_23948,N_19443,N_18744);
nand U23949 (N_23949,N_18237,N_19163);
xor U23950 (N_23950,N_19792,N_18358);
nand U23951 (N_23951,N_18748,N_18256);
xor U23952 (N_23952,N_20967,N_20884);
or U23953 (N_23953,N_20467,N_18969);
nor U23954 (N_23954,N_20125,N_18487);
xor U23955 (N_23955,N_18068,N_19293);
or U23956 (N_23956,N_19203,N_20267);
and U23957 (N_23957,N_20636,N_18045);
nor U23958 (N_23958,N_19525,N_19455);
xor U23959 (N_23959,N_19696,N_20225);
xor U23960 (N_23960,N_20263,N_19412);
nor U23961 (N_23961,N_20317,N_19112);
xnor U23962 (N_23962,N_19578,N_20525);
nor U23963 (N_23963,N_19538,N_20241);
nor U23964 (N_23964,N_20712,N_20241);
xor U23965 (N_23965,N_19349,N_19386);
or U23966 (N_23966,N_19312,N_19400);
nor U23967 (N_23967,N_19443,N_20911);
xnor U23968 (N_23968,N_20924,N_18228);
nand U23969 (N_23969,N_19408,N_18621);
nand U23970 (N_23970,N_18350,N_18820);
xnor U23971 (N_23971,N_19535,N_20437);
and U23972 (N_23972,N_19469,N_18955);
and U23973 (N_23973,N_19605,N_19879);
nand U23974 (N_23974,N_19473,N_19395);
nor U23975 (N_23975,N_18793,N_20958);
xnor U23976 (N_23976,N_18552,N_19655);
or U23977 (N_23977,N_18601,N_18847);
nor U23978 (N_23978,N_18760,N_18482);
nor U23979 (N_23979,N_18865,N_20616);
or U23980 (N_23980,N_19799,N_18105);
xnor U23981 (N_23981,N_20826,N_18878);
nor U23982 (N_23982,N_19981,N_20681);
xor U23983 (N_23983,N_19200,N_20259);
or U23984 (N_23984,N_19664,N_18385);
and U23985 (N_23985,N_20197,N_20914);
xnor U23986 (N_23986,N_20451,N_19403);
and U23987 (N_23987,N_20890,N_20041);
and U23988 (N_23988,N_20980,N_19018);
or U23989 (N_23989,N_20787,N_18316);
nor U23990 (N_23990,N_19448,N_19829);
and U23991 (N_23991,N_20512,N_20592);
xor U23992 (N_23992,N_19866,N_20156);
xor U23993 (N_23993,N_19789,N_18192);
xnor U23994 (N_23994,N_18890,N_19870);
nor U23995 (N_23995,N_18509,N_20125);
or U23996 (N_23996,N_19962,N_20076);
nand U23997 (N_23997,N_19653,N_20419);
xnor U23998 (N_23998,N_18824,N_20489);
nand U23999 (N_23999,N_20557,N_20449);
and U24000 (N_24000,N_23239,N_23474);
and U24001 (N_24001,N_21618,N_23089);
nor U24002 (N_24002,N_23749,N_22248);
nor U24003 (N_24003,N_23381,N_21730);
and U24004 (N_24004,N_21766,N_22015);
xnor U24005 (N_24005,N_23445,N_23931);
nor U24006 (N_24006,N_22932,N_23506);
and U24007 (N_24007,N_23794,N_21733);
or U24008 (N_24008,N_21617,N_21068);
xnor U24009 (N_24009,N_23156,N_21380);
nor U24010 (N_24010,N_23920,N_22483);
or U24011 (N_24011,N_23592,N_23700);
nor U24012 (N_24012,N_23973,N_21467);
or U24013 (N_24013,N_22620,N_22340);
and U24014 (N_24014,N_22025,N_23878);
or U24015 (N_24015,N_23012,N_23085);
nand U24016 (N_24016,N_22679,N_21584);
nand U24017 (N_24017,N_22956,N_21119);
xnor U24018 (N_24018,N_21966,N_22584);
and U24019 (N_24019,N_23831,N_21571);
nor U24020 (N_24020,N_23060,N_22721);
nor U24021 (N_24021,N_22580,N_22537);
or U24022 (N_24022,N_21491,N_21953);
xnor U24023 (N_24023,N_22136,N_21125);
xnor U24024 (N_24024,N_21296,N_22446);
nand U24025 (N_24025,N_22061,N_21531);
nor U24026 (N_24026,N_22065,N_22767);
xor U24027 (N_24027,N_23779,N_21422);
nor U24028 (N_24028,N_23793,N_21155);
and U24029 (N_24029,N_23271,N_21278);
nand U24030 (N_24030,N_22885,N_23660);
and U24031 (N_24031,N_22883,N_23879);
xnor U24032 (N_24032,N_22631,N_22191);
nand U24033 (N_24033,N_22059,N_22066);
or U24034 (N_24034,N_22038,N_21759);
xnor U24035 (N_24035,N_23816,N_21483);
and U24036 (N_24036,N_23753,N_21671);
and U24037 (N_24037,N_23694,N_22083);
nor U24038 (N_24038,N_22396,N_23166);
or U24039 (N_24039,N_22952,N_23511);
nand U24040 (N_24040,N_22492,N_21195);
xnor U24041 (N_24041,N_23040,N_21569);
or U24042 (N_24042,N_21056,N_21394);
nor U24043 (N_24043,N_23030,N_21309);
xnor U24044 (N_24044,N_22391,N_22953);
and U24045 (N_24045,N_23332,N_22471);
xnor U24046 (N_24046,N_23740,N_23270);
nor U24047 (N_24047,N_23672,N_22555);
xnor U24048 (N_24048,N_21346,N_23007);
and U24049 (N_24049,N_21530,N_22408);
xnor U24050 (N_24050,N_21037,N_23801);
nor U24051 (N_24051,N_22087,N_23917);
nor U24052 (N_24052,N_22001,N_23080);
or U24053 (N_24053,N_22440,N_22825);
nand U24054 (N_24054,N_22378,N_22007);
nor U24055 (N_24055,N_23743,N_23401);
xnor U24056 (N_24056,N_22520,N_21273);
nor U24057 (N_24057,N_23028,N_21414);
nor U24058 (N_24058,N_21619,N_22652);
nor U24059 (N_24059,N_21986,N_21393);
nand U24060 (N_24060,N_21222,N_21644);
nand U24061 (N_24061,N_23574,N_22216);
and U24062 (N_24062,N_22417,N_22052);
and U24063 (N_24063,N_21927,N_21866);
or U24064 (N_24064,N_22290,N_23902);
or U24065 (N_24065,N_21062,N_21433);
nand U24066 (N_24066,N_23258,N_23663);
nand U24067 (N_24067,N_23320,N_21035);
or U24068 (N_24068,N_21783,N_21769);
and U24069 (N_24069,N_21698,N_21197);
xnor U24070 (N_24070,N_21973,N_23841);
nand U24071 (N_24071,N_21622,N_23476);
xnor U24072 (N_24072,N_23921,N_23314);
and U24073 (N_24073,N_23183,N_23471);
xor U24074 (N_24074,N_21358,N_23918);
nand U24075 (N_24075,N_23750,N_23875);
xor U24076 (N_24076,N_22343,N_21282);
or U24077 (N_24077,N_23513,N_21313);
xor U24078 (N_24078,N_21824,N_22569);
or U24079 (N_24079,N_21209,N_21428);
nand U24080 (N_24080,N_22182,N_23050);
and U24081 (N_24081,N_21067,N_21147);
nor U24082 (N_24082,N_22462,N_23687);
nand U24083 (N_24083,N_23770,N_21213);
and U24084 (N_24084,N_23064,N_22848);
nor U24085 (N_24085,N_22456,N_22135);
xor U24086 (N_24086,N_22188,N_21122);
nor U24087 (N_24087,N_22639,N_23436);
and U24088 (N_24088,N_21364,N_23566);
or U24089 (N_24089,N_22246,N_21972);
or U24090 (N_24090,N_21838,N_22820);
or U24091 (N_24091,N_23097,N_21228);
nor U24092 (N_24092,N_22838,N_21573);
nand U24093 (N_24093,N_21280,N_22484);
or U24094 (N_24094,N_21686,N_22322);
or U24095 (N_24095,N_23551,N_23049);
nor U24096 (N_24096,N_22525,N_22163);
xor U24097 (N_24097,N_22844,N_23380);
xnor U24098 (N_24098,N_23107,N_21439);
or U24099 (N_24099,N_22549,N_22733);
nand U24100 (N_24100,N_23848,N_21755);
and U24101 (N_24101,N_23108,N_23941);
or U24102 (N_24102,N_23654,N_21184);
nand U24103 (N_24103,N_23544,N_21896);
or U24104 (N_24104,N_21154,N_21418);
xnor U24105 (N_24105,N_23983,N_23250);
and U24106 (N_24106,N_22117,N_22628);
or U24107 (N_24107,N_23447,N_23702);
nand U24108 (N_24108,N_21860,N_21731);
xnor U24109 (N_24109,N_23294,N_21781);
nand U24110 (N_24110,N_21989,N_22150);
or U24111 (N_24111,N_21263,N_22638);
and U24112 (N_24112,N_21203,N_21407);
and U24113 (N_24113,N_21268,N_22308);
and U24114 (N_24114,N_23913,N_22816);
nor U24115 (N_24115,N_21795,N_22164);
nand U24116 (N_24116,N_21236,N_21353);
and U24117 (N_24117,N_21942,N_21093);
and U24118 (N_24118,N_23709,N_23888);
nand U24119 (N_24119,N_23730,N_23429);
or U24120 (N_24120,N_22148,N_21980);
or U24121 (N_24121,N_23845,N_21659);
nor U24122 (N_24122,N_22239,N_22020);
nand U24123 (N_24123,N_21210,N_23729);
nand U24124 (N_24124,N_21158,N_22637);
or U24125 (N_24125,N_22728,N_21266);
nand U24126 (N_24126,N_22681,N_21620);
or U24127 (N_24127,N_21481,N_22241);
and U24128 (N_24128,N_23688,N_22818);
xnor U24129 (N_24129,N_21120,N_23982);
or U24130 (N_24130,N_21903,N_21429);
nand U24131 (N_24131,N_23019,N_21537);
xnor U24132 (N_24132,N_21649,N_22546);
and U24133 (N_24133,N_23876,N_23970);
or U24134 (N_24134,N_22923,N_21397);
or U24135 (N_24135,N_21754,N_22261);
nand U24136 (N_24136,N_22771,N_21566);
nand U24137 (N_24137,N_23833,N_23126);
xor U24138 (N_24138,N_22186,N_21727);
nor U24139 (N_24139,N_23175,N_21760);
and U24140 (N_24140,N_21319,N_22237);
nor U24141 (N_24141,N_22084,N_23919);
or U24142 (N_24142,N_23176,N_22309);
xor U24143 (N_24143,N_22807,N_23338);
xor U24144 (N_24144,N_23031,N_21128);
or U24145 (N_24145,N_22264,N_21441);
and U24146 (N_24146,N_22934,N_21322);
and U24147 (N_24147,N_23500,N_21987);
xor U24148 (N_24148,N_21066,N_22330);
xor U24149 (N_24149,N_21423,N_22392);
and U24150 (N_24150,N_23524,N_21777);
xor U24151 (N_24151,N_21857,N_22685);
and U24152 (N_24152,N_23584,N_22030);
or U24153 (N_24153,N_21765,N_23554);
xor U24154 (N_24154,N_22247,N_23881);
xnor U24155 (N_24155,N_22125,N_23890);
xor U24156 (N_24156,N_21575,N_23384);
xnor U24157 (N_24157,N_23006,N_21579);
and U24158 (N_24158,N_23449,N_22979);
xnor U24159 (N_24159,N_22010,N_21974);
xnor U24160 (N_24160,N_21142,N_23291);
xor U24161 (N_24161,N_23549,N_23783);
and U24162 (N_24162,N_21356,N_21956);
and U24163 (N_24163,N_21161,N_21643);
or U24164 (N_24164,N_23480,N_21609);
xor U24165 (N_24165,N_21241,N_23960);
and U24166 (N_24166,N_21572,N_22610);
or U24167 (N_24167,N_22947,N_23163);
or U24168 (N_24168,N_21073,N_21314);
or U24169 (N_24169,N_22332,N_23964);
or U24170 (N_24170,N_21847,N_22977);
nand U24171 (N_24171,N_21390,N_21621);
xnor U24172 (N_24172,N_21288,N_21029);
or U24173 (N_24173,N_21615,N_23977);
or U24174 (N_24174,N_21301,N_22529);
xnor U24175 (N_24175,N_23093,N_22612);
xor U24176 (N_24176,N_22832,N_21072);
nand U24177 (N_24177,N_21498,N_22600);
or U24178 (N_24178,N_23842,N_23355);
and U24179 (N_24179,N_21524,N_23228);
nor U24180 (N_24180,N_21200,N_21432);
nor U24181 (N_24181,N_22578,N_21976);
xnor U24182 (N_24182,N_22731,N_22647);
nand U24183 (N_24183,N_22381,N_21528);
nor U24184 (N_24184,N_21094,N_21276);
xor U24185 (N_24185,N_21614,N_21822);
xor U24186 (N_24186,N_23000,N_21851);
nand U24187 (N_24187,N_22716,N_22924);
nand U24188 (N_24188,N_21768,N_23665);
and U24189 (N_24189,N_23400,N_22335);
xnor U24190 (N_24190,N_22418,N_22416);
or U24191 (N_24191,N_22075,N_22984);
xor U24192 (N_24192,N_22657,N_22626);
or U24193 (N_24193,N_22576,N_23335);
or U24194 (N_24194,N_21641,N_22533);
nor U24195 (N_24195,N_23909,N_21410);
xnor U24196 (N_24196,N_22234,N_23391);
nor U24197 (N_24197,N_23748,N_21102);
and U24198 (N_24198,N_21036,N_23951);
nor U24199 (N_24199,N_21373,N_22277);
or U24200 (N_24200,N_23209,N_21914);
nor U24201 (N_24201,N_21415,N_22640);
nor U24202 (N_24202,N_21654,N_23819);
and U24203 (N_24203,N_23398,N_23304);
xor U24204 (N_24204,N_21291,N_22495);
xor U24205 (N_24205,N_23299,N_21427);
or U24206 (N_24206,N_22227,N_21389);
or U24207 (N_24207,N_21352,N_23432);
xnor U24208 (N_24208,N_21819,N_21137);
nand U24209 (N_24209,N_21006,N_21647);
nand U24210 (N_24210,N_23378,N_23178);
or U24211 (N_24211,N_21515,N_21944);
or U24212 (N_24212,N_21834,N_22215);
and U24213 (N_24213,N_22317,N_23425);
xnor U24214 (N_24214,N_21694,N_22031);
xnor U24215 (N_24215,N_22134,N_23020);
and U24216 (N_24216,N_22169,N_23457);
nor U24217 (N_24217,N_21461,N_21799);
and U24218 (N_24218,N_22987,N_22882);
nand U24219 (N_24219,N_23438,N_23356);
nor U24220 (N_24220,N_21687,N_23565);
nand U24221 (N_24221,N_21153,N_21206);
nand U24222 (N_24222,N_21794,N_23884);
or U24223 (N_24223,N_22302,N_23148);
and U24224 (N_24224,N_23764,N_23962);
and U24225 (N_24225,N_22372,N_21843);
or U24226 (N_24226,N_23388,N_23995);
and U24227 (N_24227,N_23972,N_21488);
nand U24228 (N_24228,N_23238,N_23305);
xor U24229 (N_24229,N_21684,N_23567);
xnor U24230 (N_24230,N_21541,N_22780);
xor U24231 (N_24231,N_21561,N_23319);
and U24232 (N_24232,N_21505,N_22558);
xor U24233 (N_24233,N_21281,N_21400);
xor U24234 (N_24234,N_21696,N_23346);
or U24235 (N_24235,N_23063,N_21413);
or U24236 (N_24236,N_22242,N_23069);
nor U24237 (N_24237,N_23518,N_21150);
nor U24238 (N_24238,N_21261,N_23039);
and U24239 (N_24239,N_22331,N_21229);
nor U24240 (N_24240,N_21013,N_23184);
and U24241 (N_24241,N_21040,N_23755);
nand U24242 (N_24242,N_22713,N_21875);
nor U24243 (N_24243,N_22588,N_22403);
xnor U24244 (N_24244,N_21743,N_22073);
nor U24245 (N_24245,N_23514,N_23187);
or U24246 (N_24246,N_23976,N_23067);
nor U24247 (N_24247,N_23916,N_23542);
nand U24248 (N_24248,N_21402,N_21111);
xnor U24249 (N_24249,N_22861,N_22981);
and U24250 (N_24250,N_23475,N_22579);
and U24251 (N_24251,N_22535,N_22173);
xnor U24252 (N_24252,N_23276,N_22909);
nand U24253 (N_24253,N_23034,N_22893);
or U24254 (N_24254,N_23177,N_22154);
and U24255 (N_24255,N_23010,N_23303);
or U24256 (N_24256,N_23552,N_23985);
and U24257 (N_24257,N_23136,N_23501);
xor U24258 (N_24258,N_23227,N_21806);
xor U24259 (N_24259,N_21988,N_21695);
nor U24260 (N_24260,N_22303,N_23837);
or U24261 (N_24261,N_23217,N_21836);
nor U24262 (N_24262,N_21562,N_22508);
or U24263 (N_24263,N_21658,N_23782);
nand U24264 (N_24264,N_22056,N_21164);
xor U24265 (N_24265,N_21969,N_22395);
xor U24266 (N_24266,N_23285,N_23081);
nor U24267 (N_24267,N_22361,N_23975);
and U24268 (N_24268,N_21193,N_23105);
or U24269 (N_24269,N_21300,N_23329);
nor U24270 (N_24270,N_23257,N_21014);
xor U24271 (N_24271,N_23132,N_22130);
xor U24272 (N_24272,N_22864,N_22744);
and U24273 (N_24273,N_23944,N_23843);
nor U24274 (N_24274,N_23706,N_23710);
xnor U24275 (N_24275,N_22643,N_22801);
or U24276 (N_24276,N_21770,N_23769);
and U24277 (N_24277,N_21420,N_23111);
or U24278 (N_24278,N_21060,N_23626);
nand U24279 (N_24279,N_23364,N_21199);
xnor U24280 (N_24280,N_21487,N_23751);
xor U24281 (N_24281,N_22565,N_22550);
nand U24282 (N_24282,N_21085,N_23268);
nor U24283 (N_24283,N_23150,N_22960);
nor U24284 (N_24284,N_23773,N_21290);
nand U24285 (N_24285,N_21601,N_21605);
xnor U24286 (N_24286,N_21345,N_21775);
xor U24287 (N_24287,N_21113,N_23617);
and U24288 (N_24288,N_22834,N_23033);
nor U24289 (N_24289,N_23104,N_22407);
nand U24290 (N_24290,N_22747,N_22954);
xnor U24291 (N_24291,N_23117,N_21588);
and U24292 (N_24292,N_23420,N_22473);
xnor U24293 (N_24293,N_22009,N_23677);
xor U24294 (N_24294,N_23165,N_22021);
and U24295 (N_24295,N_23042,N_22464);
nor U24296 (N_24296,N_21275,N_22739);
nor U24297 (N_24297,N_23403,N_22951);
xnor U24298 (N_24298,N_22853,N_21679);
nor U24299 (N_24299,N_21283,N_22470);
nor U24300 (N_24300,N_23267,N_21791);
xnor U24301 (N_24301,N_23247,N_22273);
and U24302 (N_24302,N_23812,N_21240);
nor U24303 (N_24303,N_22051,N_21526);
xnor U24304 (N_24304,N_23191,N_23351);
nor U24305 (N_24305,N_23823,N_22602);
xnor U24306 (N_24306,N_22755,N_23077);
nand U24307 (N_24307,N_21489,N_23171);
nor U24308 (N_24308,N_23405,N_22054);
and U24309 (N_24309,N_23018,N_23813);
and U24310 (N_24310,N_21919,N_23765);
or U24311 (N_24311,N_21933,N_22976);
nor U24312 (N_24312,N_22341,N_22459);
nand U24313 (N_24313,N_21964,N_22506);
nand U24314 (N_24314,N_22476,N_22064);
nand U24315 (N_24315,N_21326,N_21003);
nand U24316 (N_24316,N_22140,N_22870);
or U24317 (N_24317,N_23715,N_23164);
and U24318 (N_24318,N_21907,N_22692);
nand U24319 (N_24319,N_23681,N_22315);
and U24320 (N_24320,N_22365,N_21059);
nand U24321 (N_24321,N_22185,N_23644);
or U24322 (N_24322,N_21205,N_21374);
nor U24323 (N_24323,N_23468,N_22327);
nand U24324 (N_24324,N_22488,N_22604);
nand U24325 (N_24325,N_22594,N_21846);
nand U24326 (N_24326,N_23327,N_21913);
nor U24327 (N_24327,N_21930,N_23367);
and U24328 (N_24328,N_23607,N_23942);
and U24329 (N_24329,N_22841,N_23869);
nor U24330 (N_24330,N_23490,N_23434);
or U24331 (N_24331,N_23334,N_21272);
or U24332 (N_24332,N_23179,N_23302);
nand U24333 (N_24333,N_23517,N_23828);
and U24334 (N_24334,N_22259,N_22999);
xor U24335 (N_24335,N_23221,N_22386);
xnor U24336 (N_24336,N_23809,N_23900);
xor U24337 (N_24337,N_22485,N_22195);
or U24338 (N_24338,N_23426,N_22437);
nand U24339 (N_24339,N_22285,N_21547);
and U24340 (N_24340,N_21086,N_23545);
or U24341 (N_24341,N_22338,N_22852);
xnor U24342 (N_24342,N_22521,N_22581);
or U24343 (N_24343,N_22530,N_22220);
and U24344 (N_24344,N_23726,N_23846);
nor U24345 (N_24345,N_22654,N_23281);
nor U24346 (N_24346,N_23674,N_22913);
nand U24347 (N_24347,N_21665,N_21431);
xnor U24348 (N_24348,N_23989,N_23284);
and U24349 (N_24349,N_22635,N_23993);
xor U24350 (N_24350,N_22914,N_23760);
or U24351 (N_24351,N_23009,N_22701);
xor U24352 (N_24352,N_23157,N_23331);
or U24353 (N_24353,N_22063,N_23456);
nor U24354 (N_24354,N_21472,N_23313);
nand U24355 (N_24355,N_21990,N_22192);
xor U24356 (N_24356,N_23882,N_22198);
xor U24357 (N_24357,N_22871,N_23639);
nand U24358 (N_24358,N_22687,N_22175);
xor U24359 (N_24359,N_23661,N_23008);
nor U24360 (N_24360,N_21417,N_22348);
xnor U24361 (N_24361,N_22014,N_23635);
xor U24362 (N_24362,N_23253,N_21954);
nor U24363 (N_24363,N_23454,N_21295);
xor U24364 (N_24364,N_23317,N_23041);
nand U24365 (N_24365,N_21103,N_21922);
nor U24366 (N_24366,N_23658,N_22828);
or U24367 (N_24367,N_22354,N_21868);
nand U24368 (N_24368,N_23874,N_21920);
or U24369 (N_24369,N_22907,N_22350);
nor U24370 (N_24370,N_22548,N_22080);
nor U24371 (N_24371,N_22457,N_23907);
xnor U24372 (N_24372,N_21604,N_21757);
nand U24373 (N_24373,N_23261,N_22132);
xnor U24374 (N_24374,N_23120,N_22724);
or U24375 (N_24375,N_21329,N_23826);
nand U24376 (N_24376,N_23996,N_22468);
and U24377 (N_24377,N_22334,N_23458);
nand U24378 (N_24378,N_21403,N_21943);
or U24379 (N_24379,N_21902,N_23596);
or U24380 (N_24380,N_21870,N_23151);
nor U24381 (N_24381,N_21311,N_21705);
nor U24382 (N_24382,N_21112,N_21823);
and U24383 (N_24383,N_23725,N_21877);
xor U24384 (N_24384,N_22709,N_21411);
or U24385 (N_24385,N_22910,N_21438);
and U24386 (N_24386,N_23172,N_22930);
xor U24387 (N_24387,N_21267,N_21138);
nor U24388 (N_24388,N_21551,N_22887);
or U24389 (N_24389,N_22719,N_21312);
xor U24390 (N_24390,N_21269,N_22958);
xor U24391 (N_24391,N_22899,N_22275);
or U24392 (N_24392,N_21697,N_22680);
or U24393 (N_24393,N_23642,N_23885);
or U24394 (N_24394,N_23312,N_21510);
and U24395 (N_24395,N_23222,N_21758);
or U24396 (N_24396,N_23370,N_22974);
or U24397 (N_24397,N_21636,N_21091);
and U24398 (N_24398,N_22925,N_22139);
nor U24399 (N_24399,N_23419,N_22197);
nand U24400 (N_24400,N_23807,N_22211);
xor U24401 (N_24401,N_22077,N_21859);
or U24402 (N_24402,N_23195,N_21170);
xnor U24403 (N_24403,N_21054,N_22036);
nor U24404 (N_24404,N_23264,N_23371);
xor U24405 (N_24405,N_22219,N_21849);
and U24406 (N_24406,N_21114,N_21508);
xnor U24407 (N_24407,N_23047,N_21817);
nor U24408 (N_24408,N_22193,N_23959);
nor U24409 (N_24409,N_23116,N_22055);
xor U24410 (N_24410,N_23418,N_21316);
or U24411 (N_24411,N_23437,N_22337);
and U24412 (N_24412,N_21208,N_21832);
xnor U24413 (N_24413,N_22617,N_21886);
xnor U24414 (N_24414,N_23360,N_22146);
nor U24415 (N_24415,N_21334,N_21305);
or U24416 (N_24416,N_21594,N_21790);
or U24417 (N_24417,N_21858,N_23125);
or U24418 (N_24418,N_22901,N_23590);
nor U24419 (N_24419,N_21589,N_23659);
nand U24420 (N_24420,N_23657,N_21030);
nor U24421 (N_24421,N_22847,N_21399);
xnor U24422 (N_24422,N_21536,N_23936);
xor U24423 (N_24423,N_23924,N_21243);
nor U24424 (N_24424,N_23739,N_23113);
and U24425 (N_24425,N_21516,N_21406);
and U24426 (N_24426,N_22815,N_22518);
xnor U24427 (N_24427,N_21786,N_23787);
or U24428 (N_24428,N_22690,N_22043);
xnor U24429 (N_24429,N_22592,N_21645);
xor U24430 (N_24430,N_22102,N_22982);
xnor U24431 (N_24431,N_23272,N_21204);
nor U24432 (N_24432,N_22557,N_21140);
or U24433 (N_24433,N_23485,N_21404);
or U24434 (N_24434,N_21661,N_23851);
or U24435 (N_24435,N_21610,N_23987);
or U24436 (N_24436,N_23498,N_23638);
nand U24437 (N_24437,N_23208,N_21051);
xor U24438 (N_24438,N_23090,N_22991);
xnor U24439 (N_24439,N_23522,N_21355);
or U24440 (N_24440,N_21017,N_21083);
nand U24441 (N_24441,N_21978,N_21055);
and U24442 (N_24442,N_21405,N_22900);
nor U24443 (N_24443,N_22651,N_22113);
and U24444 (N_24444,N_23350,N_23139);
and U24445 (N_24445,N_21912,N_23204);
nand U24446 (N_24446,N_21734,N_21706);
and U24447 (N_24447,N_21495,N_22212);
xnor U24448 (N_24448,N_21738,N_22310);
nor U24449 (N_24449,N_22614,N_21975);
or U24450 (N_24450,N_23375,N_21118);
nand U24451 (N_24451,N_21141,N_23298);
nand U24452 (N_24452,N_23559,N_23493);
and U24453 (N_24453,N_21928,N_22624);
or U24454 (N_24454,N_21879,N_22249);
nand U24455 (N_24455,N_23992,N_21446);
or U24456 (N_24456,N_22319,N_22101);
xnor U24457 (N_24457,N_22346,N_23032);
and U24458 (N_24458,N_22256,N_23424);
nor U24459 (N_24459,N_23492,N_23859);
nand U24460 (N_24460,N_23341,N_21473);
or U24461 (N_24461,N_21340,N_22812);
nor U24462 (N_24462,N_23969,N_22857);
nor U24463 (N_24463,N_22429,N_22971);
or U24464 (N_24464,N_22489,N_21180);
or U24465 (N_24465,N_21704,N_23621);
nand U24466 (N_24466,N_22998,N_21683);
nor U24467 (N_24467,N_23101,N_21865);
and U24468 (N_24468,N_21915,N_23766);
and U24469 (N_24469,N_23800,N_21342);
nor U24470 (N_24470,N_22082,N_21265);
nand U24471 (N_24471,N_21678,N_22298);
nor U24472 (N_24472,N_22668,N_21260);
nor U24473 (N_24473,N_22004,N_21436);
nand U24474 (N_24474,N_21437,N_23218);
nand U24475 (N_24475,N_23581,N_23609);
nor U24476 (N_24476,N_21509,N_23744);
xnor U24477 (N_24477,N_22544,N_21646);
and U24478 (N_24478,N_23553,N_23442);
xnor U24479 (N_24479,N_22000,N_21507);
or U24480 (N_24480,N_22622,N_21653);
and U24481 (N_24481,N_23786,N_22441);
xor U24482 (N_24482,N_23877,N_21189);
or U24483 (N_24483,N_21298,N_22448);
or U24484 (N_24484,N_22722,N_23408);
nor U24485 (N_24485,N_22194,N_22854);
xnor U24486 (N_24486,N_23134,N_23308);
xor U24487 (N_24487,N_23200,N_21629);
nand U24488 (N_24488,N_22574,N_23255);
and U24489 (N_24489,N_21761,N_22609);
or U24490 (N_24490,N_22636,N_23452);
nand U24491 (N_24491,N_22693,N_22387);
or U24492 (N_24492,N_23713,N_21151);
nor U24493 (N_24493,N_22860,N_21689);
or U24494 (N_24494,N_22968,N_22008);
nand U24495 (N_24495,N_22349,N_23578);
xnor U24496 (N_24496,N_23194,N_23225);
and U24497 (N_24497,N_21221,N_21165);
nand U24498 (N_24498,N_21104,N_22472);
nor U24499 (N_24499,N_21248,N_21670);
or U24500 (N_24500,N_23712,N_21174);
or U24501 (N_24501,N_22865,N_22412);
nor U24502 (N_24502,N_21101,N_23955);
xor U24503 (N_24503,N_23667,N_23512);
xnor U24504 (N_24504,N_23507,N_21993);
xnor U24505 (N_24505,N_21941,N_21350);
or U24506 (N_24506,N_22933,N_22297);
nand U24507 (N_24507,N_22058,N_22218);
nand U24508 (N_24508,N_21294,N_22336);
nor U24509 (N_24509,N_21945,N_23404);
nand U24510 (N_24510,N_22867,N_21957);
nor U24511 (N_24511,N_22603,N_22373);
nor U24512 (N_24512,N_22201,N_21835);
or U24513 (N_24513,N_22515,N_22567);
or U24514 (N_24514,N_21307,N_21490);
nand U24515 (N_24515,N_23051,N_21700);
xnor U24516 (N_24516,N_21826,N_22823);
xor U24517 (N_24517,N_22627,N_22955);
xor U24518 (N_24518,N_22137,N_23190);
xnor U24519 (N_24519,N_23618,N_21845);
nand U24520 (N_24520,N_21231,N_22598);
nor U24521 (N_24521,N_23275,N_21134);
and U24522 (N_24522,N_23645,N_23417);
or U24523 (N_24523,N_21655,N_23774);
xnor U24524 (N_24524,N_22366,N_22527);
and U24525 (N_24525,N_23597,N_21286);
and U24526 (N_24526,N_21445,N_23718);
nand U24527 (N_24527,N_21233,N_22005);
xor U24528 (N_24528,N_21211,N_22666);
nor U24529 (N_24529,N_21027,N_23167);
or U24530 (N_24530,N_21194,N_23229);
or U24531 (N_24531,N_23986,N_22491);
and U24532 (N_24532,N_23593,N_22754);
or U24533 (N_24533,N_21871,N_21494);
xnor U24534 (N_24534,N_23246,N_23397);
nor U24535 (N_24535,N_23004,N_22452);
and U24536 (N_24536,N_22099,N_22496);
xnor U24537 (N_24537,N_21459,N_23614);
and U24538 (N_24538,N_21225,N_21590);
nor U24539 (N_24539,N_21063,N_23315);
nand U24540 (N_24540,N_21057,N_21812);
xnor U24541 (N_24541,N_22450,N_21201);
nor U24542 (N_24542,N_22255,N_22179);
nor U24543 (N_24543,N_23555,N_23016);
or U24544 (N_24544,N_21815,N_22370);
nor U24545 (N_24545,N_23415,N_22881);
or U24546 (N_24546,N_22545,N_23894);
and U24547 (N_24547,N_23109,N_21880);
and U24548 (N_24548,N_21793,N_21631);
or U24549 (N_24549,N_21224,N_22589);
nor U24550 (N_24550,N_23855,N_23230);
and U24551 (N_24551,N_23811,N_21821);
or U24552 (N_24552,N_23905,N_22874);
xor U24553 (N_24553,N_21457,N_22029);
xnor U24554 (N_24554,N_21009,N_23248);
and U24555 (N_24555,N_22068,N_21131);
nor U24556 (N_24556,N_21460,N_21492);
and U24557 (N_24557,N_22026,N_21578);
nand U24558 (N_24558,N_21369,N_21699);
nor U24559 (N_24559,N_22199,N_21752);
nand U24560 (N_24560,N_22725,N_22451);
or U24561 (N_24561,N_23159,N_22328);
or U24562 (N_24562,N_22100,N_21568);
xor U24563 (N_24563,N_23057,N_22689);
and U24564 (N_24564,N_23576,N_22460);
and U24565 (N_24565,N_23336,N_23464);
xor U24566 (N_24566,N_23824,N_22851);
nand U24567 (N_24567,N_23469,N_23154);
xnor U24568 (N_24568,N_22552,N_22189);
or U24569 (N_24569,N_22463,N_22568);
or U24570 (N_24570,N_21585,N_21324);
nand U24571 (N_24571,N_23279,N_23205);
and U24572 (N_24572,N_22333,N_23427);
xor U24573 (N_24573,N_22809,N_21577);
and U24574 (N_24574,N_21279,N_21099);
xnor U24575 (N_24575,N_23112,N_22203);
xnor U24576 (N_24576,N_22313,N_21999);
xnor U24577 (N_24577,N_21015,N_22512);
and U24578 (N_24578,N_22884,N_23974);
nor U24579 (N_24579,N_21202,N_21008);
nand U24580 (N_24580,N_21226,N_23673);
nor U24581 (N_24581,N_21303,N_23956);
xor U24582 (N_24582,N_23022,N_23630);
and U24583 (N_24583,N_21716,N_21183);
nand U24584 (N_24584,N_22575,N_23860);
or U24585 (N_24585,N_23605,N_21833);
and U24586 (N_24586,N_23412,N_22511);
and U24587 (N_24587,N_22547,N_22153);
xor U24588 (N_24588,N_22705,N_22128);
and U24589 (N_24589,N_23762,N_21385);
and U24590 (N_24590,N_22819,N_22254);
nand U24591 (N_24591,N_21045,N_21176);
nand U24592 (N_24592,N_21220,N_23092);
or U24593 (N_24593,N_23503,N_23076);
nor U24594 (N_24594,N_22691,N_23984);
or U24595 (N_24595,N_23348,N_21842);
nor U24596 (N_24596,N_22660,N_21480);
nand U24597 (N_24597,N_22714,N_21005);
nor U24598 (N_24598,N_22738,N_22013);
nand U24599 (N_24599,N_21274,N_21089);
or U24600 (N_24600,N_23088,N_21354);
nor U24601 (N_24601,N_23757,N_21289);
and U24602 (N_24602,N_22294,N_22122);
nor U24603 (N_24603,N_22969,N_21673);
xnor U24604 (N_24604,N_21246,N_21667);
or U24605 (N_24605,N_22079,N_23135);
or U24606 (N_24606,N_21556,N_21753);
nor U24607 (N_24607,N_22478,N_21116);
nor U24608 (N_24608,N_22006,N_21500);
and U24609 (N_24609,N_21809,N_22822);
xnor U24610 (N_24610,N_21232,N_22583);
and U24611 (N_24611,N_21763,N_21894);
nor U24612 (N_24612,N_23361,N_21692);
and U24613 (N_24613,N_21803,N_21567);
nand U24614 (N_24614,N_21612,N_23199);
and U24615 (N_24615,N_22172,N_21961);
nor U24616 (N_24616,N_23054,N_21503);
nand U24617 (N_24617,N_21901,N_22152);
nor U24618 (N_24618,N_23957,N_22616);
nand U24619 (N_24619,N_21592,N_21363);
nor U24620 (N_24620,N_21963,N_21656);
and U24621 (N_24621,N_22572,N_22435);
nor U24622 (N_24622,N_21827,N_22420);
xor U24623 (N_24623,N_21666,N_21357);
or U24624 (N_24624,N_21545,N_22623);
or U24625 (N_24625,N_21780,N_22625);
nand U24626 (N_24626,N_23486,N_22742);
nand U24627 (N_24627,N_21917,N_22481);
or U24628 (N_24628,N_22649,N_22746);
and U24629 (N_24629,N_21159,N_22353);
and U24630 (N_24630,N_21728,N_21650);
xor U24631 (N_24631,N_22621,N_22121);
nand U24632 (N_24632,N_23323,N_21124);
nand U24633 (N_24633,N_22352,N_21367);
xor U24634 (N_24634,N_23127,N_21882);
or U24635 (N_24635,N_21521,N_23689);
nand U24636 (N_24636,N_23558,N_22027);
nand U24637 (N_24637,N_23201,N_22382);
and U24638 (N_24638,N_21482,N_23895);
nand U24639 (N_24639,N_22564,N_22323);
and U24640 (N_24640,N_23953,N_21861);
xor U24641 (N_24641,N_23790,N_22662);
nand U24642 (N_24642,N_21466,N_22756);
or U24643 (N_24643,N_22675,N_21187);
nor U24644 (N_24644,N_22920,N_22040);
or U24645 (N_24645,N_22712,N_21292);
xnor U24646 (N_24646,N_21693,N_23763);
and U24647 (N_24647,N_23243,N_23925);
or U24648 (N_24648,N_23262,N_22735);
and U24649 (N_24649,N_23686,N_22240);
nor U24650 (N_24650,N_23695,N_23137);
nor U24651 (N_24651,N_21048,N_21740);
or U24652 (N_24652,N_23443,N_21895);
and U24653 (N_24653,N_23892,N_23802);
nand U24654 (N_24654,N_23224,N_21742);
and U24655 (N_24655,N_23792,N_21750);
nor U24656 (N_24656,N_21412,N_21598);
nor U24657 (N_24657,N_21109,N_21097);
nor U24658 (N_24658,N_22505,N_21909);
nand U24659 (N_24659,N_22965,N_22727);
and U24660 (N_24660,N_21096,N_23215);
xnor U24661 (N_24661,N_22720,N_21287);
nor U24662 (N_24662,N_23428,N_22563);
nor U24663 (N_24663,N_21991,N_21349);
and U24664 (N_24664,N_23839,N_23185);
nor U24665 (N_24665,N_23043,N_23098);
nor U24666 (N_24666,N_22551,N_23038);
nor U24667 (N_24667,N_22161,N_22376);
and U24668 (N_24668,N_22221,N_22664);
or U24669 (N_24669,N_23495,N_23799);
or U24670 (N_24670,N_23889,N_22942);
nand U24671 (N_24671,N_22608,N_22012);
and U24672 (N_24672,N_23505,N_23606);
nand U24673 (N_24673,N_23015,N_22090);
nor U24674 (N_24674,N_21302,N_22948);
or U24675 (N_24675,N_23535,N_22789);
or U24676 (N_24676,N_22019,N_22586);
nor U24677 (N_24677,N_22280,N_21370);
or U24678 (N_24678,N_23186,N_21042);
nor U24679 (N_24679,N_22972,N_23416);
or U24680 (N_24680,N_23594,N_22046);
nor U24681 (N_24681,N_22729,N_22560);
and U24682 (N_24682,N_23704,N_22748);
or U24683 (N_24683,N_21688,N_21544);
nand U24684 (N_24684,N_22650,N_22425);
nand U24685 (N_24685,N_23448,N_22827);
and U24686 (N_24686,N_22204,N_21365);
xor U24687 (N_24687,N_22119,N_23727);
nand U24688 (N_24688,N_21052,N_22562);
or U24689 (N_24689,N_23390,N_23528);
nor U24690 (N_24690,N_22776,N_21637);
nand U24691 (N_24691,N_21789,N_22224);
and U24692 (N_24692,N_23235,N_21565);
nand U24693 (N_24693,N_22347,N_22329);
xnor U24694 (N_24694,N_23130,N_21252);
or U24695 (N_24695,N_23805,N_22477);
nand U24696 (N_24696,N_22876,N_23908);
or U24697 (N_24697,N_23963,N_21597);
and U24698 (N_24698,N_22071,N_23316);
and U24699 (N_24699,N_22424,N_21476);
xnor U24700 (N_24700,N_22599,N_22743);
xor U24701 (N_24701,N_22994,N_23912);
nor U24702 (N_24702,N_21593,N_22050);
xor U24703 (N_24703,N_22345,N_23910);
or U24704 (N_24704,N_21157,N_21722);
or U24705 (N_24705,N_21764,N_22995);
and U24706 (N_24706,N_23887,N_21580);
or U24707 (N_24707,N_22111,N_21512);
xor U24708 (N_24708,N_21853,N_22683);
or U24709 (N_24709,N_23915,N_23721);
nor U24710 (N_24710,N_22710,N_22024);
or U24711 (N_24711,N_22783,N_23153);
nor U24712 (N_24712,N_21864,N_23048);
and U24713 (N_24713,N_22085,N_22653);
and U24714 (N_24714,N_21130,N_21076);
nand U24715 (N_24715,N_21315,N_22282);
nand U24716 (N_24716,N_22517,N_21082);
nand U24717 (N_24717,N_22260,N_21475);
nor U24718 (N_24718,N_22469,N_21525);
nand U24719 (N_24719,N_21477,N_23850);
nand U24720 (N_24720,N_23394,N_21371);
nor U24721 (N_24721,N_23515,N_21338);
and U24722 (N_24722,N_23252,N_21829);
xnor U24723 (N_24723,N_21343,N_23778);
and U24724 (N_24724,N_23741,N_23340);
xnor U24725 (N_24725,N_23058,N_22908);
or U24726 (N_24726,N_22272,N_22678);
xor U24727 (N_24727,N_22796,N_21923);
nor U24728 (N_24728,N_22480,N_21739);
and U24729 (N_24729,N_21026,N_21069);
and U24730 (N_24730,N_22133,N_21611);
nand U24731 (N_24731,N_22641,N_23547);
xor U24732 (N_24732,N_23005,N_21330);
and U24733 (N_24733,N_23326,N_22431);
nand U24734 (N_24734,N_23840,N_21726);
or U24735 (N_24735,N_21639,N_22921);
nor U24736 (N_24736,N_22205,N_23232);
and U24737 (N_24737,N_21651,N_23825);
or U24738 (N_24738,N_21084,N_23379);
and U24739 (N_24739,N_23685,N_23670);
nor U24740 (N_24740,N_22326,N_22226);
and U24741 (N_24741,N_22176,N_21186);
nor U24742 (N_24742,N_21391,N_23728);
and U24743 (N_24743,N_21946,N_22912);
nor U24744 (N_24744,N_23241,N_23182);
or U24745 (N_24745,N_22988,N_21285);
nand U24746 (N_24746,N_23352,N_22528);
nand U24747 (N_24747,N_23705,N_23021);
xor U24748 (N_24748,N_21899,N_23017);
or U24749 (N_24749,N_23240,N_22385);
and U24750 (N_24750,N_21458,N_23723);
or U24751 (N_24751,N_22532,N_23399);
nand U24752 (N_24752,N_22384,N_23168);
nand U24753 (N_24753,N_23465,N_22497);
or U24754 (N_24754,N_22078,N_23074);
and U24755 (N_24755,N_21929,N_21136);
or U24756 (N_24756,N_22606,N_21714);
xor U24757 (N_24757,N_22041,N_22873);
nor U24758 (N_24758,N_23871,N_22320);
or U24759 (N_24759,N_21863,N_22849);
and U24760 (N_24760,N_22962,N_22676);
xnor U24761 (N_24761,N_23772,N_22149);
xnor U24762 (N_24762,N_21075,N_21948);
nand U24763 (N_24763,N_22222,N_23598);
and U24764 (N_24764,N_22978,N_23068);
nor U24765 (N_24765,N_21191,N_21862);
or U24766 (N_24766,N_21306,N_22444);
nand U24767 (N_24767,N_23119,N_21627);
nand U24768 (N_24768,N_22915,N_23430);
or U24769 (N_24769,N_22276,N_21227);
nor U24770 (N_24770,N_21906,N_21452);
and U24771 (N_24771,N_23627,N_23402);
xor U24772 (N_24772,N_21050,N_21674);
nand U24773 (N_24773,N_23791,N_22611);
nor U24774 (N_24774,N_21634,N_23788);
xnor U24775 (N_24775,N_22829,N_22997);
xnor U24776 (N_24776,N_22039,N_22044);
and U24777 (N_24777,N_21361,N_22112);
and U24778 (N_24778,N_23579,N_23849);
nor U24779 (N_24779,N_23822,N_21984);
or U24780 (N_24780,N_23189,N_22230);
xnor U24781 (N_24781,N_23922,N_22371);
nand U24782 (N_24782,N_22793,N_21685);
xor U24783 (N_24783,N_21379,N_21751);
or U24784 (N_24784,N_21878,N_23330);
nor U24785 (N_24785,N_22267,N_23197);
nor U24786 (N_24786,N_21680,N_21630);
or U24787 (N_24787,N_23478,N_21800);
or U24788 (N_24788,N_22208,N_23754);
xor U24789 (N_24789,N_23287,N_21398);
nor U24790 (N_24790,N_23025,N_21626);
xnor U24791 (N_24791,N_23496,N_21396);
nor U24792 (N_24792,N_21762,N_21992);
xnor U24793 (N_24793,N_21771,N_21230);
nand U24794 (N_24794,N_22213,N_21852);
nand U24795 (N_24795,N_23883,N_22184);
xnor U24796 (N_24796,N_21681,N_22291);
or U24797 (N_24797,N_22531,N_21892);
nand U24798 (N_24798,N_23991,N_21178);
nor U24799 (N_24799,N_22037,N_22605);
nor U24800 (N_24800,N_22510,N_21392);
or U24801 (N_24801,N_21844,N_21599);
and U24802 (N_24802,N_22843,N_22736);
and U24803 (N_24803,N_23935,N_22973);
and U24804 (N_24804,N_23259,N_23724);
nor U24805 (N_24805,N_23453,N_22842);
nor U24806 (N_24806,N_23146,N_21304);
and U24807 (N_24807,N_23365,N_23059);
nor U24808 (N_24808,N_22493,N_23556);
xor U24809 (N_24809,N_23484,N_22118);
xor U24810 (N_24810,N_23343,N_22250);
or U24811 (N_24811,N_22906,N_21949);
xor U24812 (N_24812,N_22671,N_22045);
nor U24813 (N_24813,N_22772,N_23082);
xor U24814 (N_24814,N_23409,N_21796);
nor U24815 (N_24815,N_22351,N_23930);
xnor U24816 (N_24816,N_23707,N_23266);
and U24817 (N_24817,N_21339,N_22634);
or U24818 (N_24818,N_22752,N_21994);
nand U24819 (N_24819,N_21087,N_21546);
nor U24820 (N_24820,N_21181,N_22482);
and U24821 (N_24821,N_23771,N_23344);
and U24822 (N_24822,N_23014,N_23290);
xnor U24823 (N_24823,N_22028,N_21250);
nand U24824 (N_24824,N_23893,N_22158);
nor U24825 (N_24825,N_22436,N_22305);
and U24826 (N_24826,N_23676,N_23413);
and U24827 (N_24827,N_22824,N_21004);
xnor U24828 (N_24828,N_23641,N_22929);
nor U24829 (N_24829,N_23306,N_22231);
nor U24830 (N_24830,N_22400,N_22786);
xor U24831 (N_24831,N_23188,N_21216);
nor U24832 (N_24832,N_21721,N_23926);
and U24833 (N_24833,N_22682,N_21905);
nor U24834 (N_24834,N_22804,N_23529);
nor U24835 (N_24835,N_22274,N_21368);
xnor U24836 (N_24836,N_21064,N_21317);
or U24837 (N_24837,N_21767,N_21496);
and U24838 (N_24838,N_22466,N_22062);
xnor U24839 (N_24839,N_21591,N_23011);
and U24840 (N_24840,N_22142,N_21936);
or U24841 (N_24841,N_22597,N_23832);
and U24842 (N_24842,N_21251,N_21171);
and U24843 (N_24843,N_21664,N_21020);
or U24844 (N_24844,N_21271,N_21553);
and U24845 (N_24845,N_22629,N_21244);
and U24846 (N_24846,N_23891,N_22390);
and U24847 (N_24847,N_21867,N_22229);
nor U24848 (N_24848,N_22223,N_23210);
nor U24849 (N_24849,N_23516,N_23459);
or U24850 (N_24850,N_21855,N_21960);
nand U24851 (N_24851,N_22404,N_23174);
or U24852 (N_24852,N_23541,N_22601);
and U24853 (N_24853,N_22846,N_21918);
and U24854 (N_24854,N_23533,N_23311);
or U24855 (N_24855,N_22750,N_23133);
nand U24856 (N_24856,N_22318,N_23582);
xnor U24857 (N_24857,N_22766,N_22278);
nand U24858 (N_24858,N_23671,N_23206);
or U24859 (N_24859,N_21408,N_23595);
xnor U24860 (N_24860,N_21607,N_22926);
nor U24861 (N_24861,N_22917,N_23733);
xor U24862 (N_24862,N_21935,N_22661);
nor U24863 (N_24863,N_21381,N_22281);
and U24864 (N_24864,N_21965,N_21712);
xor U24865 (N_24865,N_22526,N_21497);
xnor U24866 (N_24866,N_21148,N_22596);
nand U24867 (N_24867,N_23274,N_21773);
nand U24868 (N_24868,N_22439,N_23961);
nand U24869 (N_24869,N_21959,N_21239);
nor U24870 (N_24870,N_23103,N_23277);
nor U24871 (N_24871,N_21810,N_22143);
nand U24872 (N_24872,N_23061,N_22458);
xnor U24873 (N_24873,N_21708,N_23903);
nand U24874 (N_24874,N_21748,N_22490);
nor U24875 (N_24875,N_21628,N_21890);
xnor U24876 (N_24876,N_22673,N_22094);
xor U24877 (N_24877,N_21041,N_22426);
and U24878 (N_24878,N_22422,N_22072);
or U24879 (N_24879,N_23131,N_23446);
or U24880 (N_24880,N_23144,N_21012);
nor U24881 (N_24881,N_21831,N_23037);
or U24882 (N_24882,N_22802,N_23359);
nand U24883 (N_24883,N_22210,N_22839);
nor U24884 (N_24884,N_22430,N_22170);
nand U24885 (N_24885,N_23945,N_23629);
nor U24886 (N_24886,N_23852,N_22808);
nand U24887 (N_24887,N_23233,N_23487);
nand U24888 (N_24888,N_21126,N_23722);
xnor U24889 (N_24889,N_23604,N_22949);
nor U24890 (N_24890,N_21848,N_21022);
and U24891 (N_24891,N_21596,N_23886);
or U24892 (N_24892,N_23510,N_23697);
nand U24893 (N_24893,N_21741,N_22993);
xnor U24894 (N_24894,N_22655,N_21167);
nor U24895 (N_24895,N_22286,N_23557);
and U24896 (N_24896,N_21998,N_21359);
or U24897 (N_24897,N_23075,N_23610);
or U24898 (N_24898,N_23373,N_23588);
or U24899 (N_24899,N_22301,N_21043);
or U24900 (N_24900,N_23421,N_21900);
nor U24901 (N_24901,N_22368,N_22287);
or U24902 (N_24902,N_21442,N_22749);
and U24903 (N_24903,N_22761,N_21749);
nand U24904 (N_24904,N_23333,N_22236);
nor U24905 (N_24905,N_23599,N_22145);
or U24906 (N_24906,N_23083,N_23353);
and U24907 (N_24907,N_23296,N_23387);
and U24908 (N_24908,N_22894,N_23084);
nor U24909 (N_24909,N_22536,N_21985);
or U24910 (N_24910,N_22359,N_22937);
nand U24911 (N_24911,N_21347,N_21038);
nand U24912 (N_24912,N_22033,N_22057);
nor U24913 (N_24913,N_23742,N_21624);
nor U24914 (N_24914,N_23216,N_21143);
xor U24915 (N_24915,N_21034,N_22300);
and U24916 (N_24916,N_22659,N_23937);
and U24917 (N_24917,N_22797,N_22252);
xor U24918 (N_24918,N_23322,N_22945);
or U24919 (N_24919,N_21549,N_21426);
nand U24920 (N_24920,N_22155,N_23234);
nor U24921 (N_24921,N_22507,N_23684);
xnor U24922 (N_24922,N_23719,N_22667);
nand U24923 (N_24923,N_21435,N_21574);
xor U24924 (N_24924,N_21519,N_22103);
nor U24925 (N_24925,N_22022,N_23152);
nor U24926 (N_24926,N_23180,N_21952);
nor U24927 (N_24927,N_21440,N_22067);
or U24928 (N_24928,N_23162,N_21814);
nor U24929 (N_24929,N_23836,N_21023);
nand U24930 (N_24930,N_21033,N_23114);
or U24931 (N_24931,N_21139,N_23803);
and U24932 (N_24932,N_22792,N_22397);
nand U24933 (N_24933,N_23071,N_21107);
xnor U24934 (N_24934,N_23636,N_23777);
nand U24935 (N_24935,N_23406,N_21502);
or U24936 (N_24936,N_21669,N_21811);
and U24937 (N_24937,N_21725,N_21192);
xnor U24938 (N_24938,N_22922,N_22413);
nor U24939 (N_24939,N_21785,N_23853);
and U24940 (N_24940,N_23527,N_23282);
nor U24941 (N_24941,N_23124,N_23675);
nand U24942 (N_24942,N_21711,N_23393);
or U24943 (N_24943,N_21982,N_21293);
and U24944 (N_24944,N_21873,N_23737);
nand U24945 (N_24945,N_22878,N_21310);
and U24946 (N_24946,N_23798,N_22642);
nand U24947 (N_24947,N_22342,N_21071);
or U24948 (N_24948,N_22534,N_21682);
nand U24949 (N_24949,N_23540,N_21434);
and U24950 (N_24950,N_21135,N_23820);
nand U24951 (N_24951,N_23625,N_21632);
xor U24952 (N_24952,N_21070,N_23462);
xor U24953 (N_24953,N_22423,N_23289);
nor U24954 (N_24954,N_22777,N_21893);
and U24955 (N_24955,N_23872,N_22613);
nor U24956 (N_24956,N_22665,N_21548);
nor U24957 (N_24957,N_22959,N_22244);
nand U24958 (N_24958,N_21608,N_22758);
nor U24959 (N_24959,N_23073,N_23369);
nor U24960 (N_24960,N_23971,N_22174);
nand U24961 (N_24961,N_23519,N_23170);
or U24962 (N_24962,N_22405,N_22524);
nand U24963 (N_24963,N_21538,N_23583);
nand U24964 (N_24964,N_23278,N_23223);
nor U24965 (N_24965,N_21529,N_22554);
xnor U24966 (N_24966,N_23095,N_21797);
or U24967 (N_24967,N_21190,N_22672);
or U24968 (N_24968,N_23863,N_22092);
nor U24969 (N_24969,N_23708,N_22344);
or U24970 (N_24970,N_21940,N_22393);
nor U24971 (N_24971,N_22764,N_21464);
nand U24972 (N_24972,N_23587,N_22896);
and U24973 (N_24973,N_21552,N_23602);
or U24974 (N_24974,N_21024,N_21804);
and U24975 (N_24975,N_23470,N_22964);
and U24976 (N_24976,N_22765,N_21019);
xor U24977 (N_24977,N_21215,N_22768);
and U24978 (N_24978,N_21816,N_23571);
or U24979 (N_24979,N_22811,N_21299);
or U24980 (N_24980,N_22779,N_22076);
xor U24981 (N_24981,N_21520,N_21218);
nand U24982 (N_24982,N_21484,N_22312);
xor U24983 (N_24983,N_22919,N_23978);
nand U24984 (N_24984,N_22453,N_21539);
nand U24985 (N_24985,N_22088,N_23752);
and U24986 (N_24986,N_23488,N_21720);
or U24987 (N_24987,N_23525,N_22872);
nand U24988 (N_24988,N_21550,N_21223);
xnor U24989 (N_24989,N_23696,N_23994);
and U24990 (N_24990,N_23693,N_22543);
xnor U24991 (N_24991,N_23214,N_22577);
or U24992 (N_24992,N_23455,N_21897);
or U24993 (N_24993,N_22358,N_22916);
xor U24994 (N_24994,N_21421,N_23096);
nand U24995 (N_24995,N_22114,N_22813);
or U24996 (N_24996,N_22279,N_22810);
xor U24997 (N_24997,N_21523,N_21737);
xor U24998 (N_24998,N_23509,N_21127);
and U24999 (N_24999,N_23864,N_23662);
and U25000 (N_25000,N_23904,N_22306);
or U25001 (N_25001,N_21179,N_22985);
xnor U25002 (N_25002,N_23817,N_21779);
nand U25003 (N_25003,N_23023,N_22706);
xnor U25004 (N_25004,N_21581,N_23026);
or U25005 (N_25005,N_21662,N_23366);
nor U25006 (N_25006,N_21277,N_21264);
xnor U25007 (N_25007,N_23337,N_23062);
nor U25008 (N_25008,N_23440,N_21258);
or U25009 (N_25009,N_23212,N_22374);
nand U25010 (N_25010,N_21582,N_22938);
xor U25011 (N_25011,N_23245,N_21514);
nand U25012 (N_25012,N_22670,N_22465);
nand U25013 (N_25013,N_23680,N_22138);
and U25014 (N_25014,N_22542,N_23759);
and U25015 (N_25015,N_21801,N_22011);
or U25016 (N_25016,N_22500,N_22321);
xor U25017 (N_25017,N_23868,N_22003);
and U25018 (N_25018,N_22732,N_21778);
nand U25019 (N_25019,N_22992,N_23523);
and U25020 (N_25020,N_23543,N_23283);
nand U25021 (N_25021,N_22147,N_21450);
nand U25022 (N_25022,N_21745,N_22775);
nand U25023 (N_25023,N_23537,N_23550);
and U25024 (N_25024,N_23758,N_21032);
and U25025 (N_25025,N_21284,N_22120);
xor U25026 (N_25026,N_21335,N_21623);
xor U25027 (N_25027,N_21162,N_23539);
xor U25028 (N_25028,N_23806,N_21156);
or U25029 (N_25029,N_21557,N_22553);
nor U25030 (N_25030,N_23192,N_22570);
xor U25031 (N_25031,N_21173,N_22455);
and U25032 (N_25032,N_21947,N_21123);
or U25033 (N_25033,N_22475,N_22757);
or U25034 (N_25034,N_22905,N_21238);
and U25035 (N_25035,N_21981,N_21424);
xnor U25036 (N_25036,N_21818,N_22454);
and U25037 (N_25037,N_21616,N_21002);
or U25038 (N_25038,N_22295,N_21079);
or U25039 (N_25039,N_22266,N_23668);
xor U25040 (N_25040,N_21802,N_21163);
nand U25041 (N_25041,N_23494,N_23829);
nor U25042 (N_25042,N_21874,N_21465);
and U25043 (N_25043,N_22494,N_23745);
xor U25044 (N_25044,N_22217,N_21253);
nand U25045 (N_25045,N_21657,N_22307);
xnor U25046 (N_25046,N_21448,N_23297);
and U25047 (N_25047,N_21876,N_21106);
or U25048 (N_25048,N_22034,N_22180);
or U25049 (N_25049,N_22674,N_21470);
xnor U25050 (N_25050,N_23649,N_22950);
nor U25051 (N_25051,N_23603,N_21837);
nand U25052 (N_25052,N_21921,N_21337);
and U25053 (N_25053,N_23213,N_21595);
and U25054 (N_25054,N_23613,N_23460);
or U25055 (N_25055,N_23325,N_22394);
xnor U25056 (N_25056,N_21638,N_23767);
nand U25057 (N_25057,N_22740,N_22573);
or U25058 (N_25058,N_21506,N_23775);
xnor U25059 (N_25059,N_22519,N_21175);
nor U25060 (N_25060,N_23847,N_23967);
nand U25061 (N_25061,N_23568,N_22399);
xnor U25062 (N_25062,N_22970,N_23395);
and U25063 (N_25063,N_21217,N_22726);
xor U25064 (N_25064,N_23939,N_22048);
and U25065 (N_25065,N_21603,N_23354);
nor U25066 (N_25066,N_21145,N_23526);
nor U25067 (N_25067,N_23249,N_22109);
or U25068 (N_25068,N_22879,N_21997);
nand U25069 (N_25069,N_23928,N_22292);
or U25070 (N_25070,N_22126,N_22501);
xnor U25071 (N_25071,N_22866,N_23129);
or U25072 (N_25072,N_21044,N_23198);
and U25073 (N_25073,N_23656,N_23776);
nand U25074 (N_25074,N_21444,N_21039);
or U25075 (N_25075,N_23870,N_23647);
xnor U25076 (N_25076,N_22127,N_23202);
nor U25077 (N_25077,N_21703,N_21245);
or U25078 (N_25078,N_22774,N_21576);
or U25079 (N_25079,N_21378,N_22688);
and U25080 (N_25080,N_22289,N_22897);
and U25081 (N_25081,N_22165,N_23143);
and U25082 (N_25082,N_23086,N_22243);
nor U25083 (N_25083,N_21455,N_23530);
nand U25084 (N_25084,N_22449,N_22433);
or U25085 (N_25085,N_22324,N_22814);
or U25086 (N_25086,N_22434,N_23466);
or U25087 (N_25087,N_23784,N_22238);
or U25088 (N_25088,N_21527,N_21255);
nor U25089 (N_25089,N_23732,N_21237);
and U25090 (N_25090,N_22700,N_22363);
or U25091 (N_25091,N_22585,N_23756);
xor U25092 (N_25092,N_22684,N_22785);
and U25093 (N_25093,N_23385,N_23196);
nor U25094 (N_25094,N_22053,N_23497);
nor U25095 (N_25095,N_21558,N_22795);
or U25096 (N_25096,N_22656,N_22996);
and U25097 (N_25097,N_21188,N_22943);
nand U25098 (N_25098,N_22648,N_23138);
nor U25099 (N_25099,N_21830,N_22859);
xnor U25100 (N_25100,N_23858,N_21105);
and U25101 (N_25101,N_21891,N_21977);
or U25102 (N_25102,N_23411,N_23358);
and U25103 (N_25103,N_23747,N_23534);
xor U25104 (N_25104,N_21081,N_21416);
and U25105 (N_25105,N_22251,N_23943);
xor U25106 (N_25106,N_21049,N_23382);
nor U25107 (N_25107,N_23633,N_22707);
and U25108 (N_25108,N_23789,N_21270);
and U25109 (N_25109,N_22898,N_23003);
nor U25110 (N_25110,N_22931,N_21583);
xor U25111 (N_25111,N_23102,N_23242);
or U25112 (N_25112,N_22590,N_23431);
and U25113 (N_25113,N_22356,N_22089);
and U25114 (N_25114,N_23655,N_22990);
nor U25115 (N_25115,N_21297,N_21115);
nor U25116 (N_25116,N_21675,N_21807);
nor U25117 (N_25117,N_22903,N_22669);
xor U25118 (N_25118,N_23269,N_23024);
nand U25119 (N_25119,N_22928,N_21331);
nand U25120 (N_25120,N_21660,N_22383);
nor U25121 (N_25121,N_23998,N_22311);
nor U25122 (N_25122,N_21756,N_21889);
or U25123 (N_25123,N_21185,N_21169);
nor U25124 (N_25124,N_21318,N_23643);
and U25125 (N_25125,N_23087,N_21262);
nor U25126 (N_25126,N_23698,N_22110);
nand U25127 (N_25127,N_21375,N_23934);
nor U25128 (N_25128,N_23389,N_21409);
and U25129 (N_25129,N_21932,N_23207);
nor U25130 (N_25130,N_23933,N_23147);
nand U25131 (N_25131,N_23237,N_22645);
xnor U25132 (N_25132,N_23940,N_22081);
and U25133 (N_25133,N_23508,N_22095);
xnor U25134 (N_25134,N_21884,N_21133);
nand U25135 (N_25135,N_21078,N_23220);
xor U25136 (N_25136,N_23780,N_23564);
and U25137 (N_25137,N_23929,N_23035);
xor U25138 (N_25138,N_23664,N_21332);
nor U25139 (N_25139,N_22262,N_22232);
or U25140 (N_25140,N_22989,N_21690);
nand U25141 (N_25141,N_21560,N_22697);
xor U25142 (N_25142,N_21146,N_21053);
nor U25143 (N_25143,N_21511,N_22364);
and U25144 (N_25144,N_22414,N_22632);
nand U25145 (N_25145,N_22513,N_23914);
xor U25146 (N_25146,N_23835,N_22253);
nand U25147 (N_25147,N_21018,N_22167);
nor U25148 (N_25148,N_21149,N_22967);
or U25149 (N_25149,N_23714,N_23652);
nor U25150 (N_25150,N_21881,N_22415);
and U25151 (N_25151,N_22257,N_21474);
nand U25152 (N_25152,N_21256,N_21709);
nand U25153 (N_25153,N_21885,N_21808);
nand U25154 (N_25154,N_22166,N_23901);
nor U25155 (N_25155,N_22438,N_21563);
nor U25156 (N_25156,N_21351,N_22115);
xor U25157 (N_25157,N_22516,N_23357);
or U25158 (N_25158,N_22698,N_23580);
or U25159 (N_25159,N_22918,N_21028);
or U25160 (N_25160,N_22880,N_23489);
or U25161 (N_25161,N_23044,N_21606);
and U25162 (N_25162,N_22316,N_21798);
xnor U25163 (N_25163,N_23947,N_21479);
nor U25164 (N_25164,N_21724,N_21320);
or U25165 (N_25165,N_23796,N_22983);
nand U25166 (N_25166,N_21535,N_22474);
and U25167 (N_25167,N_21934,N_23377);
and U25168 (N_25168,N_23958,N_22734);
nor U25169 (N_25169,N_23140,N_21676);
or U25170 (N_25170,N_23374,N_21493);
and U25171 (N_25171,N_21518,N_22708);
or U25172 (N_25172,N_21908,N_23433);
or U25173 (N_25173,N_21025,N_21854);
or U25174 (N_25174,N_23521,N_22803);
xnor U25175 (N_25175,N_22503,N_21784);
nor U25176 (N_25176,N_23181,N_23678);
xnor U25177 (N_25177,N_22759,N_22377);
nand U25178 (N_25178,N_22539,N_22479);
nand U25179 (N_25179,N_22157,N_21958);
nor U25180 (N_25180,N_22411,N_23738);
or U25181 (N_25181,N_21387,N_22559);
nor U25182 (N_25182,N_23444,N_22540);
or U25183 (N_25183,N_22835,N_22207);
nor U25184 (N_25184,N_23965,N_22939);
or U25185 (N_25185,N_21077,N_22737);
or U25186 (N_25186,N_23410,N_22357);
nor U25187 (N_25187,N_22156,N_22427);
and U25188 (N_25188,N_22168,N_23717);
xnor U25189 (N_25189,N_22070,N_23781);
or U25190 (N_25190,N_21152,N_21736);
nor U25191 (N_25191,N_21962,N_22104);
or U25192 (N_25192,N_22836,N_23155);
xnor U25193 (N_25193,N_21095,N_22745);
or U25194 (N_25194,N_22410,N_23736);
nand U25195 (N_25195,N_21970,N_23561);
nor U25196 (N_25196,N_21080,N_22986);
and U25197 (N_25197,N_22069,N_23070);
xnor U25198 (N_25198,N_22245,N_22401);
or U25199 (N_25199,N_22283,N_22840);
nor U25200 (N_25200,N_22904,N_23013);
nand U25201 (N_25201,N_21344,N_23637);
or U25202 (N_25202,N_21088,N_21522);
nor U25203 (N_25203,N_21663,N_21468);
xnor U25204 (N_25204,N_21384,N_23310);
nand U25205 (N_25205,N_23482,N_21454);
nand U25206 (N_25206,N_23128,N_22946);
and U25207 (N_25207,N_22902,N_21447);
xor U25208 (N_25208,N_23100,N_23295);
nand U25209 (N_25209,N_21869,N_22889);
and U25210 (N_25210,N_21534,N_23999);
xor U25211 (N_25211,N_22123,N_22541);
and U25212 (N_25212,N_21333,N_23634);
nor U25213 (N_25213,N_23640,N_23691);
or U25214 (N_25214,N_23368,N_21386);
xor U25215 (N_25215,N_23711,N_21021);
nor U25216 (N_25216,N_21257,N_21554);
nor U25217 (N_25217,N_23651,N_21463);
xor U25218 (N_25218,N_21586,N_21587);
nor U25219 (N_25219,N_21401,N_23321);
or U25220 (N_25220,N_21108,N_21485);
or U25221 (N_25221,N_23856,N_22509);
nor U25222 (N_25222,N_22830,N_21747);
or U25223 (N_25223,N_23423,N_21144);
or U25224 (N_25224,N_22753,N_22760);
xnor U25225 (N_25225,N_23631,N_23844);
nor U25226 (N_25226,N_23392,N_22911);
and U25227 (N_25227,N_23932,N_22233);
or U25228 (N_25228,N_22447,N_22375);
and U25229 (N_25229,N_23865,N_21820);
xnor U25230 (N_25230,N_21207,N_22696);
or U25231 (N_25231,N_22868,N_21955);
and U25232 (N_25232,N_22826,N_23467);
nor U25233 (N_25233,N_22177,N_22514);
nand U25234 (N_25234,N_21910,N_23532);
and U25235 (N_25235,N_23563,N_21792);
and U25236 (N_25236,N_21642,N_23309);
nor U25237 (N_25237,N_21366,N_22782);
nand U25238 (N_25238,N_23861,N_23573);
or U25239 (N_25239,N_21772,N_22060);
nor U25240 (N_25240,N_22798,N_23396);
nor U25241 (N_25241,N_23450,N_22663);
or U25242 (N_25242,N_23383,N_21362);
xor U25243 (N_25243,N_23169,N_21898);
and U25244 (N_25244,N_22178,N_22325);
nor U25245 (N_25245,N_23363,N_22271);
nor U25246 (N_25246,N_21533,N_23990);
or U25247 (N_25247,N_21701,N_23653);
xnor U25248 (N_25248,N_21007,N_21746);
nand U25249 (N_25249,N_22615,N_23569);
or U25250 (N_25250,N_21729,N_21715);
xor U25251 (N_25251,N_23036,N_22124);
xor U25252 (N_25252,N_21341,N_21336);
xnor U25253 (N_25253,N_22355,N_23461);
nand U25254 (N_25254,N_22151,N_22105);
nor U25255 (N_25255,N_21235,N_23349);
nor U25256 (N_25256,N_21325,N_23968);
nand U25257 (N_25257,N_22443,N_23263);
nor U25258 (N_25258,N_23821,N_23548);
xor U25259 (N_25259,N_23735,N_23815);
or U25260 (N_25260,N_22936,N_22214);
and U25261 (N_25261,N_23362,N_21540);
nor U25262 (N_25262,N_23954,N_22694);
nand U25263 (N_25263,N_23065,N_23952);
nand U25264 (N_25264,N_23158,N_21924);
nor U25265 (N_25265,N_21850,N_21648);
and U25266 (N_25266,N_23339,N_21100);
nand U25267 (N_25267,N_22360,N_23479);
or U25268 (N_25268,N_21377,N_21182);
nor U25269 (N_25269,N_21839,N_23118);
nand U25270 (N_25270,N_21925,N_23586);
xor U25271 (N_25271,N_21214,N_23122);
or U25272 (N_25272,N_21967,N_23854);
xnor U25273 (N_25273,N_23623,N_23254);
and U25274 (N_25274,N_21172,N_21979);
nor U25275 (N_25275,N_23260,N_21707);
or U25276 (N_25276,N_21691,N_22806);
nand U25277 (N_25277,N_21995,N_23110);
nor U25278 (N_25278,N_22032,N_22442);
nor U25279 (N_25279,N_23808,N_22895);
or U25280 (N_25280,N_23746,N_21348);
nor U25281 (N_25281,N_22891,N_23546);
and U25282 (N_25282,N_21543,N_22522);
or U25283 (N_25283,N_21242,N_21462);
xnor U25284 (N_25284,N_22686,N_22877);
or U25285 (N_25285,N_22770,N_23601);
xnor U25286 (N_25286,N_21513,N_21717);
xor U25287 (N_25287,N_23451,N_23834);
nand U25288 (N_25288,N_21813,N_23121);
or U25289 (N_25289,N_21219,N_22225);
nand U25290 (N_25290,N_23646,N_22944);
nand U25291 (N_25291,N_23830,N_23472);
nor U25292 (N_25292,N_23286,N_23768);
and U25293 (N_25293,N_23106,N_22196);
or U25294 (N_25294,N_23560,N_21327);
nand U25295 (N_25295,N_21677,N_21939);
nor U25296 (N_25296,N_22587,N_22711);
and U25297 (N_25297,N_22091,N_22131);
and U25298 (N_25298,N_22107,N_21132);
nand U25299 (N_25299,N_21047,N_21625);
and U25300 (N_25300,N_23591,N_23407);
nor U25301 (N_25301,N_22235,N_23562);
xor U25302 (N_25302,N_23231,N_23814);
nor U25303 (N_25303,N_23827,N_22162);
and U25304 (N_25304,N_22788,N_23577);
xor U25305 (N_25305,N_21058,N_23504);
or U25306 (N_25306,N_22049,N_22160);
and U25307 (N_25307,N_21321,N_21668);
nor U25308 (N_25308,N_23731,N_22106);
or U25309 (N_25309,N_23997,N_21501);
xnor U25310 (N_25310,N_21517,N_23669);
and U25311 (N_25311,N_21382,N_22718);
nand U25312 (N_25312,N_21388,N_22432);
or U25313 (N_25313,N_23720,N_21430);
xor U25314 (N_25314,N_22499,N_22582);
nor U25315 (N_25315,N_21499,N_22703);
and U25316 (N_25316,N_23600,N_22171);
nand U25317 (N_25317,N_22339,N_22855);
nor U25318 (N_25318,N_21160,N_22702);
and U25319 (N_25319,N_23307,N_22498);
or U25320 (N_25320,N_23002,N_22523);
or U25321 (N_25321,N_23619,N_23666);
nand U25322 (N_25322,N_22763,N_23692);
nand U25323 (N_25323,N_23880,N_22270);
nor U25324 (N_25324,N_22963,N_21259);
nor U25325 (N_25325,N_23145,N_23045);
nand U25326 (N_25326,N_22406,N_22741);
and U25327 (N_25327,N_22751,N_22886);
xnor U25328 (N_25328,N_23372,N_23810);
or U25329 (N_25329,N_23441,N_23292);
and U25330 (N_25330,N_23570,N_21451);
xnor U25331 (N_25331,N_23027,N_22677);
xnor U25332 (N_25332,N_21449,N_21911);
nor U25333 (N_25333,N_21938,N_21486);
or U25334 (N_25334,N_23499,N_23531);
and U25335 (N_25335,N_22502,N_23761);
xnor U25336 (N_25336,N_22773,N_23622);
nor U25337 (N_25337,N_23142,N_21360);
nand U25338 (N_25338,N_23251,N_21323);
nor U25339 (N_25339,N_22630,N_22863);
nor U25340 (N_25340,N_23804,N_23115);
and U25341 (N_25341,N_21110,N_22116);
xnor U25342 (N_25342,N_22787,N_23867);
and U25343 (N_25343,N_21856,N_21555);
or U25344 (N_25344,N_21425,N_21825);
xor U25345 (N_25345,N_21983,N_22935);
and U25346 (N_25346,N_22016,N_21061);
nand U25347 (N_25347,N_21074,N_22980);
xor U25348 (N_25348,N_23439,N_23966);
and U25349 (N_25349,N_21931,N_23538);
or U25350 (N_25350,N_22141,N_21372);
nor U25351 (N_25351,N_23703,N_21926);
nor U25352 (N_25352,N_22762,N_22369);
nand U25353 (N_25353,N_23866,N_21098);
nor U25354 (N_25354,N_22228,N_22941);
and U25355 (N_25355,N_23988,N_21774);
nor U25356 (N_25356,N_22961,N_22791);
nor U25357 (N_25357,N_22658,N_22892);
nand U25358 (N_25358,N_23679,N_23491);
or U25359 (N_25359,N_23838,N_23052);
nand U25360 (N_25360,N_23300,N_22723);
and U25361 (N_25361,N_23589,N_23615);
or U25362 (N_25362,N_21805,N_21010);
nand U25363 (N_25363,N_23273,N_21196);
xor U25364 (N_25364,N_21419,N_23616);
nand U25365 (N_25365,N_23211,N_22704);
or U25366 (N_25366,N_21735,N_21504);
nor U25367 (N_25367,N_23324,N_22699);
and U25368 (N_25368,N_23950,N_22858);
and U25369 (N_25369,N_23293,N_23422);
nor U25370 (N_25370,N_21308,N_23948);
xor U25371 (N_25371,N_22379,N_21718);
xor U25372 (N_25372,N_22800,N_23520);
xnor U25373 (N_25373,N_22209,N_23056);
nand U25374 (N_25374,N_22268,N_22206);
and U25375 (N_25375,N_21443,N_23701);
nor U25376 (N_25376,N_21968,N_23873);
or U25377 (N_25377,N_22304,N_23981);
or U25378 (N_25378,N_22957,N_22086);
nor U25379 (N_25379,N_23053,N_23226);
nor U25380 (N_25380,N_22571,N_23463);
xnor U25381 (N_25381,N_21471,N_22288);
or U25382 (N_25382,N_23288,N_21564);
and U25383 (N_25383,N_21532,N_22781);
nor U25384 (N_25384,N_22717,N_22821);
nor U25385 (N_25385,N_23898,N_22023);
nor U25386 (N_25386,N_23785,N_21788);
and U25387 (N_25387,N_22888,N_21395);
or U25388 (N_25388,N_21841,N_23938);
nand U25389 (N_25389,N_23328,N_21872);
nor U25390 (N_25390,N_22794,N_21478);
xor U25391 (N_25391,N_21168,N_23219);
nand U25392 (N_25392,N_23160,N_21121);
xnor U25393 (N_25393,N_23620,N_21904);
and U25394 (N_25394,N_21001,N_21198);
and U25395 (N_25395,N_22966,N_23979);
and U25396 (N_25396,N_23897,N_23376);
and U25397 (N_25397,N_23648,N_22790);
nor U25398 (N_25398,N_21633,N_23927);
nor U25399 (N_25399,N_23650,N_23066);
nor U25400 (N_25400,N_22421,N_23797);
xnor U25401 (N_25401,N_23923,N_22591);
and U25402 (N_25402,N_23079,N_22805);
nand U25403 (N_25403,N_22890,N_21559);
or U25404 (N_25404,N_21117,N_21782);
xor U25405 (N_25405,N_22402,N_21046);
nand U25406 (N_25406,N_22566,N_23699);
and U25407 (N_25407,N_21828,N_22561);
and U25408 (N_25408,N_22258,N_23078);
xor U25409 (N_25409,N_22183,N_21129);
nor U25410 (N_25410,N_21723,N_23345);
and U25411 (N_25411,N_22856,N_21469);
nor U25412 (N_25412,N_23624,N_23632);
nand U25413 (N_25413,N_22975,N_23149);
xnor U25414 (N_25414,N_22380,N_21996);
nand U25415 (N_25415,N_22200,N_23046);
nand U25416 (N_25416,N_22845,N_22047);
nor U25417 (N_25417,N_23473,N_23716);
and U25418 (N_25418,N_22108,N_22619);
nor U25419 (N_25419,N_22159,N_23236);
and U25420 (N_25420,N_23682,N_23265);
xor U25421 (N_25421,N_23001,N_21328);
xor U25422 (N_25422,N_23173,N_21453);
xnor U25423 (N_25423,N_23899,N_22837);
and U25424 (N_25424,N_22129,N_21166);
nor U25425 (N_25425,N_22487,N_21376);
or U25426 (N_25426,N_22850,N_21456);
and U25427 (N_25427,N_21000,N_23949);
and U25428 (N_25428,N_22017,N_22784);
nand U25429 (N_25429,N_22862,N_21640);
xor U25430 (N_25430,N_22388,N_21888);
and U25431 (N_25431,N_21065,N_21254);
or U25432 (N_25432,N_23094,N_23612);
nor U25433 (N_25433,N_23818,N_21092);
nor U25434 (N_25434,N_22769,N_22367);
or U25435 (N_25435,N_22715,N_22817);
or U25436 (N_25436,N_23896,N_21776);
and U25437 (N_25437,N_21732,N_23161);
xor U25438 (N_25438,N_21719,N_23342);
nor U25439 (N_25439,N_21177,N_23608);
or U25440 (N_25440,N_21672,N_23481);
nor U25441 (N_25441,N_21937,N_23980);
nand U25442 (N_25442,N_21744,N_22833);
and U25443 (N_25443,N_23099,N_23862);
nand U25444 (N_25444,N_22190,N_22293);
nand U25445 (N_25445,N_21570,N_21249);
xnor U25446 (N_25446,N_22299,N_23906);
nand U25447 (N_25447,N_22467,N_22644);
or U25448 (N_25448,N_22595,N_22181);
nor U25449 (N_25449,N_22035,N_23091);
xnor U25450 (N_25450,N_23141,N_23611);
xnor U25451 (N_25451,N_22927,N_22778);
or U25452 (N_25452,N_23795,N_22875);
or U25453 (N_25453,N_22409,N_22144);
xor U25454 (N_25454,N_23911,N_21031);
xnor U25455 (N_25455,N_21702,N_21212);
nor U25456 (N_25456,N_22269,N_22002);
xnor U25457 (N_25457,N_22618,N_23683);
and U25458 (N_25458,N_22486,N_22096);
xnor U25459 (N_25459,N_21916,N_23055);
or U25460 (N_25460,N_21234,N_22263);
nor U25461 (N_25461,N_22296,N_21542);
and U25462 (N_25462,N_22093,N_21247);
and U25463 (N_25463,N_23280,N_23386);
nand U25464 (N_25464,N_21600,N_22940);
nand U25465 (N_25465,N_22730,N_23628);
and U25466 (N_25466,N_22074,N_23575);
or U25467 (N_25467,N_21652,N_21011);
nor U25468 (N_25468,N_22097,N_23585);
xor U25469 (N_25469,N_22389,N_22284);
nor U25470 (N_25470,N_22607,N_23690);
nand U25471 (N_25471,N_22504,N_22428);
xor U25472 (N_25472,N_21950,N_21787);
xor U25473 (N_25473,N_23483,N_23946);
xnor U25474 (N_25474,N_23193,N_22042);
or U25475 (N_25475,N_22398,N_23347);
and U25476 (N_25476,N_21383,N_21713);
and U25477 (N_25477,N_23477,N_22869);
and U25478 (N_25478,N_22633,N_23072);
or U25479 (N_25479,N_21840,N_22556);
nand U25480 (N_25480,N_23203,N_22265);
xor U25481 (N_25481,N_23029,N_23256);
xor U25482 (N_25482,N_22202,N_23536);
xor U25483 (N_25483,N_23244,N_22646);
xor U25484 (N_25484,N_22445,N_21613);
xnor U25485 (N_25485,N_23301,N_22593);
or U25486 (N_25486,N_23572,N_22018);
and U25487 (N_25487,N_21016,N_21710);
or U25488 (N_25488,N_21090,N_22098);
xnor U25489 (N_25489,N_23502,N_22538);
and U25490 (N_25490,N_22314,N_22831);
nor U25491 (N_25491,N_21971,N_21951);
nand U25492 (N_25492,N_23435,N_21883);
nand U25493 (N_25493,N_22362,N_21635);
nor U25494 (N_25494,N_23414,N_23123);
or U25495 (N_25495,N_23318,N_23857);
nand U25496 (N_25496,N_22461,N_22799);
nor U25497 (N_25497,N_22419,N_23734);
or U25498 (N_25498,N_21887,N_21602);
xor U25499 (N_25499,N_22695,N_22187);
or U25500 (N_25500,N_23046,N_23846);
xnor U25501 (N_25501,N_21544,N_21234);
nand U25502 (N_25502,N_22256,N_21821);
and U25503 (N_25503,N_22767,N_23001);
or U25504 (N_25504,N_21968,N_23224);
or U25505 (N_25505,N_21876,N_22749);
nand U25506 (N_25506,N_21873,N_22912);
and U25507 (N_25507,N_21081,N_21209);
nand U25508 (N_25508,N_22205,N_21630);
nand U25509 (N_25509,N_22705,N_21812);
nor U25510 (N_25510,N_21752,N_21767);
or U25511 (N_25511,N_23526,N_23550);
and U25512 (N_25512,N_23596,N_23555);
and U25513 (N_25513,N_23026,N_23175);
xnor U25514 (N_25514,N_22067,N_21726);
or U25515 (N_25515,N_22420,N_23861);
nand U25516 (N_25516,N_22974,N_22129);
nand U25517 (N_25517,N_22019,N_21996);
and U25518 (N_25518,N_22203,N_21679);
nand U25519 (N_25519,N_23804,N_23784);
or U25520 (N_25520,N_23009,N_21183);
xnor U25521 (N_25521,N_22705,N_21236);
xnor U25522 (N_25522,N_21226,N_21459);
nand U25523 (N_25523,N_23835,N_22364);
nand U25524 (N_25524,N_23869,N_22114);
nor U25525 (N_25525,N_23540,N_21244);
and U25526 (N_25526,N_23931,N_22557);
xnor U25527 (N_25527,N_22377,N_23249);
xor U25528 (N_25528,N_21762,N_21445);
or U25529 (N_25529,N_21107,N_22523);
xnor U25530 (N_25530,N_23328,N_21831);
and U25531 (N_25531,N_22862,N_22782);
xor U25532 (N_25532,N_23465,N_22521);
nand U25533 (N_25533,N_21037,N_21667);
and U25534 (N_25534,N_21709,N_23056);
and U25535 (N_25535,N_22527,N_22789);
nand U25536 (N_25536,N_22454,N_23797);
and U25537 (N_25537,N_23877,N_21946);
nand U25538 (N_25538,N_22042,N_23797);
and U25539 (N_25539,N_23516,N_23588);
or U25540 (N_25540,N_23326,N_21766);
nor U25541 (N_25541,N_23906,N_21453);
xnor U25542 (N_25542,N_21146,N_21064);
or U25543 (N_25543,N_22780,N_21418);
nand U25544 (N_25544,N_22565,N_22257);
nand U25545 (N_25545,N_23727,N_22555);
xnor U25546 (N_25546,N_23815,N_22414);
and U25547 (N_25547,N_22221,N_23092);
xnor U25548 (N_25548,N_22965,N_21061);
or U25549 (N_25549,N_22845,N_23982);
and U25550 (N_25550,N_23518,N_21672);
nand U25551 (N_25551,N_21950,N_21113);
and U25552 (N_25552,N_22336,N_21426);
or U25553 (N_25553,N_21563,N_21348);
nor U25554 (N_25554,N_23886,N_23367);
xor U25555 (N_25555,N_21906,N_23728);
nand U25556 (N_25556,N_23766,N_22998);
and U25557 (N_25557,N_23191,N_23646);
nand U25558 (N_25558,N_23668,N_22581);
or U25559 (N_25559,N_22924,N_22051);
nand U25560 (N_25560,N_21322,N_22591);
nor U25561 (N_25561,N_21498,N_23879);
xor U25562 (N_25562,N_21342,N_21894);
nand U25563 (N_25563,N_23703,N_22555);
or U25564 (N_25564,N_21825,N_23521);
nand U25565 (N_25565,N_21650,N_22898);
or U25566 (N_25566,N_23566,N_21650);
xor U25567 (N_25567,N_21072,N_21600);
xnor U25568 (N_25568,N_21092,N_23145);
nand U25569 (N_25569,N_21241,N_21608);
xnor U25570 (N_25570,N_23581,N_21578);
nand U25571 (N_25571,N_22614,N_22090);
or U25572 (N_25572,N_23967,N_23838);
or U25573 (N_25573,N_23885,N_22802);
and U25574 (N_25574,N_21529,N_23448);
or U25575 (N_25575,N_21279,N_21836);
and U25576 (N_25576,N_22989,N_21450);
or U25577 (N_25577,N_21802,N_22921);
nor U25578 (N_25578,N_23712,N_22762);
or U25579 (N_25579,N_22207,N_23464);
xnor U25580 (N_25580,N_21093,N_23469);
or U25581 (N_25581,N_22982,N_21705);
xnor U25582 (N_25582,N_23101,N_22301);
nand U25583 (N_25583,N_23521,N_22343);
nand U25584 (N_25584,N_23606,N_22359);
nand U25585 (N_25585,N_22777,N_23101);
nand U25586 (N_25586,N_23690,N_23497);
or U25587 (N_25587,N_23602,N_22976);
xnor U25588 (N_25588,N_22089,N_22652);
xor U25589 (N_25589,N_21678,N_23831);
and U25590 (N_25590,N_21052,N_23046);
and U25591 (N_25591,N_21660,N_23327);
xnor U25592 (N_25592,N_21106,N_21768);
and U25593 (N_25593,N_23429,N_23499);
and U25594 (N_25594,N_22089,N_23382);
nand U25595 (N_25595,N_22574,N_21307);
nor U25596 (N_25596,N_23873,N_22490);
and U25597 (N_25597,N_23868,N_23489);
nand U25598 (N_25598,N_21290,N_22498);
or U25599 (N_25599,N_22309,N_23029);
nand U25600 (N_25600,N_23239,N_21917);
nor U25601 (N_25601,N_21287,N_23210);
xor U25602 (N_25602,N_23147,N_21670);
nor U25603 (N_25603,N_21186,N_22750);
nor U25604 (N_25604,N_21723,N_23265);
xor U25605 (N_25605,N_21896,N_22919);
nand U25606 (N_25606,N_23222,N_22935);
nor U25607 (N_25607,N_22374,N_22012);
and U25608 (N_25608,N_22562,N_22868);
xor U25609 (N_25609,N_21663,N_22308);
and U25610 (N_25610,N_22896,N_22376);
xnor U25611 (N_25611,N_22197,N_21218);
nand U25612 (N_25612,N_22823,N_23477);
nand U25613 (N_25613,N_23538,N_23450);
or U25614 (N_25614,N_21795,N_23561);
nor U25615 (N_25615,N_22288,N_22990);
nor U25616 (N_25616,N_23522,N_23211);
nand U25617 (N_25617,N_21457,N_23371);
nor U25618 (N_25618,N_22060,N_21255);
nand U25619 (N_25619,N_21400,N_23911);
nor U25620 (N_25620,N_22459,N_22885);
nand U25621 (N_25621,N_21268,N_23187);
xnor U25622 (N_25622,N_23910,N_22120);
or U25623 (N_25623,N_21664,N_21837);
nand U25624 (N_25624,N_22823,N_23615);
or U25625 (N_25625,N_21755,N_23282);
xor U25626 (N_25626,N_21866,N_21185);
nor U25627 (N_25627,N_21994,N_23857);
xor U25628 (N_25628,N_23094,N_22136);
xor U25629 (N_25629,N_22197,N_21674);
nor U25630 (N_25630,N_23093,N_22839);
or U25631 (N_25631,N_23712,N_21877);
nor U25632 (N_25632,N_21777,N_22736);
nand U25633 (N_25633,N_23873,N_21930);
or U25634 (N_25634,N_22622,N_23454);
nor U25635 (N_25635,N_22899,N_22199);
or U25636 (N_25636,N_21058,N_21032);
xor U25637 (N_25637,N_22559,N_23358);
xnor U25638 (N_25638,N_22099,N_21990);
xnor U25639 (N_25639,N_21738,N_22726);
and U25640 (N_25640,N_22579,N_23016);
xor U25641 (N_25641,N_21239,N_21073);
nor U25642 (N_25642,N_22301,N_21737);
nor U25643 (N_25643,N_22427,N_23624);
xor U25644 (N_25644,N_22571,N_22576);
and U25645 (N_25645,N_23275,N_23901);
and U25646 (N_25646,N_22914,N_21972);
or U25647 (N_25647,N_23947,N_22351);
and U25648 (N_25648,N_21290,N_23926);
and U25649 (N_25649,N_23483,N_21877);
and U25650 (N_25650,N_21643,N_21496);
xor U25651 (N_25651,N_22998,N_21362);
nor U25652 (N_25652,N_21852,N_21975);
nor U25653 (N_25653,N_21180,N_22150);
xor U25654 (N_25654,N_22285,N_22953);
nor U25655 (N_25655,N_21490,N_21047);
nor U25656 (N_25656,N_23827,N_21018);
or U25657 (N_25657,N_23282,N_21393);
nand U25658 (N_25658,N_22737,N_23848);
and U25659 (N_25659,N_23232,N_21091);
xor U25660 (N_25660,N_23996,N_23003);
or U25661 (N_25661,N_22177,N_21289);
xnor U25662 (N_25662,N_22578,N_22070);
xnor U25663 (N_25663,N_23389,N_23641);
xnor U25664 (N_25664,N_23389,N_23705);
nor U25665 (N_25665,N_21000,N_23398);
or U25666 (N_25666,N_21875,N_23749);
nand U25667 (N_25667,N_22053,N_21701);
and U25668 (N_25668,N_21853,N_22015);
nand U25669 (N_25669,N_22336,N_21552);
and U25670 (N_25670,N_22689,N_23525);
nand U25671 (N_25671,N_23695,N_23256);
nor U25672 (N_25672,N_23043,N_22807);
xnor U25673 (N_25673,N_22431,N_22031);
and U25674 (N_25674,N_21909,N_22967);
xor U25675 (N_25675,N_23775,N_23583);
xor U25676 (N_25676,N_23456,N_21986);
xnor U25677 (N_25677,N_22716,N_22087);
nand U25678 (N_25678,N_22845,N_22167);
nor U25679 (N_25679,N_22113,N_23836);
xnor U25680 (N_25680,N_22708,N_21975);
nor U25681 (N_25681,N_23852,N_23304);
and U25682 (N_25682,N_23125,N_23884);
and U25683 (N_25683,N_23033,N_23415);
or U25684 (N_25684,N_23943,N_23159);
xnor U25685 (N_25685,N_23080,N_21171);
xor U25686 (N_25686,N_21128,N_23124);
nand U25687 (N_25687,N_22676,N_22498);
and U25688 (N_25688,N_22826,N_22893);
or U25689 (N_25689,N_23517,N_21693);
nor U25690 (N_25690,N_21008,N_21759);
or U25691 (N_25691,N_22176,N_21648);
nor U25692 (N_25692,N_23135,N_21777);
nand U25693 (N_25693,N_22545,N_21515);
and U25694 (N_25694,N_22366,N_23253);
or U25695 (N_25695,N_23841,N_22594);
nor U25696 (N_25696,N_21541,N_21858);
or U25697 (N_25697,N_23567,N_21263);
or U25698 (N_25698,N_21603,N_22477);
xnor U25699 (N_25699,N_22995,N_23142);
and U25700 (N_25700,N_22013,N_21627);
xor U25701 (N_25701,N_23717,N_21621);
nand U25702 (N_25702,N_21670,N_22401);
or U25703 (N_25703,N_21204,N_21886);
or U25704 (N_25704,N_21190,N_22534);
or U25705 (N_25705,N_23790,N_23554);
xnor U25706 (N_25706,N_22237,N_21833);
and U25707 (N_25707,N_21953,N_23735);
nor U25708 (N_25708,N_21758,N_22961);
xnor U25709 (N_25709,N_22188,N_22719);
nand U25710 (N_25710,N_22032,N_22445);
xor U25711 (N_25711,N_23738,N_23168);
nor U25712 (N_25712,N_21663,N_23815);
or U25713 (N_25713,N_22971,N_22962);
nand U25714 (N_25714,N_22735,N_22451);
or U25715 (N_25715,N_22236,N_23286);
nor U25716 (N_25716,N_22754,N_22610);
and U25717 (N_25717,N_22220,N_23377);
nand U25718 (N_25718,N_22127,N_21318);
nor U25719 (N_25719,N_21308,N_22929);
nand U25720 (N_25720,N_22290,N_23000);
nand U25721 (N_25721,N_21513,N_23146);
nor U25722 (N_25722,N_22213,N_23885);
nand U25723 (N_25723,N_22454,N_23330);
and U25724 (N_25724,N_22744,N_21468);
nor U25725 (N_25725,N_22227,N_23536);
xnor U25726 (N_25726,N_22484,N_21192);
and U25727 (N_25727,N_21377,N_23022);
and U25728 (N_25728,N_22996,N_21482);
and U25729 (N_25729,N_23000,N_21541);
and U25730 (N_25730,N_22158,N_21784);
nand U25731 (N_25731,N_21861,N_21278);
nand U25732 (N_25732,N_22368,N_23697);
nor U25733 (N_25733,N_23513,N_21975);
xnor U25734 (N_25734,N_23990,N_22620);
or U25735 (N_25735,N_22062,N_21525);
or U25736 (N_25736,N_22489,N_21645);
and U25737 (N_25737,N_21093,N_22706);
or U25738 (N_25738,N_22399,N_23606);
and U25739 (N_25739,N_23772,N_22743);
or U25740 (N_25740,N_23779,N_23816);
or U25741 (N_25741,N_21897,N_22695);
xnor U25742 (N_25742,N_21977,N_23292);
and U25743 (N_25743,N_23525,N_22788);
nor U25744 (N_25744,N_22690,N_22048);
and U25745 (N_25745,N_23141,N_23180);
nor U25746 (N_25746,N_21683,N_21110);
nor U25747 (N_25747,N_23182,N_21961);
and U25748 (N_25748,N_22362,N_22246);
or U25749 (N_25749,N_21624,N_21084);
or U25750 (N_25750,N_22986,N_22865);
xnor U25751 (N_25751,N_22850,N_23539);
nand U25752 (N_25752,N_21594,N_22121);
or U25753 (N_25753,N_23000,N_23270);
xor U25754 (N_25754,N_21276,N_23306);
nand U25755 (N_25755,N_23873,N_22458);
xnor U25756 (N_25756,N_21083,N_23628);
xor U25757 (N_25757,N_21538,N_23954);
and U25758 (N_25758,N_22822,N_23919);
nor U25759 (N_25759,N_23288,N_21889);
nor U25760 (N_25760,N_23307,N_21037);
xnor U25761 (N_25761,N_21994,N_21127);
and U25762 (N_25762,N_22496,N_22485);
nand U25763 (N_25763,N_23134,N_21022);
and U25764 (N_25764,N_22545,N_23097);
nand U25765 (N_25765,N_22474,N_21984);
nor U25766 (N_25766,N_22366,N_23405);
nor U25767 (N_25767,N_22097,N_21756);
xor U25768 (N_25768,N_21346,N_23903);
xor U25769 (N_25769,N_23052,N_22814);
or U25770 (N_25770,N_22088,N_23533);
or U25771 (N_25771,N_21795,N_22086);
nand U25772 (N_25772,N_21609,N_23821);
nor U25773 (N_25773,N_22321,N_21172);
nor U25774 (N_25774,N_22863,N_21129);
xnor U25775 (N_25775,N_21359,N_22085);
or U25776 (N_25776,N_23195,N_22110);
xor U25777 (N_25777,N_23137,N_23686);
nand U25778 (N_25778,N_22681,N_23404);
or U25779 (N_25779,N_21019,N_23924);
nand U25780 (N_25780,N_22955,N_23615);
or U25781 (N_25781,N_22059,N_22015);
xnor U25782 (N_25782,N_23739,N_21516);
xnor U25783 (N_25783,N_23459,N_23234);
nor U25784 (N_25784,N_21036,N_23362);
xor U25785 (N_25785,N_22149,N_22563);
nor U25786 (N_25786,N_23503,N_23859);
nor U25787 (N_25787,N_22396,N_22924);
or U25788 (N_25788,N_23930,N_23692);
nand U25789 (N_25789,N_22376,N_21240);
nand U25790 (N_25790,N_22179,N_23870);
and U25791 (N_25791,N_23662,N_22210);
xnor U25792 (N_25792,N_22503,N_23502);
or U25793 (N_25793,N_23563,N_23217);
and U25794 (N_25794,N_21679,N_22586);
nor U25795 (N_25795,N_21898,N_21511);
nor U25796 (N_25796,N_21382,N_21841);
nand U25797 (N_25797,N_21337,N_23433);
or U25798 (N_25798,N_22188,N_23666);
nor U25799 (N_25799,N_23539,N_22680);
nor U25800 (N_25800,N_21023,N_22139);
and U25801 (N_25801,N_23240,N_21803);
nor U25802 (N_25802,N_21000,N_21787);
or U25803 (N_25803,N_21604,N_22313);
nand U25804 (N_25804,N_23770,N_22285);
xor U25805 (N_25805,N_21363,N_22432);
nor U25806 (N_25806,N_21524,N_22276);
or U25807 (N_25807,N_22966,N_22923);
and U25808 (N_25808,N_21618,N_21870);
or U25809 (N_25809,N_23721,N_21758);
and U25810 (N_25810,N_21042,N_23643);
or U25811 (N_25811,N_22390,N_22946);
and U25812 (N_25812,N_22313,N_21543);
nand U25813 (N_25813,N_21576,N_22074);
xnor U25814 (N_25814,N_21351,N_21805);
or U25815 (N_25815,N_23129,N_21681);
nand U25816 (N_25816,N_21212,N_21936);
and U25817 (N_25817,N_23502,N_23425);
or U25818 (N_25818,N_21734,N_21427);
nand U25819 (N_25819,N_22892,N_22294);
nand U25820 (N_25820,N_22636,N_22773);
or U25821 (N_25821,N_23999,N_22775);
xnor U25822 (N_25822,N_23199,N_21608);
or U25823 (N_25823,N_22776,N_22092);
nor U25824 (N_25824,N_23319,N_22282);
xor U25825 (N_25825,N_22187,N_22035);
or U25826 (N_25826,N_23253,N_23110);
xor U25827 (N_25827,N_21977,N_22173);
and U25828 (N_25828,N_23213,N_23800);
and U25829 (N_25829,N_22939,N_21234);
or U25830 (N_25830,N_22500,N_22370);
nand U25831 (N_25831,N_22155,N_21867);
nand U25832 (N_25832,N_21736,N_22420);
and U25833 (N_25833,N_23961,N_21321);
and U25834 (N_25834,N_21345,N_22301);
nor U25835 (N_25835,N_21585,N_21837);
and U25836 (N_25836,N_21728,N_21653);
xor U25837 (N_25837,N_22152,N_21365);
xnor U25838 (N_25838,N_23422,N_23775);
nand U25839 (N_25839,N_21207,N_22486);
and U25840 (N_25840,N_23878,N_21106);
or U25841 (N_25841,N_23938,N_21946);
nor U25842 (N_25842,N_22036,N_21312);
xnor U25843 (N_25843,N_22393,N_23501);
xnor U25844 (N_25844,N_23087,N_23775);
and U25845 (N_25845,N_22052,N_22530);
and U25846 (N_25846,N_22282,N_22279);
xor U25847 (N_25847,N_22296,N_23242);
nor U25848 (N_25848,N_23226,N_22170);
or U25849 (N_25849,N_21049,N_22793);
xnor U25850 (N_25850,N_22334,N_22275);
nor U25851 (N_25851,N_21516,N_22169);
nor U25852 (N_25852,N_22327,N_21622);
and U25853 (N_25853,N_22277,N_23401);
nor U25854 (N_25854,N_21739,N_22288);
or U25855 (N_25855,N_21646,N_23241);
nand U25856 (N_25856,N_22666,N_22515);
or U25857 (N_25857,N_21006,N_22589);
or U25858 (N_25858,N_21043,N_23724);
xnor U25859 (N_25859,N_22600,N_23949);
or U25860 (N_25860,N_22337,N_21819);
nor U25861 (N_25861,N_23648,N_23366);
and U25862 (N_25862,N_23577,N_21428);
nor U25863 (N_25863,N_21897,N_22520);
xor U25864 (N_25864,N_23115,N_22581);
nand U25865 (N_25865,N_21596,N_21629);
nor U25866 (N_25866,N_22244,N_22627);
nand U25867 (N_25867,N_23823,N_21506);
and U25868 (N_25868,N_22398,N_23182);
nand U25869 (N_25869,N_22703,N_22142);
nand U25870 (N_25870,N_23770,N_21044);
xnor U25871 (N_25871,N_22723,N_22581);
nand U25872 (N_25872,N_22295,N_23787);
nand U25873 (N_25873,N_23523,N_22352);
and U25874 (N_25874,N_23424,N_23446);
xnor U25875 (N_25875,N_23855,N_23288);
or U25876 (N_25876,N_21440,N_22586);
or U25877 (N_25877,N_21877,N_22803);
nor U25878 (N_25878,N_22705,N_21602);
nand U25879 (N_25879,N_22253,N_21924);
nor U25880 (N_25880,N_22531,N_22525);
nand U25881 (N_25881,N_21371,N_21356);
nor U25882 (N_25882,N_22255,N_21755);
and U25883 (N_25883,N_22673,N_21382);
and U25884 (N_25884,N_23847,N_23530);
nor U25885 (N_25885,N_21352,N_23478);
nor U25886 (N_25886,N_22291,N_22910);
nor U25887 (N_25887,N_21938,N_21653);
and U25888 (N_25888,N_22666,N_21903);
or U25889 (N_25889,N_23295,N_21942);
and U25890 (N_25890,N_21344,N_23491);
nand U25891 (N_25891,N_21589,N_21535);
nand U25892 (N_25892,N_22136,N_23089);
and U25893 (N_25893,N_22339,N_22705);
nor U25894 (N_25894,N_21773,N_22398);
nand U25895 (N_25895,N_23779,N_22642);
nor U25896 (N_25896,N_23636,N_23556);
xnor U25897 (N_25897,N_21854,N_23967);
nor U25898 (N_25898,N_21597,N_21152);
nand U25899 (N_25899,N_22662,N_23695);
nand U25900 (N_25900,N_22867,N_21596);
nor U25901 (N_25901,N_22035,N_22134);
or U25902 (N_25902,N_21124,N_23858);
xnor U25903 (N_25903,N_21189,N_22274);
xor U25904 (N_25904,N_23435,N_22445);
and U25905 (N_25905,N_21034,N_22315);
or U25906 (N_25906,N_22545,N_21259);
nor U25907 (N_25907,N_23019,N_22821);
xor U25908 (N_25908,N_23025,N_22538);
xnor U25909 (N_25909,N_21918,N_22955);
and U25910 (N_25910,N_21156,N_23893);
nor U25911 (N_25911,N_22454,N_21176);
nand U25912 (N_25912,N_22662,N_23295);
and U25913 (N_25913,N_22526,N_21114);
or U25914 (N_25914,N_23998,N_22552);
and U25915 (N_25915,N_22918,N_23729);
nand U25916 (N_25916,N_23214,N_21494);
and U25917 (N_25917,N_21464,N_22882);
and U25918 (N_25918,N_21135,N_22342);
nor U25919 (N_25919,N_21863,N_22356);
xor U25920 (N_25920,N_22146,N_22493);
xnor U25921 (N_25921,N_23951,N_23134);
nand U25922 (N_25922,N_22266,N_21534);
nor U25923 (N_25923,N_22355,N_21972);
nor U25924 (N_25924,N_22891,N_22200);
or U25925 (N_25925,N_21129,N_21634);
xor U25926 (N_25926,N_23283,N_21650);
and U25927 (N_25927,N_23424,N_21296);
xnor U25928 (N_25928,N_21409,N_23592);
xor U25929 (N_25929,N_23776,N_21440);
or U25930 (N_25930,N_23311,N_22639);
or U25931 (N_25931,N_22470,N_23502);
or U25932 (N_25932,N_22832,N_23759);
nand U25933 (N_25933,N_22023,N_23226);
or U25934 (N_25934,N_23172,N_23672);
and U25935 (N_25935,N_22579,N_23895);
nand U25936 (N_25936,N_21119,N_22256);
or U25937 (N_25937,N_22502,N_21293);
nor U25938 (N_25938,N_21206,N_22581);
and U25939 (N_25939,N_21376,N_22698);
nand U25940 (N_25940,N_21414,N_21722);
and U25941 (N_25941,N_23234,N_23323);
xor U25942 (N_25942,N_23613,N_21555);
xnor U25943 (N_25943,N_23307,N_22123);
nor U25944 (N_25944,N_23623,N_23570);
nand U25945 (N_25945,N_21600,N_21425);
nor U25946 (N_25946,N_23687,N_22196);
xnor U25947 (N_25947,N_22337,N_22022);
nor U25948 (N_25948,N_23744,N_23176);
nand U25949 (N_25949,N_22204,N_21224);
xor U25950 (N_25950,N_21839,N_21651);
nor U25951 (N_25951,N_21420,N_21238);
nand U25952 (N_25952,N_22780,N_22826);
xor U25953 (N_25953,N_23661,N_22539);
and U25954 (N_25954,N_23195,N_21822);
or U25955 (N_25955,N_21833,N_23332);
or U25956 (N_25956,N_22246,N_23966);
or U25957 (N_25957,N_21419,N_23957);
or U25958 (N_25958,N_23337,N_23204);
xor U25959 (N_25959,N_22213,N_22055);
and U25960 (N_25960,N_22829,N_22174);
and U25961 (N_25961,N_22232,N_21195);
nor U25962 (N_25962,N_23228,N_21370);
or U25963 (N_25963,N_22725,N_22528);
or U25964 (N_25964,N_23773,N_21169);
xor U25965 (N_25965,N_21096,N_22350);
and U25966 (N_25966,N_22421,N_23953);
nor U25967 (N_25967,N_22998,N_21074);
or U25968 (N_25968,N_21627,N_21502);
nor U25969 (N_25969,N_22880,N_21434);
or U25970 (N_25970,N_23813,N_23705);
or U25971 (N_25971,N_21677,N_21019);
or U25972 (N_25972,N_22622,N_21783);
and U25973 (N_25973,N_23134,N_22650);
and U25974 (N_25974,N_21143,N_22881);
and U25975 (N_25975,N_22800,N_22508);
nor U25976 (N_25976,N_23927,N_22513);
xor U25977 (N_25977,N_23411,N_23462);
or U25978 (N_25978,N_22121,N_21105);
or U25979 (N_25979,N_22397,N_23600);
or U25980 (N_25980,N_23636,N_22556);
or U25981 (N_25981,N_23457,N_23785);
or U25982 (N_25982,N_21639,N_22466);
or U25983 (N_25983,N_21055,N_21320);
nand U25984 (N_25984,N_23789,N_23721);
and U25985 (N_25985,N_23448,N_22429);
nor U25986 (N_25986,N_21222,N_23014);
nor U25987 (N_25987,N_22554,N_21759);
xnor U25988 (N_25988,N_21868,N_21071);
or U25989 (N_25989,N_22326,N_22533);
nor U25990 (N_25990,N_23814,N_22360);
and U25991 (N_25991,N_21355,N_22726);
or U25992 (N_25992,N_22271,N_21566);
nor U25993 (N_25993,N_21688,N_23936);
nand U25994 (N_25994,N_22935,N_22172);
nor U25995 (N_25995,N_22818,N_22800);
or U25996 (N_25996,N_21152,N_22757);
nand U25997 (N_25997,N_22035,N_21163);
or U25998 (N_25998,N_22992,N_23739);
nand U25999 (N_25999,N_22458,N_21710);
nor U26000 (N_26000,N_23056,N_23893);
or U26001 (N_26001,N_21286,N_21033);
nor U26002 (N_26002,N_21053,N_21355);
and U26003 (N_26003,N_22948,N_22732);
and U26004 (N_26004,N_23494,N_23690);
or U26005 (N_26005,N_22990,N_22420);
xor U26006 (N_26006,N_23187,N_21159);
nor U26007 (N_26007,N_22060,N_23644);
nand U26008 (N_26008,N_23664,N_21081);
or U26009 (N_26009,N_23115,N_21427);
nor U26010 (N_26010,N_23566,N_22892);
xnor U26011 (N_26011,N_21282,N_23432);
and U26012 (N_26012,N_21817,N_21261);
or U26013 (N_26013,N_22969,N_21646);
or U26014 (N_26014,N_22595,N_23727);
and U26015 (N_26015,N_22676,N_22519);
and U26016 (N_26016,N_21108,N_21878);
and U26017 (N_26017,N_23126,N_22448);
nor U26018 (N_26018,N_21700,N_21305);
xor U26019 (N_26019,N_22506,N_21254);
nand U26020 (N_26020,N_21358,N_22301);
nor U26021 (N_26021,N_22356,N_22834);
and U26022 (N_26022,N_21783,N_21659);
and U26023 (N_26023,N_22053,N_22035);
and U26024 (N_26024,N_23071,N_23449);
and U26025 (N_26025,N_21344,N_21889);
or U26026 (N_26026,N_23193,N_21814);
xnor U26027 (N_26027,N_23672,N_22110);
nand U26028 (N_26028,N_23950,N_23659);
or U26029 (N_26029,N_22300,N_22114);
nor U26030 (N_26030,N_22017,N_23524);
and U26031 (N_26031,N_23174,N_22792);
and U26032 (N_26032,N_22204,N_23873);
xnor U26033 (N_26033,N_21880,N_21599);
nor U26034 (N_26034,N_23893,N_23683);
xor U26035 (N_26035,N_22818,N_22736);
and U26036 (N_26036,N_21967,N_23212);
or U26037 (N_26037,N_23607,N_23288);
xor U26038 (N_26038,N_21912,N_21348);
or U26039 (N_26039,N_23388,N_22790);
or U26040 (N_26040,N_23070,N_21695);
nor U26041 (N_26041,N_22031,N_21396);
nor U26042 (N_26042,N_22444,N_21841);
nor U26043 (N_26043,N_21791,N_21771);
and U26044 (N_26044,N_22133,N_22744);
or U26045 (N_26045,N_23216,N_22070);
nor U26046 (N_26046,N_22048,N_23033);
or U26047 (N_26047,N_22909,N_23364);
xor U26048 (N_26048,N_23930,N_21802);
nor U26049 (N_26049,N_21539,N_21102);
and U26050 (N_26050,N_21567,N_22435);
or U26051 (N_26051,N_23773,N_21834);
nor U26052 (N_26052,N_22794,N_23812);
xnor U26053 (N_26053,N_21473,N_21896);
nor U26054 (N_26054,N_22492,N_23897);
or U26055 (N_26055,N_22727,N_21155);
and U26056 (N_26056,N_23390,N_21167);
nand U26057 (N_26057,N_22274,N_22843);
and U26058 (N_26058,N_22458,N_21191);
nand U26059 (N_26059,N_21643,N_23573);
nand U26060 (N_26060,N_21210,N_23947);
nor U26061 (N_26061,N_21017,N_21062);
xor U26062 (N_26062,N_23619,N_21257);
and U26063 (N_26063,N_23263,N_23279);
nor U26064 (N_26064,N_23523,N_22545);
xnor U26065 (N_26065,N_21735,N_21414);
nor U26066 (N_26066,N_22819,N_21766);
or U26067 (N_26067,N_23698,N_22424);
xnor U26068 (N_26068,N_23114,N_21785);
xnor U26069 (N_26069,N_23241,N_23475);
nor U26070 (N_26070,N_22499,N_22798);
and U26071 (N_26071,N_22351,N_23209);
nand U26072 (N_26072,N_21051,N_21009);
and U26073 (N_26073,N_23297,N_21412);
nand U26074 (N_26074,N_22916,N_23162);
xor U26075 (N_26075,N_23493,N_21053);
nor U26076 (N_26076,N_22712,N_21153);
nor U26077 (N_26077,N_23821,N_22303);
xor U26078 (N_26078,N_23972,N_22066);
nor U26079 (N_26079,N_21976,N_22163);
and U26080 (N_26080,N_22162,N_22907);
and U26081 (N_26081,N_21263,N_23289);
or U26082 (N_26082,N_23236,N_22208);
nand U26083 (N_26083,N_21839,N_23028);
nor U26084 (N_26084,N_23718,N_21550);
or U26085 (N_26085,N_21736,N_21684);
xor U26086 (N_26086,N_23138,N_21447);
nor U26087 (N_26087,N_23083,N_23548);
xor U26088 (N_26088,N_23832,N_23636);
nor U26089 (N_26089,N_23883,N_21986);
nand U26090 (N_26090,N_22442,N_21258);
nand U26091 (N_26091,N_21153,N_22964);
xor U26092 (N_26092,N_21196,N_21619);
or U26093 (N_26093,N_23089,N_21817);
nand U26094 (N_26094,N_23865,N_22345);
nand U26095 (N_26095,N_21909,N_21039);
and U26096 (N_26096,N_22072,N_23128);
xor U26097 (N_26097,N_23159,N_22221);
nor U26098 (N_26098,N_22414,N_23913);
xnor U26099 (N_26099,N_23509,N_22098);
and U26100 (N_26100,N_21711,N_21547);
or U26101 (N_26101,N_22524,N_22540);
xnor U26102 (N_26102,N_22849,N_22424);
and U26103 (N_26103,N_22268,N_22752);
and U26104 (N_26104,N_21942,N_22772);
and U26105 (N_26105,N_21909,N_21652);
nor U26106 (N_26106,N_23072,N_23685);
nor U26107 (N_26107,N_21355,N_23339);
nand U26108 (N_26108,N_22360,N_22006);
or U26109 (N_26109,N_22194,N_22827);
nor U26110 (N_26110,N_21498,N_21160);
and U26111 (N_26111,N_21442,N_21803);
or U26112 (N_26112,N_23966,N_23769);
xnor U26113 (N_26113,N_21924,N_21101);
nor U26114 (N_26114,N_22900,N_21328);
xnor U26115 (N_26115,N_21223,N_23712);
xor U26116 (N_26116,N_22032,N_22242);
or U26117 (N_26117,N_21784,N_21664);
nand U26118 (N_26118,N_23701,N_23455);
and U26119 (N_26119,N_23338,N_22304);
and U26120 (N_26120,N_22298,N_23906);
or U26121 (N_26121,N_22750,N_23915);
nand U26122 (N_26122,N_22966,N_21777);
xnor U26123 (N_26123,N_21125,N_21624);
nor U26124 (N_26124,N_22803,N_21324);
nor U26125 (N_26125,N_23029,N_23134);
nand U26126 (N_26126,N_21929,N_21715);
nand U26127 (N_26127,N_23107,N_23893);
nand U26128 (N_26128,N_22417,N_22004);
nand U26129 (N_26129,N_23983,N_22930);
nor U26130 (N_26130,N_23371,N_23909);
nand U26131 (N_26131,N_23514,N_23420);
and U26132 (N_26132,N_23999,N_22969);
and U26133 (N_26133,N_22730,N_21294);
xor U26134 (N_26134,N_21275,N_23549);
nand U26135 (N_26135,N_22068,N_22503);
nand U26136 (N_26136,N_22983,N_23311);
or U26137 (N_26137,N_23251,N_21680);
and U26138 (N_26138,N_21405,N_23515);
and U26139 (N_26139,N_22787,N_23554);
xor U26140 (N_26140,N_23937,N_21037);
and U26141 (N_26141,N_22334,N_21894);
nor U26142 (N_26142,N_23057,N_22498);
xnor U26143 (N_26143,N_23531,N_22930);
nor U26144 (N_26144,N_21334,N_21908);
xor U26145 (N_26145,N_21357,N_22759);
nor U26146 (N_26146,N_21973,N_21379);
and U26147 (N_26147,N_21380,N_22792);
and U26148 (N_26148,N_21538,N_23118);
and U26149 (N_26149,N_23534,N_22025);
or U26150 (N_26150,N_22454,N_23879);
and U26151 (N_26151,N_23251,N_22952);
and U26152 (N_26152,N_22868,N_23664);
or U26153 (N_26153,N_21564,N_23635);
nor U26154 (N_26154,N_21248,N_21127);
xor U26155 (N_26155,N_23782,N_22842);
nand U26156 (N_26156,N_22020,N_21934);
or U26157 (N_26157,N_21406,N_23633);
or U26158 (N_26158,N_22244,N_23242);
xnor U26159 (N_26159,N_23664,N_21118);
or U26160 (N_26160,N_23598,N_22632);
or U26161 (N_26161,N_21153,N_21143);
nor U26162 (N_26162,N_23208,N_22849);
or U26163 (N_26163,N_21736,N_23279);
or U26164 (N_26164,N_23596,N_22905);
xnor U26165 (N_26165,N_22486,N_21419);
and U26166 (N_26166,N_22299,N_22477);
or U26167 (N_26167,N_22422,N_22400);
nor U26168 (N_26168,N_22193,N_21443);
xor U26169 (N_26169,N_22203,N_23655);
xnor U26170 (N_26170,N_22280,N_21193);
and U26171 (N_26171,N_22485,N_21550);
xor U26172 (N_26172,N_23421,N_23444);
nor U26173 (N_26173,N_22421,N_23519);
nor U26174 (N_26174,N_22367,N_21463);
nand U26175 (N_26175,N_21439,N_21048);
or U26176 (N_26176,N_23836,N_23548);
and U26177 (N_26177,N_22153,N_23987);
nand U26178 (N_26178,N_21403,N_23288);
and U26179 (N_26179,N_22282,N_22416);
and U26180 (N_26180,N_22163,N_23430);
or U26181 (N_26181,N_21593,N_21557);
or U26182 (N_26182,N_21339,N_23259);
or U26183 (N_26183,N_21382,N_23765);
or U26184 (N_26184,N_22440,N_23465);
nand U26185 (N_26185,N_22016,N_23048);
or U26186 (N_26186,N_23000,N_21540);
and U26187 (N_26187,N_22392,N_23022);
or U26188 (N_26188,N_23656,N_21343);
xor U26189 (N_26189,N_22255,N_21908);
nand U26190 (N_26190,N_22920,N_23075);
or U26191 (N_26191,N_23427,N_22303);
nor U26192 (N_26192,N_22438,N_22795);
nor U26193 (N_26193,N_22799,N_23775);
or U26194 (N_26194,N_22879,N_21855);
or U26195 (N_26195,N_21797,N_21571);
or U26196 (N_26196,N_22700,N_23128);
nand U26197 (N_26197,N_23901,N_21434);
xor U26198 (N_26198,N_23099,N_21773);
xnor U26199 (N_26199,N_23366,N_22307);
nor U26200 (N_26200,N_21170,N_23250);
nand U26201 (N_26201,N_22141,N_23210);
xor U26202 (N_26202,N_23758,N_23436);
nand U26203 (N_26203,N_23964,N_22711);
xnor U26204 (N_26204,N_23460,N_22228);
or U26205 (N_26205,N_23957,N_23232);
xor U26206 (N_26206,N_22236,N_23931);
or U26207 (N_26207,N_22604,N_23833);
xor U26208 (N_26208,N_23604,N_21431);
nand U26209 (N_26209,N_23380,N_23700);
or U26210 (N_26210,N_21988,N_22186);
xor U26211 (N_26211,N_22732,N_23911);
or U26212 (N_26212,N_21679,N_23287);
nor U26213 (N_26213,N_22686,N_22595);
nor U26214 (N_26214,N_23945,N_22212);
nor U26215 (N_26215,N_21165,N_23876);
nor U26216 (N_26216,N_23566,N_23610);
xnor U26217 (N_26217,N_23459,N_23091);
nand U26218 (N_26218,N_23053,N_21194);
xor U26219 (N_26219,N_21590,N_23733);
xor U26220 (N_26220,N_23610,N_21729);
or U26221 (N_26221,N_22854,N_21604);
nor U26222 (N_26222,N_23547,N_22615);
nor U26223 (N_26223,N_23465,N_22491);
xnor U26224 (N_26224,N_22958,N_23576);
nand U26225 (N_26225,N_23814,N_21481);
or U26226 (N_26226,N_23197,N_22957);
xor U26227 (N_26227,N_22883,N_21737);
nor U26228 (N_26228,N_21929,N_21855);
nor U26229 (N_26229,N_21495,N_22084);
and U26230 (N_26230,N_21404,N_21897);
nand U26231 (N_26231,N_22985,N_22530);
xor U26232 (N_26232,N_23920,N_23866);
or U26233 (N_26233,N_21550,N_22114);
nor U26234 (N_26234,N_22198,N_21670);
xnor U26235 (N_26235,N_22598,N_21549);
or U26236 (N_26236,N_21268,N_22459);
or U26237 (N_26237,N_21851,N_22249);
nand U26238 (N_26238,N_23105,N_23639);
nand U26239 (N_26239,N_23298,N_22290);
nand U26240 (N_26240,N_22745,N_22448);
or U26241 (N_26241,N_21821,N_22745);
or U26242 (N_26242,N_21756,N_21682);
xor U26243 (N_26243,N_22578,N_21725);
nor U26244 (N_26244,N_22191,N_22157);
nand U26245 (N_26245,N_22028,N_23536);
nand U26246 (N_26246,N_22879,N_22059);
nand U26247 (N_26247,N_21412,N_23464);
nand U26248 (N_26248,N_22051,N_22861);
xnor U26249 (N_26249,N_23906,N_23444);
xor U26250 (N_26250,N_21500,N_23575);
nand U26251 (N_26251,N_23852,N_22194);
and U26252 (N_26252,N_23083,N_21874);
or U26253 (N_26253,N_22101,N_21879);
nor U26254 (N_26254,N_22205,N_23817);
xor U26255 (N_26255,N_22892,N_23573);
or U26256 (N_26256,N_23239,N_21518);
or U26257 (N_26257,N_22049,N_22122);
nor U26258 (N_26258,N_21720,N_23769);
xor U26259 (N_26259,N_22686,N_22620);
nand U26260 (N_26260,N_22763,N_22554);
and U26261 (N_26261,N_23855,N_23994);
nand U26262 (N_26262,N_22206,N_21907);
nor U26263 (N_26263,N_23400,N_23846);
nor U26264 (N_26264,N_23070,N_23225);
and U26265 (N_26265,N_21851,N_21497);
nor U26266 (N_26266,N_23682,N_23577);
and U26267 (N_26267,N_22244,N_23922);
xor U26268 (N_26268,N_23289,N_22164);
or U26269 (N_26269,N_22469,N_23558);
nand U26270 (N_26270,N_22743,N_22278);
nand U26271 (N_26271,N_21302,N_21205);
nor U26272 (N_26272,N_23642,N_22916);
nand U26273 (N_26273,N_21014,N_23757);
xnor U26274 (N_26274,N_23733,N_21871);
and U26275 (N_26275,N_21000,N_21936);
xor U26276 (N_26276,N_23338,N_21847);
nor U26277 (N_26277,N_23467,N_22637);
and U26278 (N_26278,N_23413,N_22228);
or U26279 (N_26279,N_23012,N_23621);
and U26280 (N_26280,N_21038,N_23131);
nor U26281 (N_26281,N_22392,N_23263);
and U26282 (N_26282,N_21967,N_22008);
nor U26283 (N_26283,N_23419,N_23119);
nand U26284 (N_26284,N_23071,N_22481);
nand U26285 (N_26285,N_22732,N_22411);
nor U26286 (N_26286,N_21944,N_22200);
or U26287 (N_26287,N_22746,N_23700);
or U26288 (N_26288,N_21722,N_21675);
nand U26289 (N_26289,N_22109,N_23403);
nor U26290 (N_26290,N_21985,N_22158);
and U26291 (N_26291,N_22345,N_22370);
and U26292 (N_26292,N_21403,N_21183);
xnor U26293 (N_26293,N_23652,N_21134);
nand U26294 (N_26294,N_21394,N_23685);
xor U26295 (N_26295,N_21445,N_23009);
xnor U26296 (N_26296,N_22860,N_21885);
and U26297 (N_26297,N_23560,N_21813);
nand U26298 (N_26298,N_22753,N_21421);
xor U26299 (N_26299,N_22237,N_21999);
nand U26300 (N_26300,N_21230,N_23939);
nand U26301 (N_26301,N_23868,N_21910);
xnor U26302 (N_26302,N_22647,N_21171);
xor U26303 (N_26303,N_21241,N_22242);
nor U26304 (N_26304,N_21143,N_22257);
nand U26305 (N_26305,N_22167,N_23076);
or U26306 (N_26306,N_23508,N_22652);
xnor U26307 (N_26307,N_21303,N_22405);
nor U26308 (N_26308,N_23220,N_21087);
or U26309 (N_26309,N_21535,N_23291);
nor U26310 (N_26310,N_23774,N_22306);
xor U26311 (N_26311,N_23753,N_23347);
nand U26312 (N_26312,N_23354,N_22313);
or U26313 (N_26313,N_21104,N_22382);
nand U26314 (N_26314,N_21369,N_23332);
and U26315 (N_26315,N_22094,N_23989);
nand U26316 (N_26316,N_21510,N_22806);
nand U26317 (N_26317,N_22472,N_22149);
and U26318 (N_26318,N_21906,N_22498);
nand U26319 (N_26319,N_22529,N_21003);
or U26320 (N_26320,N_23879,N_21782);
nand U26321 (N_26321,N_22309,N_21358);
nor U26322 (N_26322,N_21922,N_22887);
and U26323 (N_26323,N_22948,N_21058);
nor U26324 (N_26324,N_21983,N_23415);
nand U26325 (N_26325,N_23816,N_21768);
nand U26326 (N_26326,N_22332,N_22099);
nor U26327 (N_26327,N_21908,N_21032);
nor U26328 (N_26328,N_23985,N_22237);
and U26329 (N_26329,N_23197,N_23715);
or U26330 (N_26330,N_22273,N_23726);
nor U26331 (N_26331,N_22426,N_22390);
or U26332 (N_26332,N_22207,N_22669);
nor U26333 (N_26333,N_22456,N_23572);
or U26334 (N_26334,N_22328,N_21405);
or U26335 (N_26335,N_21374,N_21875);
or U26336 (N_26336,N_22518,N_22105);
or U26337 (N_26337,N_22209,N_23479);
xnor U26338 (N_26338,N_22392,N_23845);
and U26339 (N_26339,N_23598,N_21258);
or U26340 (N_26340,N_23494,N_23191);
nor U26341 (N_26341,N_21339,N_22515);
xnor U26342 (N_26342,N_22206,N_23260);
nand U26343 (N_26343,N_23135,N_23861);
nand U26344 (N_26344,N_23476,N_21477);
nand U26345 (N_26345,N_23870,N_23140);
and U26346 (N_26346,N_21863,N_21663);
xor U26347 (N_26347,N_21198,N_23740);
or U26348 (N_26348,N_22018,N_21751);
nand U26349 (N_26349,N_23297,N_21572);
nor U26350 (N_26350,N_23847,N_23199);
nor U26351 (N_26351,N_22174,N_23680);
and U26352 (N_26352,N_23273,N_21288);
xnor U26353 (N_26353,N_23322,N_23745);
and U26354 (N_26354,N_22877,N_21880);
or U26355 (N_26355,N_21529,N_21615);
xor U26356 (N_26356,N_23278,N_21289);
or U26357 (N_26357,N_23427,N_21746);
xor U26358 (N_26358,N_22309,N_21369);
nor U26359 (N_26359,N_21681,N_23250);
nor U26360 (N_26360,N_21736,N_21527);
nand U26361 (N_26361,N_21340,N_21345);
or U26362 (N_26362,N_22861,N_22521);
nor U26363 (N_26363,N_22291,N_21548);
xnor U26364 (N_26364,N_23446,N_21718);
or U26365 (N_26365,N_23349,N_22264);
nand U26366 (N_26366,N_23008,N_22412);
or U26367 (N_26367,N_21124,N_21650);
nand U26368 (N_26368,N_23128,N_22692);
nor U26369 (N_26369,N_21092,N_22970);
nor U26370 (N_26370,N_21657,N_21454);
nand U26371 (N_26371,N_23339,N_21474);
or U26372 (N_26372,N_21370,N_22313);
xor U26373 (N_26373,N_23128,N_23954);
and U26374 (N_26374,N_21803,N_23335);
or U26375 (N_26375,N_23462,N_23857);
nand U26376 (N_26376,N_22117,N_21005);
or U26377 (N_26377,N_22481,N_23044);
xor U26378 (N_26378,N_22928,N_21518);
nand U26379 (N_26379,N_23543,N_23569);
nor U26380 (N_26380,N_22523,N_23043);
nand U26381 (N_26381,N_23943,N_23257);
or U26382 (N_26382,N_21936,N_23382);
and U26383 (N_26383,N_21758,N_21219);
nor U26384 (N_26384,N_23134,N_21320);
and U26385 (N_26385,N_22415,N_22445);
nor U26386 (N_26386,N_21363,N_23238);
or U26387 (N_26387,N_22064,N_22737);
xnor U26388 (N_26388,N_23067,N_22175);
or U26389 (N_26389,N_22155,N_23770);
nor U26390 (N_26390,N_21984,N_23762);
or U26391 (N_26391,N_23428,N_21824);
nor U26392 (N_26392,N_21451,N_23954);
and U26393 (N_26393,N_21826,N_21806);
nor U26394 (N_26394,N_21765,N_22816);
and U26395 (N_26395,N_21995,N_22910);
xor U26396 (N_26396,N_21035,N_23981);
nand U26397 (N_26397,N_22485,N_21297);
nand U26398 (N_26398,N_21247,N_21971);
and U26399 (N_26399,N_22990,N_21561);
nand U26400 (N_26400,N_23077,N_22419);
and U26401 (N_26401,N_22376,N_22427);
nand U26402 (N_26402,N_22697,N_22067);
nor U26403 (N_26403,N_23179,N_21582);
nand U26404 (N_26404,N_21478,N_22566);
xor U26405 (N_26405,N_21649,N_21769);
nand U26406 (N_26406,N_23279,N_22673);
nor U26407 (N_26407,N_22411,N_23886);
xor U26408 (N_26408,N_21132,N_23153);
and U26409 (N_26409,N_23736,N_23439);
and U26410 (N_26410,N_23186,N_22161);
or U26411 (N_26411,N_23513,N_23823);
and U26412 (N_26412,N_22946,N_22114);
or U26413 (N_26413,N_23737,N_21170);
xor U26414 (N_26414,N_22663,N_23122);
xor U26415 (N_26415,N_21663,N_23613);
nor U26416 (N_26416,N_21906,N_22486);
nand U26417 (N_26417,N_22283,N_23839);
or U26418 (N_26418,N_23274,N_22220);
nor U26419 (N_26419,N_23176,N_21361);
nor U26420 (N_26420,N_21806,N_23877);
nand U26421 (N_26421,N_23367,N_23887);
xor U26422 (N_26422,N_21899,N_23869);
xor U26423 (N_26423,N_21882,N_23499);
nor U26424 (N_26424,N_21595,N_22767);
nor U26425 (N_26425,N_22811,N_22311);
nor U26426 (N_26426,N_23077,N_21281);
nand U26427 (N_26427,N_22548,N_22627);
nand U26428 (N_26428,N_21604,N_21120);
or U26429 (N_26429,N_21098,N_22043);
nor U26430 (N_26430,N_21434,N_23802);
and U26431 (N_26431,N_22787,N_21940);
xnor U26432 (N_26432,N_22957,N_21449);
nand U26433 (N_26433,N_21500,N_21162);
or U26434 (N_26434,N_22121,N_21755);
or U26435 (N_26435,N_23183,N_22072);
or U26436 (N_26436,N_23950,N_21071);
and U26437 (N_26437,N_21178,N_21087);
or U26438 (N_26438,N_23694,N_21263);
or U26439 (N_26439,N_21523,N_22411);
and U26440 (N_26440,N_22107,N_23222);
nand U26441 (N_26441,N_21188,N_21201);
nand U26442 (N_26442,N_21162,N_21564);
nand U26443 (N_26443,N_23729,N_23964);
and U26444 (N_26444,N_22466,N_21847);
and U26445 (N_26445,N_21731,N_21196);
or U26446 (N_26446,N_23158,N_22630);
or U26447 (N_26447,N_22508,N_23763);
xor U26448 (N_26448,N_23870,N_23447);
xnor U26449 (N_26449,N_21943,N_21563);
and U26450 (N_26450,N_23167,N_23482);
or U26451 (N_26451,N_23661,N_22135);
and U26452 (N_26452,N_22161,N_23678);
nand U26453 (N_26453,N_23384,N_21215);
nand U26454 (N_26454,N_21831,N_22299);
and U26455 (N_26455,N_21840,N_21813);
and U26456 (N_26456,N_22714,N_23014);
nand U26457 (N_26457,N_21193,N_23134);
or U26458 (N_26458,N_22044,N_21358);
nand U26459 (N_26459,N_21128,N_23109);
xor U26460 (N_26460,N_23589,N_23928);
or U26461 (N_26461,N_23948,N_23844);
nor U26462 (N_26462,N_21675,N_21073);
nand U26463 (N_26463,N_21043,N_22408);
or U26464 (N_26464,N_23211,N_21051);
nand U26465 (N_26465,N_22244,N_23934);
nand U26466 (N_26466,N_23442,N_23254);
xor U26467 (N_26467,N_23482,N_22395);
or U26468 (N_26468,N_21473,N_23367);
nor U26469 (N_26469,N_21934,N_21519);
and U26470 (N_26470,N_23590,N_23649);
xnor U26471 (N_26471,N_21045,N_21444);
nor U26472 (N_26472,N_23478,N_21539);
xnor U26473 (N_26473,N_22933,N_21973);
nor U26474 (N_26474,N_21113,N_22811);
or U26475 (N_26475,N_21131,N_23703);
or U26476 (N_26476,N_22000,N_21344);
and U26477 (N_26477,N_22630,N_23942);
xnor U26478 (N_26478,N_23036,N_22350);
and U26479 (N_26479,N_23699,N_22729);
and U26480 (N_26480,N_23060,N_22497);
nand U26481 (N_26481,N_23178,N_21303);
or U26482 (N_26482,N_21970,N_23392);
and U26483 (N_26483,N_22856,N_23763);
nor U26484 (N_26484,N_21001,N_23872);
nand U26485 (N_26485,N_22436,N_23315);
nand U26486 (N_26486,N_22377,N_23281);
xnor U26487 (N_26487,N_23709,N_22179);
and U26488 (N_26488,N_23990,N_22825);
and U26489 (N_26489,N_23487,N_21821);
or U26490 (N_26490,N_23802,N_21283);
or U26491 (N_26491,N_21659,N_22712);
xor U26492 (N_26492,N_23874,N_21197);
and U26493 (N_26493,N_22563,N_23103);
nor U26494 (N_26494,N_21812,N_21861);
or U26495 (N_26495,N_22203,N_22597);
nor U26496 (N_26496,N_23788,N_23478);
or U26497 (N_26497,N_21758,N_22775);
nor U26498 (N_26498,N_23426,N_21611);
xnor U26499 (N_26499,N_23560,N_22420);
nor U26500 (N_26500,N_23693,N_23251);
nand U26501 (N_26501,N_21726,N_23940);
nand U26502 (N_26502,N_22782,N_23848);
nand U26503 (N_26503,N_23599,N_23029);
and U26504 (N_26504,N_21973,N_22377);
nand U26505 (N_26505,N_21227,N_23360);
nor U26506 (N_26506,N_23253,N_23440);
xor U26507 (N_26507,N_22553,N_23813);
nor U26508 (N_26508,N_22521,N_23232);
and U26509 (N_26509,N_21548,N_22372);
nand U26510 (N_26510,N_22950,N_22129);
xor U26511 (N_26511,N_22638,N_23711);
nand U26512 (N_26512,N_23099,N_21157);
or U26513 (N_26513,N_23817,N_23028);
nand U26514 (N_26514,N_22378,N_21901);
or U26515 (N_26515,N_21076,N_23603);
and U26516 (N_26516,N_21439,N_21404);
xnor U26517 (N_26517,N_21055,N_21455);
nand U26518 (N_26518,N_21141,N_21264);
nand U26519 (N_26519,N_21871,N_21351);
nand U26520 (N_26520,N_23808,N_21798);
xnor U26521 (N_26521,N_23998,N_21428);
and U26522 (N_26522,N_21452,N_22611);
xnor U26523 (N_26523,N_21059,N_23139);
xnor U26524 (N_26524,N_23739,N_22460);
nor U26525 (N_26525,N_21036,N_21452);
xor U26526 (N_26526,N_23044,N_23708);
or U26527 (N_26527,N_22088,N_23779);
nand U26528 (N_26528,N_22743,N_21044);
nor U26529 (N_26529,N_21707,N_22749);
or U26530 (N_26530,N_22190,N_22736);
and U26531 (N_26531,N_23479,N_22815);
or U26532 (N_26532,N_23820,N_21728);
or U26533 (N_26533,N_23863,N_22720);
and U26534 (N_26534,N_23030,N_22980);
and U26535 (N_26535,N_22184,N_22733);
xor U26536 (N_26536,N_23471,N_23921);
or U26537 (N_26537,N_22289,N_21411);
nor U26538 (N_26538,N_21305,N_23603);
nand U26539 (N_26539,N_23938,N_23847);
and U26540 (N_26540,N_22133,N_21994);
xnor U26541 (N_26541,N_21062,N_23846);
or U26542 (N_26542,N_21513,N_22770);
or U26543 (N_26543,N_22590,N_21235);
nand U26544 (N_26544,N_21899,N_23635);
or U26545 (N_26545,N_22906,N_22705);
xnor U26546 (N_26546,N_22219,N_22976);
nor U26547 (N_26547,N_23450,N_23121);
xor U26548 (N_26548,N_22457,N_21169);
nor U26549 (N_26549,N_21158,N_23233);
nor U26550 (N_26550,N_22810,N_23617);
or U26551 (N_26551,N_23890,N_21612);
and U26552 (N_26552,N_23915,N_22763);
nor U26553 (N_26553,N_23518,N_21520);
xnor U26554 (N_26554,N_22177,N_23161);
and U26555 (N_26555,N_21563,N_21783);
and U26556 (N_26556,N_23805,N_21647);
or U26557 (N_26557,N_23957,N_23716);
or U26558 (N_26558,N_22567,N_22507);
xnor U26559 (N_26559,N_22126,N_22510);
and U26560 (N_26560,N_23051,N_22652);
or U26561 (N_26561,N_21013,N_23301);
xor U26562 (N_26562,N_21625,N_23385);
and U26563 (N_26563,N_21233,N_22194);
or U26564 (N_26564,N_23792,N_22286);
nor U26565 (N_26565,N_21827,N_22446);
nor U26566 (N_26566,N_23030,N_21677);
or U26567 (N_26567,N_22879,N_21962);
and U26568 (N_26568,N_23141,N_22534);
and U26569 (N_26569,N_23445,N_21332);
or U26570 (N_26570,N_22709,N_23890);
or U26571 (N_26571,N_22935,N_23182);
or U26572 (N_26572,N_22146,N_21037);
nand U26573 (N_26573,N_22385,N_21555);
and U26574 (N_26574,N_23570,N_22886);
xnor U26575 (N_26575,N_23822,N_22663);
nor U26576 (N_26576,N_21939,N_21406);
or U26577 (N_26577,N_21856,N_22527);
and U26578 (N_26578,N_21479,N_21960);
xnor U26579 (N_26579,N_21493,N_23298);
nor U26580 (N_26580,N_22645,N_21054);
nand U26581 (N_26581,N_23190,N_23441);
nand U26582 (N_26582,N_23320,N_21889);
or U26583 (N_26583,N_21099,N_22489);
xor U26584 (N_26584,N_23783,N_23747);
nand U26585 (N_26585,N_23102,N_22409);
nor U26586 (N_26586,N_23975,N_22367);
or U26587 (N_26587,N_22484,N_21628);
or U26588 (N_26588,N_22605,N_23449);
xor U26589 (N_26589,N_22844,N_23274);
or U26590 (N_26590,N_22711,N_21071);
and U26591 (N_26591,N_23208,N_21884);
and U26592 (N_26592,N_22472,N_21878);
nor U26593 (N_26593,N_22540,N_21587);
or U26594 (N_26594,N_23425,N_23262);
or U26595 (N_26595,N_22166,N_23567);
nand U26596 (N_26596,N_21297,N_22988);
nor U26597 (N_26597,N_22181,N_21708);
and U26598 (N_26598,N_21289,N_23086);
nand U26599 (N_26599,N_21191,N_21992);
nand U26600 (N_26600,N_21857,N_21951);
xnor U26601 (N_26601,N_22984,N_22009);
or U26602 (N_26602,N_22004,N_21164);
and U26603 (N_26603,N_23486,N_23985);
xnor U26604 (N_26604,N_23310,N_22427);
or U26605 (N_26605,N_23288,N_21147);
or U26606 (N_26606,N_21551,N_21211);
xnor U26607 (N_26607,N_23364,N_21231);
xor U26608 (N_26608,N_22131,N_22350);
nor U26609 (N_26609,N_23397,N_21727);
or U26610 (N_26610,N_23394,N_22234);
and U26611 (N_26611,N_23993,N_23665);
xnor U26612 (N_26612,N_22601,N_21557);
nor U26613 (N_26613,N_21317,N_21828);
and U26614 (N_26614,N_22951,N_23707);
xnor U26615 (N_26615,N_23820,N_23747);
nand U26616 (N_26616,N_21153,N_21053);
xnor U26617 (N_26617,N_22602,N_21770);
or U26618 (N_26618,N_23326,N_21695);
nor U26619 (N_26619,N_22356,N_22401);
xnor U26620 (N_26620,N_22936,N_23443);
and U26621 (N_26621,N_22308,N_21446);
and U26622 (N_26622,N_22750,N_22516);
nand U26623 (N_26623,N_22985,N_23802);
nor U26624 (N_26624,N_22421,N_21676);
xor U26625 (N_26625,N_21499,N_22198);
nor U26626 (N_26626,N_21878,N_21758);
and U26627 (N_26627,N_21297,N_21656);
and U26628 (N_26628,N_21029,N_22653);
nor U26629 (N_26629,N_23831,N_23367);
and U26630 (N_26630,N_21691,N_22614);
and U26631 (N_26631,N_21886,N_23283);
or U26632 (N_26632,N_23309,N_23553);
and U26633 (N_26633,N_21468,N_22669);
and U26634 (N_26634,N_21509,N_22979);
and U26635 (N_26635,N_22389,N_21775);
nand U26636 (N_26636,N_22813,N_22736);
and U26637 (N_26637,N_23057,N_21299);
and U26638 (N_26638,N_21818,N_22808);
xnor U26639 (N_26639,N_23546,N_23519);
nand U26640 (N_26640,N_23488,N_21222);
xor U26641 (N_26641,N_21128,N_23083);
xor U26642 (N_26642,N_23871,N_22669);
nand U26643 (N_26643,N_21431,N_21201);
xnor U26644 (N_26644,N_21273,N_23473);
or U26645 (N_26645,N_23886,N_21751);
nand U26646 (N_26646,N_21022,N_23087);
xor U26647 (N_26647,N_21105,N_21220);
and U26648 (N_26648,N_22476,N_23228);
and U26649 (N_26649,N_21742,N_21555);
nor U26650 (N_26650,N_22048,N_21418);
and U26651 (N_26651,N_23728,N_21648);
or U26652 (N_26652,N_21926,N_22204);
xnor U26653 (N_26653,N_21861,N_21934);
nand U26654 (N_26654,N_23920,N_22767);
or U26655 (N_26655,N_21108,N_23664);
nand U26656 (N_26656,N_22499,N_22514);
nand U26657 (N_26657,N_23248,N_23241);
xnor U26658 (N_26658,N_22256,N_23855);
nand U26659 (N_26659,N_23388,N_22476);
or U26660 (N_26660,N_22312,N_21914);
or U26661 (N_26661,N_22081,N_22305);
and U26662 (N_26662,N_21851,N_22667);
xnor U26663 (N_26663,N_21279,N_22455);
nor U26664 (N_26664,N_22756,N_21384);
nor U26665 (N_26665,N_21820,N_21423);
xor U26666 (N_26666,N_23842,N_21103);
nor U26667 (N_26667,N_21447,N_22056);
xnor U26668 (N_26668,N_21895,N_22551);
and U26669 (N_26669,N_21185,N_23317);
and U26670 (N_26670,N_21092,N_23444);
nor U26671 (N_26671,N_21632,N_22685);
or U26672 (N_26672,N_22733,N_22838);
xor U26673 (N_26673,N_23185,N_22905);
nand U26674 (N_26674,N_22365,N_23168);
nand U26675 (N_26675,N_21428,N_22302);
and U26676 (N_26676,N_23273,N_23896);
nor U26677 (N_26677,N_22845,N_23827);
or U26678 (N_26678,N_22087,N_21302);
xor U26679 (N_26679,N_21171,N_22788);
nand U26680 (N_26680,N_22536,N_21890);
or U26681 (N_26681,N_22692,N_23363);
xor U26682 (N_26682,N_21804,N_22980);
or U26683 (N_26683,N_22476,N_22195);
and U26684 (N_26684,N_22985,N_21059);
or U26685 (N_26685,N_22885,N_21315);
xnor U26686 (N_26686,N_22460,N_22271);
nor U26687 (N_26687,N_21511,N_23941);
or U26688 (N_26688,N_23988,N_23608);
nor U26689 (N_26689,N_21962,N_22747);
nand U26690 (N_26690,N_22057,N_22043);
nor U26691 (N_26691,N_21230,N_22315);
or U26692 (N_26692,N_23610,N_23425);
or U26693 (N_26693,N_22963,N_22852);
xor U26694 (N_26694,N_21089,N_21299);
and U26695 (N_26695,N_22934,N_23098);
xnor U26696 (N_26696,N_21433,N_23775);
nand U26697 (N_26697,N_22784,N_23158);
nor U26698 (N_26698,N_21325,N_22537);
nor U26699 (N_26699,N_21847,N_21916);
nand U26700 (N_26700,N_23170,N_23368);
nand U26701 (N_26701,N_22553,N_21182);
nand U26702 (N_26702,N_22552,N_21357);
nand U26703 (N_26703,N_21521,N_21744);
nor U26704 (N_26704,N_23667,N_22476);
nor U26705 (N_26705,N_23251,N_22589);
nand U26706 (N_26706,N_22010,N_22228);
nor U26707 (N_26707,N_23448,N_21765);
nand U26708 (N_26708,N_21682,N_23931);
nor U26709 (N_26709,N_23149,N_21887);
nand U26710 (N_26710,N_21378,N_21117);
and U26711 (N_26711,N_21149,N_23764);
nand U26712 (N_26712,N_23933,N_22336);
or U26713 (N_26713,N_21772,N_23789);
or U26714 (N_26714,N_23421,N_23954);
and U26715 (N_26715,N_23601,N_22890);
and U26716 (N_26716,N_21008,N_21887);
nand U26717 (N_26717,N_21829,N_23557);
nor U26718 (N_26718,N_23525,N_22757);
or U26719 (N_26719,N_22714,N_23783);
xnor U26720 (N_26720,N_22454,N_22925);
xor U26721 (N_26721,N_21267,N_21986);
nand U26722 (N_26722,N_22141,N_23570);
or U26723 (N_26723,N_23859,N_23216);
nand U26724 (N_26724,N_22413,N_22104);
and U26725 (N_26725,N_22484,N_22894);
and U26726 (N_26726,N_23965,N_22575);
nand U26727 (N_26727,N_21628,N_22318);
and U26728 (N_26728,N_22237,N_23863);
xnor U26729 (N_26729,N_22904,N_23280);
and U26730 (N_26730,N_22013,N_22821);
nand U26731 (N_26731,N_22897,N_21321);
or U26732 (N_26732,N_22604,N_23140);
and U26733 (N_26733,N_21486,N_23787);
xnor U26734 (N_26734,N_22361,N_22846);
xnor U26735 (N_26735,N_21542,N_23847);
and U26736 (N_26736,N_21673,N_21836);
nand U26737 (N_26737,N_21047,N_23261);
nand U26738 (N_26738,N_22271,N_22468);
and U26739 (N_26739,N_22151,N_23715);
nor U26740 (N_26740,N_22546,N_21424);
or U26741 (N_26741,N_23529,N_23304);
nand U26742 (N_26742,N_21824,N_21280);
or U26743 (N_26743,N_22169,N_23360);
nor U26744 (N_26744,N_23504,N_21955);
xor U26745 (N_26745,N_23626,N_23781);
or U26746 (N_26746,N_22197,N_23303);
or U26747 (N_26747,N_23250,N_21811);
nor U26748 (N_26748,N_21632,N_22070);
or U26749 (N_26749,N_21305,N_22463);
nand U26750 (N_26750,N_22157,N_21029);
nor U26751 (N_26751,N_22215,N_23228);
xor U26752 (N_26752,N_23096,N_22825);
and U26753 (N_26753,N_22578,N_22437);
xnor U26754 (N_26754,N_21363,N_21656);
and U26755 (N_26755,N_21282,N_23347);
nand U26756 (N_26756,N_21736,N_22267);
and U26757 (N_26757,N_22790,N_23313);
nor U26758 (N_26758,N_22544,N_21812);
nor U26759 (N_26759,N_21510,N_23379);
or U26760 (N_26760,N_21642,N_22308);
or U26761 (N_26761,N_21408,N_22637);
and U26762 (N_26762,N_22982,N_22707);
or U26763 (N_26763,N_21623,N_21747);
nor U26764 (N_26764,N_22266,N_23280);
nand U26765 (N_26765,N_22186,N_23879);
and U26766 (N_26766,N_22877,N_21440);
nand U26767 (N_26767,N_22498,N_22726);
nand U26768 (N_26768,N_23214,N_22869);
nor U26769 (N_26769,N_22222,N_23919);
and U26770 (N_26770,N_22576,N_23857);
or U26771 (N_26771,N_21747,N_21853);
nand U26772 (N_26772,N_23758,N_22313);
nor U26773 (N_26773,N_23426,N_21300);
nand U26774 (N_26774,N_22151,N_22538);
and U26775 (N_26775,N_22752,N_21119);
nand U26776 (N_26776,N_23556,N_23367);
or U26777 (N_26777,N_22385,N_22988);
or U26778 (N_26778,N_22398,N_21676);
xor U26779 (N_26779,N_21768,N_21302);
and U26780 (N_26780,N_22780,N_23844);
and U26781 (N_26781,N_22913,N_21988);
nand U26782 (N_26782,N_23958,N_22721);
and U26783 (N_26783,N_21785,N_22045);
nor U26784 (N_26784,N_23996,N_22121);
and U26785 (N_26785,N_22916,N_21026);
and U26786 (N_26786,N_21602,N_23294);
xnor U26787 (N_26787,N_23104,N_21549);
xnor U26788 (N_26788,N_23373,N_21135);
or U26789 (N_26789,N_21886,N_22081);
xor U26790 (N_26790,N_23116,N_22368);
or U26791 (N_26791,N_23991,N_23424);
nand U26792 (N_26792,N_22425,N_21869);
nand U26793 (N_26793,N_23290,N_23898);
nand U26794 (N_26794,N_23667,N_21854);
or U26795 (N_26795,N_22486,N_23580);
or U26796 (N_26796,N_22471,N_22530);
or U26797 (N_26797,N_23300,N_23428);
nor U26798 (N_26798,N_21237,N_22095);
or U26799 (N_26799,N_22637,N_21528);
or U26800 (N_26800,N_22040,N_22104);
or U26801 (N_26801,N_21488,N_23181);
and U26802 (N_26802,N_22036,N_22730);
nor U26803 (N_26803,N_23755,N_21121);
nor U26804 (N_26804,N_22337,N_23444);
xor U26805 (N_26805,N_22434,N_21693);
or U26806 (N_26806,N_23263,N_21366);
or U26807 (N_26807,N_22410,N_22373);
xnor U26808 (N_26808,N_22505,N_23286);
nand U26809 (N_26809,N_23228,N_23776);
or U26810 (N_26810,N_22070,N_23045);
nand U26811 (N_26811,N_23561,N_22891);
nor U26812 (N_26812,N_22244,N_21253);
or U26813 (N_26813,N_21537,N_21916);
and U26814 (N_26814,N_23903,N_23409);
and U26815 (N_26815,N_23243,N_22143);
xnor U26816 (N_26816,N_21386,N_22807);
nor U26817 (N_26817,N_23326,N_22952);
or U26818 (N_26818,N_21455,N_21940);
nand U26819 (N_26819,N_21408,N_23928);
xnor U26820 (N_26820,N_23439,N_23608);
and U26821 (N_26821,N_23809,N_23014);
or U26822 (N_26822,N_23960,N_22205);
xor U26823 (N_26823,N_22072,N_21988);
xor U26824 (N_26824,N_22320,N_22942);
and U26825 (N_26825,N_21417,N_21679);
nand U26826 (N_26826,N_21319,N_23931);
xnor U26827 (N_26827,N_22934,N_23911);
xor U26828 (N_26828,N_22706,N_22041);
or U26829 (N_26829,N_21718,N_22398);
and U26830 (N_26830,N_21030,N_21905);
nor U26831 (N_26831,N_22888,N_23665);
xor U26832 (N_26832,N_22029,N_21687);
or U26833 (N_26833,N_21598,N_23156);
nor U26834 (N_26834,N_22926,N_21046);
and U26835 (N_26835,N_22015,N_23550);
xor U26836 (N_26836,N_23703,N_21700);
nand U26837 (N_26837,N_22932,N_22527);
and U26838 (N_26838,N_22839,N_22286);
nor U26839 (N_26839,N_23670,N_22017);
nand U26840 (N_26840,N_22099,N_21238);
and U26841 (N_26841,N_21765,N_23165);
nor U26842 (N_26842,N_22278,N_23949);
and U26843 (N_26843,N_22668,N_21074);
nand U26844 (N_26844,N_22947,N_22593);
nor U26845 (N_26845,N_21274,N_21618);
nand U26846 (N_26846,N_21971,N_22235);
nand U26847 (N_26847,N_23360,N_23254);
nor U26848 (N_26848,N_22757,N_22138);
nor U26849 (N_26849,N_21619,N_23614);
xnor U26850 (N_26850,N_21395,N_22708);
nor U26851 (N_26851,N_22224,N_21815);
xnor U26852 (N_26852,N_22684,N_21920);
xnor U26853 (N_26853,N_22162,N_23015);
and U26854 (N_26854,N_22168,N_21370);
or U26855 (N_26855,N_21590,N_22235);
xnor U26856 (N_26856,N_23577,N_22383);
xor U26857 (N_26857,N_21044,N_23826);
nor U26858 (N_26858,N_22825,N_22508);
xor U26859 (N_26859,N_23571,N_23392);
and U26860 (N_26860,N_23458,N_22758);
nand U26861 (N_26861,N_21207,N_22222);
or U26862 (N_26862,N_21871,N_23918);
or U26863 (N_26863,N_21814,N_21965);
nand U26864 (N_26864,N_22659,N_23744);
or U26865 (N_26865,N_21460,N_23698);
xnor U26866 (N_26866,N_22936,N_22271);
nor U26867 (N_26867,N_23792,N_22158);
or U26868 (N_26868,N_23757,N_22944);
and U26869 (N_26869,N_23007,N_21475);
xnor U26870 (N_26870,N_21510,N_23851);
or U26871 (N_26871,N_22961,N_23720);
or U26872 (N_26872,N_23058,N_23285);
nand U26873 (N_26873,N_21075,N_22919);
nand U26874 (N_26874,N_22812,N_21207);
nand U26875 (N_26875,N_23864,N_21503);
or U26876 (N_26876,N_22189,N_21676);
nand U26877 (N_26877,N_23616,N_23672);
xnor U26878 (N_26878,N_22010,N_22106);
or U26879 (N_26879,N_23275,N_22815);
nor U26880 (N_26880,N_21807,N_23231);
nor U26881 (N_26881,N_23781,N_23431);
or U26882 (N_26882,N_22757,N_21331);
or U26883 (N_26883,N_21722,N_21036);
nor U26884 (N_26884,N_23321,N_22464);
xnor U26885 (N_26885,N_23391,N_21560);
or U26886 (N_26886,N_21008,N_22946);
xnor U26887 (N_26887,N_22216,N_21733);
and U26888 (N_26888,N_22823,N_23176);
or U26889 (N_26889,N_21109,N_23341);
xor U26890 (N_26890,N_21560,N_23865);
or U26891 (N_26891,N_22702,N_23602);
and U26892 (N_26892,N_23131,N_23653);
nand U26893 (N_26893,N_21783,N_23951);
nand U26894 (N_26894,N_21534,N_21448);
or U26895 (N_26895,N_22526,N_23026);
nor U26896 (N_26896,N_21168,N_21224);
xor U26897 (N_26897,N_21637,N_21758);
and U26898 (N_26898,N_23305,N_22135);
nor U26899 (N_26899,N_22731,N_22676);
nor U26900 (N_26900,N_21471,N_23480);
nand U26901 (N_26901,N_23472,N_22614);
nor U26902 (N_26902,N_22844,N_22938);
xor U26903 (N_26903,N_22455,N_23586);
nor U26904 (N_26904,N_22478,N_21394);
or U26905 (N_26905,N_23199,N_21818);
xnor U26906 (N_26906,N_23628,N_21986);
or U26907 (N_26907,N_22255,N_21838);
xnor U26908 (N_26908,N_21637,N_22655);
nand U26909 (N_26909,N_23713,N_22042);
nor U26910 (N_26910,N_22759,N_21920);
nor U26911 (N_26911,N_22745,N_23341);
or U26912 (N_26912,N_23143,N_23076);
and U26913 (N_26913,N_21143,N_23614);
nor U26914 (N_26914,N_21242,N_21253);
nand U26915 (N_26915,N_21682,N_22612);
xor U26916 (N_26916,N_22784,N_21677);
nand U26917 (N_26917,N_21488,N_21876);
nor U26918 (N_26918,N_22008,N_22974);
nand U26919 (N_26919,N_21305,N_22992);
nand U26920 (N_26920,N_21503,N_22602);
and U26921 (N_26921,N_23365,N_23475);
nand U26922 (N_26922,N_23025,N_21492);
or U26923 (N_26923,N_21846,N_22535);
nand U26924 (N_26924,N_21817,N_23481);
xnor U26925 (N_26925,N_23955,N_22541);
nand U26926 (N_26926,N_21359,N_23040);
or U26927 (N_26927,N_21107,N_23076);
xor U26928 (N_26928,N_21173,N_22742);
or U26929 (N_26929,N_21087,N_23504);
nand U26930 (N_26930,N_21374,N_23034);
and U26931 (N_26931,N_21603,N_21602);
and U26932 (N_26932,N_21134,N_23609);
and U26933 (N_26933,N_23757,N_23984);
xor U26934 (N_26934,N_23329,N_22268);
and U26935 (N_26935,N_23086,N_21310);
and U26936 (N_26936,N_23924,N_23711);
and U26937 (N_26937,N_21181,N_22837);
nand U26938 (N_26938,N_21230,N_22932);
nor U26939 (N_26939,N_22330,N_23893);
or U26940 (N_26940,N_23786,N_23788);
nor U26941 (N_26941,N_23066,N_21922);
and U26942 (N_26942,N_23934,N_23105);
xor U26943 (N_26943,N_23479,N_23326);
nor U26944 (N_26944,N_21974,N_23417);
nand U26945 (N_26945,N_22407,N_22144);
and U26946 (N_26946,N_22727,N_23012);
xnor U26947 (N_26947,N_23499,N_23455);
or U26948 (N_26948,N_23377,N_23559);
and U26949 (N_26949,N_22781,N_21157);
nand U26950 (N_26950,N_22543,N_23599);
and U26951 (N_26951,N_23072,N_22526);
nor U26952 (N_26952,N_21833,N_22138);
nor U26953 (N_26953,N_22195,N_23076);
nand U26954 (N_26954,N_23040,N_22747);
nor U26955 (N_26955,N_23289,N_22956);
xnor U26956 (N_26956,N_22170,N_22317);
nand U26957 (N_26957,N_21905,N_23948);
nor U26958 (N_26958,N_23551,N_23933);
or U26959 (N_26959,N_22598,N_22449);
xnor U26960 (N_26960,N_22618,N_23959);
or U26961 (N_26961,N_22164,N_22679);
nor U26962 (N_26962,N_21284,N_23883);
or U26963 (N_26963,N_21540,N_22245);
or U26964 (N_26964,N_22895,N_22884);
nor U26965 (N_26965,N_21424,N_22021);
xnor U26966 (N_26966,N_21009,N_21896);
or U26967 (N_26967,N_21220,N_21610);
xnor U26968 (N_26968,N_22341,N_23442);
or U26969 (N_26969,N_23928,N_23031);
nand U26970 (N_26970,N_22465,N_22784);
and U26971 (N_26971,N_22958,N_23509);
nor U26972 (N_26972,N_21029,N_22312);
nand U26973 (N_26973,N_23178,N_22124);
xor U26974 (N_26974,N_23662,N_23617);
xnor U26975 (N_26975,N_21854,N_23124);
or U26976 (N_26976,N_22764,N_22390);
xnor U26977 (N_26977,N_22899,N_21788);
or U26978 (N_26978,N_22897,N_21625);
and U26979 (N_26979,N_23138,N_21336);
nand U26980 (N_26980,N_21125,N_23186);
nor U26981 (N_26981,N_22079,N_23009);
or U26982 (N_26982,N_23538,N_22278);
or U26983 (N_26983,N_21460,N_22003);
and U26984 (N_26984,N_23088,N_21610);
nor U26985 (N_26985,N_23796,N_21829);
nand U26986 (N_26986,N_23976,N_21985);
nand U26987 (N_26987,N_22532,N_22533);
or U26988 (N_26988,N_23734,N_21498);
xnor U26989 (N_26989,N_22692,N_23224);
and U26990 (N_26990,N_21292,N_22045);
nand U26991 (N_26991,N_23984,N_21872);
xnor U26992 (N_26992,N_23267,N_23044);
xnor U26993 (N_26993,N_23453,N_23009);
xnor U26994 (N_26994,N_22918,N_22131);
nor U26995 (N_26995,N_22095,N_22990);
and U26996 (N_26996,N_21565,N_23071);
nand U26997 (N_26997,N_22289,N_21421);
nor U26998 (N_26998,N_22020,N_21135);
and U26999 (N_26999,N_22611,N_21740);
and U27000 (N_27000,N_24542,N_24499);
and U27001 (N_27001,N_24620,N_26017);
and U27002 (N_27002,N_26129,N_25285);
xor U27003 (N_27003,N_26839,N_26429);
or U27004 (N_27004,N_26148,N_25834);
xnor U27005 (N_27005,N_26569,N_25944);
and U27006 (N_27006,N_26145,N_25626);
xor U27007 (N_27007,N_26547,N_24365);
nor U27008 (N_27008,N_26557,N_26906);
nor U27009 (N_27009,N_26920,N_26486);
nand U27010 (N_27010,N_24064,N_26771);
nor U27011 (N_27011,N_26413,N_25686);
and U27012 (N_27012,N_25935,N_25102);
nand U27013 (N_27013,N_25151,N_25144);
nand U27014 (N_27014,N_25128,N_25331);
or U27015 (N_27015,N_24356,N_24908);
xnor U27016 (N_27016,N_24801,N_24077);
nor U27017 (N_27017,N_26855,N_26253);
nor U27018 (N_27018,N_25130,N_25039);
nand U27019 (N_27019,N_26312,N_26690);
or U27020 (N_27020,N_26924,N_25399);
nor U27021 (N_27021,N_25545,N_24661);
xnor U27022 (N_27022,N_25550,N_25630);
and U27023 (N_27023,N_26386,N_25057);
or U27024 (N_27024,N_25607,N_24385);
and U27025 (N_27025,N_24872,N_26729);
and U27026 (N_27026,N_24191,N_24979);
nand U27027 (N_27027,N_26764,N_25249);
or U27028 (N_27028,N_25147,N_26317);
and U27029 (N_27029,N_26914,N_24183);
or U27030 (N_27030,N_24949,N_25354);
or U27031 (N_27031,N_25581,N_25235);
nor U27032 (N_27032,N_24472,N_25127);
or U27033 (N_27033,N_25802,N_25831);
nand U27034 (N_27034,N_24273,N_24474);
nand U27035 (N_27035,N_26388,N_25899);
or U27036 (N_27036,N_26096,N_26268);
nor U27037 (N_27037,N_25692,N_25044);
or U27038 (N_27038,N_25906,N_25685);
xor U27039 (N_27039,N_26768,N_26738);
and U27040 (N_27040,N_26825,N_24337);
or U27041 (N_27041,N_25483,N_25111);
or U27042 (N_27042,N_25073,N_24343);
and U27043 (N_27043,N_25972,N_26634);
xnor U27044 (N_27044,N_25827,N_26907);
nor U27045 (N_27045,N_24274,N_25306);
or U27046 (N_27046,N_24126,N_24044);
and U27047 (N_27047,N_25442,N_25293);
and U27048 (N_27048,N_25311,N_26524);
and U27049 (N_27049,N_25360,N_24798);
xor U27050 (N_27050,N_26435,N_24732);
xnor U27051 (N_27051,N_25245,N_26896);
or U27052 (N_27052,N_25560,N_25475);
nand U27053 (N_27053,N_25992,N_26337);
or U27054 (N_27054,N_26610,N_25003);
or U27055 (N_27055,N_25749,N_24362);
or U27056 (N_27056,N_26329,N_25782);
or U27057 (N_27057,N_25759,N_25175);
nor U27058 (N_27058,N_25850,N_26284);
nor U27059 (N_27059,N_26490,N_25923);
and U27060 (N_27060,N_24649,N_25845);
xor U27061 (N_27061,N_25417,N_26482);
nor U27062 (N_27062,N_24617,N_26876);
xor U27063 (N_27063,N_26058,N_25933);
or U27064 (N_27064,N_24079,N_26628);
nand U27065 (N_27065,N_25366,N_26892);
nand U27066 (N_27066,N_24935,N_26846);
nor U27067 (N_27067,N_24958,N_26843);
nand U27068 (N_27068,N_25484,N_26326);
or U27069 (N_27069,N_25148,N_24639);
and U27070 (N_27070,N_24648,N_25884);
or U27071 (N_27071,N_24111,N_25324);
and U27072 (N_27072,N_24293,N_24720);
nor U27073 (N_27073,N_24626,N_25321);
xnor U27074 (N_27074,N_26452,N_26278);
nor U27075 (N_27075,N_25784,N_24058);
and U27076 (N_27076,N_25317,N_25573);
nand U27077 (N_27077,N_24084,N_25721);
or U27078 (N_27078,N_26277,N_25490);
or U27079 (N_27079,N_26471,N_25553);
nor U27080 (N_27080,N_26689,N_25722);
nand U27081 (N_27081,N_24432,N_25453);
or U27082 (N_27082,N_26667,N_26020);
nand U27083 (N_27083,N_25520,N_25726);
or U27084 (N_27084,N_25569,N_26643);
nand U27085 (N_27085,N_24063,N_24262);
nand U27086 (N_27086,N_24242,N_25835);
xor U27087 (N_27087,N_26320,N_25281);
nor U27088 (N_27088,N_25514,N_25267);
or U27089 (N_27089,N_25880,N_26402);
nor U27090 (N_27090,N_24226,N_25107);
xnor U27091 (N_27091,N_24896,N_26179);
or U27092 (N_27092,N_24690,N_25555);
xnor U27093 (N_27093,N_25392,N_26727);
nand U27094 (N_27094,N_25305,N_26731);
or U27095 (N_27095,N_24139,N_25903);
or U27096 (N_27096,N_26522,N_25762);
and U27097 (N_27097,N_24651,N_26872);
or U27098 (N_27098,N_25084,N_24995);
and U27099 (N_27099,N_24934,N_25589);
or U27100 (N_27100,N_24937,N_25499);
nor U27101 (N_27101,N_24818,N_25866);
xnor U27102 (N_27102,N_24445,N_24624);
xor U27103 (N_27103,N_24714,N_26543);
xnor U27104 (N_27104,N_25382,N_24718);
xor U27105 (N_27105,N_24227,N_26897);
nand U27106 (N_27106,N_24839,N_26871);
and U27107 (N_27107,N_25604,N_24879);
nor U27108 (N_27108,N_25590,N_25715);
nand U27109 (N_27109,N_24590,N_24909);
xor U27110 (N_27110,N_24860,N_26963);
or U27111 (N_27111,N_25415,N_26696);
xor U27112 (N_27112,N_26883,N_24660);
and U27113 (N_27113,N_26523,N_24820);
xnor U27114 (N_27114,N_24278,N_24987);
or U27115 (N_27115,N_24291,N_24476);
or U27116 (N_27116,N_25945,N_26874);
and U27117 (N_27117,N_26160,N_26588);
nand U27118 (N_27118,N_26292,N_25074);
or U27119 (N_27119,N_26219,N_25250);
or U27120 (N_27120,N_25450,N_26507);
nand U27121 (N_27121,N_26712,N_25817);
nand U27122 (N_27122,N_24912,N_25928);
xnor U27123 (N_27123,N_25800,N_24730);
xor U27124 (N_27124,N_25004,N_26308);
or U27125 (N_27125,N_25952,N_25606);
nor U27126 (N_27126,N_25342,N_26080);
nor U27127 (N_27127,N_26021,N_26010);
nor U27128 (N_27128,N_24192,N_25209);
nor U27129 (N_27129,N_25428,N_25507);
or U27130 (N_27130,N_24880,N_25385);
xnor U27131 (N_27131,N_25363,N_26181);
nand U27132 (N_27132,N_25007,N_24994);
and U27133 (N_27133,N_24026,N_24706);
or U27134 (N_27134,N_26953,N_24536);
xnor U27135 (N_27135,N_26314,N_25167);
xnor U27136 (N_27136,N_26587,N_24727);
and U27137 (N_27137,N_26755,N_24859);
or U27138 (N_27138,N_24329,N_26197);
nor U27139 (N_27139,N_26614,N_25296);
or U27140 (N_27140,N_24037,N_24414);
xnor U27141 (N_27141,N_24986,N_26745);
or U27142 (N_27142,N_26209,N_25008);
xor U27143 (N_27143,N_24376,N_26296);
nand U27144 (N_27144,N_24253,N_24216);
nor U27145 (N_27145,N_25830,N_24409);
or U27146 (N_27146,N_26552,N_26695);
or U27147 (N_27147,N_24157,N_26321);
nor U27148 (N_27148,N_26147,N_26332);
or U27149 (N_27149,N_25271,N_24106);
nand U27150 (N_27150,N_26791,N_24604);
and U27151 (N_27151,N_26662,N_24245);
xor U27152 (N_27152,N_25467,N_26997);
and U27153 (N_27153,N_26974,N_26918);
xor U27154 (N_27154,N_26477,N_26468);
nand U27155 (N_27155,N_24777,N_25913);
or U27156 (N_27156,N_25395,N_24711);
nor U27157 (N_27157,N_25757,N_25705);
nor U27158 (N_27158,N_26378,N_25885);
nand U27159 (N_27159,N_24892,N_26844);
nand U27160 (N_27160,N_25254,N_24688);
xnor U27161 (N_27161,N_24076,N_24311);
xor U27162 (N_27162,N_25423,N_24004);
xor U27163 (N_27163,N_25896,N_25414);
or U27164 (N_27164,N_24315,N_26748);
nor U27165 (N_27165,N_24121,N_25904);
and U27166 (N_27166,N_26707,N_25977);
nand U27167 (N_27167,N_25954,N_24665);
xor U27168 (N_27168,N_25124,N_24965);
nor U27169 (N_27169,N_26813,N_25825);
and U27170 (N_27170,N_26891,N_25709);
and U27171 (N_27171,N_24533,N_26701);
xnor U27172 (N_27172,N_26367,N_26819);
or U27173 (N_27173,N_25248,N_24712);
nand U27174 (N_27174,N_24047,N_25469);
nor U27175 (N_27175,N_24259,N_26315);
xnor U27176 (N_27176,N_24486,N_24438);
xor U27177 (N_27177,N_24940,N_24426);
nor U27178 (N_27178,N_24043,N_25289);
xor U27179 (N_27179,N_25698,N_25905);
xor U27180 (N_27180,N_24941,N_25165);
nor U27181 (N_27181,N_24155,N_25265);
nor U27182 (N_27182,N_26105,N_24846);
and U27183 (N_27183,N_25822,N_24007);
nand U27184 (N_27184,N_24855,N_25302);
nand U27185 (N_27185,N_26014,N_24478);
and U27186 (N_27186,N_24538,N_26608);
nor U27187 (N_27187,N_26306,N_25857);
nor U27188 (N_27188,N_25451,N_25040);
nor U27189 (N_27189,N_24930,N_25205);
nand U27190 (N_27190,N_26762,N_26788);
nand U27191 (N_27191,N_24381,N_24924);
or U27192 (N_27192,N_24557,N_25925);
or U27193 (N_27193,N_24147,N_24372);
or U27194 (N_27194,N_24049,N_25194);
or U27195 (N_27195,N_26808,N_26538);
nand U27196 (N_27196,N_25159,N_24917);
nor U27197 (N_27197,N_25595,N_24596);
nor U27198 (N_27198,N_26946,N_25878);
and U27199 (N_27199,N_25547,N_25063);
nor U27200 (N_27200,N_24593,N_25129);
or U27201 (N_27201,N_24821,N_25751);
nand U27202 (N_27202,N_26840,N_24124);
nor U27203 (N_27203,N_26514,N_25276);
or U27204 (N_27204,N_25110,N_24387);
or U27205 (N_27205,N_26101,N_26816);
nor U27206 (N_27206,N_24320,N_25892);
and U27207 (N_27207,N_26900,N_26463);
nor U27208 (N_27208,N_25558,N_24889);
nand U27209 (N_27209,N_24401,N_24375);
xor U27210 (N_27210,N_24524,N_24422);
and U27211 (N_27211,N_24104,N_24899);
and U27212 (N_27212,N_24333,N_25051);
nand U27213 (N_27213,N_24150,N_24276);
xnor U27214 (N_27214,N_24922,N_24440);
or U27215 (N_27215,N_26870,N_25731);
nand U27216 (N_27216,N_24747,N_25523);
or U27217 (N_27217,N_24360,N_25234);
nand U27218 (N_27218,N_25199,N_25663);
nand U27219 (N_27219,N_25023,N_24645);
nor U27220 (N_27220,N_26940,N_25844);
and U27221 (N_27221,N_25990,N_26602);
and U27222 (N_27222,N_26051,N_24471);
nand U27223 (N_27223,N_25037,N_25656);
nand U27224 (N_27224,N_25020,N_26409);
and U27225 (N_27225,N_25158,N_25678);
nor U27226 (N_27226,N_25410,N_26563);
and U27227 (N_27227,N_24662,N_25744);
and U27228 (N_27228,N_26678,N_24161);
xnor U27229 (N_27229,N_26687,N_26991);
xor U27230 (N_27230,N_26323,N_26998);
nand U27231 (N_27231,N_26521,N_26030);
nand U27232 (N_27232,N_24769,N_26747);
nor U27233 (N_27233,N_25501,N_26240);
or U27234 (N_27234,N_24984,N_25443);
xnor U27235 (N_27235,N_25869,N_24721);
or U27236 (N_27236,N_25379,N_25900);
nand U27237 (N_27237,N_26214,N_24804);
nor U27238 (N_27238,N_25773,N_24016);
and U27239 (N_27239,N_24489,N_24850);
or U27240 (N_27240,N_25812,N_25761);
and U27241 (N_27241,N_26289,N_26439);
or U27242 (N_27242,N_26448,N_26453);
xor U27243 (N_27243,N_24193,N_26192);
and U27244 (N_27244,N_25618,N_24803);
nand U27245 (N_27245,N_24316,N_25966);
or U27246 (N_27246,N_25401,N_26078);
and U27247 (N_27247,N_26324,N_26369);
and U27248 (N_27248,N_26350,N_26631);
or U27249 (N_27249,N_24963,N_24285);
and U27250 (N_27250,N_25367,N_26269);
nand U27251 (N_27251,N_26737,N_24545);
and U27252 (N_27252,N_24384,N_26121);
xor U27253 (N_27253,N_24511,N_25349);
or U27254 (N_27254,N_26024,N_24715);
or U27255 (N_27255,N_25251,N_25372);
and U27256 (N_27256,N_26646,N_25700);
or U27257 (N_27257,N_25587,N_24921);
nor U27258 (N_27258,N_25103,N_25202);
nor U27259 (N_27259,N_24345,N_25099);
nor U27260 (N_27260,N_26142,N_26651);
or U27261 (N_27261,N_26090,N_26176);
nand U27262 (N_27262,N_24723,N_25754);
nor U27263 (N_27263,N_26591,N_26603);
nand U27264 (N_27264,N_25651,N_24097);
nor U27265 (N_27265,N_25921,N_24882);
xor U27266 (N_27266,N_26812,N_26194);
and U27267 (N_27267,N_25815,N_25434);
nand U27268 (N_27268,N_25162,N_24092);
nor U27269 (N_27269,N_26815,N_24287);
nor U27270 (N_27270,N_26178,N_26141);
xnor U27271 (N_27271,N_25783,N_24030);
nand U27272 (N_27272,N_25619,N_26195);
nand U27273 (N_27273,N_25340,N_26267);
nand U27274 (N_27274,N_26499,N_25764);
nor U27275 (N_27275,N_24326,N_25294);
or U27276 (N_27276,N_26912,N_25807);
xnor U27277 (N_27277,N_24089,N_25986);
xor U27278 (N_27278,N_25088,N_24606);
nor U27279 (N_27279,N_26880,N_24854);
nor U27280 (N_27280,N_24607,N_24558);
nor U27281 (N_27281,N_24647,N_26984);
or U27282 (N_27282,N_26919,N_25776);
nand U27283 (N_27283,N_26211,N_24110);
nor U27284 (N_27284,N_25351,N_25516);
or U27285 (N_27285,N_24523,N_25593);
nor U27286 (N_27286,N_24100,N_26879);
xnor U27287 (N_27287,N_25201,N_26119);
and U27288 (N_27288,N_24289,N_26140);
nor U27289 (N_27289,N_26705,N_25531);
or U27290 (N_27290,N_26611,N_26793);
nand U27291 (N_27291,N_24074,N_25243);
and U27292 (N_27292,N_24166,N_25492);
or U27293 (N_27293,N_24065,N_26057);
nor U27294 (N_27294,N_26780,N_24865);
or U27295 (N_27295,N_24988,N_25237);
and U27296 (N_27296,N_26795,N_24307);
xor U27297 (N_27297,N_25756,N_25498);
or U27298 (N_27298,N_24194,N_26124);
nor U27299 (N_27299,N_26743,N_25960);
nor U27300 (N_27300,N_24415,N_24477);
nor U27301 (N_27301,N_25582,N_25384);
and U27302 (N_27302,N_26827,N_26134);
or U27303 (N_27303,N_26999,N_24109);
and U27304 (N_27304,N_26358,N_24927);
or U27305 (N_27305,N_24789,N_26261);
or U27306 (N_27306,N_24546,N_25238);
xnor U27307 (N_27307,N_24842,N_24613);
or U27308 (N_27308,N_25309,N_25098);
nand U27309 (N_27309,N_24666,N_24819);
and U27310 (N_27310,N_26878,N_24456);
nor U27311 (N_27311,N_26962,N_24689);
or U27312 (N_27312,N_24099,N_26375);
and U27313 (N_27313,N_24981,N_24412);
and U27314 (N_27314,N_25454,N_26070);
xor U27315 (N_27315,N_24070,N_24770);
nand U27316 (N_27316,N_24378,N_24449);
nand U27317 (N_27317,N_24504,N_26865);
nand U27318 (N_27318,N_25432,N_25022);
or U27319 (N_27319,N_25228,N_26424);
and U27320 (N_27320,N_26995,N_26288);
nand U27321 (N_27321,N_25120,N_24083);
xnor U27322 (N_27322,N_26043,N_26183);
and U27323 (N_27323,N_25479,N_26174);
xnor U27324 (N_27324,N_26652,N_25070);
nand U27325 (N_27325,N_24851,N_24141);
nand U27326 (N_27326,N_24013,N_26244);
nand U27327 (N_27327,N_24982,N_24996);
xnor U27328 (N_27328,N_25509,N_26670);
nand U27329 (N_27329,N_26076,N_24469);
or U27330 (N_27330,N_25393,N_24530);
nor U27331 (N_27331,N_26540,N_26927);
and U27332 (N_27332,N_24323,N_24067);
nor U27333 (N_27333,N_25180,N_25045);
nor U27334 (N_27334,N_26884,N_26492);
xnor U27335 (N_27335,N_25769,N_25771);
nand U27336 (N_27336,N_25343,N_24705);
and U27337 (N_27337,N_25203,N_25424);
and U27338 (N_27338,N_26437,N_25968);
xnor U27339 (N_27339,N_24010,N_24252);
and U27340 (N_27340,N_25053,N_25583);
and U27341 (N_27341,N_26389,N_25131);
nand U27342 (N_27342,N_25233,N_25240);
nand U27343 (N_27343,N_24210,N_26451);
or U27344 (N_27344,N_25031,N_26868);
and U27345 (N_27345,N_26126,N_25940);
nor U27346 (N_27346,N_24642,N_24122);
or U27347 (N_27347,N_25580,N_24778);
nor U27348 (N_27348,N_24266,N_24496);
xor U27349 (N_27349,N_25313,N_26774);
xnor U27350 (N_27350,N_25862,N_26640);
nand U27351 (N_27351,N_25075,N_26433);
or U27352 (N_27352,N_25801,N_24295);
xnor U27353 (N_27353,N_24383,N_24061);
and U27354 (N_27354,N_25221,N_26352);
nor U27355 (N_27355,N_24313,N_26742);
nor U27356 (N_27356,N_25461,N_25611);
or U27357 (N_27357,N_25189,N_25792);
nand U27358 (N_27358,N_25310,N_26222);
nand U27359 (N_27359,N_25763,N_25563);
xnor U27360 (N_27360,N_26525,N_25474);
xnor U27361 (N_27361,N_25222,N_26889);
or U27362 (N_27362,N_24591,N_26110);
or U27363 (N_27363,N_26954,N_25303);
and U27364 (N_27364,N_24583,N_26506);
nand U27365 (N_27365,N_26069,N_26806);
nor U27366 (N_27366,N_25543,N_24142);
nor U27367 (N_27367,N_26188,N_26952);
xnor U27368 (N_27368,N_26237,N_26909);
nor U27369 (N_27369,N_24627,N_24454);
and U27370 (N_27370,N_24348,N_24429);
xor U27371 (N_27371,N_25460,N_26103);
nor U27372 (N_27372,N_24485,N_24260);
nand U27373 (N_27373,N_24925,N_25781);
or U27374 (N_27374,N_24239,N_26710);
nand U27375 (N_27375,N_24431,N_26766);
nor U27376 (N_27376,N_26527,N_26282);
nand U27377 (N_27377,N_24231,N_24615);
nand U27378 (N_27378,N_26849,N_26075);
or U27379 (N_27379,N_26445,N_24336);
or U27380 (N_27380,N_26725,N_24780);
and U27381 (N_27381,N_25380,N_24840);
nor U27382 (N_27382,N_26833,N_26852);
or U27383 (N_27383,N_26342,N_24670);
xnor U27384 (N_27384,N_25999,N_26407);
nor U27385 (N_27385,N_25049,N_24073);
nor U27386 (N_27386,N_24202,N_26660);
nand U27387 (N_27387,N_24494,N_26048);
or U27388 (N_27388,N_24197,N_24340);
or U27389 (N_27389,N_26144,N_24579);
and U27390 (N_27390,N_25655,N_24971);
or U27391 (N_27391,N_25123,N_24829);
xnor U27392 (N_27392,N_24933,N_25297);
or U27393 (N_27393,N_24806,N_25316);
and U27394 (N_27394,N_24355,N_24450);
and U27395 (N_27395,N_24363,N_24785);
nor U27396 (N_27396,N_24584,N_26474);
nor U27397 (N_27397,N_26325,N_25574);
nand U27398 (N_27398,N_26724,N_26656);
or U27399 (N_27399,N_26544,N_26036);
xnor U27400 (N_27400,N_24005,N_26894);
and U27401 (N_27401,N_25050,N_25562);
nand U27402 (N_27402,N_25347,N_24271);
or U27403 (N_27403,N_26081,N_26639);
nand U27404 (N_27404,N_25732,N_24021);
or U27405 (N_27405,N_25983,N_24997);
and U27406 (N_27406,N_26580,N_26354);
nand U27407 (N_27407,N_25279,N_26503);
or U27408 (N_27408,N_24327,N_25671);
xor U27409 (N_27409,N_24024,N_26818);
nor U27410 (N_27410,N_25006,N_26049);
xor U27411 (N_27411,N_26302,N_25811);
nand U27412 (N_27412,N_25266,N_26227);
nor U27413 (N_27413,N_26489,N_26559);
nand U27414 (N_27414,N_24731,N_26012);
and U27415 (N_27415,N_25466,N_25299);
nor U27416 (N_27416,N_24938,N_26297);
nor U27417 (N_27417,N_24565,N_24163);
and U27418 (N_27418,N_26488,N_26693);
xnor U27419 (N_27419,N_24212,N_24328);
or U27420 (N_27420,N_25694,N_24824);
and U27421 (N_27421,N_24175,N_24640);
nor U27422 (N_27422,N_26853,N_26931);
nand U27423 (N_27423,N_26777,N_26595);
and U27424 (N_27424,N_26309,N_25932);
nand U27425 (N_27425,N_24926,N_26597);
nand U27426 (N_27426,N_24011,N_26403);
nand U27427 (N_27427,N_26415,N_24547);
nand U27428 (N_27428,N_24170,N_24900);
xnor U27429 (N_27429,N_26348,N_24875);
and U27430 (N_27430,N_24960,N_24039);
and U27431 (N_27431,N_26162,N_26960);
and U27432 (N_27432,N_25344,N_24796);
nand U27433 (N_27433,N_24575,N_24783);
or U27434 (N_27434,N_24200,N_26895);
nor U27435 (N_27435,N_24208,N_24521);
or U27436 (N_27436,N_26387,N_25609);
and U27437 (N_27437,N_25758,N_24148);
nor U27438 (N_27438,N_24448,N_26034);
nor U27439 (N_27439,N_25090,N_24129);
and U27440 (N_27440,N_26985,N_24167);
or U27441 (N_27441,N_26581,N_26467);
xnor U27442 (N_27442,N_24434,N_25134);
and U27443 (N_27443,N_26382,N_24754);
nor U27444 (N_27444,N_25258,N_24868);
xor U27445 (N_27445,N_26845,N_26166);
or U27446 (N_27446,N_26254,N_25370);
and U27447 (N_27447,N_26405,N_26246);
or U27448 (N_27448,N_24916,N_26592);
and U27449 (N_27449,N_24862,N_26376);
and U27450 (N_27450,N_25988,N_25522);
or U27451 (N_27451,N_24439,N_24417);
nand U27452 (N_27452,N_25462,N_25533);
and U27453 (N_27453,N_26050,N_26223);
nand U27454 (N_27454,N_25413,N_24177);
xor U27455 (N_27455,N_26787,N_24402);
xor U27456 (N_27456,N_26466,N_25868);
and U27457 (N_27457,N_26861,N_24768);
and U27458 (N_27458,N_25101,N_25768);
nand U27459 (N_27459,N_24867,N_25377);
or U27460 (N_27460,N_25922,N_26113);
nand U27461 (N_27461,N_26831,N_26007);
or U27462 (N_27462,N_26986,N_26590);
and U27463 (N_27463,N_26401,N_25642);
xor U27464 (N_27464,N_26399,N_24369);
or U27465 (N_27465,N_24817,N_25019);
and U27466 (N_27466,N_26374,N_25799);
nand U27467 (N_27467,N_24683,N_25605);
nand U27468 (N_27468,N_26599,N_24246);
nand U27469 (N_27469,N_24279,N_24403);
nand U27470 (N_27470,N_24568,N_26131);
nor U27471 (N_27471,N_26447,N_24599);
nand U27472 (N_27472,N_25624,N_24339);
or U27473 (N_27473,N_25602,N_25214);
nand U27474 (N_27474,N_26882,N_25216);
nand U27475 (N_27475,N_24275,N_24676);
or U27476 (N_27476,N_24374,N_24220);
nor U27477 (N_27477,N_25264,N_24972);
or U27478 (N_27478,N_24667,N_26485);
xor U27479 (N_27479,N_25502,N_26534);
and U27480 (N_27480,N_25673,N_25330);
or U27481 (N_27481,N_24929,N_26573);
and U27482 (N_27482,N_26455,N_25860);
and U27483 (N_27483,N_25959,N_24696);
and U27484 (N_27484,N_24713,N_24869);
or U27485 (N_27485,N_26015,N_26941);
or U27486 (N_27486,N_26629,N_25269);
and U27487 (N_27487,N_24240,N_26200);
or U27488 (N_27488,N_25976,N_26657);
and U27489 (N_27489,N_25946,N_24603);
and U27490 (N_27490,N_25375,N_25867);
and U27491 (N_27491,N_26836,N_25736);
xnor U27492 (N_27492,N_25468,N_25005);
and U27493 (N_27493,N_24810,N_26976);
or U27494 (N_27494,N_26130,N_25080);
nor U27495 (N_27495,N_26410,N_25252);
or U27496 (N_27496,N_24605,N_24587);
or U27497 (N_27497,N_26063,N_24512);
or U27498 (N_27498,N_26630,N_25298);
and U27499 (N_27499,N_25421,N_25654);
nor U27500 (N_27500,N_25823,N_26098);
and U27501 (N_27501,N_24219,N_24634);
or U27502 (N_27502,N_25661,N_26760);
nor U27503 (N_27503,N_24009,N_25083);
nor U27504 (N_27504,N_24708,N_25629);
or U27505 (N_27505,N_26336,N_24693);
nor U27506 (N_27506,N_26802,N_24022);
or U27507 (N_27507,N_26135,N_24497);
and U27508 (N_27508,N_26146,N_25188);
nor U27509 (N_27509,N_25755,N_25069);
nand U27510 (N_27510,N_25106,N_24728);
nor U27511 (N_27511,N_26225,N_24578);
nand U27512 (N_27512,N_26182,N_24790);
nor U27513 (N_27513,N_24541,N_25963);
and U27514 (N_27514,N_24703,N_25920);
or U27515 (N_27515,N_26797,N_24350);
or U27516 (N_27516,N_24843,N_26505);
and U27517 (N_27517,N_25119,N_24028);
nor U27518 (N_27518,N_25197,N_26589);
nor U27519 (N_27519,N_26715,N_26905);
nand U27520 (N_27520,N_24792,N_24787);
nand U27521 (N_27521,N_25614,N_25236);
or U27522 (N_27522,N_25962,N_24205);
nor U27523 (N_27523,N_25332,N_25819);
xor U27524 (N_27524,N_26177,N_26184);
and U27525 (N_27525,N_26832,N_24744);
and U27526 (N_27526,N_26553,N_26968);
nand U27527 (N_27527,N_25931,N_24592);
or U27528 (N_27528,N_24550,N_26769);
or U27529 (N_27529,N_24108,N_25601);
nor U27530 (N_27530,N_24098,N_26851);
nor U27531 (N_27531,N_25325,N_26420);
xnor U27532 (N_27532,N_24179,N_26528);
or U27533 (N_27533,N_24299,N_25280);
nor U27534 (N_27534,N_24894,N_26163);
nand U27535 (N_27535,N_25383,N_24405);
or U27536 (N_27536,N_24614,N_25791);
xor U27537 (N_27537,N_26251,N_24646);
nor U27538 (N_27538,N_25985,N_26086);
nor U27539 (N_27539,N_25032,N_26293);
xor U27540 (N_27540,N_24493,N_26272);
nand U27541 (N_27541,N_24131,N_26763);
nor U27542 (N_27542,N_24535,N_25695);
and U27543 (N_27543,N_26746,N_24919);
nor U27544 (N_27544,N_25138,N_24211);
nand U27545 (N_27545,N_24040,N_25472);
nand U27546 (N_27546,N_24825,N_24424);
or U27547 (N_27547,N_25054,N_25849);
or U27548 (N_27548,N_24091,N_24729);
nor U27549 (N_27549,N_26432,N_25471);
and U27550 (N_27550,N_26085,N_25882);
nor U27551 (N_27551,N_26838,N_25312);
xor U27552 (N_27552,N_25435,N_26770);
nand U27553 (N_27553,N_26377,N_24539);
nand U27554 (N_27554,N_25510,N_26005);
and U27555 (N_27555,N_25727,N_25320);
nand U27556 (N_27556,N_24571,N_26741);
or U27557 (N_27557,N_25873,N_24664);
and U27558 (N_27558,N_26975,N_24059);
or U27559 (N_27559,N_24481,N_26226);
or U27560 (N_27560,N_24594,N_24382);
xnor U27561 (N_27561,N_25517,N_25198);
xor U27562 (N_27562,N_25314,N_24989);
or U27563 (N_27563,N_26438,N_24096);
xnor U27564 (N_27564,N_24118,N_26837);
xor U27565 (N_27565,N_24701,N_24413);
xor U27566 (N_27566,N_24506,N_26231);
or U27567 (N_27567,N_24870,N_26680);
nor U27568 (N_27568,N_24045,N_24373);
nor U27569 (N_27569,N_26046,N_25575);
nor U27570 (N_27570,N_26708,N_24410);
or U27571 (N_27571,N_26561,N_25011);
xnor U27572 (N_27572,N_24288,N_24213);
or U27573 (N_27573,N_24446,N_25538);
nor U27574 (N_27574,N_24297,N_25613);
nand U27575 (N_27575,N_24898,N_24822);
xor U27576 (N_27576,N_26773,N_26565);
or U27577 (N_27577,N_25095,N_24229);
or U27578 (N_27578,N_24983,N_24903);
nor U27579 (N_27579,N_25577,N_24856);
xnor U27580 (N_27580,N_25406,N_25217);
nor U27581 (N_27581,N_26009,N_25072);
and U27582 (N_27582,N_25291,N_24272);
xnor U27583 (N_27583,N_24399,N_26890);
nand U27584 (N_27584,N_26801,N_25091);
and U27585 (N_27585,N_24172,N_24761);
nand U27586 (N_27586,N_26805,N_26460);
xor U27587 (N_27587,N_24095,N_26068);
xnor U27588 (N_27588,N_26294,N_24283);
nor U27589 (N_27589,N_26798,N_24577);
nand U27590 (N_27590,N_25872,N_25820);
nand U27591 (N_27591,N_24420,N_24020);
and U27592 (N_27592,N_26804,N_26383);
and U27593 (N_27593,N_25186,N_24514);
nand U27594 (N_27594,N_26366,N_25919);
and U27595 (N_27595,N_25052,N_26979);
xor U27596 (N_27596,N_26274,N_26362);
or U27597 (N_27597,N_26965,N_24957);
and U27598 (N_27598,N_24421,N_25114);
and U27599 (N_27599,N_26841,N_25009);
nand U27600 (N_27600,N_25263,N_24786);
xor U27601 (N_27601,N_24400,N_24159);
or U27602 (N_27602,N_26235,N_24697);
or U27603 (N_27603,N_25974,N_26546);
nand U27604 (N_27604,N_25436,N_26665);
nor U27605 (N_27605,N_25404,N_26792);
xnor U27606 (N_27606,N_26556,N_26648);
xor U27607 (N_27607,N_24874,N_25301);
xnor U27608 (N_27608,N_25402,N_24716);
nor U27609 (N_27609,N_24094,N_24528);
xnor U27610 (N_27610,N_25893,N_24764);
or U27611 (N_27611,N_25173,N_26228);
and U27612 (N_27612,N_26734,N_24338);
and U27613 (N_27613,N_24572,N_26395);
or U27614 (N_27614,N_26345,N_25975);
nor U27615 (N_27615,N_25918,N_26981);
or U27616 (N_27616,N_25458,N_24832);
nor U27617 (N_27617,N_24143,N_25681);
and U27618 (N_27618,N_26079,N_25419);
xnor U27619 (N_27619,N_24527,N_25910);
nand U27620 (N_27620,N_26404,N_26616);
or U27621 (N_27621,N_26716,N_25969);
nand U27622 (N_27622,N_25308,N_24544);
nor U27623 (N_27623,N_24158,N_26154);
nor U27624 (N_27624,N_24668,N_24884);
nor U27625 (N_27625,N_24331,N_25431);
nand U27626 (N_27626,N_26679,N_26346);
or U27627 (N_27627,N_25658,N_24335);
or U27628 (N_27628,N_26022,N_24015);
nand U27629 (N_27629,N_24187,N_26800);
or U27630 (N_27630,N_25141,N_26242);
or U27631 (N_27631,N_26982,N_24491);
xnor U27632 (N_27632,N_25559,N_26035);
nor U27633 (N_27633,N_25223,N_26697);
nor U27634 (N_27634,N_25871,N_24954);
or U27635 (N_27635,N_25741,N_26444);
nor U27636 (N_27636,N_24990,N_25441);
xnor U27637 (N_27637,N_25551,N_25979);
nand U27638 (N_27638,N_25062,N_25033);
nand U27639 (N_27639,N_24132,N_26199);
nor U27640 (N_27640,N_26548,N_24657);
nor U27641 (N_27641,N_25163,N_25025);
nand U27642 (N_27642,N_24595,N_26571);
nor U27643 (N_27643,N_24695,N_26564);
xor U27644 (N_27644,N_25584,N_24243);
nor U27645 (N_27645,N_24130,N_24698);
and U27646 (N_27646,N_26752,N_25981);
nand U27647 (N_27647,N_24324,N_24848);
and U27648 (N_27648,N_26704,N_26055);
or U27649 (N_27649,N_24811,N_24967);
xnor U27650 (N_27650,N_25579,N_25737);
and U27651 (N_27651,N_24222,N_25341);
and U27652 (N_27652,N_26220,N_25172);
or U27653 (N_27653,N_25373,N_26339);
nor U27654 (N_27654,N_25728,N_24265);
xnor U27655 (N_27655,N_25427,N_26649);
nand U27656 (N_27656,N_26391,N_26138);
or U27657 (N_27657,N_26167,N_26411);
and U27658 (N_27658,N_24280,N_25646);
nand U27659 (N_27659,N_25337,N_26504);
nand U27660 (N_27660,N_25570,N_26783);
xor U27661 (N_27661,N_26781,N_24447);
and U27662 (N_27662,N_25687,N_24891);
nand U27663 (N_27663,N_24835,N_24444);
nand U27664 (N_27664,N_25534,N_24951);
nor U27665 (N_27665,N_26842,N_26191);
xnor U27666 (N_27666,N_25622,N_26915);
nand U27667 (N_27667,N_24330,N_26969);
or U27668 (N_27668,N_25068,N_25504);
xnor U27669 (N_27669,N_25887,N_25400);
nand U27670 (N_27670,N_26252,N_25143);
or U27671 (N_27671,N_25042,N_24377);
or U27672 (N_27672,N_24105,N_26193);
nand U27673 (N_27673,N_26379,N_25898);
and U27674 (N_27674,N_24513,N_25018);
xor U27675 (N_27675,N_24371,N_25505);
nand U27676 (N_27676,N_25693,N_25038);
or U27677 (N_27677,N_24757,N_25641);
or U27678 (N_27678,N_26751,N_25295);
nor U27679 (N_27679,N_26273,N_25470);
and U27680 (N_27680,N_24309,N_24247);
xnor U27681 (N_27681,N_25833,N_24364);
or U27682 (N_27682,N_26108,N_24379);
or U27683 (N_27683,N_24956,N_26461);
or U27684 (N_27684,N_24069,N_26137);
or U27685 (N_27685,N_24739,N_24014);
xor U27686 (N_27686,N_25512,N_24653);
nand U27687 (N_27687,N_26218,N_24224);
nor U27688 (N_27688,N_26186,N_25339);
or U27689 (N_27689,N_25420,N_25934);
nand U27690 (N_27690,N_25770,N_24964);
xnor U27691 (N_27691,N_25557,N_25561);
and U27692 (N_27692,N_25676,N_25408);
or U27693 (N_27693,N_24230,N_24828);
xor U27694 (N_27694,N_26713,N_25916);
or U27695 (N_27695,N_25714,N_26932);
xnor U27696 (N_27696,N_25598,N_26786);
xnor U27697 (N_27697,N_25998,N_25506);
nand U27698 (N_27698,N_25638,N_26243);
nand U27699 (N_27699,N_24518,N_25270);
and U27700 (N_27700,N_26885,N_25497);
or U27701 (N_27701,N_25422,N_25836);
nor U27702 (N_27702,N_25917,N_24610);
or U27703 (N_27703,N_24140,N_25081);
xnor U27704 (N_27704,N_25982,N_25193);
nor U27705 (N_27705,N_25886,N_24128);
nand U27706 (N_27706,N_25077,N_24508);
nand U27707 (N_27707,N_26672,N_24034);
xnor U27708 (N_27708,N_24251,N_26215);
xor U27709 (N_27709,N_25683,N_24113);
nand U27710 (N_27710,N_25515,N_24628);
xnor U27711 (N_27711,N_26661,N_26776);
xor U27712 (N_27712,N_24062,N_24629);
or U27713 (N_27713,N_24404,N_25789);
nand U27714 (N_27714,N_24581,N_24038);
or U27715 (N_27715,N_25632,N_26380);
and U27716 (N_27716,N_26877,N_24763);
nor U27717 (N_27717,N_26340,N_24841);
nor U27718 (N_27718,N_25283,N_25444);
nor U27719 (N_27719,N_26123,N_24625);
nor U27720 (N_27720,N_25674,N_24419);
xor U27721 (N_27721,N_25338,N_24522);
nor U27722 (N_27722,N_26887,N_24249);
or U27723 (N_27723,N_26908,N_26473);
and U27724 (N_27724,N_25670,N_24978);
nor U27725 (N_27725,N_26784,N_24188);
nand U27726 (N_27726,N_26740,N_24771);
xnor U27727 (N_27727,N_24300,N_24586);
or U27728 (N_27728,N_24945,N_25459);
xor U27729 (N_27729,N_24928,N_26767);
nor U27730 (N_27730,N_25086,N_25473);
or U27731 (N_27731,N_24914,N_26360);
or U27732 (N_27732,N_25495,N_25927);
or U27733 (N_27733,N_24724,N_26519);
xor U27734 (N_27734,N_26371,N_26245);
nand U27735 (N_27735,N_25552,N_26921);
or U27736 (N_27736,N_24351,N_25766);
nand U27737 (N_27737,N_24888,N_24347);
nand U27738 (N_27738,N_26901,N_26241);
nand U27739 (N_27739,N_25542,N_26609);
and U27740 (N_27740,N_25486,N_26726);
nand U27741 (N_27741,N_25600,N_24248);
nand U27742 (N_27742,N_24762,N_25227);
and U27743 (N_27743,N_26255,N_25476);
and U27744 (N_27744,N_24133,N_26152);
nor U27745 (N_27745,N_25096,N_25864);
or U27746 (N_27746,N_26650,N_26212);
and U27747 (N_27747,N_26778,N_24509);
or U27748 (N_27748,N_26626,N_26093);
nand U27749 (N_27749,N_24023,N_25631);
xor U27750 (N_27750,N_26216,N_26699);
or U27751 (N_27751,N_26691,N_24502);
and U27752 (N_27752,N_25571,N_25785);
or U27753 (N_27753,N_25682,N_24503);
nor U27754 (N_27754,N_25196,N_24501);
nand U27755 (N_27755,N_26809,N_25149);
xnor U27756 (N_27756,N_26972,N_24310);
or U27757 (N_27757,N_26600,N_25544);
nor U27758 (N_27758,N_24425,N_24164);
nor U27759 (N_27759,N_25411,N_25566);
xnor U27760 (N_27760,N_25665,N_26207);
nor U27761 (N_27761,N_25939,N_24116);
nor U27762 (N_27762,N_25014,N_26898);
nand U27763 (N_27763,N_26088,N_24864);
xnor U27764 (N_27764,N_24075,N_24598);
nor U27765 (N_27765,N_25061,N_25041);
nor U27766 (N_27766,N_25115,N_25691);
nand U27767 (N_27767,N_25941,N_24082);
xor U27768 (N_27768,N_24725,N_26577);
nand U27769 (N_27769,N_24286,N_26280);
nor U27770 (N_27770,N_26938,N_24234);
nor U27771 (N_27771,N_26572,N_26706);
and U27772 (N_27772,N_24858,N_25213);
nor U27773 (N_27773,N_26937,N_26606);
nor U27774 (N_27774,N_26298,N_25518);
nand U27775 (N_27775,N_25717,N_25637);
and U27776 (N_27776,N_25991,N_24574);
nand U27777 (N_27777,N_26537,N_24970);
or U27778 (N_27778,N_25540,N_26728);
nand U27779 (N_27779,N_26313,N_25286);
nand U27780 (N_27780,N_26248,N_26641);
and U27781 (N_27781,N_24947,N_24250);
and U27782 (N_27782,N_24427,N_26234);
or U27783 (N_27783,N_24318,N_26685);
xor U27784 (N_27784,N_26933,N_25405);
nand U27785 (N_27785,N_25247,N_26698);
xnor U27786 (N_27786,N_25644,N_25529);
or U27787 (N_27787,N_25150,N_25089);
nor U27788 (N_27788,N_24221,N_24507);
or U27789 (N_27789,N_24752,N_26187);
nor U27790 (N_27790,N_25627,N_25290);
nor U27791 (N_27791,N_25924,N_24537);
nor U27792 (N_27792,N_26338,N_25284);
xnor U27793 (N_27793,N_24735,N_26970);
and U27794 (N_27794,N_26295,N_24918);
xor U27795 (N_27795,N_26281,N_26331);
nand U27796 (N_27796,N_24103,N_24774);
nand U27797 (N_27797,N_24389,N_26257);
or U27798 (N_27798,N_26423,N_26469);
nor U27799 (N_27799,N_24361,N_25346);
nand U27800 (N_27800,N_24797,N_26478);
and U27801 (N_27801,N_25879,N_25358);
nor U27802 (N_27802,N_25195,N_24057);
xnor U27803 (N_27803,N_24319,N_25046);
nand U27804 (N_27804,N_24050,N_25463);
and U27805 (N_27805,N_24018,N_26421);
xnor U27806 (N_27806,N_25164,N_25723);
or U27807 (N_27807,N_26006,N_26735);
and U27808 (N_27808,N_26155,N_24526);
nor U27809 (N_27809,N_26517,N_25356);
nor U27810 (N_27810,N_26867,N_26814);
xnor U27811 (N_27811,N_25649,N_26621);
and U27812 (N_27812,N_25711,N_24566);
and U27813 (N_27813,N_24218,N_25359);
xnor U27814 (N_27814,N_24733,N_25212);
or U27815 (N_27815,N_25650,N_25725);
nor U27816 (N_27816,N_26185,N_25112);
or U27817 (N_27817,N_24029,N_25355);
or U27818 (N_27818,N_25191,N_24102);
nor U27819 (N_27819,N_25122,N_25669);
and U27820 (N_27820,N_24663,N_26221);
nor U27821 (N_27821,N_24162,N_24041);
nor U27822 (N_27822,N_24442,N_25936);
nand U27823 (N_27823,N_26122,N_26862);
nor U27824 (N_27824,N_26917,N_25664);
and U27825 (N_27825,N_25208,N_25908);
xor U27826 (N_27826,N_24630,N_26025);
xnor U27827 (N_27827,N_24631,N_26496);
nand U27828 (N_27828,N_25076,N_26000);
and U27829 (N_27829,N_25734,N_24802);
and U27830 (N_27830,N_25742,N_24980);
nand U27831 (N_27831,N_25667,N_26635);
xnor U27832 (N_27832,N_26111,N_24033);
nor U27833 (N_27833,N_24805,N_26446);
nand U27834 (N_27834,N_24254,N_26663);
nor U27835 (N_27835,N_24680,N_26956);
nor U27836 (N_27836,N_26654,N_26618);
and U27837 (N_27837,N_26584,N_25440);
and U27838 (N_27838,N_26671,N_24895);
nor U27839 (N_27839,N_25888,N_25775);
nor U27840 (N_27840,N_26087,N_25858);
nand U27841 (N_27841,N_26826,N_25387);
xnor U27842 (N_27842,N_24236,N_24408);
or U27843 (N_27843,N_24671,N_26266);
nand U27844 (N_27844,N_26502,N_26967);
and U27845 (N_27845,N_24500,N_25889);
nand U27846 (N_27846,N_26532,N_24117);
nor U27847 (N_27847,N_25398,N_26992);
xnor U27848 (N_27848,N_26576,N_24775);
nor U27849 (N_27849,N_25079,N_24144);
nand U27850 (N_27850,N_26061,N_26638);
or U27851 (N_27851,N_25092,N_24101);
and U27852 (N_27852,N_25645,N_26759);
nor U27853 (N_27853,N_24321,N_26136);
nor U27854 (N_27854,N_25909,N_26688);
xor U27855 (N_27855,N_25839,N_24146);
nor U27856 (N_27856,N_24042,N_25105);
nand U27857 (N_27857,N_24952,N_24465);
xnor U27858 (N_27858,N_25636,N_24644);
nand U27859 (N_27859,N_24863,N_25790);
and U27860 (N_27860,N_26622,N_25716);
nor U27861 (N_27861,N_26799,N_26396);
nor U27862 (N_27862,N_24800,N_26757);
xor U27863 (N_27863,N_25021,N_24959);
nand U27864 (N_27864,N_24685,N_26615);
or U27865 (N_27865,N_25368,N_26579);
xor U27866 (N_27866,N_25588,N_25948);
nand U27867 (N_27867,N_25219,N_26305);
nand U27868 (N_27868,N_26041,N_26761);
nor U27869 (N_27869,N_26810,N_24455);
and U27870 (N_27870,N_24151,N_24053);
or U27871 (N_27871,N_26988,N_26094);
xor U27872 (N_27872,N_26092,N_25161);
and U27873 (N_27873,N_25712,N_25412);
nor U27874 (N_27874,N_25287,N_25818);
nor U27875 (N_27875,N_25190,N_26196);
nor U27876 (N_27876,N_25938,N_26300);
and U27877 (N_27877,N_25793,N_26568);
and U27878 (N_27878,N_24341,N_26161);
nor U27879 (N_27879,N_25719,N_24153);
nand U27880 (N_27880,N_26442,N_25788);
xnor U27881 (N_27881,N_24437,N_25876);
xor U27882 (N_27882,N_24480,N_26322);
or U27883 (N_27883,N_26493,N_24263);
and U27884 (N_27884,N_24931,N_26971);
or U27885 (N_27885,N_25272,N_24261);
xnor U27886 (N_27886,N_24619,N_24641);
xor U27887 (N_27887,N_25017,N_26381);
and U27888 (N_27888,N_26004,N_24601);
xnor U27889 (N_27889,N_25735,N_24658);
nor U27890 (N_27890,N_26318,N_25275);
and U27891 (N_27891,N_25621,N_26700);
or U27892 (N_27892,N_25743,N_25292);
and U27893 (N_27893,N_25861,N_24452);
xnor U27894 (N_27894,N_26658,N_26583);
or U27895 (N_27895,N_24852,N_25798);
and U27896 (N_27896,N_24388,N_26542);
nor U27897 (N_27897,N_25947,N_24515);
nand U27898 (N_27898,N_25635,N_25956);
and U27899 (N_27899,N_26074,N_25058);
or U27900 (N_27900,N_26511,N_24582);
or U27901 (N_27901,N_24552,N_24031);
nor U27902 (N_27902,N_26594,N_25870);
nand U27903 (N_27903,N_25030,N_26132);
and U27904 (N_27904,N_25684,N_25429);
nor U27905 (N_27905,N_25688,N_26203);
nor U27906 (N_27906,N_25851,N_24830);
and U27907 (N_27907,N_25390,N_26431);
nand U27908 (N_27908,N_24650,N_24001);
or U27909 (N_27909,N_24611,N_24397);
or U27910 (N_27910,N_25152,N_25554);
and U27911 (N_27911,N_26925,N_26450);
nor U27912 (N_27912,N_26961,N_25617);
and U27913 (N_27913,N_25615,N_25381);
or U27914 (N_27914,N_26343,N_26355);
nor U27915 (N_27915,N_25388,N_25482);
nor U27916 (N_27916,N_26359,N_26263);
or U27917 (N_27917,N_26531,N_24621);
nand U27918 (N_27918,N_25035,N_25132);
xnor U27919 (N_27919,N_25511,N_26456);
or U27920 (N_27920,N_25277,N_25100);
nor U27921 (N_27921,N_26264,N_26428);
nor U27922 (N_27922,N_26586,N_25526);
xor U27923 (N_27923,N_25174,N_26045);
nand U27924 (N_27924,N_25690,N_25326);
nor U27925 (N_27925,N_25318,N_24195);
nand U27926 (N_27926,N_25274,N_26850);
xnor U27927 (N_27927,N_25513,N_26549);
or U27928 (N_27928,N_25528,N_25508);
and U27929 (N_27929,N_24317,N_24681);
and U27930 (N_27930,N_25026,N_25546);
and U27931 (N_27931,N_25480,N_26911);
nand U27932 (N_27932,N_26903,N_25549);
nand U27933 (N_27933,N_25797,N_26422);
xor U27934 (N_27934,N_26011,N_26089);
and U27935 (N_27935,N_26392,N_24652);
or U27936 (N_27936,N_26091,N_24178);
nor U27937 (N_27937,N_25015,N_26158);
xor U27938 (N_27938,N_24529,N_24684);
and U27939 (N_27939,N_26107,N_25980);
xor U27940 (N_27940,N_25333,N_24495);
xor U27941 (N_27941,N_24655,N_25335);
and U27942 (N_27942,N_26230,N_24782);
nand U27943 (N_27943,N_25226,N_24993);
or U27944 (N_27944,N_24567,N_24087);
nand U27945 (N_27945,N_25211,N_25950);
nor U27946 (N_27946,N_25536,N_26239);
and U27947 (N_27947,N_26673,N_25679);
xor U27948 (N_27948,N_25964,N_26686);
and U27949 (N_27949,N_25838,N_25530);
and U27950 (N_27950,N_24156,N_24505);
nor U27951 (N_27951,N_26518,N_25995);
and U27952 (N_27952,N_26929,N_24883);
and U27953 (N_27953,N_25000,N_25353);
and U27954 (N_27954,N_25082,N_25365);
xor U27955 (N_27955,N_26541,N_25087);
nand U27956 (N_27956,N_25437,N_25953);
and U27957 (N_27957,N_26311,N_24974);
nand U27958 (N_27958,N_25826,N_24853);
nand U27959 (N_27959,N_26910,N_25718);
xor U27960 (N_27960,N_25137,N_26328);
or U27961 (N_27961,N_25378,N_24332);
and U27962 (N_27962,N_25425,N_25182);
or U27963 (N_27963,N_26633,N_25795);
or U27964 (N_27964,N_25065,N_24561);
and U27965 (N_27965,N_25171,N_25949);
nor U27966 (N_27966,N_25154,N_25336);
or U27967 (N_27967,N_26018,N_25160);
nand U27968 (N_27968,N_24687,N_24939);
nand U27969 (N_27969,N_24998,N_24461);
nor U27970 (N_27970,N_24992,N_26723);
nand U27971 (N_27971,N_25433,N_26283);
nor U27972 (N_27972,N_26714,N_26835);
xnor U27973 (N_27973,N_24588,N_26899);
and U27974 (N_27974,N_24749,N_25804);
nor U27975 (N_27975,N_25109,N_26775);
nor U27976 (N_27976,N_26250,N_25478);
nor U27977 (N_27977,N_24055,N_24149);
nand U27978 (N_27978,N_24169,N_25166);
or U27979 (N_27979,N_24831,N_26659);
nor U27980 (N_27980,N_24633,N_26566);
or U27981 (N_27981,N_25824,N_24359);
and U27982 (N_27982,N_24793,N_26416);
xnor U27983 (N_27983,N_25720,N_25746);
nand U27984 (N_27984,N_26149,N_26562);
xnor U27985 (N_27985,N_26664,N_24296);
and U27986 (N_27986,N_26520,N_25599);
and U27987 (N_27987,N_24269,N_26668);
and U27988 (N_27988,N_26229,N_26623);
or U27989 (N_27989,N_25085,N_24277);
and U27990 (N_27990,N_24392,N_25984);
nand U27991 (N_27991,N_25814,N_26530);
and U27992 (N_27992,N_24911,N_25779);
and U27993 (N_27993,N_24532,N_25288);
xnor U27994 (N_27994,N_26683,N_26604);
nand U27995 (N_27995,N_24396,N_26102);
and U27996 (N_27996,N_26987,N_25487);
and U27997 (N_27997,N_24235,N_24897);
nand U27998 (N_27998,N_25955,N_24845);
and U27999 (N_27999,N_25890,N_24492);
or U28000 (N_28000,N_26750,N_26736);
xor U28001 (N_28001,N_24753,N_25912);
and U28002 (N_28002,N_24767,N_26692);
nand U28003 (N_28003,N_25449,N_25610);
xnor U28004 (N_28004,N_26205,N_24585);
nand U28005 (N_28005,N_25765,N_24462);
or U28006 (N_28006,N_25586,N_25750);
xnor U28007 (N_28007,N_25178,N_25064);
nor U28008 (N_28008,N_26830,N_26365);
nand U28009 (N_28009,N_25133,N_26419);
or U28010 (N_28010,N_24207,N_26099);
and U28011 (N_28011,N_25971,N_26636);
xnor U28012 (N_28012,N_25328,N_25877);
nor U28013 (N_28013,N_24325,N_26624);
or U28014 (N_28014,N_24256,N_26619);
xnor U28015 (N_28015,N_26232,N_25055);
or U28016 (N_28016,N_25772,N_26694);
nor U28017 (N_28017,N_25591,N_25747);
and U28018 (N_28018,N_26959,N_26536);
nand U28019 (N_28019,N_25672,N_25989);
and U28020 (N_28020,N_26408,N_26732);
nand U28021 (N_28021,N_24160,N_26598);
xnor U28022 (N_28022,N_25200,N_25391);
nor U28023 (N_28023,N_24543,N_25875);
or U28024 (N_28024,N_26217,N_25578);
nor U28025 (N_28025,N_25585,N_26236);
nor U28026 (N_28026,N_25322,N_25118);
xnor U28027 (N_28027,N_25142,N_24019);
or U28028 (N_28028,N_26436,N_24206);
nor U28029 (N_28029,N_25997,N_25662);
nand U28030 (N_28030,N_26551,N_26150);
or U28031 (N_28031,N_26817,N_26739);
xnor U28032 (N_28032,N_24357,N_24923);
nand U28033 (N_28033,N_26100,N_26682);
nor U28034 (N_28034,N_25699,N_26270);
or U28035 (N_28035,N_26782,N_26430);
and U28036 (N_28036,N_25832,N_24112);
and U28037 (N_28037,N_25556,N_25852);
and U28038 (N_28038,N_25481,N_24873);
xnor U28039 (N_28039,N_26066,N_25837);
nand U28040 (N_28040,N_26983,N_24878);
xor U28041 (N_28041,N_25125,N_25093);
and U28042 (N_28042,N_26412,N_25056);
and U28043 (N_28043,N_24977,N_26056);
nor U28044 (N_28044,N_25796,N_24198);
xor U28045 (N_28045,N_26943,N_24966);
nand U28046 (N_28046,N_25168,N_24549);
or U28047 (N_28047,N_26172,N_26441);
nor U28048 (N_28048,N_24354,N_26875);
nor U28049 (N_28049,N_24134,N_25048);
or U28050 (N_28050,N_24334,N_24738);
nor U28051 (N_28051,N_25724,N_25350);
or U28052 (N_28052,N_26276,N_25145);
nand U28053 (N_28053,N_26720,N_26427);
or U28054 (N_28054,N_25386,N_24460);
or U28055 (N_28055,N_24008,N_24214);
nand U28056 (N_28056,N_24196,N_24710);
nor U28057 (N_28057,N_25567,N_26394);
and U28058 (N_28058,N_26040,N_25396);
nand U28059 (N_28059,N_26866,N_24773);
xor U28060 (N_28060,N_25680,N_26980);
and U28061 (N_28061,N_24766,N_24719);
or U28062 (N_28062,N_24622,N_26669);
and U28063 (N_28063,N_24398,N_24290);
nor U28064 (N_28064,N_24808,N_24443);
nor U28065 (N_28065,N_24756,N_24861);
xnor U28066 (N_28066,N_24081,N_24225);
or U28067 (N_28067,N_25307,N_25369);
nand U28068 (N_28068,N_26676,N_25739);
nand U28069 (N_28069,N_26785,N_26479);
xor U28070 (N_28070,N_26032,N_24837);
xor U28071 (N_28071,N_25539,N_24961);
or U28072 (N_28072,N_24072,N_26744);
nor U28073 (N_28073,N_24740,N_26027);
xor U28074 (N_28074,N_26361,N_25521);
nor U28075 (N_28075,N_26632,N_25261);
and U28076 (N_28076,N_26038,N_24136);
or U28077 (N_28077,N_25996,N_25639);
nor U28078 (N_28078,N_25215,N_26120);
or U28079 (N_28079,N_25895,N_26811);
xor U28080 (N_28080,N_25126,N_26535);
or U28081 (N_28081,N_26449,N_24093);
or U28082 (N_28082,N_25183,N_24025);
or U28083 (N_28083,N_24284,N_24258);
nand U28084 (N_28084,N_25527,N_25067);
nand U28085 (N_28085,N_25242,N_24138);
nand U28086 (N_28086,N_24673,N_24826);
and U28087 (N_28087,N_25786,N_24844);
nand U28088 (N_28088,N_24746,N_24612);
nand U28089 (N_28089,N_26425,N_24185);
and U28090 (N_28090,N_24743,N_25371);
nand U28091 (N_28091,N_25537,N_24784);
xnor U28092 (N_28092,N_25967,N_25094);
xor U28093 (N_28093,N_26260,N_26645);
nor U28094 (N_28094,N_24562,N_24836);
xnor U28095 (N_28095,N_25345,N_26902);
nand U28096 (N_28096,N_26019,N_26258);
nor U28097 (N_28097,N_24060,N_25943);
nor U28098 (N_28098,N_25816,N_25787);
or U28099 (N_28099,N_25951,N_26790);
and U28100 (N_28100,N_24580,N_24312);
xnor U28101 (N_28101,N_24540,N_25192);
and U28102 (N_28102,N_26655,N_26607);
xnor U28103 (N_28103,N_26204,N_25493);
nand U28104 (N_28104,N_26820,N_25809);
or U28105 (N_28105,N_24301,N_25300);
xnor U28106 (N_28106,N_26013,N_26515);
and U28107 (N_28107,N_24686,N_25155);
or U28108 (N_28108,N_25323,N_26059);
or U28109 (N_28109,N_26279,N_24692);
xor U28110 (N_28110,N_25597,N_26803);
xnor U28111 (N_28111,N_24962,N_26501);
nand U28112 (N_28112,N_25348,N_25821);
nor U28113 (N_28113,N_26977,N_26434);
xnor U28114 (N_28114,N_26095,N_24490);
xor U28115 (N_28115,N_24654,N_24048);
nand U28116 (N_28116,N_26711,N_25001);
or U28117 (N_28117,N_25806,N_24517);
xor U28118 (N_28118,N_25246,N_24395);
or U28119 (N_28119,N_24675,N_24969);
nor U28120 (N_28120,N_24268,N_25496);
nor U28121 (N_28121,N_24035,N_26307);
nand U28122 (N_28122,N_24618,N_25643);
xor U28123 (N_28123,N_26955,N_26171);
or U28124 (N_28124,N_25232,N_25013);
nor U28125 (N_28125,N_24012,N_25426);
xor U28126 (N_28126,N_26224,N_26037);
or U28127 (N_28127,N_25881,N_26916);
and U28128 (N_28128,N_26003,N_24901);
and U28129 (N_28129,N_26400,N_25256);
or U28130 (N_28130,N_25625,N_26494);
nor U28131 (N_28131,N_24416,N_26973);
xnor U28132 (N_28132,N_24085,N_26353);
nand U28133 (N_28133,N_26854,N_24352);
and U28134 (N_28134,N_24223,N_26341);
and U28135 (N_28135,N_24816,N_24520);
nor U28136 (N_28136,N_24525,N_26316);
or U28137 (N_28137,N_26848,N_24181);
nor U28138 (N_28138,N_24887,N_25930);
xnor U28139 (N_28139,N_25701,N_26159);
xor U28140 (N_28140,N_26824,N_24294);
nand U28141 (N_28141,N_24407,N_24736);
xor U28142 (N_28142,N_24815,N_25846);
and U28143 (N_28143,N_25108,N_25907);
xor U28144 (N_28144,N_24638,N_25457);
and U28145 (N_28145,N_24027,N_24904);
nand U28146 (N_28146,N_24406,N_24847);
xnor U28147 (N_28147,N_24717,N_24674);
nor U28148 (N_28148,N_26935,N_24267);
nor U28149 (N_28149,N_26481,N_26303);
xnor U28150 (N_28150,N_25220,N_25957);
and U28151 (N_28151,N_25706,N_25012);
nand U28152 (N_28152,N_26718,N_26873);
or U28153 (N_28153,N_26500,N_24702);
or U28154 (N_28154,N_26116,N_26484);
and U28155 (N_28155,N_26275,N_26290);
nand U28156 (N_28156,N_25978,N_26363);
and U28157 (N_28157,N_25730,N_26008);
or U28158 (N_28158,N_25648,N_26385);
or U28159 (N_28159,N_24344,N_25060);
and U28160 (N_28160,N_25113,N_25863);
and U28161 (N_28161,N_25937,N_26994);
nand U28162 (N_28162,N_24292,N_25926);
xor U28163 (N_28163,N_26052,N_25389);
nor U28164 (N_28164,N_26860,N_26989);
nand U28165 (N_28165,N_24451,N_24991);
or U28166 (N_28166,N_25278,N_26417);
and U28167 (N_28167,N_24906,N_25689);
and U28168 (N_28168,N_26575,N_24257);
and U28169 (N_28169,N_25576,N_25633);
nand U28170 (N_28170,N_25596,N_24563);
nand U28171 (N_28171,N_24741,N_25902);
nor U28172 (N_28172,N_24342,N_24677);
or U28173 (N_28173,N_26157,N_25657);
xnor U28174 (N_28174,N_24609,N_24051);
nor U28175 (N_28175,N_26847,N_26189);
and U28176 (N_28176,N_25760,N_25117);
or U28177 (N_28177,N_24125,N_25146);
xnor U28178 (N_28178,N_26001,N_26031);
xnor U28179 (N_28179,N_26772,N_24119);
xnor U28180 (N_28180,N_25668,N_25352);
xnor U28181 (N_28181,N_26498,N_24441);
xnor U28182 (N_28182,N_24393,N_25503);
nand U28183 (N_28183,N_26238,N_26397);
and U28184 (N_28184,N_24616,N_26966);
nor U28185 (N_28185,N_26828,N_26990);
nor U28186 (N_28186,N_26578,N_26384);
and U28187 (N_28187,N_25374,N_24600);
and U28188 (N_28188,N_26926,N_24189);
and U28189 (N_28189,N_25738,N_25666);
nand U28190 (N_28190,N_25456,N_24699);
nand U28191 (N_28191,N_26016,N_24765);
and U28192 (N_28192,N_26106,N_25702);
or U28193 (N_28193,N_25157,N_24217);
nor U28194 (N_28194,N_24032,N_24090);
or U28195 (N_28195,N_26863,N_25675);
nor U28196 (N_28196,N_25696,N_24704);
nor U28197 (N_28197,N_25612,N_24168);
or U28198 (N_28198,N_25327,N_26570);
nor U28199 (N_28199,N_24368,N_24458);
xnor U28200 (N_28200,N_24165,N_25047);
and U28201 (N_28201,N_24948,N_25016);
and U28202 (N_28202,N_24080,N_26165);
or U28203 (N_28203,N_26083,N_24726);
and U28204 (N_28204,N_26567,N_24955);
nand U28205 (N_28205,N_24722,N_24322);
or U28206 (N_28206,N_25653,N_25843);
xnor U28207 (N_28207,N_26978,N_26529);
xor U28208 (N_28208,N_25229,N_24679);
xnor U28209 (N_28209,N_25315,N_24745);
nand U28210 (N_28210,N_24017,N_26625);
nand U28211 (N_28211,N_26613,N_26928);
and U28212 (N_28212,N_26198,N_24180);
nor U28213 (N_28213,N_26286,N_26356);
or U28214 (N_28214,N_26393,N_24682);
nand U28215 (N_28215,N_25156,N_26082);
and U28216 (N_28216,N_26789,N_24659);
and U28217 (N_28217,N_24468,N_26190);
xor U28218 (N_28218,N_24554,N_26996);
or U28219 (N_28219,N_25260,N_24759);
or U28220 (N_28220,N_24046,N_25329);
and U28221 (N_28221,N_26807,N_26779);
xor U28222 (N_28222,N_26077,N_26054);
or U28223 (N_28223,N_25808,N_24241);
nor U28224 (N_28224,N_26859,N_26913);
or U28225 (N_28225,N_26653,N_26508);
xor U28226 (N_28226,N_24573,N_25623);
nand U28227 (N_28227,N_24470,N_26513);
and U28228 (N_28228,N_26605,N_26904);
nand U28229 (N_28229,N_26958,N_24487);
and U28230 (N_28230,N_25987,N_24907);
xor U28231 (N_28231,N_26291,N_24510);
xor U28232 (N_28232,N_25029,N_26256);
nand U28233 (N_28233,N_26758,N_26117);
and U28234 (N_28234,N_24849,N_24182);
and U28235 (N_28235,N_25697,N_25210);
or U28236 (N_28236,N_26084,N_26357);
xnor U28237 (N_28237,N_24201,N_24556);
nor U28238 (N_28238,N_25901,N_26582);
nand U28239 (N_28239,N_24794,N_25704);
and U28240 (N_28240,N_24788,N_26344);
nand U28241 (N_28241,N_24608,N_25071);
xnor U28242 (N_28242,N_24823,N_26247);
or U28243 (N_28243,N_26104,N_24700);
or U28244 (N_28244,N_26864,N_24298);
nand U28245 (N_28245,N_25477,N_26857);
and U28246 (N_28246,N_26869,N_24435);
and U28247 (N_28247,N_25207,N_25855);
and U28248 (N_28248,N_24795,N_24120);
and U28249 (N_28249,N_25828,N_24123);
xnor U28250 (N_28250,N_24758,N_25652);
nand U28251 (N_28251,N_24390,N_25519);
xor U28252 (N_28252,N_24750,N_24857);
xor U28253 (N_28253,N_24386,N_26033);
or U28254 (N_28254,N_26475,N_24483);
and U28255 (N_28255,N_25767,N_26753);
nand U28256 (N_28256,N_24464,N_24643);
and U28257 (N_28257,N_25362,N_25397);
nor U28258 (N_28258,N_26398,N_25361);
or U28259 (N_28259,N_25859,N_24107);
nor U28260 (N_28260,N_26249,N_26721);
or U28261 (N_28261,N_24453,N_26042);
or U28262 (N_28262,N_26349,N_25066);
nor U28263 (N_28263,N_24281,N_25253);
or U28264 (N_28264,N_25894,N_26951);
or U28265 (N_28265,N_24154,N_25043);
nor U28266 (N_28266,N_26944,N_24881);
and U28267 (N_28267,N_24555,N_24920);
nand U28268 (N_28268,N_25407,N_25620);
and U28269 (N_28269,N_26539,N_25805);
nor U28270 (N_28270,N_26574,N_26443);
and U28271 (N_28271,N_25028,N_24799);
xnor U28272 (N_28272,N_25929,N_24635);
nand U28273 (N_28273,N_24078,N_25206);
and U28274 (N_28274,N_25409,N_26065);
xnor U28275 (N_28275,N_26039,N_24807);
nor U28276 (N_28276,N_24760,N_26373);
nor U28277 (N_28277,N_25181,N_26125);
or U28278 (N_28278,N_26071,N_26330);
or U28279 (N_28279,N_26169,N_26585);
and U28280 (N_28280,N_24358,N_26168);
or U28281 (N_28281,N_25097,N_26310);
nor U28282 (N_28282,N_25255,N_24430);
nor U28283 (N_28283,N_24597,N_26627);
or U28284 (N_28284,N_24463,N_26265);
or U28285 (N_28285,N_26023,N_25179);
xnor U28286 (N_28286,N_25958,N_25777);
and U28287 (N_28287,N_24066,N_26957);
or U28288 (N_28288,N_25304,N_24570);
nor U28289 (N_28289,N_26487,N_24560);
xnor U28290 (N_28290,N_25364,N_26319);
nand U28291 (N_28291,N_26156,N_24174);
or U28292 (N_28292,N_24137,N_25185);
and U28293 (N_28293,N_25452,N_24380);
nor U28294 (N_28294,N_26480,N_26922);
or U28295 (N_28295,N_25169,N_25394);
xor U28296 (N_28296,N_24233,N_26702);
and U28297 (N_28297,N_24833,N_25565);
and U28298 (N_28298,N_25177,N_25002);
xor U28299 (N_28299,N_26593,N_26271);
or U28300 (N_28300,N_25010,N_25525);
xnor U28301 (N_28301,N_26472,N_25568);
and U28302 (N_28302,N_26044,N_26202);
or U28303 (N_28303,N_24871,N_25856);
and U28304 (N_28304,N_24975,N_24976);
or U28305 (N_28305,N_24519,N_24135);
nand U28306 (N_28306,N_26118,N_25244);
and U28307 (N_28307,N_24199,N_25225);
nor U28308 (N_28308,N_25813,N_24071);
nand U28309 (N_28309,N_24936,N_25334);
or U28310 (N_28310,N_26114,N_24459);
xor U28311 (N_28311,N_25489,N_24186);
nor U28312 (N_28312,N_26677,N_24457);
nor U28313 (N_28313,N_25708,N_25572);
xnor U28314 (N_28314,N_25973,N_26097);
or U28315 (N_28315,N_24781,N_26333);
nand U28316 (N_28316,N_26418,N_24418);
and U28317 (N_28317,N_26335,N_25865);
xnor U28318 (N_28318,N_24127,N_24176);
and U28319 (N_28319,N_24428,N_24531);
or U28320 (N_28320,N_25911,N_25485);
or U28321 (N_28321,N_26612,N_24270);
and U28322 (N_28322,N_24003,N_24473);
nor U28323 (N_28323,N_25854,N_26601);
nor U28324 (N_28324,N_24088,N_26210);
nor U28325 (N_28325,N_26709,N_26881);
and U28326 (N_28326,N_26406,N_24171);
nor U28327 (N_28327,N_25282,N_25965);
nor U28328 (N_28328,N_25774,N_26703);
or U28329 (N_28329,N_26028,N_24264);
and U28330 (N_28330,N_26465,N_24190);
nand U28331 (N_28331,N_26351,N_26285);
nand U28332 (N_28332,N_24308,N_26893);
nand U28333 (N_28333,N_25116,N_26558);
nand U28334 (N_28334,N_25803,N_26213);
nand U28335 (N_28335,N_24068,N_25059);
xor U28336 (N_28336,N_25842,N_25660);
and U28337 (N_28337,N_25262,N_24999);
nor U28338 (N_28338,N_24056,N_26533);
or U28339 (N_28339,N_25239,N_26304);
or U28340 (N_28340,N_26823,N_25616);
or U28341 (N_28341,N_25438,N_26555);
nand U28342 (N_28342,N_25416,N_24036);
nor U28343 (N_28343,N_24751,N_24636);
nand U28344 (N_28344,N_25993,N_26647);
nor U28345 (N_28345,N_24052,N_26834);
or U28346 (N_28346,N_24953,N_25036);
nand U28347 (N_28347,N_26109,N_26440);
nand U28348 (N_28348,N_26942,N_26112);
or U28349 (N_28349,N_26796,N_24282);
nor U28350 (N_28350,N_25187,N_24306);
nand U28351 (N_28351,N_24346,N_25603);
and U28352 (N_28352,N_24423,N_25659);
xor U28353 (N_28353,N_26170,N_26139);
and U28354 (N_28354,N_25677,N_26510);
and U28355 (N_28355,N_26327,N_26923);
or U28356 (N_28356,N_26262,N_24394);
nor U28357 (N_28357,N_26201,N_26173);
nand U28358 (N_28358,N_25078,N_24086);
or U28359 (N_28359,N_25564,N_24209);
nor U28360 (N_28360,N_25135,N_24944);
and U28361 (N_28361,N_25748,N_26765);
nand U28362 (N_28362,N_26681,N_24152);
and U28363 (N_28363,N_24173,N_25994);
xnor U28364 (N_28364,N_24755,N_24589);
xnor U28365 (N_28365,N_24482,N_24776);
and U28366 (N_28366,N_25541,N_24569);
xnor U28367 (N_28367,N_26143,N_24742);
and U28368 (N_28368,N_25121,N_26208);
and U28369 (N_28369,N_24436,N_25810);
and U28370 (N_28370,N_24791,N_24813);
nor U28371 (N_28371,N_26950,N_26675);
and U28372 (N_28372,N_25430,N_26299);
nand U28373 (N_28373,N_25729,N_25204);
xor U28374 (N_28374,N_25840,N_26516);
or U28375 (N_28375,N_24932,N_25376);
and U28376 (N_28376,N_26233,N_24812);
xnor U28377 (N_28377,N_24238,N_24366);
nand U28378 (N_28378,N_25535,N_26560);
xnor U28379 (N_28379,N_24314,N_26164);
and U28380 (N_28380,N_25608,N_25224);
nor U28381 (N_28381,N_25915,N_26948);
nor U28382 (N_28382,N_24467,N_24370);
or U28383 (N_28383,N_25532,N_24054);
nand U28384 (N_28384,N_24827,N_24838);
and U28385 (N_28385,N_24002,N_25970);
nor U28386 (N_28386,N_24973,N_25439);
or U28387 (N_28387,N_25257,N_25640);
and U28388 (N_28388,N_24656,N_26939);
nand U28389 (N_28389,N_26062,N_24942);
or U28390 (N_28390,N_26930,N_25853);
nor U28391 (N_28391,N_24215,N_24303);
nand U28392 (N_28392,N_26936,N_24913);
and U28393 (N_28393,N_25136,N_24204);
and U28394 (N_28394,N_26545,N_26756);
xor U28395 (N_28395,N_25241,N_26993);
xnor U28396 (N_28396,N_25745,N_26390);
xnor U28397 (N_28397,N_24748,N_26666);
or U28398 (N_28398,N_26749,N_26414);
nor U28399 (N_28399,N_24876,N_24576);
or U28400 (N_28400,N_26550,N_24946);
and U28401 (N_28401,N_24488,N_24866);
and U28402 (N_28402,N_24623,N_26512);
nor U28403 (N_28403,N_24391,N_24902);
and U28404 (N_28404,N_24184,N_25494);
and U28405 (N_28405,N_24349,N_25548);
and U28406 (N_28406,N_26454,N_24950);
and U28407 (N_28407,N_24772,N_24877);
xnor U28408 (N_28408,N_25874,N_24602);
or U28409 (N_28409,N_25231,N_24893);
or U28410 (N_28410,N_24302,N_26458);
xnor U28411 (N_28411,N_25153,N_25710);
nor U28412 (N_28412,N_26026,N_26301);
nand U28413 (N_28413,N_24304,N_24632);
nor U28414 (N_28414,N_26886,N_25447);
or U28415 (N_28415,N_24255,N_26730);
or U28416 (N_28416,N_26949,N_25707);
or U28417 (N_28417,N_26002,N_24115);
and U28418 (N_28418,N_24145,N_26497);
nor U28419 (N_28419,N_26053,N_25524);
or U28420 (N_28420,N_26128,N_24516);
and U28421 (N_28421,N_24669,N_25273);
nor U28422 (N_28422,N_24548,N_25488);
or U28423 (N_28423,N_26642,N_26072);
or U28424 (N_28424,N_25592,N_26684);
nor U28425 (N_28425,N_26794,N_24411);
and U28426 (N_28426,N_24637,N_26067);
nor U28427 (N_28427,N_26153,N_25847);
and U28428 (N_28428,N_26822,N_25753);
nand U28429 (N_28429,N_25024,N_26733);
or U28430 (N_28430,N_25491,N_26858);
nand U28431 (N_28431,N_26133,N_24691);
xor U28432 (N_28432,N_26596,N_26462);
xnor U28433 (N_28433,N_25883,N_25914);
and U28434 (N_28434,N_26717,N_25259);
or U28435 (N_28435,N_24367,N_26459);
xor U28436 (N_28436,N_26064,N_24694);
and U28437 (N_28437,N_25139,N_24466);
nand U28438 (N_28438,N_25446,N_24814);
and U28439 (N_28439,N_26347,N_24237);
nand U28440 (N_28440,N_25445,N_26483);
or U28441 (N_28441,N_26175,N_24834);
or U28442 (N_28442,N_25752,N_24244);
nand U28443 (N_28443,N_26856,N_24910);
or U28444 (N_28444,N_24353,N_26491);
nand U28445 (N_28445,N_26206,N_24305);
and U28446 (N_28446,N_24114,N_25713);
xnor U28447 (N_28447,N_24006,N_26617);
nand U28448 (N_28448,N_25794,N_25897);
or U28449 (N_28449,N_26047,N_24707);
nand U28450 (N_28450,N_25733,N_24228);
nand U28451 (N_28451,N_24809,N_24905);
xor U28452 (N_28452,N_24484,N_24553);
and U28453 (N_28453,N_24672,N_24968);
or U28454 (N_28454,N_24534,N_25140);
nand U28455 (N_28455,N_25594,N_26754);
xnor U28456 (N_28456,N_26287,N_24433);
xnor U28457 (N_28457,N_26829,N_25780);
nand U28458 (N_28458,N_25455,N_25104);
nor U28459 (N_28459,N_25170,N_25027);
nor U28460 (N_28460,N_25891,N_25703);
and U28461 (N_28461,N_26821,N_26509);
or U28462 (N_28462,N_26370,N_25841);
nor U28463 (N_28463,N_26364,N_26029);
nand U28464 (N_28464,N_26888,N_24000);
or U28465 (N_28465,N_26495,N_25268);
nand U28466 (N_28466,N_24734,N_26526);
and U28467 (N_28467,N_26945,N_25403);
nand U28468 (N_28468,N_25319,N_26719);
or U28469 (N_28469,N_26259,N_26947);
nor U28470 (N_28470,N_25961,N_25218);
or U28471 (N_28471,N_25848,N_25448);
xnor U28472 (N_28472,N_24885,N_25778);
xnor U28473 (N_28473,N_26674,N_24985);
and U28474 (N_28474,N_26620,N_25942);
or U28475 (N_28475,N_26127,N_26115);
nand U28476 (N_28476,N_25034,N_25500);
or U28477 (N_28477,N_25357,N_26151);
nor U28478 (N_28478,N_24203,N_26476);
or U28479 (N_28479,N_26073,N_25184);
nor U28480 (N_28480,N_26554,N_24564);
xor U28481 (N_28481,N_24559,N_24678);
nand U28482 (N_28482,N_25634,N_26470);
and U28483 (N_28483,N_24475,N_26368);
nor U28484 (N_28484,N_26426,N_25740);
nor U28485 (N_28485,N_26637,N_26464);
and U28486 (N_28486,N_26722,N_24779);
nand U28487 (N_28487,N_26644,N_24737);
nand U28488 (N_28488,N_24886,N_26934);
nand U28489 (N_28489,N_26457,N_26334);
nor U28490 (N_28490,N_25230,N_25418);
xor U28491 (N_28491,N_25829,N_24479);
xor U28492 (N_28492,N_25465,N_24915);
or U28493 (N_28493,N_24551,N_26964);
xnor U28494 (N_28494,N_24890,N_25628);
nor U28495 (N_28495,N_24943,N_25647);
or U28496 (N_28496,N_24498,N_24232);
and U28497 (N_28497,N_26180,N_24709);
and U28498 (N_28498,N_25464,N_26372);
or U28499 (N_28499,N_26060,N_25176);
nand U28500 (N_28500,N_24462,N_25255);
or U28501 (N_28501,N_26104,N_25304);
xnor U28502 (N_28502,N_25797,N_26495);
nand U28503 (N_28503,N_24191,N_26560);
xnor U28504 (N_28504,N_24692,N_24781);
nand U28505 (N_28505,N_25629,N_26002);
nor U28506 (N_28506,N_25089,N_26782);
and U28507 (N_28507,N_26636,N_24851);
nor U28508 (N_28508,N_26242,N_26193);
nor U28509 (N_28509,N_26861,N_26531);
and U28510 (N_28510,N_26311,N_25890);
nor U28511 (N_28511,N_24572,N_24720);
xnor U28512 (N_28512,N_25152,N_26478);
nor U28513 (N_28513,N_25058,N_24396);
nand U28514 (N_28514,N_24021,N_24647);
and U28515 (N_28515,N_25251,N_26142);
nand U28516 (N_28516,N_26842,N_24691);
xnor U28517 (N_28517,N_25790,N_25164);
xor U28518 (N_28518,N_26864,N_24653);
nand U28519 (N_28519,N_24083,N_25685);
nand U28520 (N_28520,N_26281,N_26289);
xor U28521 (N_28521,N_26942,N_24044);
nand U28522 (N_28522,N_24203,N_26182);
nor U28523 (N_28523,N_24459,N_25497);
nand U28524 (N_28524,N_24812,N_25118);
and U28525 (N_28525,N_24347,N_26431);
nand U28526 (N_28526,N_25473,N_26449);
xor U28527 (N_28527,N_25782,N_26337);
and U28528 (N_28528,N_25926,N_26503);
or U28529 (N_28529,N_25553,N_24810);
or U28530 (N_28530,N_26123,N_25797);
and U28531 (N_28531,N_24891,N_25374);
xor U28532 (N_28532,N_26600,N_25617);
and U28533 (N_28533,N_25531,N_24090);
nor U28534 (N_28534,N_26447,N_25496);
nor U28535 (N_28535,N_25714,N_24563);
nand U28536 (N_28536,N_26557,N_24547);
xnor U28537 (N_28537,N_25095,N_26489);
xnor U28538 (N_28538,N_24691,N_24614);
or U28539 (N_28539,N_24558,N_26994);
xnor U28540 (N_28540,N_26099,N_26566);
or U28541 (N_28541,N_24426,N_25729);
nor U28542 (N_28542,N_24284,N_24819);
xor U28543 (N_28543,N_26795,N_26892);
and U28544 (N_28544,N_26055,N_25610);
xnor U28545 (N_28545,N_24560,N_25359);
nand U28546 (N_28546,N_26190,N_26786);
xor U28547 (N_28547,N_25496,N_24697);
and U28548 (N_28548,N_25323,N_25876);
nor U28549 (N_28549,N_24101,N_25335);
and U28550 (N_28550,N_24705,N_25667);
or U28551 (N_28551,N_25213,N_25487);
xnor U28552 (N_28552,N_26217,N_26482);
or U28553 (N_28553,N_25618,N_26134);
and U28554 (N_28554,N_26056,N_25970);
nand U28555 (N_28555,N_26222,N_24730);
xnor U28556 (N_28556,N_24400,N_26411);
xor U28557 (N_28557,N_26138,N_26010);
xor U28558 (N_28558,N_25650,N_25250);
xnor U28559 (N_28559,N_24048,N_25982);
and U28560 (N_28560,N_25886,N_26677);
nand U28561 (N_28561,N_25412,N_24606);
nor U28562 (N_28562,N_26570,N_25216);
or U28563 (N_28563,N_24201,N_26644);
or U28564 (N_28564,N_24244,N_25224);
or U28565 (N_28565,N_25706,N_24909);
xnor U28566 (N_28566,N_25310,N_24191);
and U28567 (N_28567,N_24862,N_25371);
nor U28568 (N_28568,N_25450,N_25518);
or U28569 (N_28569,N_24073,N_25043);
or U28570 (N_28570,N_26425,N_24492);
nor U28571 (N_28571,N_24308,N_26176);
or U28572 (N_28572,N_24939,N_25303);
and U28573 (N_28573,N_24145,N_25595);
xor U28574 (N_28574,N_24000,N_25497);
nand U28575 (N_28575,N_24792,N_24662);
and U28576 (N_28576,N_25132,N_24027);
nand U28577 (N_28577,N_26286,N_24156);
nand U28578 (N_28578,N_24541,N_25365);
xor U28579 (N_28579,N_24290,N_25811);
nor U28580 (N_28580,N_26185,N_26217);
nor U28581 (N_28581,N_26983,N_26222);
xnor U28582 (N_28582,N_24710,N_24668);
nand U28583 (N_28583,N_25609,N_24487);
nand U28584 (N_28584,N_24236,N_26761);
and U28585 (N_28585,N_24993,N_26729);
and U28586 (N_28586,N_25755,N_24583);
xor U28587 (N_28587,N_24883,N_26172);
nand U28588 (N_28588,N_26529,N_24853);
or U28589 (N_28589,N_26498,N_24709);
or U28590 (N_28590,N_26720,N_25286);
and U28591 (N_28591,N_26631,N_26822);
xor U28592 (N_28592,N_25294,N_24858);
and U28593 (N_28593,N_24926,N_26645);
nand U28594 (N_28594,N_26741,N_24123);
nand U28595 (N_28595,N_25018,N_26418);
nor U28596 (N_28596,N_25730,N_24584);
nand U28597 (N_28597,N_24746,N_26823);
or U28598 (N_28598,N_24745,N_24128);
nor U28599 (N_28599,N_25538,N_26554);
nor U28600 (N_28600,N_25789,N_24638);
or U28601 (N_28601,N_26177,N_26062);
and U28602 (N_28602,N_25308,N_25647);
xor U28603 (N_28603,N_26343,N_24251);
nand U28604 (N_28604,N_26642,N_24804);
xor U28605 (N_28605,N_25364,N_26502);
or U28606 (N_28606,N_24124,N_24490);
or U28607 (N_28607,N_26373,N_25056);
nor U28608 (N_28608,N_25724,N_25465);
or U28609 (N_28609,N_26168,N_25606);
nor U28610 (N_28610,N_24443,N_24654);
or U28611 (N_28611,N_24396,N_24207);
nand U28612 (N_28612,N_24202,N_25291);
or U28613 (N_28613,N_24714,N_24964);
or U28614 (N_28614,N_24864,N_26618);
nor U28615 (N_28615,N_24111,N_26793);
xnor U28616 (N_28616,N_24265,N_26627);
xor U28617 (N_28617,N_24390,N_26234);
and U28618 (N_28618,N_24991,N_26815);
or U28619 (N_28619,N_26674,N_26234);
xor U28620 (N_28620,N_26787,N_24191);
xor U28621 (N_28621,N_25030,N_25246);
or U28622 (N_28622,N_24187,N_26996);
nor U28623 (N_28623,N_26221,N_24744);
nor U28624 (N_28624,N_25507,N_24869);
or U28625 (N_28625,N_25490,N_25826);
and U28626 (N_28626,N_24824,N_26245);
nor U28627 (N_28627,N_26797,N_24196);
xor U28628 (N_28628,N_24439,N_25471);
xor U28629 (N_28629,N_24342,N_25635);
nor U28630 (N_28630,N_26056,N_26545);
nand U28631 (N_28631,N_25530,N_25388);
and U28632 (N_28632,N_24607,N_26142);
xor U28633 (N_28633,N_24962,N_24905);
or U28634 (N_28634,N_25482,N_26430);
and U28635 (N_28635,N_24288,N_25792);
nand U28636 (N_28636,N_25030,N_25895);
xnor U28637 (N_28637,N_24723,N_25809);
xnor U28638 (N_28638,N_26713,N_25459);
or U28639 (N_28639,N_26547,N_26252);
or U28640 (N_28640,N_24642,N_26388);
and U28641 (N_28641,N_26195,N_26387);
and U28642 (N_28642,N_25469,N_24318);
or U28643 (N_28643,N_24958,N_26639);
and U28644 (N_28644,N_25728,N_24211);
or U28645 (N_28645,N_25752,N_24199);
and U28646 (N_28646,N_25521,N_24112);
or U28647 (N_28647,N_26229,N_25945);
nand U28648 (N_28648,N_25249,N_24671);
nor U28649 (N_28649,N_24279,N_25248);
nor U28650 (N_28650,N_26989,N_24897);
nand U28651 (N_28651,N_26976,N_26563);
nand U28652 (N_28652,N_26383,N_25975);
and U28653 (N_28653,N_25989,N_26269);
and U28654 (N_28654,N_26657,N_26674);
and U28655 (N_28655,N_24236,N_26509);
and U28656 (N_28656,N_26773,N_26711);
or U28657 (N_28657,N_24725,N_25097);
nor U28658 (N_28658,N_25067,N_24128);
or U28659 (N_28659,N_24870,N_24111);
and U28660 (N_28660,N_26872,N_24578);
and U28661 (N_28661,N_25800,N_26844);
or U28662 (N_28662,N_26712,N_24469);
nand U28663 (N_28663,N_26970,N_26969);
xor U28664 (N_28664,N_24588,N_24611);
nor U28665 (N_28665,N_26195,N_25308);
or U28666 (N_28666,N_25353,N_24092);
nand U28667 (N_28667,N_25032,N_24485);
or U28668 (N_28668,N_25041,N_25849);
nor U28669 (N_28669,N_26926,N_24220);
xor U28670 (N_28670,N_25061,N_25478);
or U28671 (N_28671,N_25821,N_26500);
and U28672 (N_28672,N_26877,N_24711);
nor U28673 (N_28673,N_25468,N_26056);
and U28674 (N_28674,N_25696,N_25413);
xor U28675 (N_28675,N_26242,N_24604);
and U28676 (N_28676,N_26921,N_24861);
and U28677 (N_28677,N_24039,N_25588);
nand U28678 (N_28678,N_26022,N_25424);
nand U28679 (N_28679,N_26246,N_26810);
xor U28680 (N_28680,N_26809,N_26761);
nor U28681 (N_28681,N_25124,N_24919);
nand U28682 (N_28682,N_24698,N_24657);
nor U28683 (N_28683,N_25093,N_24970);
and U28684 (N_28684,N_26498,N_24696);
nand U28685 (N_28685,N_24733,N_26633);
nand U28686 (N_28686,N_25849,N_25466);
or U28687 (N_28687,N_25229,N_26559);
or U28688 (N_28688,N_25962,N_24239);
or U28689 (N_28689,N_26964,N_25376);
xnor U28690 (N_28690,N_26651,N_24370);
and U28691 (N_28691,N_26669,N_26124);
nand U28692 (N_28692,N_26469,N_26273);
nor U28693 (N_28693,N_26674,N_24253);
and U28694 (N_28694,N_26040,N_26892);
xnor U28695 (N_28695,N_25110,N_24932);
xor U28696 (N_28696,N_25421,N_25473);
and U28697 (N_28697,N_25705,N_24777);
nand U28698 (N_28698,N_25945,N_25816);
and U28699 (N_28699,N_26989,N_25592);
xor U28700 (N_28700,N_26663,N_26320);
or U28701 (N_28701,N_26117,N_26967);
nand U28702 (N_28702,N_26658,N_26459);
xor U28703 (N_28703,N_25659,N_24390);
or U28704 (N_28704,N_24158,N_26792);
xor U28705 (N_28705,N_25734,N_24206);
and U28706 (N_28706,N_24959,N_26748);
nand U28707 (N_28707,N_26568,N_24037);
xnor U28708 (N_28708,N_26408,N_25491);
nor U28709 (N_28709,N_25912,N_26517);
xnor U28710 (N_28710,N_26042,N_25775);
or U28711 (N_28711,N_25633,N_26870);
or U28712 (N_28712,N_25953,N_25747);
or U28713 (N_28713,N_26930,N_24341);
or U28714 (N_28714,N_26404,N_24919);
or U28715 (N_28715,N_24972,N_24537);
nand U28716 (N_28716,N_26015,N_25402);
xor U28717 (N_28717,N_24373,N_24682);
or U28718 (N_28718,N_25307,N_24406);
and U28719 (N_28719,N_26556,N_25023);
and U28720 (N_28720,N_24786,N_24920);
and U28721 (N_28721,N_24728,N_26096);
xnor U28722 (N_28722,N_25042,N_26229);
nor U28723 (N_28723,N_26858,N_25797);
xnor U28724 (N_28724,N_26977,N_26616);
nand U28725 (N_28725,N_24252,N_24125);
xor U28726 (N_28726,N_24282,N_24838);
or U28727 (N_28727,N_24016,N_24159);
or U28728 (N_28728,N_24016,N_25621);
nor U28729 (N_28729,N_26222,N_25170);
nand U28730 (N_28730,N_26095,N_26542);
and U28731 (N_28731,N_24860,N_25156);
nand U28732 (N_28732,N_24517,N_25413);
nor U28733 (N_28733,N_25132,N_24103);
xnor U28734 (N_28734,N_24933,N_25985);
xor U28735 (N_28735,N_24654,N_25048);
or U28736 (N_28736,N_24227,N_25454);
and U28737 (N_28737,N_26582,N_25402);
nand U28738 (N_28738,N_26006,N_26737);
or U28739 (N_28739,N_25913,N_26683);
xor U28740 (N_28740,N_25723,N_24805);
nand U28741 (N_28741,N_25226,N_24258);
nand U28742 (N_28742,N_25995,N_26443);
or U28743 (N_28743,N_24473,N_24446);
xnor U28744 (N_28744,N_24451,N_26108);
nor U28745 (N_28745,N_24662,N_24770);
nor U28746 (N_28746,N_26428,N_26403);
and U28747 (N_28747,N_25609,N_24532);
or U28748 (N_28748,N_24946,N_24534);
or U28749 (N_28749,N_24120,N_24127);
nand U28750 (N_28750,N_26303,N_24493);
or U28751 (N_28751,N_26889,N_25640);
and U28752 (N_28752,N_26839,N_24175);
nand U28753 (N_28753,N_25765,N_26270);
and U28754 (N_28754,N_25368,N_25615);
and U28755 (N_28755,N_25136,N_26220);
nor U28756 (N_28756,N_26399,N_25772);
or U28757 (N_28757,N_25213,N_25096);
and U28758 (N_28758,N_24550,N_26687);
nand U28759 (N_28759,N_25856,N_26036);
or U28760 (N_28760,N_26531,N_25262);
or U28761 (N_28761,N_26314,N_25667);
or U28762 (N_28762,N_25616,N_26784);
xnor U28763 (N_28763,N_25390,N_26399);
or U28764 (N_28764,N_24413,N_26998);
nand U28765 (N_28765,N_25795,N_24472);
or U28766 (N_28766,N_26546,N_24379);
and U28767 (N_28767,N_26442,N_25522);
nand U28768 (N_28768,N_25019,N_26760);
nand U28769 (N_28769,N_24950,N_25247);
nor U28770 (N_28770,N_26308,N_26394);
nand U28771 (N_28771,N_25275,N_24327);
nor U28772 (N_28772,N_24027,N_25025);
xnor U28773 (N_28773,N_26503,N_26268);
xor U28774 (N_28774,N_25994,N_25752);
nand U28775 (N_28775,N_26444,N_25248);
and U28776 (N_28776,N_25707,N_25635);
xnor U28777 (N_28777,N_26125,N_24193);
nor U28778 (N_28778,N_26083,N_26528);
and U28779 (N_28779,N_25279,N_24312);
and U28780 (N_28780,N_25104,N_25207);
or U28781 (N_28781,N_25782,N_25190);
nor U28782 (N_28782,N_26626,N_25586);
or U28783 (N_28783,N_26675,N_24075);
nand U28784 (N_28784,N_25806,N_24433);
xnor U28785 (N_28785,N_24274,N_24437);
nor U28786 (N_28786,N_24140,N_24421);
nor U28787 (N_28787,N_26528,N_24835);
nand U28788 (N_28788,N_24993,N_25388);
nor U28789 (N_28789,N_24147,N_25757);
nor U28790 (N_28790,N_25852,N_24042);
or U28791 (N_28791,N_25724,N_24532);
xor U28792 (N_28792,N_26529,N_24019);
and U28793 (N_28793,N_24839,N_26952);
nor U28794 (N_28794,N_25387,N_25936);
nor U28795 (N_28795,N_24034,N_25189);
and U28796 (N_28796,N_25063,N_24307);
or U28797 (N_28797,N_26229,N_25310);
nor U28798 (N_28798,N_24159,N_24855);
nand U28799 (N_28799,N_24489,N_25264);
xor U28800 (N_28800,N_24236,N_26395);
xnor U28801 (N_28801,N_24965,N_26505);
or U28802 (N_28802,N_25969,N_25911);
nand U28803 (N_28803,N_25541,N_24891);
or U28804 (N_28804,N_25845,N_26132);
xor U28805 (N_28805,N_26987,N_26857);
nor U28806 (N_28806,N_25521,N_25289);
xor U28807 (N_28807,N_25049,N_24778);
nor U28808 (N_28808,N_25550,N_24152);
xor U28809 (N_28809,N_26147,N_25864);
or U28810 (N_28810,N_26395,N_24641);
or U28811 (N_28811,N_24660,N_24485);
nand U28812 (N_28812,N_26355,N_24134);
xnor U28813 (N_28813,N_25181,N_25071);
nand U28814 (N_28814,N_26681,N_24690);
xnor U28815 (N_28815,N_24477,N_25125);
and U28816 (N_28816,N_24131,N_24538);
or U28817 (N_28817,N_24182,N_26839);
and U28818 (N_28818,N_24587,N_24859);
and U28819 (N_28819,N_24462,N_25814);
xnor U28820 (N_28820,N_25503,N_24703);
nand U28821 (N_28821,N_25127,N_24967);
or U28822 (N_28822,N_26276,N_26741);
xnor U28823 (N_28823,N_26731,N_26596);
xnor U28824 (N_28824,N_25685,N_24087);
nor U28825 (N_28825,N_25648,N_24575);
nand U28826 (N_28826,N_25738,N_24951);
xor U28827 (N_28827,N_24944,N_24008);
or U28828 (N_28828,N_24773,N_25247);
and U28829 (N_28829,N_25549,N_24838);
nor U28830 (N_28830,N_26470,N_25046);
nor U28831 (N_28831,N_25599,N_26315);
nor U28832 (N_28832,N_25357,N_26109);
and U28833 (N_28833,N_26810,N_24045);
nand U28834 (N_28834,N_25246,N_24192);
or U28835 (N_28835,N_24613,N_26338);
or U28836 (N_28836,N_24614,N_25605);
nor U28837 (N_28837,N_26280,N_24055);
xnor U28838 (N_28838,N_24942,N_25981);
and U28839 (N_28839,N_24853,N_26759);
nand U28840 (N_28840,N_25595,N_26560);
nor U28841 (N_28841,N_24639,N_24808);
nor U28842 (N_28842,N_24263,N_26520);
nand U28843 (N_28843,N_25636,N_26551);
or U28844 (N_28844,N_25572,N_26956);
and U28845 (N_28845,N_26661,N_26659);
nor U28846 (N_28846,N_25475,N_24710);
xnor U28847 (N_28847,N_24879,N_24171);
nand U28848 (N_28848,N_26493,N_26582);
and U28849 (N_28849,N_24660,N_26101);
xnor U28850 (N_28850,N_24140,N_26662);
or U28851 (N_28851,N_25121,N_26960);
xor U28852 (N_28852,N_25443,N_25663);
xnor U28853 (N_28853,N_25860,N_26581);
nor U28854 (N_28854,N_24962,N_24103);
or U28855 (N_28855,N_26853,N_24953);
nor U28856 (N_28856,N_24294,N_25092);
and U28857 (N_28857,N_24663,N_25184);
nor U28858 (N_28858,N_24961,N_26225);
or U28859 (N_28859,N_25925,N_24692);
nor U28860 (N_28860,N_24538,N_25677);
and U28861 (N_28861,N_24004,N_25763);
xor U28862 (N_28862,N_26614,N_25022);
nand U28863 (N_28863,N_25872,N_24715);
or U28864 (N_28864,N_24337,N_25229);
nand U28865 (N_28865,N_24289,N_25871);
nand U28866 (N_28866,N_25946,N_26096);
or U28867 (N_28867,N_24059,N_24126);
nand U28868 (N_28868,N_25804,N_26334);
nand U28869 (N_28869,N_24369,N_26012);
and U28870 (N_28870,N_24763,N_25938);
or U28871 (N_28871,N_24359,N_26326);
or U28872 (N_28872,N_26697,N_24277);
nand U28873 (N_28873,N_25787,N_24024);
xnor U28874 (N_28874,N_24416,N_26441);
or U28875 (N_28875,N_24145,N_25317);
and U28876 (N_28876,N_26209,N_26765);
or U28877 (N_28877,N_24269,N_24722);
nor U28878 (N_28878,N_25020,N_25939);
and U28879 (N_28879,N_24381,N_25881);
nor U28880 (N_28880,N_26712,N_26767);
and U28881 (N_28881,N_26772,N_25240);
nand U28882 (N_28882,N_26098,N_25193);
nand U28883 (N_28883,N_24384,N_24005);
nor U28884 (N_28884,N_24298,N_26393);
and U28885 (N_28885,N_24857,N_26031);
nor U28886 (N_28886,N_26502,N_25197);
and U28887 (N_28887,N_25117,N_24905);
and U28888 (N_28888,N_26184,N_26979);
or U28889 (N_28889,N_24997,N_26166);
nor U28890 (N_28890,N_25746,N_24683);
and U28891 (N_28891,N_26488,N_25338);
and U28892 (N_28892,N_24651,N_25160);
nor U28893 (N_28893,N_26270,N_25693);
nand U28894 (N_28894,N_25793,N_26980);
or U28895 (N_28895,N_26934,N_24086);
nor U28896 (N_28896,N_24946,N_26825);
and U28897 (N_28897,N_26975,N_25078);
xor U28898 (N_28898,N_26008,N_26869);
nand U28899 (N_28899,N_25509,N_25151);
or U28900 (N_28900,N_26204,N_24442);
and U28901 (N_28901,N_26918,N_25780);
and U28902 (N_28902,N_26952,N_26715);
or U28903 (N_28903,N_25104,N_24668);
or U28904 (N_28904,N_25003,N_26181);
or U28905 (N_28905,N_24489,N_25003);
and U28906 (N_28906,N_26893,N_24070);
nand U28907 (N_28907,N_24179,N_24338);
xor U28908 (N_28908,N_24563,N_26796);
xnor U28909 (N_28909,N_25135,N_26110);
or U28910 (N_28910,N_26685,N_24092);
xor U28911 (N_28911,N_26049,N_24794);
and U28912 (N_28912,N_25865,N_24822);
nand U28913 (N_28913,N_26263,N_25481);
nor U28914 (N_28914,N_24599,N_26158);
nor U28915 (N_28915,N_24933,N_24858);
nor U28916 (N_28916,N_24640,N_26972);
nor U28917 (N_28917,N_26738,N_25651);
and U28918 (N_28918,N_25335,N_24387);
and U28919 (N_28919,N_25379,N_24828);
xor U28920 (N_28920,N_24343,N_24597);
nor U28921 (N_28921,N_26194,N_24092);
and U28922 (N_28922,N_25769,N_25601);
or U28923 (N_28923,N_25085,N_25521);
and U28924 (N_28924,N_24996,N_25688);
nand U28925 (N_28925,N_25655,N_24279);
nor U28926 (N_28926,N_26200,N_24081);
or U28927 (N_28927,N_26832,N_26736);
or U28928 (N_28928,N_24773,N_25269);
nor U28929 (N_28929,N_26732,N_25208);
nor U28930 (N_28930,N_26871,N_25995);
nor U28931 (N_28931,N_24478,N_26709);
and U28932 (N_28932,N_24057,N_26790);
nor U28933 (N_28933,N_24240,N_25359);
and U28934 (N_28934,N_26265,N_26801);
nor U28935 (N_28935,N_25315,N_25432);
nand U28936 (N_28936,N_26622,N_24750);
xnor U28937 (N_28937,N_25762,N_26652);
or U28938 (N_28938,N_25573,N_25373);
xor U28939 (N_28939,N_26012,N_24503);
or U28940 (N_28940,N_25085,N_26373);
or U28941 (N_28941,N_25630,N_25985);
nand U28942 (N_28942,N_25718,N_26215);
and U28943 (N_28943,N_25467,N_25301);
or U28944 (N_28944,N_26550,N_24506);
nand U28945 (N_28945,N_26167,N_25340);
and U28946 (N_28946,N_25886,N_26525);
and U28947 (N_28947,N_26729,N_26096);
nand U28948 (N_28948,N_26835,N_25838);
or U28949 (N_28949,N_25211,N_24347);
and U28950 (N_28950,N_26728,N_26752);
or U28951 (N_28951,N_24662,N_26935);
nor U28952 (N_28952,N_25569,N_25797);
nor U28953 (N_28953,N_24860,N_26442);
xor U28954 (N_28954,N_26320,N_26364);
and U28955 (N_28955,N_24090,N_24140);
nor U28956 (N_28956,N_24762,N_26362);
nor U28957 (N_28957,N_25957,N_26883);
and U28958 (N_28958,N_24284,N_24277);
and U28959 (N_28959,N_25431,N_24821);
nand U28960 (N_28960,N_26609,N_24161);
and U28961 (N_28961,N_25253,N_26331);
nand U28962 (N_28962,N_24191,N_26763);
nor U28963 (N_28963,N_26052,N_25010);
nand U28964 (N_28964,N_26828,N_24647);
xnor U28965 (N_28965,N_25071,N_25142);
nor U28966 (N_28966,N_25143,N_26981);
xnor U28967 (N_28967,N_25933,N_25143);
nor U28968 (N_28968,N_24067,N_25091);
and U28969 (N_28969,N_24694,N_25784);
and U28970 (N_28970,N_24832,N_24561);
or U28971 (N_28971,N_24726,N_26351);
and U28972 (N_28972,N_25323,N_25848);
nor U28973 (N_28973,N_25695,N_26167);
nand U28974 (N_28974,N_25746,N_25204);
nor U28975 (N_28975,N_25120,N_25379);
nand U28976 (N_28976,N_25502,N_24341);
nor U28977 (N_28977,N_25747,N_25714);
nand U28978 (N_28978,N_24805,N_25627);
xor U28979 (N_28979,N_25919,N_25816);
or U28980 (N_28980,N_24566,N_24312);
nor U28981 (N_28981,N_24394,N_25910);
xnor U28982 (N_28982,N_26385,N_25920);
or U28983 (N_28983,N_26394,N_24797);
nand U28984 (N_28984,N_26249,N_26385);
nand U28985 (N_28985,N_24350,N_24850);
or U28986 (N_28986,N_25559,N_26063);
or U28987 (N_28987,N_24248,N_24736);
nand U28988 (N_28988,N_24931,N_24439);
nor U28989 (N_28989,N_26252,N_25603);
xor U28990 (N_28990,N_26855,N_24304);
and U28991 (N_28991,N_25402,N_24946);
nor U28992 (N_28992,N_25916,N_24124);
nor U28993 (N_28993,N_25999,N_24709);
nand U28994 (N_28994,N_24320,N_24829);
xnor U28995 (N_28995,N_24807,N_26805);
xor U28996 (N_28996,N_26867,N_24438);
xnor U28997 (N_28997,N_24997,N_24778);
or U28998 (N_28998,N_24443,N_26889);
and U28999 (N_28999,N_25016,N_26561);
nand U29000 (N_29000,N_26227,N_25017);
nand U29001 (N_29001,N_25036,N_26501);
and U29002 (N_29002,N_26687,N_25006);
or U29003 (N_29003,N_25688,N_24724);
nor U29004 (N_29004,N_24048,N_25867);
nor U29005 (N_29005,N_24071,N_24745);
and U29006 (N_29006,N_24572,N_25157);
xnor U29007 (N_29007,N_26037,N_26809);
and U29008 (N_29008,N_26267,N_24600);
nand U29009 (N_29009,N_25310,N_26501);
or U29010 (N_29010,N_25728,N_24435);
nor U29011 (N_29011,N_24550,N_26878);
nand U29012 (N_29012,N_24853,N_26087);
nand U29013 (N_29013,N_26830,N_25788);
and U29014 (N_29014,N_26029,N_26901);
and U29015 (N_29015,N_24568,N_25766);
or U29016 (N_29016,N_26038,N_24661);
and U29017 (N_29017,N_25610,N_24161);
and U29018 (N_29018,N_25347,N_25502);
or U29019 (N_29019,N_25791,N_24411);
xnor U29020 (N_29020,N_25436,N_25330);
xnor U29021 (N_29021,N_25419,N_26118);
xor U29022 (N_29022,N_25954,N_24324);
and U29023 (N_29023,N_25473,N_26878);
or U29024 (N_29024,N_24225,N_25780);
or U29025 (N_29025,N_25360,N_26850);
nand U29026 (N_29026,N_25809,N_26850);
nor U29027 (N_29027,N_26424,N_26837);
nand U29028 (N_29028,N_24619,N_25732);
and U29029 (N_29029,N_24893,N_24424);
or U29030 (N_29030,N_24903,N_26609);
and U29031 (N_29031,N_24030,N_25018);
or U29032 (N_29032,N_24541,N_24296);
nand U29033 (N_29033,N_26825,N_26339);
and U29034 (N_29034,N_25073,N_25711);
xnor U29035 (N_29035,N_25358,N_25437);
xnor U29036 (N_29036,N_25670,N_25133);
nand U29037 (N_29037,N_24422,N_25941);
xor U29038 (N_29038,N_26844,N_25721);
and U29039 (N_29039,N_26237,N_25582);
and U29040 (N_29040,N_26940,N_24667);
or U29041 (N_29041,N_26832,N_26869);
nand U29042 (N_29042,N_24920,N_24597);
nor U29043 (N_29043,N_25433,N_24468);
nor U29044 (N_29044,N_25074,N_24627);
or U29045 (N_29045,N_24783,N_25094);
or U29046 (N_29046,N_25122,N_26956);
and U29047 (N_29047,N_25698,N_26205);
and U29048 (N_29048,N_25697,N_25569);
nor U29049 (N_29049,N_26529,N_26344);
or U29050 (N_29050,N_26321,N_26979);
nand U29051 (N_29051,N_26460,N_26580);
or U29052 (N_29052,N_25093,N_26552);
and U29053 (N_29053,N_24999,N_24993);
xor U29054 (N_29054,N_24139,N_26781);
xnor U29055 (N_29055,N_25557,N_26608);
nor U29056 (N_29056,N_25284,N_25474);
xnor U29057 (N_29057,N_26656,N_24314);
nand U29058 (N_29058,N_26435,N_24697);
and U29059 (N_29059,N_25955,N_24869);
and U29060 (N_29060,N_26602,N_24300);
nor U29061 (N_29061,N_26947,N_25899);
xor U29062 (N_29062,N_24738,N_25040);
nand U29063 (N_29063,N_25022,N_24013);
xnor U29064 (N_29064,N_26033,N_25521);
xnor U29065 (N_29065,N_24788,N_26494);
xor U29066 (N_29066,N_25192,N_26602);
nand U29067 (N_29067,N_24403,N_26218);
xor U29068 (N_29068,N_26651,N_25645);
nor U29069 (N_29069,N_26406,N_26461);
or U29070 (N_29070,N_26187,N_24330);
nor U29071 (N_29071,N_26542,N_25382);
xor U29072 (N_29072,N_24908,N_24507);
or U29073 (N_29073,N_25557,N_24151);
nor U29074 (N_29074,N_26314,N_24819);
and U29075 (N_29075,N_24300,N_25487);
or U29076 (N_29076,N_25942,N_25810);
nor U29077 (N_29077,N_25069,N_24545);
nand U29078 (N_29078,N_26255,N_24892);
nor U29079 (N_29079,N_24965,N_24196);
xor U29080 (N_29080,N_24112,N_25692);
nand U29081 (N_29081,N_24968,N_25074);
and U29082 (N_29082,N_26928,N_25878);
xor U29083 (N_29083,N_25854,N_25015);
nor U29084 (N_29084,N_25922,N_24105);
nor U29085 (N_29085,N_26663,N_24776);
nand U29086 (N_29086,N_26176,N_25059);
or U29087 (N_29087,N_26110,N_24250);
nand U29088 (N_29088,N_24195,N_25242);
and U29089 (N_29089,N_25075,N_24569);
xnor U29090 (N_29090,N_24856,N_25117);
and U29091 (N_29091,N_26007,N_24544);
nor U29092 (N_29092,N_25446,N_24424);
nand U29093 (N_29093,N_25104,N_26330);
xor U29094 (N_29094,N_25762,N_25033);
nand U29095 (N_29095,N_25972,N_25092);
nand U29096 (N_29096,N_24800,N_26266);
nand U29097 (N_29097,N_26292,N_25425);
and U29098 (N_29098,N_24975,N_25149);
xnor U29099 (N_29099,N_24255,N_24056);
or U29100 (N_29100,N_24584,N_26548);
nand U29101 (N_29101,N_26044,N_25105);
nor U29102 (N_29102,N_26864,N_26645);
and U29103 (N_29103,N_25780,N_24610);
xnor U29104 (N_29104,N_24092,N_24783);
nand U29105 (N_29105,N_24879,N_24072);
or U29106 (N_29106,N_26279,N_24391);
and U29107 (N_29107,N_24595,N_24664);
or U29108 (N_29108,N_26593,N_26608);
nor U29109 (N_29109,N_24154,N_24803);
or U29110 (N_29110,N_25546,N_24945);
xnor U29111 (N_29111,N_24198,N_26355);
or U29112 (N_29112,N_24410,N_25043);
nand U29113 (N_29113,N_26558,N_25247);
nand U29114 (N_29114,N_26607,N_25915);
and U29115 (N_29115,N_26756,N_25467);
and U29116 (N_29116,N_26698,N_25885);
or U29117 (N_29117,N_26331,N_25318);
and U29118 (N_29118,N_25410,N_26068);
or U29119 (N_29119,N_24421,N_24994);
xor U29120 (N_29120,N_25622,N_24332);
or U29121 (N_29121,N_24936,N_25379);
xnor U29122 (N_29122,N_24480,N_25677);
xnor U29123 (N_29123,N_24685,N_25033);
nand U29124 (N_29124,N_26454,N_24121);
nor U29125 (N_29125,N_24032,N_24677);
nand U29126 (N_29126,N_25856,N_24847);
or U29127 (N_29127,N_25869,N_26069);
nor U29128 (N_29128,N_24465,N_26080);
nor U29129 (N_29129,N_26146,N_25215);
xor U29130 (N_29130,N_24166,N_25615);
nand U29131 (N_29131,N_25366,N_25745);
nand U29132 (N_29132,N_24152,N_26683);
xnor U29133 (N_29133,N_26447,N_26504);
nand U29134 (N_29134,N_25194,N_24470);
nor U29135 (N_29135,N_24434,N_26338);
and U29136 (N_29136,N_26252,N_24173);
xnor U29137 (N_29137,N_26739,N_26983);
nor U29138 (N_29138,N_26490,N_26894);
nand U29139 (N_29139,N_25030,N_25898);
nand U29140 (N_29140,N_24390,N_25772);
xnor U29141 (N_29141,N_24330,N_26565);
or U29142 (N_29142,N_24070,N_25372);
nand U29143 (N_29143,N_25930,N_24443);
nand U29144 (N_29144,N_24342,N_26022);
nand U29145 (N_29145,N_25957,N_25271);
nand U29146 (N_29146,N_26155,N_26293);
or U29147 (N_29147,N_25811,N_24422);
and U29148 (N_29148,N_26090,N_26021);
nor U29149 (N_29149,N_25869,N_24416);
or U29150 (N_29150,N_25132,N_25463);
xor U29151 (N_29151,N_26007,N_25639);
and U29152 (N_29152,N_26065,N_25495);
or U29153 (N_29153,N_26103,N_24323);
nor U29154 (N_29154,N_25116,N_26307);
nor U29155 (N_29155,N_25672,N_25407);
and U29156 (N_29156,N_24618,N_25740);
nor U29157 (N_29157,N_26524,N_25968);
nand U29158 (N_29158,N_26878,N_26531);
nand U29159 (N_29159,N_25251,N_24044);
or U29160 (N_29160,N_26300,N_25806);
and U29161 (N_29161,N_25464,N_24565);
nand U29162 (N_29162,N_24601,N_25822);
nand U29163 (N_29163,N_26674,N_25848);
xor U29164 (N_29164,N_26232,N_25754);
nand U29165 (N_29165,N_25707,N_25463);
xnor U29166 (N_29166,N_26676,N_25683);
nand U29167 (N_29167,N_24571,N_25112);
nand U29168 (N_29168,N_26177,N_24206);
or U29169 (N_29169,N_25192,N_26586);
or U29170 (N_29170,N_25292,N_26428);
xor U29171 (N_29171,N_26284,N_25089);
or U29172 (N_29172,N_26532,N_26145);
and U29173 (N_29173,N_25706,N_24142);
xnor U29174 (N_29174,N_26334,N_24333);
nor U29175 (N_29175,N_24962,N_24751);
nand U29176 (N_29176,N_25132,N_26454);
or U29177 (N_29177,N_24319,N_24105);
nand U29178 (N_29178,N_24913,N_26959);
and U29179 (N_29179,N_24868,N_25093);
nand U29180 (N_29180,N_26739,N_24931);
nand U29181 (N_29181,N_24144,N_26124);
xor U29182 (N_29182,N_26902,N_24180);
nand U29183 (N_29183,N_24255,N_24646);
xnor U29184 (N_29184,N_24426,N_24613);
or U29185 (N_29185,N_25406,N_26298);
and U29186 (N_29186,N_26836,N_24383);
and U29187 (N_29187,N_24307,N_24490);
xor U29188 (N_29188,N_26112,N_24561);
nor U29189 (N_29189,N_26471,N_26961);
xor U29190 (N_29190,N_25188,N_24326);
xor U29191 (N_29191,N_25001,N_24708);
xor U29192 (N_29192,N_24965,N_25307);
or U29193 (N_29193,N_26684,N_25946);
or U29194 (N_29194,N_26336,N_25631);
nor U29195 (N_29195,N_25736,N_25958);
or U29196 (N_29196,N_25179,N_24594);
xor U29197 (N_29197,N_26695,N_25730);
or U29198 (N_29198,N_25535,N_24967);
and U29199 (N_29199,N_26496,N_26562);
nand U29200 (N_29200,N_25618,N_24427);
nand U29201 (N_29201,N_25273,N_24244);
xnor U29202 (N_29202,N_25882,N_25286);
nor U29203 (N_29203,N_26106,N_24626);
nor U29204 (N_29204,N_24791,N_24878);
xnor U29205 (N_29205,N_24678,N_24212);
nand U29206 (N_29206,N_24490,N_24219);
or U29207 (N_29207,N_25109,N_24829);
xnor U29208 (N_29208,N_24369,N_25720);
nor U29209 (N_29209,N_24186,N_25246);
and U29210 (N_29210,N_24084,N_25596);
nor U29211 (N_29211,N_25664,N_24009);
nand U29212 (N_29212,N_26128,N_25057);
nor U29213 (N_29213,N_26191,N_26173);
nand U29214 (N_29214,N_26743,N_24009);
xor U29215 (N_29215,N_26061,N_24480);
nor U29216 (N_29216,N_25159,N_24037);
and U29217 (N_29217,N_26598,N_25089);
or U29218 (N_29218,N_24696,N_26269);
or U29219 (N_29219,N_26627,N_26725);
xnor U29220 (N_29220,N_25478,N_24374);
and U29221 (N_29221,N_24860,N_25710);
nor U29222 (N_29222,N_26370,N_25858);
nand U29223 (N_29223,N_24100,N_26444);
nand U29224 (N_29224,N_24413,N_26467);
and U29225 (N_29225,N_24704,N_24523);
xnor U29226 (N_29226,N_26467,N_26119);
nand U29227 (N_29227,N_24881,N_24691);
and U29228 (N_29228,N_25158,N_24239);
nand U29229 (N_29229,N_26587,N_25065);
or U29230 (N_29230,N_25271,N_25991);
nor U29231 (N_29231,N_25169,N_25823);
and U29232 (N_29232,N_24813,N_24278);
xor U29233 (N_29233,N_26367,N_24010);
nand U29234 (N_29234,N_24308,N_25513);
or U29235 (N_29235,N_24459,N_24914);
and U29236 (N_29236,N_25802,N_24282);
or U29237 (N_29237,N_26154,N_24576);
nand U29238 (N_29238,N_24333,N_24234);
and U29239 (N_29239,N_24293,N_24301);
nand U29240 (N_29240,N_26468,N_25689);
xor U29241 (N_29241,N_26959,N_24318);
nand U29242 (N_29242,N_26148,N_24938);
nor U29243 (N_29243,N_24655,N_24980);
or U29244 (N_29244,N_25468,N_24030);
or U29245 (N_29245,N_26825,N_25014);
nand U29246 (N_29246,N_26140,N_25504);
xor U29247 (N_29247,N_24784,N_25672);
or U29248 (N_29248,N_24993,N_24347);
and U29249 (N_29249,N_24393,N_24021);
nor U29250 (N_29250,N_24590,N_26295);
and U29251 (N_29251,N_24951,N_24826);
xnor U29252 (N_29252,N_24108,N_24755);
xnor U29253 (N_29253,N_25840,N_25248);
or U29254 (N_29254,N_25328,N_25909);
and U29255 (N_29255,N_24243,N_25667);
or U29256 (N_29256,N_26883,N_25548);
xnor U29257 (N_29257,N_25678,N_24632);
nor U29258 (N_29258,N_26793,N_26107);
xnor U29259 (N_29259,N_26434,N_26960);
nor U29260 (N_29260,N_25368,N_26783);
nor U29261 (N_29261,N_26661,N_24777);
xnor U29262 (N_29262,N_24531,N_25312);
xor U29263 (N_29263,N_26156,N_24655);
or U29264 (N_29264,N_26116,N_24930);
nor U29265 (N_29265,N_26327,N_26982);
nand U29266 (N_29266,N_24080,N_26473);
nor U29267 (N_29267,N_26534,N_25637);
xor U29268 (N_29268,N_24649,N_26699);
nand U29269 (N_29269,N_25780,N_25445);
or U29270 (N_29270,N_26416,N_24931);
and U29271 (N_29271,N_25794,N_26534);
and U29272 (N_29272,N_25787,N_24877);
or U29273 (N_29273,N_24865,N_26708);
xor U29274 (N_29274,N_25439,N_25561);
xor U29275 (N_29275,N_26105,N_24645);
or U29276 (N_29276,N_26926,N_24100);
xor U29277 (N_29277,N_24852,N_26143);
xor U29278 (N_29278,N_25873,N_26801);
or U29279 (N_29279,N_24937,N_25854);
and U29280 (N_29280,N_26777,N_25762);
or U29281 (N_29281,N_24455,N_25019);
nor U29282 (N_29282,N_26276,N_24006);
and U29283 (N_29283,N_24667,N_25552);
nand U29284 (N_29284,N_25208,N_26445);
nand U29285 (N_29285,N_24764,N_26444);
nand U29286 (N_29286,N_25610,N_25163);
or U29287 (N_29287,N_24151,N_24626);
and U29288 (N_29288,N_25170,N_24240);
or U29289 (N_29289,N_26512,N_24532);
xor U29290 (N_29290,N_24060,N_25674);
nand U29291 (N_29291,N_25259,N_24939);
nand U29292 (N_29292,N_24184,N_25751);
and U29293 (N_29293,N_25608,N_26531);
xnor U29294 (N_29294,N_24173,N_26376);
xnor U29295 (N_29295,N_26719,N_24737);
nand U29296 (N_29296,N_24513,N_24718);
xnor U29297 (N_29297,N_26902,N_25144);
nor U29298 (N_29298,N_26409,N_25528);
nand U29299 (N_29299,N_26907,N_24416);
and U29300 (N_29300,N_24279,N_24654);
xnor U29301 (N_29301,N_26110,N_25523);
nand U29302 (N_29302,N_24033,N_26533);
and U29303 (N_29303,N_25204,N_25295);
nand U29304 (N_29304,N_25949,N_25876);
nand U29305 (N_29305,N_26378,N_24476);
or U29306 (N_29306,N_26712,N_24664);
nor U29307 (N_29307,N_25807,N_24089);
or U29308 (N_29308,N_25192,N_25896);
xnor U29309 (N_29309,N_26435,N_25972);
nand U29310 (N_29310,N_26443,N_26548);
and U29311 (N_29311,N_24664,N_25092);
nor U29312 (N_29312,N_26341,N_26193);
or U29313 (N_29313,N_25728,N_25251);
or U29314 (N_29314,N_24004,N_26552);
nand U29315 (N_29315,N_26318,N_25463);
xor U29316 (N_29316,N_24281,N_26413);
nor U29317 (N_29317,N_25271,N_25652);
xnor U29318 (N_29318,N_24992,N_26973);
xnor U29319 (N_29319,N_26560,N_25727);
or U29320 (N_29320,N_25534,N_24956);
nor U29321 (N_29321,N_25578,N_26901);
nand U29322 (N_29322,N_25160,N_25546);
or U29323 (N_29323,N_26698,N_26076);
nor U29324 (N_29324,N_26020,N_24965);
nor U29325 (N_29325,N_26689,N_24499);
nor U29326 (N_29326,N_25549,N_26321);
and U29327 (N_29327,N_24346,N_26727);
nor U29328 (N_29328,N_26966,N_24146);
nor U29329 (N_29329,N_24880,N_25070);
or U29330 (N_29330,N_24842,N_24450);
nor U29331 (N_29331,N_24125,N_26430);
xnor U29332 (N_29332,N_25846,N_26608);
and U29333 (N_29333,N_26678,N_25199);
nand U29334 (N_29334,N_24233,N_24668);
nand U29335 (N_29335,N_24272,N_26729);
nor U29336 (N_29336,N_26504,N_24195);
and U29337 (N_29337,N_26860,N_24130);
nor U29338 (N_29338,N_26637,N_26509);
nand U29339 (N_29339,N_24999,N_26571);
and U29340 (N_29340,N_26607,N_24988);
or U29341 (N_29341,N_24100,N_24936);
and U29342 (N_29342,N_25954,N_25453);
and U29343 (N_29343,N_25758,N_26505);
and U29344 (N_29344,N_24026,N_26090);
and U29345 (N_29345,N_24996,N_26846);
xnor U29346 (N_29346,N_26390,N_25018);
nand U29347 (N_29347,N_24121,N_26484);
and U29348 (N_29348,N_25654,N_24474);
or U29349 (N_29349,N_25818,N_24017);
nor U29350 (N_29350,N_25024,N_25839);
and U29351 (N_29351,N_26996,N_26826);
and U29352 (N_29352,N_26409,N_25992);
nor U29353 (N_29353,N_26748,N_25626);
or U29354 (N_29354,N_26312,N_25909);
or U29355 (N_29355,N_24729,N_26373);
nand U29356 (N_29356,N_25763,N_26140);
xnor U29357 (N_29357,N_24442,N_26555);
or U29358 (N_29358,N_25997,N_25850);
and U29359 (N_29359,N_26910,N_24376);
nor U29360 (N_29360,N_25509,N_24390);
xnor U29361 (N_29361,N_26849,N_25288);
and U29362 (N_29362,N_24071,N_24506);
nand U29363 (N_29363,N_26462,N_24519);
xnor U29364 (N_29364,N_26167,N_26692);
nand U29365 (N_29365,N_24783,N_26400);
nor U29366 (N_29366,N_24898,N_24464);
and U29367 (N_29367,N_24623,N_24642);
nand U29368 (N_29368,N_26086,N_24424);
nand U29369 (N_29369,N_25194,N_25499);
nor U29370 (N_29370,N_25970,N_26692);
xnor U29371 (N_29371,N_24768,N_26757);
nor U29372 (N_29372,N_25598,N_25949);
nand U29373 (N_29373,N_25048,N_25616);
and U29374 (N_29374,N_26914,N_25051);
nor U29375 (N_29375,N_25968,N_26592);
nor U29376 (N_29376,N_25138,N_25218);
or U29377 (N_29377,N_25306,N_26814);
nand U29378 (N_29378,N_26839,N_26950);
or U29379 (N_29379,N_26018,N_24530);
nand U29380 (N_29380,N_24830,N_25317);
nand U29381 (N_29381,N_25185,N_25478);
or U29382 (N_29382,N_24482,N_26781);
xnor U29383 (N_29383,N_24414,N_26409);
or U29384 (N_29384,N_26551,N_25929);
nor U29385 (N_29385,N_24824,N_24892);
nor U29386 (N_29386,N_24488,N_26815);
or U29387 (N_29387,N_24968,N_26527);
and U29388 (N_29388,N_24906,N_25082);
and U29389 (N_29389,N_26151,N_24466);
or U29390 (N_29390,N_25797,N_24322);
and U29391 (N_29391,N_25358,N_26054);
and U29392 (N_29392,N_26143,N_26038);
xnor U29393 (N_29393,N_25339,N_26595);
xnor U29394 (N_29394,N_26446,N_26065);
and U29395 (N_29395,N_25730,N_24508);
or U29396 (N_29396,N_26725,N_26327);
nor U29397 (N_29397,N_26462,N_25378);
nand U29398 (N_29398,N_24710,N_24963);
nand U29399 (N_29399,N_25004,N_26163);
nor U29400 (N_29400,N_24123,N_26492);
nor U29401 (N_29401,N_24621,N_25719);
xnor U29402 (N_29402,N_24794,N_26722);
nor U29403 (N_29403,N_24867,N_26467);
and U29404 (N_29404,N_24410,N_26820);
nand U29405 (N_29405,N_25090,N_24939);
or U29406 (N_29406,N_25922,N_25000);
xnor U29407 (N_29407,N_26026,N_25064);
or U29408 (N_29408,N_26088,N_26027);
and U29409 (N_29409,N_24877,N_24940);
or U29410 (N_29410,N_25138,N_26919);
xnor U29411 (N_29411,N_24842,N_25987);
nor U29412 (N_29412,N_24703,N_24152);
nand U29413 (N_29413,N_26306,N_26296);
and U29414 (N_29414,N_26384,N_24403);
xor U29415 (N_29415,N_24785,N_25222);
or U29416 (N_29416,N_25538,N_25438);
or U29417 (N_29417,N_26448,N_26714);
nand U29418 (N_29418,N_26346,N_26937);
or U29419 (N_29419,N_26094,N_25087);
xor U29420 (N_29420,N_25205,N_25477);
nand U29421 (N_29421,N_24074,N_24380);
nor U29422 (N_29422,N_26590,N_26264);
nand U29423 (N_29423,N_25822,N_25670);
nand U29424 (N_29424,N_26276,N_24255);
nor U29425 (N_29425,N_25480,N_26904);
and U29426 (N_29426,N_26700,N_26061);
nor U29427 (N_29427,N_25174,N_25967);
xor U29428 (N_29428,N_25604,N_25840);
or U29429 (N_29429,N_25790,N_26067);
and U29430 (N_29430,N_25957,N_26950);
nor U29431 (N_29431,N_25773,N_26277);
xnor U29432 (N_29432,N_26250,N_25777);
nor U29433 (N_29433,N_26687,N_25863);
nor U29434 (N_29434,N_24762,N_26778);
nand U29435 (N_29435,N_24328,N_24078);
and U29436 (N_29436,N_26813,N_25993);
xor U29437 (N_29437,N_24048,N_25274);
nor U29438 (N_29438,N_26760,N_25491);
or U29439 (N_29439,N_25268,N_24520);
xor U29440 (N_29440,N_24524,N_25520);
or U29441 (N_29441,N_24954,N_26613);
or U29442 (N_29442,N_25347,N_25708);
nor U29443 (N_29443,N_26288,N_24013);
and U29444 (N_29444,N_25607,N_24301);
xnor U29445 (N_29445,N_26136,N_25130);
nand U29446 (N_29446,N_26891,N_26879);
or U29447 (N_29447,N_26712,N_24832);
or U29448 (N_29448,N_26806,N_25559);
nor U29449 (N_29449,N_24140,N_26141);
nand U29450 (N_29450,N_26958,N_25807);
nand U29451 (N_29451,N_26756,N_26821);
and U29452 (N_29452,N_24961,N_25312);
or U29453 (N_29453,N_26857,N_24919);
and U29454 (N_29454,N_26675,N_25647);
nor U29455 (N_29455,N_24995,N_26299);
xor U29456 (N_29456,N_26404,N_25728);
or U29457 (N_29457,N_24031,N_25664);
nor U29458 (N_29458,N_24385,N_25840);
xnor U29459 (N_29459,N_25883,N_25431);
and U29460 (N_29460,N_26112,N_25194);
nand U29461 (N_29461,N_24428,N_25182);
and U29462 (N_29462,N_24790,N_26746);
xor U29463 (N_29463,N_24775,N_25200);
xor U29464 (N_29464,N_26912,N_26992);
or U29465 (N_29465,N_26344,N_25981);
and U29466 (N_29466,N_24355,N_24177);
or U29467 (N_29467,N_25899,N_26820);
nor U29468 (N_29468,N_25997,N_24885);
xnor U29469 (N_29469,N_25514,N_25596);
or U29470 (N_29470,N_25600,N_24784);
nor U29471 (N_29471,N_24965,N_25266);
nand U29472 (N_29472,N_25215,N_24056);
nor U29473 (N_29473,N_25402,N_25898);
or U29474 (N_29474,N_25488,N_26973);
nand U29475 (N_29475,N_26971,N_24471);
or U29476 (N_29476,N_25661,N_25043);
nor U29477 (N_29477,N_24533,N_24625);
xor U29478 (N_29478,N_24590,N_24260);
nor U29479 (N_29479,N_26052,N_24360);
xnor U29480 (N_29480,N_26921,N_25182);
or U29481 (N_29481,N_25192,N_26963);
nor U29482 (N_29482,N_26945,N_25148);
and U29483 (N_29483,N_24767,N_26590);
or U29484 (N_29484,N_25844,N_26469);
xnor U29485 (N_29485,N_24501,N_26007);
nor U29486 (N_29486,N_26367,N_25903);
xor U29487 (N_29487,N_26819,N_24432);
nor U29488 (N_29488,N_25178,N_25116);
or U29489 (N_29489,N_26418,N_25631);
and U29490 (N_29490,N_25242,N_24163);
xnor U29491 (N_29491,N_25721,N_26204);
and U29492 (N_29492,N_26459,N_24799);
xnor U29493 (N_29493,N_26585,N_24928);
or U29494 (N_29494,N_26499,N_26752);
or U29495 (N_29495,N_25102,N_24084);
xnor U29496 (N_29496,N_25475,N_25264);
and U29497 (N_29497,N_25317,N_25636);
nand U29498 (N_29498,N_26874,N_24012);
nor U29499 (N_29499,N_26248,N_25250);
and U29500 (N_29500,N_24630,N_25053);
or U29501 (N_29501,N_25668,N_25799);
nand U29502 (N_29502,N_24312,N_26081);
and U29503 (N_29503,N_25883,N_25044);
or U29504 (N_29504,N_26470,N_25177);
and U29505 (N_29505,N_25331,N_25582);
xnor U29506 (N_29506,N_26818,N_26582);
xor U29507 (N_29507,N_25456,N_26705);
xor U29508 (N_29508,N_24293,N_24149);
and U29509 (N_29509,N_25084,N_24449);
or U29510 (N_29510,N_24582,N_26804);
or U29511 (N_29511,N_26977,N_24416);
nor U29512 (N_29512,N_26251,N_25099);
and U29513 (N_29513,N_25930,N_26559);
nor U29514 (N_29514,N_25267,N_25282);
nor U29515 (N_29515,N_26119,N_24992);
nor U29516 (N_29516,N_25642,N_25076);
and U29517 (N_29517,N_24856,N_26788);
or U29518 (N_29518,N_24694,N_24451);
nand U29519 (N_29519,N_26268,N_26995);
xnor U29520 (N_29520,N_24986,N_24927);
nand U29521 (N_29521,N_24243,N_24658);
nand U29522 (N_29522,N_24861,N_25058);
nand U29523 (N_29523,N_25590,N_24223);
nand U29524 (N_29524,N_25513,N_26547);
nand U29525 (N_29525,N_24780,N_26949);
nor U29526 (N_29526,N_24962,N_26244);
and U29527 (N_29527,N_26454,N_25557);
xnor U29528 (N_29528,N_26053,N_24710);
or U29529 (N_29529,N_24176,N_24095);
xor U29530 (N_29530,N_26813,N_25874);
or U29531 (N_29531,N_26300,N_24573);
nand U29532 (N_29532,N_25226,N_24205);
nand U29533 (N_29533,N_25208,N_25348);
or U29534 (N_29534,N_24096,N_26655);
or U29535 (N_29535,N_24649,N_24262);
or U29536 (N_29536,N_24668,N_25541);
nor U29537 (N_29537,N_24932,N_24524);
nor U29538 (N_29538,N_25603,N_25507);
nor U29539 (N_29539,N_24858,N_24849);
or U29540 (N_29540,N_26189,N_26227);
nor U29541 (N_29541,N_25443,N_24351);
nand U29542 (N_29542,N_26195,N_26865);
or U29543 (N_29543,N_25377,N_25601);
and U29544 (N_29544,N_25529,N_26771);
or U29545 (N_29545,N_24473,N_24622);
or U29546 (N_29546,N_26478,N_25240);
or U29547 (N_29547,N_25274,N_24425);
and U29548 (N_29548,N_26185,N_26747);
and U29549 (N_29549,N_24179,N_26985);
nor U29550 (N_29550,N_24246,N_26133);
nand U29551 (N_29551,N_24579,N_24985);
nor U29552 (N_29552,N_25037,N_25020);
and U29553 (N_29553,N_24839,N_26117);
or U29554 (N_29554,N_25174,N_25121);
and U29555 (N_29555,N_25909,N_25928);
and U29556 (N_29556,N_24166,N_25514);
nor U29557 (N_29557,N_25913,N_24177);
and U29558 (N_29558,N_26454,N_25883);
xnor U29559 (N_29559,N_24552,N_25995);
xor U29560 (N_29560,N_26414,N_26208);
or U29561 (N_29561,N_25227,N_24460);
xor U29562 (N_29562,N_25343,N_25084);
nand U29563 (N_29563,N_26070,N_25792);
or U29564 (N_29564,N_24830,N_24467);
or U29565 (N_29565,N_26697,N_25386);
or U29566 (N_29566,N_25053,N_25305);
xor U29567 (N_29567,N_24301,N_24406);
nor U29568 (N_29568,N_26905,N_24118);
nand U29569 (N_29569,N_24306,N_25323);
and U29570 (N_29570,N_26246,N_24678);
xor U29571 (N_29571,N_25111,N_26218);
or U29572 (N_29572,N_24702,N_26925);
nor U29573 (N_29573,N_24930,N_24719);
or U29574 (N_29574,N_26641,N_25728);
xnor U29575 (N_29575,N_24643,N_26260);
or U29576 (N_29576,N_26844,N_26360);
nor U29577 (N_29577,N_25226,N_26359);
nand U29578 (N_29578,N_24118,N_25148);
nand U29579 (N_29579,N_25435,N_25897);
or U29580 (N_29580,N_25397,N_25151);
or U29581 (N_29581,N_25613,N_24038);
nor U29582 (N_29582,N_26546,N_25124);
nor U29583 (N_29583,N_24196,N_26393);
nor U29584 (N_29584,N_26657,N_24129);
nand U29585 (N_29585,N_24671,N_25963);
xor U29586 (N_29586,N_24394,N_24779);
nand U29587 (N_29587,N_25608,N_26694);
nor U29588 (N_29588,N_26129,N_25559);
xor U29589 (N_29589,N_26599,N_25116);
xnor U29590 (N_29590,N_24306,N_26986);
nor U29591 (N_29591,N_26094,N_24904);
nor U29592 (N_29592,N_25448,N_24527);
or U29593 (N_29593,N_26254,N_24690);
or U29594 (N_29594,N_24150,N_25688);
nor U29595 (N_29595,N_24290,N_24190);
xor U29596 (N_29596,N_25714,N_26929);
and U29597 (N_29597,N_25568,N_26735);
or U29598 (N_29598,N_25236,N_26145);
and U29599 (N_29599,N_25814,N_26867);
xnor U29600 (N_29600,N_25808,N_25231);
or U29601 (N_29601,N_24132,N_25356);
nand U29602 (N_29602,N_25819,N_26311);
or U29603 (N_29603,N_26803,N_26521);
nor U29604 (N_29604,N_25532,N_24835);
nor U29605 (N_29605,N_25018,N_26852);
or U29606 (N_29606,N_24823,N_25226);
nand U29607 (N_29607,N_26064,N_24999);
xor U29608 (N_29608,N_26684,N_25537);
xor U29609 (N_29609,N_26034,N_24217);
nor U29610 (N_29610,N_25980,N_24668);
xor U29611 (N_29611,N_26333,N_25378);
and U29612 (N_29612,N_25843,N_24049);
nand U29613 (N_29613,N_25441,N_25861);
nor U29614 (N_29614,N_25195,N_25078);
nand U29615 (N_29615,N_25107,N_24567);
or U29616 (N_29616,N_25414,N_24444);
nor U29617 (N_29617,N_25749,N_26723);
nand U29618 (N_29618,N_25084,N_25719);
nor U29619 (N_29619,N_24018,N_25527);
nor U29620 (N_29620,N_26780,N_25102);
nor U29621 (N_29621,N_25408,N_25519);
nand U29622 (N_29622,N_24942,N_25515);
nor U29623 (N_29623,N_26209,N_26821);
xor U29624 (N_29624,N_26536,N_25969);
nand U29625 (N_29625,N_26659,N_24854);
xnor U29626 (N_29626,N_24354,N_26551);
nor U29627 (N_29627,N_25908,N_24432);
and U29628 (N_29628,N_25688,N_24156);
nor U29629 (N_29629,N_26791,N_25061);
or U29630 (N_29630,N_26237,N_26894);
and U29631 (N_29631,N_25236,N_24812);
nand U29632 (N_29632,N_25534,N_26755);
or U29633 (N_29633,N_26889,N_24181);
or U29634 (N_29634,N_25666,N_26405);
nand U29635 (N_29635,N_26493,N_25702);
or U29636 (N_29636,N_26753,N_24153);
and U29637 (N_29637,N_26793,N_26284);
xor U29638 (N_29638,N_25906,N_24002);
and U29639 (N_29639,N_25016,N_26020);
nand U29640 (N_29640,N_24632,N_25046);
and U29641 (N_29641,N_26952,N_26430);
xor U29642 (N_29642,N_25145,N_24642);
xor U29643 (N_29643,N_26863,N_26455);
nand U29644 (N_29644,N_26118,N_24987);
or U29645 (N_29645,N_24379,N_24908);
or U29646 (N_29646,N_26437,N_25030);
nand U29647 (N_29647,N_24975,N_26735);
xnor U29648 (N_29648,N_24594,N_25744);
or U29649 (N_29649,N_26637,N_25974);
xnor U29650 (N_29650,N_25072,N_26112);
nor U29651 (N_29651,N_26319,N_24894);
nand U29652 (N_29652,N_24790,N_25496);
nor U29653 (N_29653,N_25297,N_26572);
xnor U29654 (N_29654,N_26108,N_26010);
nand U29655 (N_29655,N_25589,N_26239);
xor U29656 (N_29656,N_26462,N_24032);
and U29657 (N_29657,N_26527,N_25446);
nor U29658 (N_29658,N_26731,N_24950);
nor U29659 (N_29659,N_24432,N_26993);
and U29660 (N_29660,N_26123,N_26697);
or U29661 (N_29661,N_25833,N_25716);
nor U29662 (N_29662,N_25332,N_25478);
xor U29663 (N_29663,N_25323,N_25625);
or U29664 (N_29664,N_26295,N_25282);
nor U29665 (N_29665,N_26568,N_24161);
or U29666 (N_29666,N_24716,N_26717);
nand U29667 (N_29667,N_24953,N_25029);
and U29668 (N_29668,N_24225,N_25875);
nor U29669 (N_29669,N_24016,N_25216);
nand U29670 (N_29670,N_26718,N_24975);
or U29671 (N_29671,N_24915,N_26050);
nor U29672 (N_29672,N_24774,N_26404);
nand U29673 (N_29673,N_24166,N_26580);
nor U29674 (N_29674,N_25685,N_26873);
xor U29675 (N_29675,N_24909,N_25904);
nand U29676 (N_29676,N_26855,N_24609);
nand U29677 (N_29677,N_26242,N_24374);
xnor U29678 (N_29678,N_26726,N_25339);
xor U29679 (N_29679,N_26290,N_26695);
xnor U29680 (N_29680,N_24920,N_25372);
and U29681 (N_29681,N_24765,N_25011);
or U29682 (N_29682,N_26838,N_26078);
nand U29683 (N_29683,N_26022,N_24575);
xnor U29684 (N_29684,N_26939,N_25708);
nand U29685 (N_29685,N_26967,N_25784);
and U29686 (N_29686,N_26109,N_24922);
or U29687 (N_29687,N_26789,N_25186);
and U29688 (N_29688,N_25677,N_25691);
or U29689 (N_29689,N_25248,N_26502);
nand U29690 (N_29690,N_24000,N_25021);
and U29691 (N_29691,N_26010,N_24909);
xor U29692 (N_29692,N_24878,N_25445);
nor U29693 (N_29693,N_25548,N_25738);
or U29694 (N_29694,N_26292,N_24746);
nor U29695 (N_29695,N_26468,N_25630);
xnor U29696 (N_29696,N_25252,N_25837);
xor U29697 (N_29697,N_24707,N_26738);
and U29698 (N_29698,N_26000,N_25646);
xor U29699 (N_29699,N_25984,N_24167);
or U29700 (N_29700,N_25878,N_26217);
xor U29701 (N_29701,N_25528,N_25872);
nand U29702 (N_29702,N_25935,N_25049);
or U29703 (N_29703,N_26320,N_24950);
or U29704 (N_29704,N_26186,N_24150);
and U29705 (N_29705,N_25436,N_26023);
nor U29706 (N_29706,N_25329,N_25957);
and U29707 (N_29707,N_25624,N_26030);
nor U29708 (N_29708,N_24248,N_25954);
xnor U29709 (N_29709,N_25115,N_24144);
or U29710 (N_29710,N_25002,N_24373);
or U29711 (N_29711,N_24667,N_25360);
or U29712 (N_29712,N_26695,N_26189);
nor U29713 (N_29713,N_26769,N_26701);
nand U29714 (N_29714,N_26476,N_26976);
nand U29715 (N_29715,N_25499,N_25160);
nand U29716 (N_29716,N_24450,N_26688);
and U29717 (N_29717,N_25920,N_26512);
nand U29718 (N_29718,N_26227,N_24856);
xor U29719 (N_29719,N_25225,N_24964);
nand U29720 (N_29720,N_24716,N_24163);
xnor U29721 (N_29721,N_25380,N_24374);
or U29722 (N_29722,N_24368,N_25925);
or U29723 (N_29723,N_26390,N_26953);
nand U29724 (N_29724,N_26236,N_26994);
and U29725 (N_29725,N_24220,N_24593);
and U29726 (N_29726,N_25025,N_26032);
nor U29727 (N_29727,N_25987,N_25048);
xnor U29728 (N_29728,N_25030,N_26093);
or U29729 (N_29729,N_26353,N_24066);
nand U29730 (N_29730,N_24471,N_24567);
or U29731 (N_29731,N_25500,N_26181);
or U29732 (N_29732,N_26426,N_26256);
and U29733 (N_29733,N_24809,N_24951);
xnor U29734 (N_29734,N_26759,N_25553);
nor U29735 (N_29735,N_25069,N_25649);
nor U29736 (N_29736,N_26974,N_25793);
xnor U29737 (N_29737,N_24618,N_24135);
nand U29738 (N_29738,N_25090,N_25848);
nand U29739 (N_29739,N_24433,N_26150);
or U29740 (N_29740,N_25370,N_24276);
nor U29741 (N_29741,N_24735,N_26134);
and U29742 (N_29742,N_26345,N_24268);
nand U29743 (N_29743,N_24222,N_26363);
and U29744 (N_29744,N_25695,N_24591);
nand U29745 (N_29745,N_24591,N_26394);
xor U29746 (N_29746,N_25595,N_25514);
and U29747 (N_29747,N_26215,N_26927);
nor U29748 (N_29748,N_24372,N_25386);
or U29749 (N_29749,N_26367,N_26891);
nand U29750 (N_29750,N_25483,N_26269);
xor U29751 (N_29751,N_24334,N_24113);
or U29752 (N_29752,N_24924,N_24449);
or U29753 (N_29753,N_25015,N_24927);
nor U29754 (N_29754,N_25139,N_25068);
nand U29755 (N_29755,N_25360,N_24084);
xor U29756 (N_29756,N_25219,N_26509);
and U29757 (N_29757,N_24869,N_26302);
and U29758 (N_29758,N_26231,N_26438);
or U29759 (N_29759,N_26620,N_25717);
nor U29760 (N_29760,N_25564,N_26261);
xnor U29761 (N_29761,N_24608,N_26021);
and U29762 (N_29762,N_25065,N_26909);
xor U29763 (N_29763,N_26758,N_26375);
and U29764 (N_29764,N_25567,N_26886);
xor U29765 (N_29765,N_25001,N_24270);
and U29766 (N_29766,N_26658,N_26133);
nand U29767 (N_29767,N_24549,N_26988);
nand U29768 (N_29768,N_24463,N_24660);
or U29769 (N_29769,N_25509,N_24967);
and U29770 (N_29770,N_26340,N_24778);
xnor U29771 (N_29771,N_25601,N_24885);
nand U29772 (N_29772,N_25332,N_24758);
xor U29773 (N_29773,N_26548,N_26603);
nor U29774 (N_29774,N_25355,N_25934);
nand U29775 (N_29775,N_24546,N_25154);
and U29776 (N_29776,N_25998,N_25250);
or U29777 (N_29777,N_26524,N_25905);
nand U29778 (N_29778,N_25960,N_25444);
or U29779 (N_29779,N_25349,N_24536);
or U29780 (N_29780,N_25421,N_26702);
nor U29781 (N_29781,N_24314,N_25293);
and U29782 (N_29782,N_25780,N_24467);
nor U29783 (N_29783,N_25053,N_25711);
nand U29784 (N_29784,N_24995,N_25924);
nand U29785 (N_29785,N_26952,N_25222);
nor U29786 (N_29786,N_26189,N_26698);
nand U29787 (N_29787,N_25330,N_25116);
nor U29788 (N_29788,N_25276,N_25717);
nand U29789 (N_29789,N_26056,N_25046);
and U29790 (N_29790,N_26538,N_25909);
or U29791 (N_29791,N_24485,N_26241);
xnor U29792 (N_29792,N_25158,N_24120);
and U29793 (N_29793,N_25922,N_26151);
nand U29794 (N_29794,N_26701,N_26007);
xor U29795 (N_29795,N_26211,N_26711);
nand U29796 (N_29796,N_26980,N_26964);
xnor U29797 (N_29797,N_24006,N_26858);
and U29798 (N_29798,N_26797,N_26531);
and U29799 (N_29799,N_26064,N_25523);
and U29800 (N_29800,N_26953,N_26115);
nor U29801 (N_29801,N_26125,N_26050);
nand U29802 (N_29802,N_24020,N_25521);
nor U29803 (N_29803,N_24805,N_24176);
nor U29804 (N_29804,N_26208,N_26191);
and U29805 (N_29805,N_25628,N_24651);
and U29806 (N_29806,N_24572,N_26077);
or U29807 (N_29807,N_26562,N_25366);
or U29808 (N_29808,N_26736,N_26003);
and U29809 (N_29809,N_25385,N_25030);
xnor U29810 (N_29810,N_25698,N_25256);
xnor U29811 (N_29811,N_24326,N_25981);
and U29812 (N_29812,N_26500,N_26124);
and U29813 (N_29813,N_25597,N_25210);
xnor U29814 (N_29814,N_26160,N_25911);
nor U29815 (N_29815,N_25249,N_24592);
nand U29816 (N_29816,N_24397,N_24688);
nand U29817 (N_29817,N_25489,N_24052);
xor U29818 (N_29818,N_26463,N_25314);
xor U29819 (N_29819,N_25865,N_26127);
xnor U29820 (N_29820,N_26968,N_24289);
or U29821 (N_29821,N_24836,N_25710);
and U29822 (N_29822,N_26160,N_24173);
nand U29823 (N_29823,N_25277,N_25252);
and U29824 (N_29824,N_25538,N_24933);
nor U29825 (N_29825,N_25539,N_24908);
xnor U29826 (N_29826,N_26701,N_24778);
nor U29827 (N_29827,N_25427,N_25961);
nand U29828 (N_29828,N_24645,N_26889);
nand U29829 (N_29829,N_25284,N_24006);
nor U29830 (N_29830,N_25659,N_26371);
and U29831 (N_29831,N_26569,N_25534);
and U29832 (N_29832,N_24694,N_26620);
xnor U29833 (N_29833,N_25299,N_26904);
xnor U29834 (N_29834,N_24760,N_25009);
nor U29835 (N_29835,N_26733,N_24502);
nor U29836 (N_29836,N_24227,N_25123);
xnor U29837 (N_29837,N_26178,N_25747);
nand U29838 (N_29838,N_24624,N_26212);
xor U29839 (N_29839,N_26400,N_26344);
nand U29840 (N_29840,N_25846,N_24172);
nor U29841 (N_29841,N_25291,N_25544);
or U29842 (N_29842,N_24133,N_25028);
and U29843 (N_29843,N_25462,N_24125);
and U29844 (N_29844,N_24891,N_26872);
nand U29845 (N_29845,N_26049,N_25342);
nor U29846 (N_29846,N_24027,N_26360);
or U29847 (N_29847,N_24204,N_25399);
nand U29848 (N_29848,N_26886,N_24897);
and U29849 (N_29849,N_24234,N_26327);
nor U29850 (N_29850,N_24792,N_26860);
and U29851 (N_29851,N_25796,N_24664);
or U29852 (N_29852,N_26017,N_24984);
and U29853 (N_29853,N_24914,N_24952);
nor U29854 (N_29854,N_26922,N_25648);
nand U29855 (N_29855,N_24504,N_25698);
and U29856 (N_29856,N_26994,N_25963);
or U29857 (N_29857,N_24468,N_26107);
and U29858 (N_29858,N_25667,N_24985);
xor U29859 (N_29859,N_26701,N_26509);
xnor U29860 (N_29860,N_26978,N_25051);
nand U29861 (N_29861,N_24168,N_24856);
nand U29862 (N_29862,N_24131,N_26863);
nand U29863 (N_29863,N_25148,N_26069);
nor U29864 (N_29864,N_26482,N_24699);
nand U29865 (N_29865,N_26296,N_26039);
nand U29866 (N_29866,N_25719,N_26078);
and U29867 (N_29867,N_26903,N_25483);
nor U29868 (N_29868,N_26469,N_26834);
and U29869 (N_29869,N_25403,N_26765);
xnor U29870 (N_29870,N_26502,N_24804);
nor U29871 (N_29871,N_25068,N_26635);
and U29872 (N_29872,N_25960,N_24385);
and U29873 (N_29873,N_24592,N_26099);
nor U29874 (N_29874,N_26905,N_25706);
xor U29875 (N_29875,N_24386,N_26810);
nor U29876 (N_29876,N_26296,N_24062);
xor U29877 (N_29877,N_25610,N_25584);
or U29878 (N_29878,N_25537,N_26430);
nand U29879 (N_29879,N_25706,N_25785);
nand U29880 (N_29880,N_26871,N_26318);
nand U29881 (N_29881,N_25598,N_25701);
or U29882 (N_29882,N_25465,N_24601);
nand U29883 (N_29883,N_24740,N_25578);
xnor U29884 (N_29884,N_26956,N_25332);
nor U29885 (N_29885,N_26108,N_24362);
xnor U29886 (N_29886,N_26666,N_25574);
nor U29887 (N_29887,N_24784,N_24114);
nand U29888 (N_29888,N_24048,N_26668);
or U29889 (N_29889,N_24277,N_26412);
nor U29890 (N_29890,N_26632,N_24539);
xor U29891 (N_29891,N_24566,N_25474);
and U29892 (N_29892,N_26791,N_26801);
or U29893 (N_29893,N_26961,N_25598);
or U29894 (N_29894,N_24110,N_24029);
or U29895 (N_29895,N_24277,N_26349);
and U29896 (N_29896,N_25770,N_25756);
nand U29897 (N_29897,N_26934,N_25406);
xnor U29898 (N_29898,N_24103,N_26467);
and U29899 (N_29899,N_24444,N_26381);
or U29900 (N_29900,N_26395,N_25203);
or U29901 (N_29901,N_24076,N_26734);
nand U29902 (N_29902,N_25656,N_25821);
nand U29903 (N_29903,N_25313,N_26556);
nor U29904 (N_29904,N_24918,N_26442);
or U29905 (N_29905,N_24828,N_24488);
nand U29906 (N_29906,N_26581,N_25178);
xnor U29907 (N_29907,N_25035,N_25694);
nand U29908 (N_29908,N_24305,N_24049);
nor U29909 (N_29909,N_25416,N_24750);
nor U29910 (N_29910,N_25331,N_26825);
nor U29911 (N_29911,N_26184,N_24871);
nor U29912 (N_29912,N_24282,N_26227);
and U29913 (N_29913,N_26608,N_26759);
xnor U29914 (N_29914,N_25897,N_24469);
xnor U29915 (N_29915,N_26634,N_26829);
or U29916 (N_29916,N_25369,N_25502);
and U29917 (N_29917,N_25763,N_24590);
xor U29918 (N_29918,N_24556,N_26610);
and U29919 (N_29919,N_26034,N_24463);
nor U29920 (N_29920,N_25603,N_26946);
nand U29921 (N_29921,N_25255,N_25969);
nor U29922 (N_29922,N_26643,N_26788);
xnor U29923 (N_29923,N_25409,N_26550);
nor U29924 (N_29924,N_26716,N_26562);
nand U29925 (N_29925,N_25057,N_26255);
nor U29926 (N_29926,N_24347,N_26058);
and U29927 (N_29927,N_25107,N_26306);
xor U29928 (N_29928,N_25503,N_24007);
nor U29929 (N_29929,N_26501,N_24896);
nand U29930 (N_29930,N_25186,N_26241);
xnor U29931 (N_29931,N_24803,N_26636);
or U29932 (N_29932,N_26831,N_25026);
or U29933 (N_29933,N_26016,N_26424);
and U29934 (N_29934,N_26748,N_24756);
and U29935 (N_29935,N_26284,N_24323);
or U29936 (N_29936,N_26538,N_25505);
or U29937 (N_29937,N_25621,N_25825);
or U29938 (N_29938,N_24958,N_24625);
nor U29939 (N_29939,N_26291,N_25817);
nor U29940 (N_29940,N_24150,N_25827);
nor U29941 (N_29941,N_26187,N_26815);
or U29942 (N_29942,N_25223,N_25915);
nand U29943 (N_29943,N_25091,N_26526);
xor U29944 (N_29944,N_26014,N_24626);
and U29945 (N_29945,N_25310,N_26132);
xnor U29946 (N_29946,N_25243,N_25372);
nor U29947 (N_29947,N_24616,N_24508);
nand U29948 (N_29948,N_24852,N_26203);
nand U29949 (N_29949,N_24034,N_26570);
and U29950 (N_29950,N_25737,N_25374);
nand U29951 (N_29951,N_25966,N_26877);
or U29952 (N_29952,N_26492,N_26956);
nand U29953 (N_29953,N_24691,N_26381);
nand U29954 (N_29954,N_26360,N_25704);
nand U29955 (N_29955,N_24620,N_26126);
or U29956 (N_29956,N_24055,N_26343);
and U29957 (N_29957,N_26974,N_26087);
nand U29958 (N_29958,N_26634,N_24699);
and U29959 (N_29959,N_26462,N_26108);
xor U29960 (N_29960,N_25251,N_26309);
nand U29961 (N_29961,N_25946,N_24106);
nand U29962 (N_29962,N_24159,N_24404);
or U29963 (N_29963,N_24418,N_24041);
or U29964 (N_29964,N_25269,N_24537);
and U29965 (N_29965,N_24945,N_25343);
or U29966 (N_29966,N_24510,N_25368);
nand U29967 (N_29967,N_24883,N_24271);
nor U29968 (N_29968,N_24282,N_26223);
xnor U29969 (N_29969,N_24075,N_25348);
or U29970 (N_29970,N_24815,N_25039);
nor U29971 (N_29971,N_24320,N_26486);
xnor U29972 (N_29972,N_25261,N_25770);
xor U29973 (N_29973,N_25602,N_26065);
nand U29974 (N_29974,N_24272,N_26324);
or U29975 (N_29975,N_25911,N_24333);
xor U29976 (N_29976,N_25709,N_26910);
nor U29977 (N_29977,N_25420,N_26902);
nand U29978 (N_29978,N_24774,N_25558);
nand U29979 (N_29979,N_26540,N_26661);
nand U29980 (N_29980,N_24667,N_25515);
xnor U29981 (N_29981,N_26684,N_26381);
or U29982 (N_29982,N_26641,N_25654);
and U29983 (N_29983,N_26299,N_25390);
or U29984 (N_29984,N_25535,N_25615);
or U29985 (N_29985,N_25385,N_26546);
and U29986 (N_29986,N_26788,N_25991);
or U29987 (N_29987,N_24146,N_25406);
nand U29988 (N_29988,N_26281,N_24380);
nor U29989 (N_29989,N_26109,N_26782);
or U29990 (N_29990,N_25552,N_25706);
or U29991 (N_29991,N_26461,N_26921);
nand U29992 (N_29992,N_26249,N_24842);
nand U29993 (N_29993,N_25871,N_26868);
nor U29994 (N_29994,N_25726,N_24605);
nor U29995 (N_29995,N_24162,N_24935);
xor U29996 (N_29996,N_26375,N_26340);
or U29997 (N_29997,N_26983,N_24100);
nand U29998 (N_29998,N_24067,N_26695);
nand U29999 (N_29999,N_25625,N_24991);
xnor UO_0 (O_0,N_27570,N_27727);
nor UO_1 (O_1,N_28671,N_29805);
nand UO_2 (O_2,N_29964,N_27989);
and UO_3 (O_3,N_29660,N_28923);
and UO_4 (O_4,N_29701,N_29896);
nor UO_5 (O_5,N_27765,N_27962);
nand UO_6 (O_6,N_27612,N_28900);
and UO_7 (O_7,N_27928,N_27457);
nand UO_8 (O_8,N_28562,N_28784);
or UO_9 (O_9,N_29295,N_29301);
nand UO_10 (O_10,N_29387,N_27029);
and UO_11 (O_11,N_27346,N_27538);
or UO_12 (O_12,N_29210,N_27609);
and UO_13 (O_13,N_27806,N_28928);
and UO_14 (O_14,N_29405,N_29793);
xnor UO_15 (O_15,N_29895,N_27582);
or UO_16 (O_16,N_27172,N_28228);
and UO_17 (O_17,N_27317,N_28772);
and UO_18 (O_18,N_28131,N_27975);
nor UO_19 (O_19,N_28764,N_28181);
or UO_20 (O_20,N_29399,N_29417);
nand UO_21 (O_21,N_29316,N_27551);
xor UO_22 (O_22,N_28031,N_27639);
nand UO_23 (O_23,N_29476,N_29891);
and UO_24 (O_24,N_27914,N_28028);
or UO_25 (O_25,N_27658,N_27284);
or UO_26 (O_26,N_28263,N_28492);
or UO_27 (O_27,N_28761,N_28596);
or UO_28 (O_28,N_28939,N_28849);
or UO_29 (O_29,N_28269,N_28201);
xnor UO_30 (O_30,N_28896,N_28411);
nor UO_31 (O_31,N_29211,N_29470);
or UO_32 (O_32,N_29328,N_29058);
xor UO_33 (O_33,N_28553,N_29702);
nor UO_34 (O_34,N_28817,N_27348);
or UO_35 (O_35,N_27643,N_28262);
xor UO_36 (O_36,N_28264,N_29952);
xor UO_37 (O_37,N_29081,N_29449);
or UO_38 (O_38,N_27498,N_27752);
and UO_39 (O_39,N_28978,N_28888);
or UO_40 (O_40,N_27456,N_27180);
nor UO_41 (O_41,N_28558,N_29086);
or UO_42 (O_42,N_27473,N_28815);
and UO_43 (O_43,N_28357,N_29483);
and UO_44 (O_44,N_27329,N_28027);
nand UO_45 (O_45,N_28977,N_29382);
xor UO_46 (O_46,N_27065,N_27364);
xor UO_47 (O_47,N_27949,N_27145);
nor UO_48 (O_48,N_29471,N_29718);
or UO_49 (O_49,N_27548,N_28997);
and UO_50 (O_50,N_28628,N_29107);
and UO_51 (O_51,N_29951,N_27585);
or UO_52 (O_52,N_27462,N_27615);
and UO_53 (O_53,N_27124,N_27061);
or UO_54 (O_54,N_29593,N_29053);
nor UO_55 (O_55,N_29267,N_29216);
or UO_56 (O_56,N_29713,N_29361);
nand UO_57 (O_57,N_29428,N_29584);
or UO_58 (O_58,N_27851,N_27020);
xnor UO_59 (O_59,N_28491,N_29826);
and UO_60 (O_60,N_29598,N_29446);
or UO_61 (O_61,N_29240,N_27229);
nor UO_62 (O_62,N_28616,N_27074);
nor UO_63 (O_63,N_27453,N_29563);
xnor UO_64 (O_64,N_29078,N_27628);
nor UO_65 (O_65,N_29359,N_28069);
or UO_66 (O_66,N_28347,N_28349);
nor UO_67 (O_67,N_28305,N_27597);
nor UO_68 (O_68,N_29924,N_28052);
and UO_69 (O_69,N_28276,N_28319);
or UO_70 (O_70,N_28698,N_28531);
and UO_71 (O_71,N_29151,N_27645);
nor UO_72 (O_72,N_27552,N_28499);
nor UO_73 (O_73,N_27505,N_27897);
and UO_74 (O_74,N_28890,N_29903);
and UO_75 (O_75,N_28431,N_29221);
nand UO_76 (O_76,N_28162,N_27719);
nand UO_77 (O_77,N_29422,N_28718);
nand UO_78 (O_78,N_29234,N_27671);
nor UO_79 (O_79,N_29651,N_28451);
and UO_80 (O_80,N_28078,N_29653);
xnor UO_81 (O_81,N_28344,N_28641);
and UO_82 (O_82,N_29372,N_27500);
xnor UO_83 (O_83,N_27856,N_27848);
nand UO_84 (O_84,N_28476,N_29438);
nor UO_85 (O_85,N_28871,N_28992);
xnor UO_86 (O_86,N_27011,N_29126);
xnor UO_87 (O_87,N_28404,N_27748);
or UO_88 (O_88,N_29768,N_27063);
nor UO_89 (O_89,N_29735,N_27702);
xnor UO_90 (O_90,N_28296,N_29818);
nand UO_91 (O_91,N_28642,N_28017);
nand UO_92 (O_92,N_27472,N_29279);
xor UO_93 (O_93,N_28299,N_29925);
xor UO_94 (O_94,N_29520,N_28412);
or UO_95 (O_95,N_27427,N_28643);
or UO_96 (O_96,N_28086,N_27711);
nand UO_97 (O_97,N_29259,N_28521);
xnor UO_98 (O_98,N_27019,N_27474);
xnor UO_99 (O_99,N_28223,N_28571);
nor UO_100 (O_100,N_28824,N_27313);
nand UO_101 (O_101,N_27660,N_29159);
xnor UO_102 (O_102,N_29670,N_28705);
nor UO_103 (O_103,N_27194,N_29066);
and UO_104 (O_104,N_27789,N_29000);
and UO_105 (O_105,N_28000,N_28530);
and UO_106 (O_106,N_29332,N_28420);
nor UO_107 (O_107,N_29753,N_27423);
or UO_108 (O_108,N_29043,N_29353);
or UO_109 (O_109,N_29282,N_29723);
or UO_110 (O_110,N_28044,N_28875);
xor UO_111 (O_111,N_27139,N_27735);
xnor UO_112 (O_112,N_28753,N_27361);
nor UO_113 (O_113,N_27535,N_29919);
nor UO_114 (O_114,N_27439,N_29215);
nor UO_115 (O_115,N_28683,N_27657);
nand UO_116 (O_116,N_29338,N_29588);
nand UO_117 (O_117,N_29070,N_27118);
and UO_118 (O_118,N_27630,N_27683);
and UO_119 (O_119,N_29406,N_27314);
nand UO_120 (O_120,N_29906,N_27526);
xor UO_121 (O_121,N_28182,N_29764);
xnor UO_122 (O_122,N_28667,N_27146);
nand UO_123 (O_123,N_28238,N_29715);
nor UO_124 (O_124,N_29902,N_29934);
nand UO_125 (O_125,N_29423,N_28979);
xor UO_126 (O_126,N_27874,N_27753);
and UO_127 (O_127,N_28438,N_28147);
xnor UO_128 (O_128,N_27843,N_29778);
nand UO_129 (O_129,N_29163,N_29694);
nor UO_130 (O_130,N_28260,N_27808);
and UO_131 (O_131,N_29067,N_27008);
xor UO_132 (O_132,N_28533,N_27939);
or UO_133 (O_133,N_28676,N_27906);
and UO_134 (O_134,N_29590,N_27771);
nand UO_135 (O_135,N_28777,N_28161);
nor UO_136 (O_136,N_28934,N_29466);
xor UO_137 (O_137,N_29655,N_27050);
nor UO_138 (O_138,N_29810,N_28141);
nand UO_139 (O_139,N_29512,N_27680);
nand UO_140 (O_140,N_27149,N_27318);
or UO_141 (O_141,N_28774,N_29671);
nor UO_142 (O_142,N_28517,N_27129);
nor UO_143 (O_143,N_28072,N_27704);
or UO_144 (O_144,N_27530,N_27103);
or UO_145 (O_145,N_29122,N_28436);
nor UO_146 (O_146,N_27106,N_28919);
or UO_147 (O_147,N_29138,N_28423);
xor UO_148 (O_148,N_27446,N_27432);
xor UO_149 (O_149,N_27688,N_28732);
or UO_150 (O_150,N_27007,N_28703);
or UO_151 (O_151,N_29418,N_27824);
nor UO_152 (O_152,N_27220,N_29401);
and UO_153 (O_153,N_29500,N_27088);
nand UO_154 (O_154,N_28687,N_28883);
nand UO_155 (O_155,N_28605,N_29668);
nor UO_156 (O_156,N_27076,N_28457);
or UO_157 (O_157,N_27811,N_28821);
or UO_158 (O_158,N_27413,N_29909);
nor UO_159 (O_159,N_29928,N_29089);
nand UO_160 (O_160,N_28367,N_29275);
nand UO_161 (O_161,N_27160,N_29343);
nand UO_162 (O_162,N_28982,N_28425);
or UO_163 (O_163,N_27070,N_29614);
nor UO_164 (O_164,N_28623,N_29369);
xor UO_165 (O_165,N_29965,N_27945);
or UO_166 (O_166,N_28448,N_27754);
and UO_167 (O_167,N_29543,N_27434);
xor UO_168 (O_168,N_27039,N_29371);
nand UO_169 (O_169,N_28070,N_27232);
or UO_170 (O_170,N_29542,N_27218);
nor UO_171 (O_171,N_27522,N_28102);
or UO_172 (O_172,N_29530,N_28608);
nor UO_173 (O_173,N_28866,N_29348);
nand UO_174 (O_174,N_28833,N_28422);
nor UO_175 (O_175,N_28502,N_27721);
or UO_176 (O_176,N_29276,N_29324);
xor UO_177 (O_177,N_27210,N_28631);
and UO_178 (O_178,N_27828,N_29879);
or UO_179 (O_179,N_28011,N_27470);
xor UO_180 (O_180,N_29124,N_27844);
nor UO_181 (O_181,N_28130,N_28635);
nor UO_182 (O_182,N_27780,N_27835);
and UO_183 (O_183,N_29561,N_27234);
nor UO_184 (O_184,N_28666,N_29088);
nor UO_185 (O_185,N_28284,N_27100);
or UO_186 (O_186,N_27540,N_27875);
nor UO_187 (O_187,N_28439,N_29734);
nand UO_188 (O_188,N_27511,N_29189);
nor UO_189 (O_189,N_29101,N_27681);
xnor UO_190 (O_190,N_29959,N_28967);
or UO_191 (O_191,N_28770,N_29747);
or UO_192 (O_192,N_28787,N_29569);
or UO_193 (O_193,N_28337,N_27972);
nand UO_194 (O_194,N_28668,N_28306);
and UO_195 (O_195,N_28512,N_28094);
or UO_196 (O_196,N_28681,N_28803);
nand UO_197 (O_197,N_29468,N_27695);
nand UO_198 (O_198,N_29991,N_27991);
xnor UO_199 (O_199,N_29609,N_29686);
xor UO_200 (O_200,N_28286,N_28012);
xnor UO_201 (O_201,N_29586,N_28931);
or UO_202 (O_202,N_27770,N_28677);
or UO_203 (O_203,N_27443,N_28843);
or UO_204 (O_204,N_27974,N_29344);
nand UO_205 (O_205,N_29678,N_28617);
nand UO_206 (O_206,N_27521,N_28552);
and UO_207 (O_207,N_27254,N_29013);
nor UO_208 (O_208,N_29626,N_27613);
xnor UO_209 (O_209,N_29885,N_28200);
and UO_210 (O_210,N_27487,N_29935);
nand UO_211 (O_211,N_28889,N_28901);
nor UO_212 (O_212,N_28758,N_28719);
xnor UO_213 (O_213,N_27256,N_29631);
xor UO_214 (O_214,N_28509,N_28852);
nand UO_215 (O_215,N_29444,N_29581);
xnor UO_216 (O_216,N_28154,N_29001);
nor UO_217 (O_217,N_28085,N_29378);
nor UO_218 (O_218,N_27805,N_27121);
nor UO_219 (O_219,N_27560,N_29862);
and UO_220 (O_220,N_28893,N_29624);
or UO_221 (O_221,N_27831,N_28316);
or UO_222 (O_222,N_27214,N_28092);
or UO_223 (O_223,N_28213,N_28107);
nand UO_224 (O_224,N_28996,N_28932);
or UO_225 (O_225,N_29289,N_28272);
nand UO_226 (O_226,N_28462,N_29535);
nor UO_227 (O_227,N_28725,N_27280);
xor UO_228 (O_228,N_27801,N_29900);
nor UO_229 (O_229,N_29308,N_27827);
or UO_230 (O_230,N_27839,N_27921);
or UO_231 (O_231,N_27116,N_28727);
nand UO_232 (O_232,N_29238,N_28449);
or UO_233 (O_233,N_27374,N_28661);
xor UO_234 (O_234,N_27449,N_27266);
nor UO_235 (O_235,N_27901,N_27541);
nand UO_236 (O_236,N_27454,N_29710);
or UO_237 (O_237,N_29085,N_27415);
xor UO_238 (O_238,N_28482,N_29123);
and UO_239 (O_239,N_28734,N_27113);
and UO_240 (O_240,N_29523,N_27764);
nand UO_241 (O_241,N_29179,N_29011);
xor UO_242 (O_242,N_29209,N_28744);
nand UO_243 (O_243,N_28249,N_27114);
and UO_244 (O_244,N_29983,N_27502);
nor UO_245 (O_245,N_27442,N_28183);
nor UO_246 (O_246,N_29203,N_29776);
nand UO_247 (O_247,N_28090,N_28595);
xnor UO_248 (O_248,N_29673,N_29491);
nand UO_249 (O_249,N_28779,N_28087);
xnor UO_250 (O_250,N_29800,N_28970);
or UO_251 (O_251,N_29068,N_27590);
and UO_252 (O_252,N_29882,N_28909);
and UO_253 (O_253,N_27016,N_27594);
xor UO_254 (O_254,N_27954,N_28535);
or UO_255 (O_255,N_28168,N_28322);
xnor UO_256 (O_256,N_28990,N_29821);
nand UO_257 (O_257,N_29941,N_28298);
xnor UO_258 (O_258,N_27757,N_29802);
nor UO_259 (O_259,N_29017,N_27325);
xnor UO_260 (O_260,N_29766,N_28902);
and UO_261 (O_261,N_27793,N_28807);
and UO_262 (O_262,N_29813,N_29060);
nor UO_263 (O_263,N_27004,N_27304);
or UO_264 (O_264,N_28569,N_28184);
nand UO_265 (O_265,N_27923,N_29849);
nor UO_266 (O_266,N_27352,N_29222);
xnor UO_267 (O_267,N_28164,N_27638);
xnor UO_268 (O_268,N_28678,N_29330);
and UO_269 (O_269,N_27572,N_27048);
or UO_270 (O_270,N_29415,N_28211);
xor UO_271 (O_271,N_27565,N_29097);
or UO_272 (O_272,N_28981,N_28537);
nor UO_273 (O_273,N_29135,N_28860);
and UO_274 (O_274,N_28606,N_29443);
or UO_275 (O_275,N_27403,N_29726);
or UO_276 (O_276,N_27850,N_28124);
xnor UO_277 (O_277,N_28007,N_27075);
nand UO_278 (O_278,N_29914,N_28494);
and UO_279 (O_279,N_29229,N_29398);
and UO_280 (O_280,N_29908,N_28785);
nor UO_281 (O_281,N_27444,N_29567);
nand UO_282 (O_282,N_29918,N_28508);
and UO_283 (O_283,N_27097,N_28040);
and UO_284 (O_284,N_28755,N_27216);
and UO_285 (O_285,N_27316,N_29811);
nor UO_286 (O_286,N_27903,N_29219);
or UO_287 (O_287,N_28385,N_29019);
nor UO_288 (O_288,N_27323,N_27494);
and UO_289 (O_289,N_27815,N_28143);
or UO_290 (O_290,N_27133,N_28954);
xor UO_291 (O_291,N_28861,N_29806);
nand UO_292 (O_292,N_28020,N_28892);
nor UO_293 (O_293,N_27108,N_27606);
xor UO_294 (O_294,N_27913,N_27938);
xor UO_295 (O_295,N_29386,N_27199);
and UO_296 (O_296,N_29357,N_28520);
xnor UO_297 (O_297,N_29319,N_29358);
or UO_298 (O_298,N_29707,N_27136);
xor UO_299 (O_299,N_28484,N_29192);
nor UO_300 (O_300,N_29178,N_27942);
nand UO_301 (O_301,N_27246,N_27722);
and UO_302 (O_302,N_27476,N_27288);
nor UO_303 (O_303,N_29208,N_29575);
xnor UO_304 (O_304,N_28874,N_27320);
and UO_305 (O_305,N_29193,N_28334);
nor UO_306 (O_306,N_28534,N_29455);
and UO_307 (O_307,N_29474,N_27337);
and UO_308 (O_308,N_28644,N_28601);
nand UO_309 (O_309,N_28196,N_27094);
nor UO_310 (O_310,N_28818,N_28749);
nand UO_311 (O_311,N_28704,N_27896);
nand UO_312 (O_312,N_28016,N_29478);
nor UO_313 (O_313,N_28064,N_29910);
nor UO_314 (O_314,N_27948,N_28663);
and UO_315 (O_315,N_29880,N_28947);
nor UO_316 (O_316,N_27983,N_27508);
xnor UO_317 (O_317,N_27576,N_29341);
and UO_318 (O_318,N_27148,N_28495);
nand UO_319 (O_319,N_29460,N_28490);
or UO_320 (O_320,N_27743,N_29197);
and UO_321 (O_321,N_27188,N_27900);
or UO_322 (O_322,N_29082,N_27177);
and UO_323 (O_323,N_28878,N_29247);
nand UO_324 (O_324,N_28971,N_27137);
xor UO_325 (O_325,N_28307,N_28540);
nor UO_326 (O_326,N_28999,N_27099);
and UO_327 (O_327,N_27045,N_28415);
or UO_328 (O_328,N_29286,N_29489);
xnor UO_329 (O_329,N_29205,N_29505);
xor UO_330 (O_330,N_28426,N_28342);
or UO_331 (O_331,N_27790,N_29224);
xnor UO_332 (O_332,N_27049,N_27359);
and UO_333 (O_333,N_29785,N_27968);
and UO_334 (O_334,N_28034,N_29127);
nand UO_335 (O_335,N_29187,N_28479);
and UO_336 (O_336,N_29027,N_28315);
or UO_337 (O_337,N_29878,N_28578);
xnor UO_338 (O_338,N_29704,N_27212);
nand UO_339 (O_339,N_27278,N_27525);
nand UO_340 (O_340,N_28116,N_27608);
xnor UO_341 (O_341,N_28962,N_29913);
and UO_342 (O_342,N_27916,N_28811);
nand UO_343 (O_343,N_28022,N_27534);
xor UO_344 (O_344,N_28897,N_28268);
nand UO_345 (O_345,N_29158,N_27703);
and UO_346 (O_346,N_28099,N_28145);
or UO_347 (O_347,N_29022,N_28049);
nor UO_348 (O_348,N_29967,N_27055);
nor UO_349 (O_349,N_28949,N_28194);
xor UO_350 (O_350,N_27464,N_27621);
xor UO_351 (O_351,N_27080,N_28039);
or UO_352 (O_352,N_29527,N_27271);
nand UO_353 (O_353,N_27819,N_28593);
nor UO_354 (O_354,N_29699,N_27886);
xnor UO_355 (O_355,N_28801,N_28882);
nor UO_356 (O_356,N_29160,N_27959);
nand UO_357 (O_357,N_29741,N_28619);
or UO_358 (O_358,N_29585,N_27539);
nor UO_359 (O_359,N_27377,N_29038);
or UO_360 (O_360,N_27184,N_27395);
nand UO_361 (O_361,N_29258,N_29789);
or UO_362 (O_362,N_28081,N_29596);
and UO_363 (O_363,N_27512,N_28345);
xor UO_364 (O_364,N_27169,N_29389);
and UO_365 (O_365,N_29248,N_28056);
nand UO_366 (O_366,N_28246,N_27718);
xnor UO_367 (O_367,N_27797,N_27773);
or UO_368 (O_368,N_28670,N_28244);
and UO_369 (O_369,N_27884,N_28432);
or UO_370 (O_370,N_28325,N_27396);
nand UO_371 (O_371,N_29946,N_27410);
and UO_372 (O_372,N_28318,N_29080);
nand UO_373 (O_373,N_29533,N_29749);
nand UO_374 (O_374,N_28477,N_29287);
or UO_375 (O_375,N_28273,N_29521);
xnor UO_376 (O_376,N_27190,N_27341);
and UO_377 (O_377,N_27119,N_27784);
nor UO_378 (O_378,N_27109,N_29613);
nand UO_379 (O_379,N_28123,N_28946);
xnor UO_380 (O_380,N_27372,N_29497);
and UO_381 (O_381,N_29758,N_27622);
or UO_382 (O_382,N_29752,N_29524);
nand UO_383 (O_383,N_29300,N_29808);
xnor UO_384 (O_384,N_27458,N_28691);
xor UO_385 (O_385,N_29181,N_27386);
and UO_386 (O_386,N_27385,N_29182);
nor UO_387 (O_387,N_28500,N_27072);
or UO_388 (O_388,N_28831,N_27079);
or UO_389 (O_389,N_27600,N_29379);
nor UO_390 (O_390,N_27544,N_27774);
nand UO_391 (O_391,N_28115,N_29577);
or UO_392 (O_392,N_28783,N_27290);
xnor UO_393 (O_393,N_27746,N_29150);
nor UO_394 (O_394,N_28146,N_28454);
xnor UO_395 (O_395,N_27616,N_28441);
xor UO_396 (O_396,N_29206,N_28215);
nor UO_397 (O_397,N_29393,N_27005);
xor UO_398 (O_398,N_27733,N_28752);
nand UO_399 (O_399,N_29922,N_29616);
nor UO_400 (O_400,N_27175,N_27173);
or UO_401 (O_401,N_29644,N_29939);
nand UO_402 (O_402,N_27854,N_28062);
xor UO_403 (O_403,N_28865,N_29729);
nor UO_404 (O_404,N_27816,N_29095);
and UO_405 (O_405,N_28096,N_27475);
nor UO_406 (O_406,N_28554,N_28247);
xnor UO_407 (O_407,N_29973,N_29213);
or UO_408 (O_408,N_29562,N_27849);
xnor UO_409 (O_409,N_28583,N_29439);
xor UO_410 (O_410,N_27373,N_28279);
xor UO_411 (O_411,N_27969,N_27391);
nand UO_412 (O_412,N_27744,N_27101);
or UO_413 (O_413,N_28030,N_28125);
nand UO_414 (O_414,N_29069,N_28132);
or UO_415 (O_415,N_28084,N_28708);
or UO_416 (O_416,N_27489,N_27224);
nand UO_417 (O_417,N_28149,N_27672);
nor UO_418 (O_418,N_27618,N_28602);
and UO_419 (O_419,N_28859,N_28455);
xnor UO_420 (O_420,N_28952,N_29604);
or UO_421 (O_421,N_28624,N_28195);
nand UO_422 (O_422,N_28235,N_29075);
and UO_423 (O_423,N_27687,N_28109);
or UO_424 (O_424,N_29177,N_28739);
nor UO_425 (O_425,N_27370,N_28814);
nor UO_426 (O_426,N_28187,N_27052);
nor UO_427 (O_427,N_29241,N_28074);
nor UO_428 (O_428,N_29893,N_27082);
xnor UO_429 (O_429,N_29787,N_29312);
nand UO_430 (O_430,N_29829,N_27251);
xnor UO_431 (O_431,N_29133,N_27971);
nor UO_432 (O_432,N_27918,N_27637);
nor UO_433 (O_433,N_29815,N_28290);
nand UO_434 (O_434,N_28684,N_27492);
and UO_435 (O_435,N_29031,N_28392);
or UO_436 (O_436,N_28937,N_28217);
or UO_437 (O_437,N_27296,N_27555);
or UO_438 (O_438,N_27862,N_29669);
and UO_439 (O_439,N_28098,N_27632);
xor UO_440 (O_440,N_29271,N_29071);
nor UO_441 (O_441,N_28768,N_29599);
and UO_442 (O_442,N_27509,N_28710);
xor UO_443 (O_443,N_28802,N_28516);
nor UO_444 (O_444,N_28459,N_28353);
xnor UO_445 (O_445,N_28538,N_29858);
or UO_446 (O_446,N_27159,N_29290);
nor UO_447 (O_447,N_27932,N_28277);
or UO_448 (O_448,N_29976,N_28498);
and UO_449 (O_449,N_28969,N_28778);
and UO_450 (O_450,N_28383,N_27795);
nand UO_451 (O_451,N_27040,N_27347);
nor UO_452 (O_452,N_27664,N_29730);
and UO_453 (O_453,N_29564,N_27245);
xor UO_454 (O_454,N_28864,N_28075);
or UO_455 (O_455,N_28523,N_29283);
nor UO_456 (O_456,N_29998,N_27355);
xor UO_457 (O_457,N_29465,N_29658);
or UO_458 (O_458,N_29457,N_29050);
xnor UO_459 (O_459,N_29875,N_28461);
and UO_460 (O_460,N_29549,N_27567);
or UO_461 (O_461,N_28626,N_28697);
nor UO_462 (O_462,N_29469,N_28837);
and UO_463 (O_463,N_28372,N_28178);
nor UO_464 (O_464,N_27559,N_28757);
or UO_465 (O_465,N_27178,N_29846);
and UO_466 (O_466,N_29106,N_29498);
nand UO_467 (O_467,N_27532,N_27400);
and UO_468 (O_468,N_27984,N_29881);
and UO_469 (O_469,N_28408,N_28799);
nand UO_470 (O_470,N_28812,N_29518);
xnor UO_471 (O_471,N_29534,N_27707);
xor UO_472 (O_472,N_28063,N_27527);
and UO_473 (O_473,N_29641,N_28715);
nor UO_474 (O_474,N_27388,N_27956);
and UO_475 (O_475,N_27605,N_29266);
xor UO_476 (O_476,N_29748,N_27580);
and UO_477 (O_477,N_29394,N_29169);
or UO_478 (O_478,N_29664,N_27406);
nor UO_479 (O_479,N_29061,N_28776);
or UO_480 (O_480,N_27322,N_28250);
or UO_481 (O_481,N_29696,N_28735);
or UO_482 (O_482,N_28169,N_27228);
and UO_483 (O_483,N_28113,N_28014);
xor UO_484 (O_484,N_28060,N_28114);
nor UO_485 (O_485,N_27556,N_28689);
and UO_486 (O_486,N_29963,N_29514);
nor UO_487 (O_487,N_28489,N_29490);
xnor UO_488 (O_488,N_27717,N_28980);
nor UO_489 (O_489,N_29850,N_27581);
nor UO_490 (O_490,N_27759,N_29350);
xnor UO_491 (O_491,N_28907,N_29176);
nor UO_492 (O_492,N_28542,N_27147);
xor UO_493 (O_493,N_28924,N_29486);
and UO_494 (O_494,N_28227,N_28790);
or UO_495 (O_495,N_28314,N_28001);
xor UO_496 (O_496,N_28471,N_29077);
nor UO_497 (O_497,N_28252,N_29780);
xnor UO_498 (O_498,N_29601,N_27157);
or UO_499 (O_499,N_29953,N_29296);
nand UO_500 (O_500,N_28926,N_28948);
nor UO_501 (O_501,N_28816,N_29949);
nand UO_502 (O_502,N_28651,N_29617);
nand UO_503 (O_503,N_27634,N_29366);
nor UO_504 (O_504,N_29650,N_28368);
and UO_505 (O_505,N_29062,N_28118);
and UO_506 (O_506,N_28150,N_28629);
nand UO_507 (O_507,N_29175,N_27593);
and UO_508 (O_508,N_27652,N_29397);
and UO_509 (O_509,N_28045,N_28328);
or UO_510 (O_510,N_27673,N_29014);
nand UO_511 (O_511,N_27006,N_29636);
nor UO_512 (O_512,N_27046,N_27531);
nor UO_513 (O_513,N_29602,N_28203);
nand UO_514 (O_514,N_27908,N_27761);
nand UO_515 (O_515,N_27000,N_29989);
or UO_516 (O_516,N_28138,N_29996);
and UO_517 (O_517,N_29975,N_28912);
and UO_518 (O_518,N_27223,N_27987);
nor UO_519 (O_519,N_28632,N_27818);
or UO_520 (O_520,N_28577,N_29659);
nand UO_521 (O_521,N_29844,N_29746);
nor UO_522 (O_522,N_29083,N_28589);
nand UO_523 (O_523,N_28618,N_29728);
nand UO_524 (O_524,N_28539,N_27293);
xnor UO_525 (O_525,N_27941,N_27203);
and UO_526 (O_526,N_28329,N_29691);
nand UO_527 (O_527,N_28288,N_29084);
or UO_528 (O_528,N_29024,N_27692);
and UO_529 (O_529,N_27015,N_29732);
or UO_530 (O_530,N_28615,N_29035);
nor UO_531 (O_531,N_29755,N_29923);
and UO_532 (O_532,N_27303,N_27781);
and UO_533 (O_533,N_28650,N_29560);
and UO_534 (O_534,N_27741,N_29452);
and UO_535 (O_535,N_29190,N_28604);
nand UO_536 (O_536,N_29522,N_28857);
and UO_537 (O_537,N_28702,N_29873);
xor UO_538 (O_538,N_27233,N_28613);
and UO_539 (O_539,N_28136,N_27724);
nand UO_540 (O_540,N_29110,N_27356);
nor UO_541 (O_541,N_29199,N_29637);
or UO_542 (O_542,N_28822,N_28460);
nand UO_543 (O_543,N_28076,N_29684);
nand UO_544 (O_544,N_28467,N_28762);
nand UO_545 (O_545,N_29409,N_27257);
nand UO_546 (O_546,N_29304,N_28566);
nor UO_547 (O_547,N_27678,N_29784);
or UO_548 (O_548,N_28366,N_27200);
xor UO_549 (O_549,N_27846,N_28963);
or UO_550 (O_550,N_29305,N_27219);
and UO_551 (O_551,N_28218,N_27128);
nand UO_552 (O_552,N_28877,N_27351);
xor UO_553 (O_553,N_28041,N_28111);
and UO_554 (O_554,N_29194,N_29306);
xnor UO_555 (O_555,N_29867,N_27550);
nand UO_556 (O_556,N_29459,N_27301);
or UO_557 (O_557,N_27591,N_28033);
xor UO_558 (O_558,N_27419,N_28407);
and UO_559 (O_559,N_27662,N_27098);
nand UO_560 (O_560,N_29587,N_29508);
or UO_561 (O_561,N_27888,N_28598);
nor UO_562 (O_562,N_27191,N_29757);
or UO_563 (O_563,N_28664,N_28134);
nand UO_564 (O_564,N_27768,N_29712);
nor UO_565 (O_565,N_29252,N_28271);
and UO_566 (O_566,N_27078,N_27420);
xnor UO_567 (O_567,N_27155,N_27588);
or UO_568 (O_568,N_27363,N_27587);
nor UO_569 (O_569,N_28863,N_27737);
xor UO_570 (O_570,N_28782,N_29733);
nor UO_571 (O_571,N_28518,N_27650);
xnor UO_572 (O_572,N_27732,N_29098);
xor UO_573 (O_573,N_28544,N_29597);
nand UO_574 (O_574,N_28133,N_28358);
xnor UO_575 (O_575,N_28835,N_28853);
xor UO_576 (O_576,N_27873,N_27796);
xor UO_577 (O_577,N_27275,N_28160);
or UO_578 (O_578,N_29244,N_27999);
and UO_579 (O_579,N_28015,N_29643);
nor UO_580 (O_580,N_28192,N_27091);
and UO_581 (O_581,N_27710,N_27877);
nor UO_582 (O_582,N_28071,N_27852);
or UO_583 (O_583,N_29705,N_28302);
nand UO_584 (O_584,N_27243,N_28151);
and UO_585 (O_585,N_28998,N_29503);
and UO_586 (O_586,N_28265,N_27171);
and UO_587 (O_587,N_28582,N_29700);
nand UO_588 (O_588,N_27651,N_28019);
or UO_589 (O_589,N_28452,N_27927);
nand UO_590 (O_590,N_28335,N_27669);
or UO_591 (O_591,N_29072,N_27362);
and UO_592 (O_592,N_29679,N_29168);
nor UO_593 (O_593,N_29482,N_28795);
and UO_594 (O_594,N_27132,N_27350);
and UO_595 (O_595,N_29843,N_28410);
xnor UO_596 (O_596,N_27714,N_27261);
nor UO_597 (O_597,N_28117,N_27021);
or UO_598 (O_598,N_27196,N_28694);
nand UO_599 (O_599,N_29087,N_27817);
and UO_600 (O_600,N_27111,N_27421);
or UO_601 (O_601,N_29281,N_28198);
xnor UO_602 (O_602,N_28464,N_27653);
nor UO_603 (O_603,N_28522,N_27336);
nand UO_604 (O_604,N_27766,N_29656);
and UO_605 (O_605,N_28830,N_27785);
nand UO_606 (O_606,N_28916,N_27343);
and UO_607 (O_607,N_27095,N_28396);
and UO_608 (O_608,N_28724,N_28445);
nand UO_609 (O_609,N_29385,N_29703);
nand UO_610 (O_610,N_27239,N_29759);
and UO_611 (O_611,N_27952,N_29847);
or UO_612 (O_612,N_29396,N_28560);
nand UO_613 (O_613,N_29529,N_29739);
xnor UO_614 (O_614,N_28486,N_29988);
nand UO_615 (O_615,N_29129,N_28258);
or UO_616 (O_616,N_29956,N_28148);
or UO_617 (O_617,N_28382,N_28079);
and UO_618 (O_618,N_28870,N_27425);
or UO_619 (O_619,N_29680,N_27910);
xnor UO_620 (O_620,N_29904,N_29582);
xnor UO_621 (O_621,N_28189,N_29837);
xnor UO_622 (O_622,N_27977,N_29570);
nand UO_623 (O_623,N_27206,N_27919);
nand UO_624 (O_624,N_28005,N_28326);
nor UO_625 (O_625,N_29580,N_29539);
nand UO_626 (O_626,N_27131,N_29819);
nand UO_627 (O_627,N_27167,N_28819);
xnor UO_628 (O_628,N_27950,N_29121);
xnor UO_629 (O_629,N_29118,N_27066);
and UO_630 (O_630,N_27647,N_28805);
and UO_631 (O_631,N_29367,N_29868);
nand UO_632 (O_632,N_28023,N_29744);
nor UO_633 (O_633,N_27170,N_27151);
or UO_634 (O_634,N_29364,N_28640);
and UO_635 (O_635,N_27665,N_29246);
xor UO_636 (O_636,N_29188,N_28929);
nor UO_637 (O_637,N_28966,N_29492);
and UO_638 (O_638,N_27235,N_28157);
or UO_639 (O_639,N_29105,N_27772);
nand UO_640 (O_640,N_28573,N_29303);
and UO_641 (O_641,N_28846,N_28941);
nand UO_642 (O_642,N_27092,N_29481);
nand UO_643 (O_643,N_28446,N_27682);
nand UO_644 (O_644,N_29464,N_27944);
nor UO_645 (O_645,N_29310,N_28394);
and UO_646 (O_646,N_29861,N_27127);
or UO_647 (O_647,N_29472,N_28741);
or UO_648 (O_648,N_28548,N_28536);
and UO_649 (O_649,N_29288,N_27625);
and UO_650 (O_650,N_28140,N_27705);
nand UO_651 (O_651,N_28568,N_28733);
nand UO_652 (O_652,N_27144,N_27996);
and UO_653 (O_653,N_27340,N_29487);
or UO_654 (O_654,N_28301,N_27001);
nor UO_655 (O_655,N_29897,N_28010);
and UO_656 (O_656,N_27272,N_27936);
xnor UO_657 (O_657,N_29100,N_29547);
and UO_658 (O_658,N_27310,N_28289);
xnor UO_659 (O_659,N_29932,N_28750);
or UO_660 (O_660,N_28903,N_29864);
nand UO_661 (O_661,N_29770,N_29342);
and UO_662 (O_662,N_27607,N_27750);
nand UO_663 (O_663,N_27154,N_29742);
or UO_664 (O_664,N_27448,N_27547);
nor UO_665 (O_665,N_28885,N_28003);
nor UO_666 (O_666,N_27459,N_29727);
and UO_667 (O_667,N_28620,N_28364);
nand UO_668 (O_668,N_28630,N_29509);
xnor UO_669 (O_669,N_29384,N_29957);
xor UO_670 (O_670,N_27107,N_27038);
xor UO_671 (O_671,N_29041,N_28820);
and UO_672 (O_672,N_27249,N_27438);
or UO_673 (O_673,N_29437,N_27577);
nand UO_674 (O_674,N_29894,N_27349);
xor UO_675 (O_675,N_27656,N_29920);
or UO_676 (O_676,N_28391,N_29981);
nand UO_677 (O_677,N_27876,N_28323);
nor UO_678 (O_678,N_27463,N_29915);
or UO_679 (O_679,N_29475,N_29851);
nor UO_680 (O_680,N_28574,N_28343);
nand UO_681 (O_681,N_27696,N_27562);
nand UO_682 (O_682,N_28444,N_27998);
or UO_683 (O_683,N_28059,N_29901);
nor UO_684 (O_684,N_29052,N_27533);
or UO_685 (O_685,N_29298,N_28868);
and UO_686 (O_686,N_28406,N_27367);
nand UO_687 (O_687,N_28514,N_27241);
nand UO_688 (O_688,N_27633,N_29557);
xor UO_689 (O_689,N_29830,N_29532);
nor UO_690 (O_690,N_27982,N_27418);
xor UO_691 (O_691,N_29134,N_27461);
nor UO_692 (O_692,N_29235,N_29883);
nand UO_693 (O_693,N_29839,N_27958);
nand UO_694 (O_694,N_28515,N_29646);
nand UO_695 (O_695,N_27466,N_29318);
xor UO_696 (O_696,N_27417,N_28951);
nand UO_697 (O_697,N_27514,N_29986);
nand UO_698 (O_698,N_28155,N_28210);
nand UO_699 (O_699,N_29931,N_27315);
xnor UO_700 (O_700,N_29972,N_27031);
and UO_701 (O_701,N_28592,N_27592);
and UO_702 (O_702,N_28035,N_28266);
nand UO_703 (O_703,N_29842,N_29420);
and UO_704 (O_704,N_28957,N_27501);
and UO_705 (O_705,N_27837,N_27546);
or UO_706 (O_706,N_28827,N_28809);
nor UO_707 (O_707,N_28443,N_29494);
xnor UO_708 (O_708,N_29430,N_28336);
nor UO_709 (O_709,N_29511,N_29039);
nor UO_710 (O_710,N_28371,N_28647);
nand UO_711 (O_711,N_27207,N_27558);
and UO_712 (O_712,N_28622,N_28170);
or UO_713 (O_713,N_27933,N_27483);
nand UO_714 (O_714,N_28915,N_29250);
xnor UO_715 (O_715,N_29132,N_27433);
nand UO_716 (O_716,N_27644,N_29109);
nand UO_717 (O_717,N_27519,N_27611);
nor UO_718 (O_718,N_29899,N_27345);
nand UO_719 (O_719,N_29202,N_27965);
and UO_720 (O_720,N_28173,N_27429);
nand UO_721 (O_721,N_29317,N_28904);
nor UO_722 (O_722,N_27891,N_27493);
or UO_723 (O_723,N_28736,N_28165);
or UO_724 (O_724,N_28197,N_28714);
nor UO_725 (O_725,N_29788,N_27339);
nor UO_726 (O_726,N_27868,N_29756);
nand UO_727 (O_727,N_28363,N_29933);
and UO_728 (O_728,N_28379,N_29950);
and UO_729 (O_729,N_29840,N_27230);
and UO_730 (O_730,N_29392,N_28053);
xor UO_731 (O_731,N_28740,N_28458);
nor UO_732 (O_732,N_27782,N_27185);
and UO_733 (O_733,N_27518,N_28338);
and UO_734 (O_734,N_28834,N_28693);
nor UO_735 (O_735,N_28401,N_29997);
or UO_736 (O_736,N_28480,N_28378);
xor UO_737 (O_737,N_27564,N_27163);
nor UO_738 (O_738,N_29823,N_29092);
and UO_739 (O_739,N_27027,N_29419);
nor UO_740 (O_740,N_29608,N_27504);
xor UO_741 (O_741,N_27834,N_29223);
xor UO_742 (O_742,N_27858,N_27569);
or UO_743 (O_743,N_28695,N_27777);
nand UO_744 (O_744,N_28549,N_28242);
or UO_745 (O_745,N_29773,N_27698);
nor UO_746 (O_746,N_29424,N_29360);
xor UO_747 (O_747,N_27543,N_28983);
or UO_748 (O_748,N_29365,N_29458);
or UO_749 (O_749,N_28100,N_29531);
and UO_750 (O_750,N_29023,N_29334);
xor UO_751 (O_751,N_28842,N_29036);
and UO_752 (O_752,N_27515,N_29201);
nor UO_753 (O_753,N_27820,N_29642);
xnor UO_754 (O_754,N_29725,N_28960);
and UO_755 (O_755,N_28106,N_28965);
nand UO_756 (O_756,N_27060,N_27117);
xor UO_757 (O_757,N_28191,N_29033);
nor UO_758 (O_758,N_28886,N_29681);
nor UO_759 (O_759,N_28281,N_27596);
or UO_760 (O_760,N_28856,N_29940);
and UO_761 (O_761,N_28519,N_28222);
nand UO_762 (O_762,N_29499,N_29161);
or UO_763 (O_763,N_27328,N_28586);
nor UO_764 (O_764,N_27745,N_29363);
nor UO_765 (O_765,N_28791,N_28918);
nand UO_766 (O_766,N_27684,N_28850);
xor UO_767 (O_767,N_29877,N_27990);
and UO_768 (O_768,N_28280,N_27378);
and UO_769 (O_769,N_27299,N_29907);
nor UO_770 (O_770,N_29099,N_29771);
and UO_771 (O_771,N_28585,N_29128);
nor UO_772 (O_772,N_28310,N_28935);
nor UO_773 (O_773,N_28638,N_27507);
and UO_774 (O_774,N_28662,N_27394);
or UO_775 (O_775,N_29473,N_27110);
xnor UO_776 (O_776,N_27264,N_28362);
nor UO_777 (O_777,N_29196,N_29898);
or UO_778 (O_778,N_28751,N_27619);
or UO_779 (O_779,N_28097,N_27701);
nand UO_780 (O_780,N_28780,N_27730);
xor UO_781 (O_781,N_27387,N_29634);
xnor UO_782 (O_782,N_29111,N_27477);
xnor UO_783 (O_783,N_27156,N_28135);
nand UO_784 (O_784,N_29352,N_28876);
xor UO_785 (O_785,N_29104,N_27994);
nand UO_786 (O_786,N_27383,N_28251);
or UO_787 (O_787,N_29857,N_28665);
or UO_788 (O_788,N_29325,N_29125);
or UO_789 (O_789,N_27751,N_29751);
or UO_790 (O_790,N_29738,N_27822);
xnor UO_791 (O_791,N_29926,N_29006);
nand UO_792 (O_792,N_29803,N_29184);
or UO_793 (O_793,N_29346,N_29217);
nor UO_794 (O_794,N_28088,N_29693);
or UO_795 (O_795,N_29754,N_28950);
xor UO_796 (O_796,N_27047,N_28065);
and UO_797 (O_797,N_29251,N_29141);
nand UO_798 (O_798,N_28331,N_29044);
or UO_799 (O_799,N_27740,N_28254);
and UO_800 (O_800,N_28938,N_29630);
nor UO_801 (O_801,N_27749,N_28082);
and UO_802 (O_802,N_28359,N_27953);
or UO_803 (O_803,N_27833,N_28895);
nor UO_804 (O_804,N_29146,N_27488);
and UO_805 (O_805,N_29007,N_28769);
xnor UO_806 (O_806,N_28255,N_27291);
and UO_807 (O_807,N_27804,N_28648);
and UO_808 (O_808,N_27469,N_27840);
and UO_809 (O_809,N_28711,N_29794);
nor UO_810 (O_810,N_28324,N_28418);
nand UO_811 (O_811,N_29695,N_27617);
nand UO_812 (O_812,N_29320,N_27176);
nand UO_813 (O_813,N_27864,N_28267);
and UO_814 (O_814,N_29954,N_27321);
or UO_815 (O_815,N_27691,N_29657);
and UO_816 (O_816,N_29115,N_27017);
nand UO_817 (O_817,N_28933,N_28395);
and UO_818 (O_818,N_27338,N_29971);
and UO_819 (O_819,N_29760,N_28179);
nor UO_820 (O_820,N_27416,N_28346);
nor UO_821 (O_821,N_28731,N_28881);
or UO_822 (O_822,N_27723,N_28506);
and UO_823 (O_823,N_27503,N_29307);
nand UO_824 (O_824,N_27013,N_27058);
or UO_825 (O_825,N_29938,N_27287);
xor UO_826 (O_826,N_27179,N_28465);
nand UO_827 (O_827,N_28101,N_28636);
xnor UO_828 (O_828,N_27282,N_27880);
nand UO_829 (O_829,N_28543,N_29165);
nor UO_830 (O_830,N_27215,N_27360);
nand UO_831 (O_831,N_28825,N_29838);
and UO_832 (O_832,N_29480,N_28057);
or UO_833 (O_833,N_29554,N_28729);
xnor UO_834 (O_834,N_28229,N_27760);
nand UO_835 (O_835,N_29467,N_27032);
or UO_836 (O_836,N_28706,N_28887);
xor UO_837 (O_837,N_29195,N_28994);
nor UO_838 (O_838,N_29889,N_27878);
or UO_839 (O_839,N_28447,N_29555);
or UO_840 (O_840,N_28584,N_29425);
xnor UO_841 (O_841,N_28555,N_27115);
nand UO_842 (O_842,N_29390,N_28456);
or UO_843 (O_843,N_29147,N_28657);
or UO_844 (O_844,N_29736,N_28914);
xnor UO_845 (O_845,N_29102,N_27857);
or UO_846 (O_846,N_28297,N_29717);
nand UO_847 (O_847,N_28321,N_28652);
xnor UO_848 (O_848,N_29860,N_29375);
or UO_849 (O_849,N_27152,N_29204);
or UO_850 (O_850,N_27431,N_29854);
nor UO_851 (O_851,N_27197,N_27408);
or UO_852 (O_852,N_28158,N_27465);
and UO_853 (O_853,N_28955,N_28541);
nand UO_854 (O_854,N_27887,N_29144);
or UO_855 (O_855,N_27250,N_29351);
or UO_856 (O_856,N_27479,N_29559);
nor UO_857 (O_857,N_28806,N_27836);
nand UO_858 (O_858,N_28701,N_28221);
and UO_859 (O_859,N_29783,N_28611);
or UO_860 (O_860,N_28174,N_27940);
and UO_861 (O_861,N_28561,N_27237);
and UO_862 (O_862,N_29945,N_28745);
nor UO_863 (O_863,N_27667,N_28973);
and UO_864 (O_864,N_28872,N_29937);
xnor UO_865 (O_865,N_29049,N_29982);
and UO_866 (O_866,N_27211,N_27165);
nor UO_867 (O_867,N_27973,N_29541);
nand UO_868 (O_868,N_29987,N_27389);
and UO_869 (O_869,N_27285,N_29403);
or UO_870 (O_870,N_28559,N_27093);
nor UO_871 (O_871,N_29853,N_27979);
xor UO_872 (O_872,N_28655,N_27455);
xnor UO_873 (O_873,N_28171,N_29721);
nand UO_874 (O_874,N_29395,N_28156);
nand UO_875 (O_875,N_28575,N_28348);
and UO_876 (O_876,N_29647,N_28603);
nand UO_877 (O_877,N_29822,N_28417);
nand UO_878 (O_878,N_28985,N_29504);
and UO_879 (O_879,N_27480,N_27451);
xor UO_880 (O_880,N_27073,N_29615);
nand UO_881 (O_881,N_27033,N_29091);
or UO_882 (O_882,N_29545,N_27468);
or UO_883 (O_883,N_29362,N_28804);
and UO_884 (O_884,N_29373,N_28524);
nand UO_885 (O_885,N_27297,N_27126);
nand UO_886 (O_886,N_29230,N_27084);
nand UO_887 (O_887,N_27392,N_29170);
nor UO_888 (O_888,N_27578,N_29576);
and UO_889 (O_889,N_27368,N_28440);
nor UO_890 (O_890,N_27071,N_29021);
nor UO_891 (O_891,N_27135,N_28529);
nand UO_892 (O_892,N_27579,N_27274);
or UO_893 (O_893,N_27676,N_27189);
and UO_894 (O_894,N_27599,N_27424);
nor UO_895 (O_895,N_27143,N_28202);
or UO_896 (O_896,N_29076,N_27247);
nor UO_897 (O_897,N_27202,N_28927);
and UO_898 (O_898,N_27947,N_27904);
or UO_899 (O_899,N_29552,N_28497);
and UO_900 (O_900,N_29136,N_29414);
nor UO_901 (O_901,N_29434,N_29689);
and UO_902 (O_902,N_28389,N_29697);
or UO_903 (O_903,N_27042,N_27861);
and UO_904 (O_904,N_27478,N_28692);
nor UO_905 (O_905,N_28993,N_27882);
nor UO_906 (O_906,N_29153,N_28673);
nor UO_907 (O_907,N_27853,N_28836);
or UO_908 (O_908,N_29645,N_29714);
and UO_909 (O_909,N_28421,N_29948);
and UO_910 (O_910,N_28122,N_28414);
nand UO_911 (O_911,N_29029,N_28066);
or UO_912 (O_912,N_27085,N_28737);
and UO_913 (O_913,N_29516,N_28340);
or UO_914 (O_914,N_27955,N_28225);
nor UO_915 (O_915,N_29032,N_28278);
and UO_916 (O_916,N_27830,N_27332);
or UO_917 (O_917,N_27838,N_27034);
xnor UO_918 (O_918,N_27758,N_28239);
nand UO_919 (O_919,N_28940,N_29692);
xor UO_920 (O_920,N_28920,N_27168);
or UO_921 (O_921,N_27729,N_29866);
nor UO_922 (O_922,N_28172,N_29073);
nand UO_923 (O_923,N_29648,N_29454);
xor UO_924 (O_924,N_29326,N_27646);
nand UO_925 (O_925,N_29553,N_29261);
nand UO_926 (O_926,N_28720,N_28285);
nor UO_927 (O_927,N_29892,N_29550);
or UO_928 (O_928,N_28036,N_28126);
nand UO_929 (O_929,N_29025,N_28026);
and UO_930 (O_930,N_29612,N_27915);
nor UO_931 (O_931,N_29724,N_28528);
xor UO_932 (O_932,N_29556,N_28002);
nor UO_933 (O_933,N_27426,N_28600);
nand UO_934 (O_934,N_29876,N_27269);
nand UO_935 (O_935,N_27557,N_27829);
nand UO_936 (O_936,N_29270,N_27414);
and UO_937 (O_937,N_27988,N_28067);
and UO_938 (O_938,N_28550,N_29661);
nor UO_939 (O_939,N_27659,N_28419);
nor UO_940 (O_940,N_27964,N_27018);
and UO_941 (O_941,N_27666,N_28207);
and UO_942 (O_942,N_27041,N_29628);
nand UO_943 (O_943,N_28093,N_29528);
or UO_944 (O_944,N_28808,N_29040);
or UO_945 (O_945,N_27841,N_27802);
xnor UO_946 (O_946,N_28716,N_29510);
nand UO_947 (O_947,N_27883,N_27879);
or UO_948 (O_948,N_28304,N_28570);
nor UO_949 (O_949,N_29479,N_27067);
nand UO_950 (O_950,N_28527,N_28089);
xnor UO_951 (O_951,N_28361,N_27225);
nor UO_952 (O_952,N_27123,N_29314);
xor UO_953 (O_953,N_28327,N_29551);
and UO_954 (O_954,N_27384,N_29790);
nor UO_955 (O_955,N_29649,N_28398);
or UO_956 (O_956,N_27125,N_28838);
and UO_957 (O_957,N_29618,N_27236);
nand UO_958 (O_958,N_28354,N_29322);
nor UO_959 (O_959,N_28891,N_27860);
and UO_960 (O_960,N_28854,N_28579);
nand UO_961 (O_961,N_28956,N_29047);
nand UO_962 (O_962,N_28726,N_29572);
and UO_963 (O_963,N_29186,N_27986);
and UO_964 (O_964,N_27404,N_29627);
nor UO_965 (O_965,N_28551,N_27648);
nor UO_966 (O_966,N_28545,N_29992);
nand UO_967 (O_967,N_27482,N_29743);
and UO_968 (O_968,N_28660,N_28798);
nor UO_969 (O_969,N_27051,N_27726);
or UO_970 (O_970,N_27258,N_29672);
xnor UO_971 (O_971,N_27024,N_29321);
or UO_972 (O_972,N_29519,N_28759);
and UO_973 (O_973,N_28654,N_27326);
nand UO_974 (O_974,N_27405,N_27161);
nand UO_975 (O_975,N_28826,N_27690);
nand UO_976 (O_976,N_29496,N_29848);
and UO_977 (O_977,N_28637,N_28152);
nand UO_978 (O_978,N_27675,N_27778);
and UO_979 (O_979,N_27598,N_29619);
nand UO_980 (O_980,N_29930,N_28754);
nor UO_981 (O_981,N_29763,N_28050);
xor UO_982 (O_982,N_28858,N_28453);
nor UO_983 (O_983,N_28793,N_28567);
xor UO_984 (O_984,N_27747,N_27411);
and UO_985 (O_985,N_27221,N_27087);
nor UO_986 (O_986,N_27823,N_29432);
and UO_987 (O_987,N_29149,N_27595);
or UO_988 (O_988,N_28216,N_27309);
xnor UO_989 (O_989,N_27890,N_29632);
nand UO_990 (O_990,N_29028,N_27674);
and UO_991 (O_991,N_28061,N_27376);
nor UO_992 (O_992,N_28840,N_29016);
nor UO_993 (O_993,N_29355,N_27268);
xor UO_994 (O_994,N_29824,N_27863);
nand UO_995 (O_995,N_28332,N_29871);
and UO_996 (O_996,N_29253,N_29633);
nor UO_997 (O_997,N_28763,N_27490);
nor UO_998 (O_998,N_27294,N_29331);
and UO_999 (O_999,N_27222,N_28953);
or UO_1000 (O_1000,N_29057,N_27090);
and UO_1001 (O_1001,N_29172,N_29239);
nor UO_1002 (O_1002,N_27762,N_29708);
xnor UO_1003 (O_1003,N_29629,N_28513);
and UO_1004 (O_1004,N_28646,N_28430);
or UO_1005 (O_1005,N_28908,N_28481);
nand UO_1006 (O_1006,N_27641,N_27244);
nor UO_1007 (O_1007,N_29269,N_27832);
nand UO_1008 (O_1008,N_27150,N_28526);
nand UO_1009 (O_1009,N_29263,N_28649);
or UO_1010 (O_1010,N_29383,N_27966);
nor UO_1011 (O_1011,N_28046,N_28505);
or UO_1012 (O_1012,N_29820,N_27926);
or UO_1013 (O_1013,N_28240,N_28682);
and UO_1014 (O_1014,N_29792,N_27985);
nor UO_1015 (O_1015,N_28658,N_28054);
nand UO_1016 (O_1016,N_28922,N_27467);
xnor UO_1017 (O_1017,N_28199,N_27308);
xnor UO_1018 (O_1018,N_29463,N_29337);
and UO_1019 (O_1019,N_27183,N_28121);
nor UO_1020 (O_1020,N_29595,N_28633);
nor UO_1021 (O_1021,N_28862,N_27997);
or UO_1022 (O_1022,N_29456,N_28722);
xor UO_1023 (O_1023,N_28365,N_27788);
nor UO_1024 (O_1024,N_27276,N_29433);
or UO_1025 (O_1025,N_29809,N_28442);
xor UO_1026 (O_1026,N_29978,N_27917);
nand UO_1027 (O_1027,N_27604,N_27407);
or UO_1028 (O_1028,N_28917,N_29441);
xnor UO_1029 (O_1029,N_29218,N_27153);
and UO_1030 (O_1030,N_27626,N_27693);
or UO_1031 (O_1031,N_29833,N_27573);
and UO_1032 (O_1032,N_28696,N_29436);
and UO_1033 (O_1033,N_28995,N_29045);
nand UO_1034 (O_1034,N_28237,N_27976);
xnor UO_1035 (O_1035,N_29183,N_28813);
nor UO_1036 (O_1036,N_28869,N_28679);
nor UO_1037 (O_1037,N_28839,N_27992);
nand UO_1038 (O_1038,N_29426,N_28468);
and UO_1039 (O_1039,N_27354,N_28746);
xnor UO_1040 (O_1040,N_29442,N_28021);
xnor UO_1041 (O_1041,N_29376,N_29791);
nor UO_1042 (O_1042,N_29114,N_28341);
nand UO_1043 (O_1043,N_27614,N_28166);
and UO_1044 (O_1044,N_29140,N_29488);
nor UO_1045 (O_1045,N_28964,N_29578);
nor UO_1046 (O_1046,N_29280,N_27265);
and UO_1047 (O_1047,N_27141,N_29484);
nor UO_1048 (O_1048,N_27677,N_29814);
and UO_1049 (O_1049,N_27402,N_28159);
or UO_1050 (O_1050,N_29037,N_28976);
nor UO_1051 (O_1051,N_27428,N_27471);
xnor UO_1052 (O_1052,N_27800,N_28435);
and UO_1053 (O_1053,N_28587,N_28188);
and UO_1054 (O_1054,N_28127,N_27907);
xnor UO_1055 (O_1055,N_28029,N_27763);
and UO_1056 (O_1056,N_27450,N_29863);
and UO_1057 (O_1057,N_29769,N_29356);
or UO_1058 (O_1058,N_28634,N_27775);
xnor UO_1059 (O_1059,N_29719,N_29034);
nand UO_1060 (O_1060,N_27679,N_27182);
nor UO_1061 (O_1061,N_29558,N_29277);
nor UO_1062 (O_1062,N_27912,N_29059);
xor UO_1063 (O_1063,N_27186,N_27198);
xor UO_1064 (O_1064,N_29762,N_28723);
and UO_1065 (O_1065,N_27629,N_29589);
nand UO_1066 (O_1066,N_28721,N_29349);
nor UO_1067 (O_1067,N_27499,N_28317);
nand UO_1068 (O_1068,N_28845,N_27731);
nor UO_1069 (O_1069,N_27825,N_28275);
or UO_1070 (O_1070,N_28095,N_28339);
or UO_1071 (O_1071,N_29030,N_28073);
nand UO_1072 (O_1072,N_28612,N_29113);
xnor UO_1073 (O_1073,N_27516,N_29574);
xor UO_1074 (O_1074,N_29603,N_27213);
and UO_1075 (O_1075,N_28256,N_27192);
or UO_1076 (O_1076,N_28627,N_28936);
and UO_1077 (O_1077,N_28220,N_27931);
xnor UO_1078 (O_1078,N_27053,N_28707);
and UO_1079 (O_1079,N_28108,N_29005);
nor UO_1080 (O_1080,N_28083,N_28756);
and UO_1081 (O_1081,N_28303,N_27902);
nor UO_1082 (O_1082,N_29493,N_28645);
nor UO_1083 (O_1083,N_29055,N_28230);
nor UO_1084 (O_1084,N_27742,N_29737);
xor UO_1085 (O_1085,N_27010,N_27924);
or UO_1086 (O_1086,N_28433,N_28004);
nor UO_1087 (O_1087,N_28104,N_27935);
nor UO_1088 (O_1088,N_27187,N_28110);
or UO_1089 (O_1089,N_28728,N_27756);
nor UO_1090 (O_1090,N_29315,N_27122);
xnor UO_1091 (O_1091,N_27327,N_28103);
and UO_1092 (O_1092,N_27713,N_27603);
nand UO_1093 (O_1093,N_29622,N_28376);
and UO_1094 (O_1094,N_29245,N_27870);
and UO_1095 (O_1095,N_29566,N_29272);
nor UO_1096 (O_1096,N_29625,N_27893);
xor UO_1097 (O_1097,N_27302,N_28594);
nor UO_1098 (O_1098,N_29621,N_29870);
nand UO_1099 (O_1099,N_28294,N_28055);
xnor UO_1100 (O_1100,N_27553,N_27685);
or UO_1101 (O_1101,N_27231,N_29711);
xnor UO_1102 (O_1102,N_27706,N_27929);
nor UO_1103 (O_1103,N_27357,N_29804);
nand UO_1104 (O_1104,N_28475,N_27068);
nor UO_1105 (O_1105,N_29154,N_27755);
or UO_1106 (O_1106,N_27120,N_27792);
nand UO_1107 (O_1107,N_29226,N_27542);
or UO_1108 (O_1108,N_28283,N_27201);
and UO_1109 (O_1109,N_28474,N_27059);
nand UO_1110 (O_1110,N_28841,N_29777);
or UO_1111 (O_1111,N_29200,N_27716);
nand UO_1112 (O_1112,N_28413,N_29620);
or UO_1113 (O_1113,N_28942,N_28686);
xnor UO_1114 (O_1114,N_29869,N_29795);
nand UO_1115 (O_1115,N_29255,N_28429);
nor UO_1116 (O_1116,N_27708,N_28142);
nand UO_1117 (O_1117,N_27398,N_29990);
nand UO_1118 (O_1118,N_28792,N_27445);
and UO_1119 (O_1119,N_29268,N_29782);
xnor UO_1120 (O_1120,N_29970,N_27545);
nand UO_1121 (O_1121,N_29311,N_29662);
nor UO_1122 (O_1122,N_28153,N_28625);
or UO_1123 (O_1123,N_27259,N_28789);
xnor UO_1124 (O_1124,N_27728,N_28037);
nor UO_1125 (O_1125,N_29517,N_29606);
nand UO_1126 (O_1126,N_28355,N_27390);
nor UO_1127 (O_1127,N_28747,N_27810);
nand UO_1128 (O_1128,N_29143,N_28470);
and UO_1129 (O_1129,N_29506,N_27023);
nor UO_1130 (O_1130,N_27335,N_28472);
or UO_1131 (O_1131,N_28851,N_28013);
nor UO_1132 (O_1132,N_27174,N_28399);
and UO_1133 (O_1133,N_28008,N_29236);
nor UO_1134 (O_1134,N_29845,N_29688);
and UO_1135 (O_1135,N_28282,N_27963);
and UO_1136 (O_1136,N_27610,N_27670);
and UO_1137 (O_1137,N_29816,N_28669);
and UO_1138 (O_1138,N_27524,N_29273);
nand UO_1139 (O_1139,N_27709,N_29666);
or UO_1140 (O_1140,N_27905,N_27937);
or UO_1141 (O_1141,N_29292,N_27623);
xor UO_1142 (O_1142,N_28224,N_28501);
nor UO_1143 (O_1143,N_28350,N_29961);
nor UO_1144 (O_1144,N_29663,N_28989);
or UO_1145 (O_1145,N_27911,N_27510);
and UO_1146 (O_1146,N_29402,N_29225);
or UO_1147 (O_1147,N_29745,N_28546);
xor UO_1148 (O_1148,N_27208,N_27536);
xnor UO_1149 (O_1149,N_27978,N_28193);
xor UO_1150 (O_1150,N_29048,N_29515);
nand UO_1151 (O_1151,N_29391,N_29191);
and UO_1152 (O_1152,N_28974,N_27158);
xnor UO_1153 (O_1153,N_29605,N_27561);
nor UO_1154 (O_1154,N_29852,N_29329);
nor UO_1155 (O_1155,N_28511,N_28921);
xor UO_1156 (O_1156,N_27371,N_29257);
nor UO_1157 (O_1157,N_29888,N_28219);
and UO_1158 (O_1158,N_27452,N_28847);
nand UO_1159 (O_1159,N_28313,N_28311);
xor UO_1160 (O_1160,N_29600,N_27009);
nand UO_1161 (O_1161,N_27030,N_29836);
and UO_1162 (O_1162,N_27440,N_27529);
and UO_1163 (O_1163,N_29388,N_28588);
nor UO_1164 (O_1164,N_28185,N_28796);
or UO_1165 (O_1165,N_28766,N_28248);
xor UO_1166 (O_1166,N_28388,N_28058);
xor UO_1167 (O_1167,N_27286,N_27289);
and UO_1168 (O_1168,N_29103,N_29683);
or UO_1169 (O_1169,N_29354,N_28525);
xor UO_1170 (O_1170,N_28503,N_28867);
or UO_1171 (O_1171,N_27281,N_28959);
and UO_1172 (O_1172,N_29690,N_29156);
nand UO_1173 (O_1173,N_29054,N_27563);
xor UO_1174 (O_1174,N_27635,N_29152);
xor UO_1175 (O_1175,N_27700,N_28374);
xnor UO_1176 (O_1176,N_28234,N_29265);
nor UO_1177 (O_1177,N_29652,N_27807);
or UO_1178 (O_1178,N_28496,N_27697);
nor UO_1179 (O_1179,N_29228,N_28400);
nor UO_1180 (O_1180,N_28105,N_27142);
nor UO_1181 (O_1181,N_29676,N_28730);
and UO_1182 (O_1182,N_28599,N_28607);
xnor UO_1183 (O_1183,N_27584,N_27104);
or UO_1184 (O_1184,N_27686,N_27319);
xor UO_1185 (O_1185,N_27715,N_28384);
nor UO_1186 (O_1186,N_29313,N_29968);
nand UO_1187 (O_1187,N_27574,N_27025);
nand UO_1188 (O_1188,N_28261,N_27627);
and UO_1189 (O_1189,N_27855,N_28119);
nor UO_1190 (O_1190,N_27899,N_28945);
nand UO_1191 (O_1191,N_27872,N_27311);
or UO_1192 (O_1192,N_29009,N_29339);
and UO_1193 (O_1193,N_28351,N_29297);
xor UO_1194 (O_1194,N_29065,N_29064);
xor UO_1195 (O_1195,N_28614,N_28913);
nor UO_1196 (O_1196,N_28352,N_28972);
and UO_1197 (O_1197,N_28243,N_28572);
nand UO_1198 (O_1198,N_28884,N_27081);
and UO_1199 (O_1199,N_28786,N_29828);
nor UO_1200 (O_1200,N_29094,N_28828);
or UO_1201 (O_1201,N_29682,N_28760);
or UO_1202 (O_1202,N_27655,N_27447);
and UO_1203 (O_1203,N_29675,N_27865);
nand UO_1204 (O_1204,N_27248,N_29461);
xor UO_1205 (O_1205,N_28944,N_27885);
xor UO_1206 (O_1206,N_27164,N_29400);
or UO_1207 (O_1207,N_29750,N_28564);
or UO_1208 (O_1208,N_28397,N_29995);
or UO_1209 (O_1209,N_27571,N_28137);
or UO_1210 (O_1210,N_28930,N_29018);
nor UO_1211 (O_1211,N_27712,N_29131);
nor UO_1212 (O_1212,N_27779,N_29323);
xnor UO_1213 (O_1213,N_29167,N_28610);
xnor UO_1214 (O_1214,N_29374,N_27002);
nand UO_1215 (O_1215,N_29548,N_29278);
nor UO_1216 (O_1216,N_29886,N_28208);
nor UO_1217 (O_1217,N_27602,N_28580);
and UO_1218 (O_1218,N_28381,N_28205);
or UO_1219 (O_1219,N_28375,N_29166);
or UO_1220 (O_1220,N_29427,N_28186);
xnor UO_1221 (O_1221,N_27057,N_27689);
and UO_1222 (O_1222,N_29404,N_29916);
nand UO_1223 (O_1223,N_29056,N_27620);
xor UO_1224 (O_1224,N_29450,N_27306);
nand UO_1225 (O_1225,N_29546,N_27393);
nand UO_1226 (O_1226,N_29051,N_29984);
or UO_1227 (O_1227,N_27809,N_28832);
and UO_1228 (O_1228,N_27734,N_28986);
nand UO_1229 (O_1229,N_27485,N_27435);
nand UO_1230 (O_1230,N_28270,N_29731);
nand UO_1231 (O_1231,N_27195,N_28330);
and UO_1232 (O_1232,N_28167,N_29477);
nand UO_1233 (O_1233,N_28009,N_29798);
xnor UO_1234 (O_1234,N_29969,N_29765);
nor UO_1235 (O_1235,N_28675,N_29859);
nor UO_1236 (O_1236,N_27204,N_29157);
nand UO_1237 (O_1237,N_28274,N_28911);
and UO_1238 (O_1238,N_28748,N_28473);
nand UO_1239 (O_1239,N_29429,N_28773);
nor UO_1240 (O_1240,N_29977,N_29774);
nand UO_1241 (O_1241,N_29917,N_28309);
and UO_1242 (O_1242,N_27253,N_29740);
nand UO_1243 (O_1243,N_27209,N_27995);
or UO_1244 (O_1244,N_29198,N_29232);
or UO_1245 (O_1245,N_28532,N_27920);
and UO_1246 (O_1246,N_29538,N_28176);
or UO_1247 (O_1247,N_29453,N_29807);
and UO_1248 (O_1248,N_29410,N_27295);
and UO_1249 (O_1249,N_27813,N_29408);
and UO_1250 (O_1250,N_29579,N_27821);
nand UO_1251 (O_1251,N_29623,N_27636);
nand UO_1252 (O_1252,N_29377,N_28291);
and UO_1253 (O_1253,N_27794,N_29974);
xnor UO_1254 (O_1254,N_28639,N_29309);
or UO_1255 (O_1255,N_27895,N_27401);
and UO_1256 (O_1256,N_27044,N_28360);
and UO_1257 (O_1257,N_29171,N_27381);
and UO_1258 (O_1258,N_27566,N_28292);
xor UO_1259 (O_1259,N_29445,N_28006);
or UO_1260 (O_1260,N_28879,N_29262);
or UO_1261 (O_1261,N_28910,N_28469);
and UO_1262 (O_1262,N_28080,N_27263);
and UO_1263 (O_1263,N_29501,N_29571);
xor UO_1264 (O_1264,N_29139,N_27961);
and UO_1265 (O_1265,N_27575,N_28463);
nor UO_1266 (O_1266,N_28848,N_29779);
xnor UO_1267 (O_1267,N_28557,N_27273);
nor UO_1268 (O_1268,N_27803,N_28402);
xor UO_1269 (O_1269,N_28112,N_27365);
or UO_1270 (O_1270,N_28018,N_29173);
and UO_1271 (O_1271,N_29026,N_27640);
xnor UO_1272 (O_1272,N_28688,N_27412);
and UO_1273 (O_1273,N_28905,N_29416);
nand UO_1274 (O_1274,N_28975,N_28690);
xnor UO_1275 (O_1275,N_29130,N_28245);
xor UO_1276 (O_1276,N_29544,N_29042);
nand UO_1277 (O_1277,N_29537,N_29831);
or UO_1278 (O_1278,N_27369,N_29706);
nor UO_1279 (O_1279,N_29993,N_27967);
nor UO_1280 (O_1280,N_29761,N_29540);
nor UO_1281 (O_1281,N_28047,N_28450);
nor UO_1282 (O_1282,N_27814,N_27422);
xnor UO_1283 (O_1283,N_29116,N_28797);
nand UO_1284 (O_1284,N_28032,N_29855);
nand UO_1285 (O_1285,N_28713,N_27397);
nor UO_1286 (O_1286,N_28810,N_28232);
nand UO_1287 (O_1287,N_27382,N_29929);
nand UO_1288 (O_1288,N_28709,N_29220);
or UO_1289 (O_1289,N_29874,N_27460);
nand UO_1290 (O_1290,N_28487,N_27869);
xor UO_1291 (O_1291,N_29431,N_29002);
nand UO_1292 (O_1292,N_28504,N_27035);
xnor UO_1293 (O_1293,N_28128,N_27240);
xor UO_1294 (O_1294,N_27430,N_29583);
and UO_1295 (O_1295,N_27484,N_27331);
nor UO_1296 (O_1296,N_27086,N_27513);
nand UO_1297 (O_1297,N_29640,N_28231);
nor UO_1298 (O_1298,N_28387,N_29835);
or UO_1299 (O_1299,N_28742,N_27089);
xor UO_1300 (O_1300,N_28437,N_29507);
xor UO_1301 (O_1301,N_27934,N_28403);
and UO_1302 (O_1302,N_27776,N_27379);
and UO_1303 (O_1303,N_28386,N_27003);
or UO_1304 (O_1304,N_28590,N_29010);
nor UO_1305 (O_1305,N_28943,N_29801);
or UO_1306 (O_1306,N_28493,N_29285);
and UO_1307 (O_1307,N_28485,N_28300);
nor UO_1308 (O_1308,N_27668,N_29451);
xor UO_1309 (O_1309,N_28712,N_27436);
nor UO_1310 (O_1310,N_29610,N_28214);
xnor UO_1311 (O_1311,N_29999,N_29591);
nand UO_1312 (O_1312,N_28393,N_29958);
nor UO_1313 (O_1313,N_27798,N_27537);
and UO_1314 (O_1314,N_29665,N_27481);
and UO_1315 (O_1315,N_29327,N_27305);
xnor UO_1316 (O_1316,N_27960,N_28038);
and UO_1317 (O_1317,N_27867,N_28259);
nand UO_1318 (O_1318,N_29264,N_28241);
or UO_1319 (O_1319,N_27300,N_27014);
and UO_1320 (O_1320,N_27437,N_28233);
nand UO_1321 (O_1321,N_28591,N_29093);
nor UO_1322 (O_1322,N_29639,N_27334);
nor UO_1323 (O_1323,N_29674,N_27062);
nor UO_1324 (O_1324,N_29960,N_29832);
nor UO_1325 (O_1325,N_28547,N_27166);
xnor UO_1326 (O_1326,N_29212,N_27866);
xor UO_1327 (O_1327,N_28253,N_29412);
xnor UO_1328 (O_1328,N_27826,N_29180);
and UO_1329 (O_1329,N_27739,N_29825);
or UO_1330 (O_1330,N_29340,N_28043);
xnor UO_1331 (O_1331,N_29207,N_28987);
and UO_1332 (O_1332,N_27720,N_29421);
or UO_1333 (O_1333,N_29607,N_27270);
nand UO_1334 (O_1334,N_27791,N_27767);
nand UO_1335 (O_1335,N_29817,N_29936);
nor UO_1336 (O_1336,N_29079,N_29148);
and UO_1337 (O_1337,N_27642,N_27366);
xor UO_1338 (O_1338,N_29233,N_29812);
nor UO_1339 (O_1339,N_27787,N_29112);
and UO_1340 (O_1340,N_27654,N_28576);
or UO_1341 (O_1341,N_29775,N_29856);
nand UO_1342 (O_1342,N_28899,N_28855);
nor UO_1343 (O_1343,N_29865,N_28416);
nand UO_1344 (O_1344,N_28680,N_27922);
or UO_1345 (O_1345,N_27589,N_27262);
and UO_1346 (O_1346,N_27725,N_27491);
xnor UO_1347 (O_1347,N_27523,N_27898);
xor UO_1348 (O_1348,N_28597,N_29090);
nand UO_1349 (O_1349,N_27738,N_27399);
and UO_1350 (O_1350,N_27847,N_29336);
or UO_1351 (O_1351,N_27283,N_28988);
nor UO_1352 (O_1352,N_28483,N_29772);
nand UO_1353 (O_1353,N_27012,N_27649);
nand UO_1354 (O_1354,N_29781,N_28781);
and UO_1355 (O_1355,N_28898,N_27624);
nor UO_1356 (O_1356,N_27227,N_29943);
nand UO_1357 (O_1357,N_27134,N_28829);
or UO_1358 (O_1358,N_27036,N_29120);
or UO_1359 (O_1359,N_29004,N_28308);
or UO_1360 (O_1360,N_28775,N_28925);
xor UO_1361 (O_1361,N_28717,N_28048);
or UO_1362 (O_1362,N_27130,N_29890);
or UO_1363 (O_1363,N_29495,N_29003);
xnor UO_1364 (O_1364,N_28428,N_27267);
nand UO_1365 (O_1365,N_27056,N_29145);
nor UO_1366 (O_1366,N_27495,N_27568);
nor UO_1367 (O_1367,N_29955,N_27980);
nand UO_1368 (O_1368,N_27226,N_28765);
nor UO_1369 (O_1369,N_27312,N_29635);
or UO_1370 (O_1370,N_29568,N_28180);
nor UO_1371 (O_1371,N_27353,N_29980);
xor UO_1372 (O_1372,N_29284,N_28880);
and UO_1373 (O_1373,N_29447,N_29256);
nand UO_1374 (O_1374,N_29485,N_27344);
xnor UO_1375 (O_1375,N_29709,N_28894);
nor UO_1376 (O_1376,N_29687,N_27520);
or UO_1377 (O_1377,N_28068,N_28563);
and UO_1378 (O_1378,N_27957,N_28488);
nand UO_1379 (O_1379,N_29841,N_28163);
nand UO_1380 (O_1380,N_27554,N_29526);
and UO_1381 (O_1381,N_29677,N_27497);
nand UO_1382 (O_1382,N_28051,N_29368);
nand UO_1383 (O_1383,N_29370,N_29108);
nand UO_1384 (O_1384,N_27217,N_28984);
nor UO_1385 (O_1385,N_29291,N_28609);
xor UO_1386 (O_1386,N_29119,N_29407);
nor UO_1387 (O_1387,N_27077,N_27943);
or UO_1388 (O_1388,N_29834,N_28177);
nand UO_1389 (O_1389,N_27298,N_27699);
nand UO_1390 (O_1390,N_28672,N_28209);
or UO_1391 (O_1391,N_28700,N_29015);
and UO_1392 (O_1392,N_29294,N_28293);
nor UO_1393 (O_1393,N_29592,N_27324);
nand UO_1394 (O_1394,N_29243,N_29927);
and UO_1395 (O_1395,N_27799,N_29994);
or UO_1396 (O_1396,N_29448,N_28204);
xor UO_1397 (O_1397,N_27330,N_27894);
nand UO_1398 (O_1398,N_27026,N_27736);
nand UO_1399 (O_1399,N_28427,N_27694);
xnor UO_1400 (O_1400,N_27112,N_29720);
or UO_1401 (O_1401,N_29921,N_27028);
nor UO_1402 (O_1402,N_27292,N_28373);
nor UO_1403 (O_1403,N_29912,N_27022);
xnor UO_1404 (O_1404,N_27889,N_28190);
and UO_1405 (O_1405,N_29137,N_29164);
or UO_1406 (O_1406,N_29162,N_27140);
or UO_1407 (O_1407,N_29962,N_29698);
and UO_1408 (O_1408,N_28409,N_29413);
nand UO_1409 (O_1409,N_28380,N_29411);
and UO_1410 (O_1410,N_27069,N_27260);
xor UO_1411 (O_1411,N_27993,N_28024);
nand UO_1412 (O_1412,N_29796,N_29063);
or UO_1413 (O_1413,N_27951,N_29716);
and UO_1414 (O_1414,N_28823,N_28958);
and UO_1415 (O_1415,N_28206,N_27054);
nand UO_1416 (O_1416,N_27037,N_29799);
xor UO_1417 (O_1417,N_28377,N_27783);
xnor UO_1418 (O_1418,N_29012,N_29237);
nand UO_1419 (O_1419,N_29872,N_28844);
xor UO_1420 (O_1420,N_29565,N_27549);
nand UO_1421 (O_1421,N_29884,N_27255);
nor UO_1422 (O_1422,N_27583,N_29214);
nor UO_1423 (O_1423,N_29462,N_28699);
nand UO_1424 (O_1424,N_28674,N_27786);
or UO_1425 (O_1425,N_28144,N_27441);
or UO_1426 (O_1426,N_28788,N_28873);
nand UO_1427 (O_1427,N_27845,N_28236);
or UO_1428 (O_1428,N_27663,N_28621);
and UO_1429 (O_1429,N_27496,N_28120);
nor UO_1430 (O_1430,N_29638,N_27486);
nand UO_1431 (O_1431,N_28139,N_27909);
or UO_1432 (O_1432,N_29074,N_27064);
nor UO_1433 (O_1433,N_29347,N_27333);
nand UO_1434 (O_1434,N_29227,N_29020);
xor UO_1435 (O_1435,N_28906,N_29231);
xnor UO_1436 (O_1436,N_28794,N_28320);
nand UO_1437 (O_1437,N_28287,N_27358);
xnor UO_1438 (O_1438,N_29797,N_29302);
or UO_1439 (O_1439,N_29654,N_29142);
and UO_1440 (O_1440,N_29435,N_29117);
and UO_1441 (O_1441,N_29827,N_29513);
xor UO_1442 (O_1442,N_28961,N_28312);
xor UO_1443 (O_1443,N_28466,N_29944);
nor UO_1444 (O_1444,N_29254,N_27375);
and UO_1445 (O_1445,N_29380,N_29685);
nor UO_1446 (O_1446,N_28565,N_29242);
nand UO_1447 (O_1447,N_27409,N_29174);
and UO_1448 (O_1448,N_29525,N_28369);
nor UO_1449 (O_1449,N_29299,N_28581);
nand UO_1450 (O_1450,N_27238,N_27307);
xnor UO_1451 (O_1451,N_29594,N_29611);
xor UO_1452 (O_1452,N_29345,N_27631);
and UO_1453 (O_1453,N_27812,N_29008);
nor UO_1454 (O_1454,N_28405,N_27181);
and UO_1455 (O_1455,N_27769,N_27842);
nand UO_1456 (O_1456,N_27930,N_27661);
or UO_1457 (O_1457,N_29887,N_29293);
and UO_1458 (O_1458,N_27981,N_28042);
xnor UO_1459 (O_1459,N_28226,N_27102);
or UO_1460 (O_1460,N_29333,N_27242);
or UO_1461 (O_1461,N_29942,N_28212);
xnor UO_1462 (O_1462,N_27506,N_27043);
nand UO_1463 (O_1463,N_28478,N_29947);
nor UO_1464 (O_1464,N_27586,N_29502);
and UO_1465 (O_1465,N_28333,N_28025);
xor UO_1466 (O_1466,N_28424,N_27205);
or UO_1467 (O_1467,N_28659,N_28653);
or UO_1468 (O_1468,N_28800,N_27871);
nor UO_1469 (O_1469,N_28091,N_28257);
and UO_1470 (O_1470,N_29905,N_27517);
or UO_1471 (O_1471,N_27528,N_28738);
nand UO_1472 (O_1472,N_28370,N_29274);
and UO_1473 (O_1473,N_29985,N_29185);
nor UO_1474 (O_1474,N_27279,N_28510);
nor UO_1475 (O_1475,N_27096,N_29979);
nand UO_1476 (O_1476,N_27859,N_28507);
and UO_1477 (O_1477,N_27892,N_29966);
xor UO_1478 (O_1478,N_27946,N_28434);
or UO_1479 (O_1479,N_28556,N_27970);
nand UO_1480 (O_1480,N_29911,N_27925);
xor UO_1481 (O_1481,N_29786,N_27252);
xnor UO_1482 (O_1482,N_27162,N_29260);
xor UO_1483 (O_1483,N_27193,N_27105);
and UO_1484 (O_1484,N_28743,N_29573);
and UO_1485 (O_1485,N_28968,N_27881);
xor UO_1486 (O_1486,N_27083,N_28771);
xor UO_1487 (O_1487,N_27342,N_28390);
nor UO_1488 (O_1488,N_28356,N_27601);
nand UO_1489 (O_1489,N_29536,N_29249);
nand UO_1490 (O_1490,N_29667,N_29155);
nor UO_1491 (O_1491,N_28175,N_27138);
and UO_1492 (O_1492,N_28077,N_27277);
nor UO_1493 (O_1493,N_29767,N_29096);
and UO_1494 (O_1494,N_29335,N_29381);
xor UO_1495 (O_1495,N_28991,N_28685);
nor UO_1496 (O_1496,N_29046,N_28295);
and UO_1497 (O_1497,N_28129,N_28767);
or UO_1498 (O_1498,N_29440,N_28656);
and UO_1499 (O_1499,N_29722,N_27380);
or UO_1500 (O_1500,N_28603,N_27740);
xnor UO_1501 (O_1501,N_27578,N_27066);
nand UO_1502 (O_1502,N_28618,N_28265);
xor UO_1503 (O_1503,N_29806,N_28478);
and UO_1504 (O_1504,N_29515,N_29362);
xor UO_1505 (O_1505,N_28846,N_29802);
and UO_1506 (O_1506,N_28909,N_27245);
and UO_1507 (O_1507,N_29537,N_29809);
nand UO_1508 (O_1508,N_28885,N_29186);
and UO_1509 (O_1509,N_27415,N_27279);
or UO_1510 (O_1510,N_29105,N_27517);
or UO_1511 (O_1511,N_27205,N_27923);
and UO_1512 (O_1512,N_27496,N_28269);
or UO_1513 (O_1513,N_29031,N_29069);
nand UO_1514 (O_1514,N_28316,N_28657);
xnor UO_1515 (O_1515,N_27065,N_28501);
xor UO_1516 (O_1516,N_29063,N_28236);
xnor UO_1517 (O_1517,N_28754,N_27752);
xor UO_1518 (O_1518,N_27602,N_28937);
nor UO_1519 (O_1519,N_27994,N_28019);
or UO_1520 (O_1520,N_28893,N_28359);
xnor UO_1521 (O_1521,N_28394,N_29212);
nor UO_1522 (O_1522,N_27987,N_28961);
nor UO_1523 (O_1523,N_29312,N_29666);
xnor UO_1524 (O_1524,N_27952,N_29352);
nand UO_1525 (O_1525,N_27131,N_28694);
or UO_1526 (O_1526,N_27598,N_28483);
nor UO_1527 (O_1527,N_28530,N_28823);
nand UO_1528 (O_1528,N_28788,N_28891);
and UO_1529 (O_1529,N_29305,N_29920);
nand UO_1530 (O_1530,N_29620,N_28332);
xor UO_1531 (O_1531,N_29481,N_29224);
and UO_1532 (O_1532,N_28631,N_29276);
or UO_1533 (O_1533,N_28983,N_28743);
or UO_1534 (O_1534,N_28598,N_27857);
or UO_1535 (O_1535,N_29104,N_27670);
or UO_1536 (O_1536,N_27191,N_27818);
xor UO_1537 (O_1537,N_27546,N_29201);
or UO_1538 (O_1538,N_28767,N_28686);
nor UO_1539 (O_1539,N_29997,N_27038);
or UO_1540 (O_1540,N_28000,N_27241);
and UO_1541 (O_1541,N_29357,N_27209);
and UO_1542 (O_1542,N_28822,N_29145);
nor UO_1543 (O_1543,N_27823,N_29139);
xnor UO_1544 (O_1544,N_27318,N_28874);
or UO_1545 (O_1545,N_27447,N_29128);
xnor UO_1546 (O_1546,N_28034,N_28721);
nand UO_1547 (O_1547,N_27095,N_27353);
and UO_1548 (O_1548,N_29850,N_29887);
nor UO_1549 (O_1549,N_27467,N_29961);
and UO_1550 (O_1550,N_27112,N_29012);
or UO_1551 (O_1551,N_27435,N_28218);
or UO_1552 (O_1552,N_29725,N_29578);
nand UO_1553 (O_1553,N_27243,N_27563);
nand UO_1554 (O_1554,N_27727,N_27174);
nor UO_1555 (O_1555,N_29218,N_28512);
nor UO_1556 (O_1556,N_28758,N_29241);
nor UO_1557 (O_1557,N_28510,N_29779);
nor UO_1558 (O_1558,N_27194,N_27647);
xnor UO_1559 (O_1559,N_28369,N_29708);
nand UO_1560 (O_1560,N_27903,N_29280);
and UO_1561 (O_1561,N_29971,N_29767);
nor UO_1562 (O_1562,N_28784,N_27842);
or UO_1563 (O_1563,N_29575,N_28896);
nand UO_1564 (O_1564,N_28337,N_29515);
and UO_1565 (O_1565,N_29940,N_28390);
nand UO_1566 (O_1566,N_28548,N_27643);
nand UO_1567 (O_1567,N_27602,N_29128);
and UO_1568 (O_1568,N_28345,N_28493);
or UO_1569 (O_1569,N_28860,N_27701);
nand UO_1570 (O_1570,N_27317,N_29476);
xor UO_1571 (O_1571,N_28513,N_29201);
xor UO_1572 (O_1572,N_27146,N_29847);
and UO_1573 (O_1573,N_29833,N_28382);
nor UO_1574 (O_1574,N_29014,N_27940);
xnor UO_1575 (O_1575,N_28636,N_29715);
and UO_1576 (O_1576,N_27704,N_28406);
or UO_1577 (O_1577,N_29986,N_29398);
nand UO_1578 (O_1578,N_29989,N_27014);
xnor UO_1579 (O_1579,N_29845,N_28784);
xor UO_1580 (O_1580,N_29105,N_28826);
and UO_1581 (O_1581,N_29979,N_28387);
xnor UO_1582 (O_1582,N_29692,N_29390);
nand UO_1583 (O_1583,N_28321,N_29089);
and UO_1584 (O_1584,N_29268,N_28944);
or UO_1585 (O_1585,N_29967,N_28363);
or UO_1586 (O_1586,N_28662,N_28431);
xor UO_1587 (O_1587,N_28662,N_27416);
or UO_1588 (O_1588,N_27197,N_29327);
and UO_1589 (O_1589,N_29027,N_28537);
or UO_1590 (O_1590,N_29354,N_28995);
xnor UO_1591 (O_1591,N_27258,N_29575);
nor UO_1592 (O_1592,N_27612,N_27112);
xnor UO_1593 (O_1593,N_29263,N_28563);
or UO_1594 (O_1594,N_27460,N_28806);
xor UO_1595 (O_1595,N_28608,N_27590);
and UO_1596 (O_1596,N_28149,N_27235);
nor UO_1597 (O_1597,N_29562,N_27986);
or UO_1598 (O_1598,N_29011,N_29475);
and UO_1599 (O_1599,N_28054,N_29337);
nand UO_1600 (O_1600,N_29642,N_29846);
and UO_1601 (O_1601,N_28577,N_27193);
xor UO_1602 (O_1602,N_28124,N_27547);
and UO_1603 (O_1603,N_29577,N_27308);
xor UO_1604 (O_1604,N_27384,N_29165);
or UO_1605 (O_1605,N_28084,N_28789);
and UO_1606 (O_1606,N_28226,N_27303);
and UO_1607 (O_1607,N_27857,N_29586);
xnor UO_1608 (O_1608,N_27277,N_28116);
nor UO_1609 (O_1609,N_29704,N_28402);
xnor UO_1610 (O_1610,N_29532,N_28439);
xnor UO_1611 (O_1611,N_27698,N_29442);
nand UO_1612 (O_1612,N_28638,N_27903);
or UO_1613 (O_1613,N_29368,N_27481);
xor UO_1614 (O_1614,N_27298,N_27801);
nor UO_1615 (O_1615,N_29618,N_28657);
nand UO_1616 (O_1616,N_28065,N_28844);
or UO_1617 (O_1617,N_27884,N_27438);
or UO_1618 (O_1618,N_28221,N_27235);
xor UO_1619 (O_1619,N_27969,N_27474);
or UO_1620 (O_1620,N_28873,N_29927);
and UO_1621 (O_1621,N_28952,N_29402);
and UO_1622 (O_1622,N_28965,N_28233);
or UO_1623 (O_1623,N_29214,N_28425);
and UO_1624 (O_1624,N_28025,N_29451);
or UO_1625 (O_1625,N_28207,N_29386);
nor UO_1626 (O_1626,N_29717,N_29429);
and UO_1627 (O_1627,N_29064,N_29767);
and UO_1628 (O_1628,N_28071,N_27481);
nor UO_1629 (O_1629,N_29506,N_29743);
nor UO_1630 (O_1630,N_29460,N_28933);
and UO_1631 (O_1631,N_27425,N_27413);
nor UO_1632 (O_1632,N_28607,N_28444);
nor UO_1633 (O_1633,N_27666,N_29776);
and UO_1634 (O_1634,N_27836,N_28730);
nand UO_1635 (O_1635,N_29141,N_29726);
and UO_1636 (O_1636,N_28003,N_27902);
xor UO_1637 (O_1637,N_28803,N_28671);
nand UO_1638 (O_1638,N_28501,N_28887);
nor UO_1639 (O_1639,N_29443,N_29243);
or UO_1640 (O_1640,N_27014,N_28655);
xnor UO_1641 (O_1641,N_28301,N_29246);
and UO_1642 (O_1642,N_29673,N_27809);
or UO_1643 (O_1643,N_29938,N_28102);
or UO_1644 (O_1644,N_29366,N_28971);
or UO_1645 (O_1645,N_28138,N_29683);
and UO_1646 (O_1646,N_28135,N_27715);
and UO_1647 (O_1647,N_28160,N_27396);
and UO_1648 (O_1648,N_29067,N_28065);
or UO_1649 (O_1649,N_27382,N_28608);
or UO_1650 (O_1650,N_28392,N_29734);
nor UO_1651 (O_1651,N_28037,N_27296);
xnor UO_1652 (O_1652,N_27230,N_27136);
nand UO_1653 (O_1653,N_29402,N_28652);
nand UO_1654 (O_1654,N_28984,N_27116);
or UO_1655 (O_1655,N_28699,N_29569);
and UO_1656 (O_1656,N_29467,N_29607);
nand UO_1657 (O_1657,N_27875,N_27302);
xnor UO_1658 (O_1658,N_27715,N_27143);
nand UO_1659 (O_1659,N_29285,N_27536);
xor UO_1660 (O_1660,N_28540,N_29000);
nand UO_1661 (O_1661,N_27564,N_27241);
nor UO_1662 (O_1662,N_28806,N_27660);
or UO_1663 (O_1663,N_29380,N_28787);
xnor UO_1664 (O_1664,N_27790,N_27734);
or UO_1665 (O_1665,N_27019,N_28184);
nor UO_1666 (O_1666,N_28326,N_27829);
and UO_1667 (O_1667,N_28823,N_28944);
nor UO_1668 (O_1668,N_29712,N_27663);
xnor UO_1669 (O_1669,N_29495,N_28531);
nand UO_1670 (O_1670,N_27670,N_28506);
nand UO_1671 (O_1671,N_27471,N_27299);
nand UO_1672 (O_1672,N_28460,N_27502);
xor UO_1673 (O_1673,N_28123,N_28825);
xnor UO_1674 (O_1674,N_28718,N_29319);
and UO_1675 (O_1675,N_29552,N_28153);
or UO_1676 (O_1676,N_27952,N_28433);
nand UO_1677 (O_1677,N_28916,N_29585);
xor UO_1678 (O_1678,N_29940,N_28531);
or UO_1679 (O_1679,N_27461,N_27556);
or UO_1680 (O_1680,N_27160,N_28438);
nor UO_1681 (O_1681,N_28549,N_28556);
and UO_1682 (O_1682,N_27929,N_27268);
xnor UO_1683 (O_1683,N_28006,N_28365);
or UO_1684 (O_1684,N_29244,N_28053);
xor UO_1685 (O_1685,N_27202,N_27773);
or UO_1686 (O_1686,N_27896,N_29548);
nor UO_1687 (O_1687,N_28440,N_27529);
or UO_1688 (O_1688,N_29713,N_28238);
xor UO_1689 (O_1689,N_27828,N_27633);
nor UO_1690 (O_1690,N_29851,N_28475);
or UO_1691 (O_1691,N_28870,N_29168);
nor UO_1692 (O_1692,N_29522,N_27928);
xnor UO_1693 (O_1693,N_27658,N_28066);
or UO_1694 (O_1694,N_28528,N_28896);
or UO_1695 (O_1695,N_27664,N_28382);
nand UO_1696 (O_1696,N_29559,N_29059);
nor UO_1697 (O_1697,N_28504,N_29047);
and UO_1698 (O_1698,N_27981,N_28706);
nand UO_1699 (O_1699,N_27727,N_28467);
or UO_1700 (O_1700,N_28283,N_29743);
or UO_1701 (O_1701,N_29259,N_29921);
nor UO_1702 (O_1702,N_29899,N_29069);
xnor UO_1703 (O_1703,N_29520,N_29544);
nand UO_1704 (O_1704,N_29527,N_29290);
xnor UO_1705 (O_1705,N_27906,N_27539);
nand UO_1706 (O_1706,N_27313,N_28755);
nand UO_1707 (O_1707,N_29415,N_29536);
nor UO_1708 (O_1708,N_28815,N_27863);
nand UO_1709 (O_1709,N_27067,N_28933);
or UO_1710 (O_1710,N_28179,N_29841);
and UO_1711 (O_1711,N_27256,N_28319);
and UO_1712 (O_1712,N_28478,N_29647);
nand UO_1713 (O_1713,N_27375,N_29424);
nand UO_1714 (O_1714,N_27201,N_28231);
nand UO_1715 (O_1715,N_28058,N_28254);
or UO_1716 (O_1716,N_27147,N_27695);
nor UO_1717 (O_1717,N_27711,N_27408);
xor UO_1718 (O_1718,N_28107,N_28462);
or UO_1719 (O_1719,N_29413,N_28526);
or UO_1720 (O_1720,N_27787,N_29831);
or UO_1721 (O_1721,N_27239,N_29227);
nand UO_1722 (O_1722,N_28167,N_29196);
xnor UO_1723 (O_1723,N_28739,N_29625);
nand UO_1724 (O_1724,N_28042,N_29034);
nand UO_1725 (O_1725,N_29581,N_27338);
nand UO_1726 (O_1726,N_28766,N_27673);
nand UO_1727 (O_1727,N_29273,N_27893);
or UO_1728 (O_1728,N_29741,N_27560);
xor UO_1729 (O_1729,N_29389,N_28360);
xor UO_1730 (O_1730,N_27244,N_29136);
and UO_1731 (O_1731,N_29057,N_28962);
nand UO_1732 (O_1732,N_29272,N_27906);
and UO_1733 (O_1733,N_27518,N_29696);
nand UO_1734 (O_1734,N_28402,N_29553);
or UO_1735 (O_1735,N_29551,N_28820);
xnor UO_1736 (O_1736,N_28251,N_27846);
nor UO_1737 (O_1737,N_29182,N_27855);
or UO_1738 (O_1738,N_29925,N_27693);
nand UO_1739 (O_1739,N_27092,N_27898);
or UO_1740 (O_1740,N_29920,N_28548);
or UO_1741 (O_1741,N_28644,N_27938);
and UO_1742 (O_1742,N_29509,N_28728);
and UO_1743 (O_1743,N_28803,N_28497);
nand UO_1744 (O_1744,N_28405,N_27732);
nand UO_1745 (O_1745,N_28328,N_28648);
nand UO_1746 (O_1746,N_27989,N_27891);
nor UO_1747 (O_1747,N_29730,N_28077);
nand UO_1748 (O_1748,N_29755,N_27479);
or UO_1749 (O_1749,N_28225,N_28412);
or UO_1750 (O_1750,N_28304,N_29316);
or UO_1751 (O_1751,N_27975,N_27343);
xnor UO_1752 (O_1752,N_29491,N_28724);
or UO_1753 (O_1753,N_27639,N_29417);
xnor UO_1754 (O_1754,N_27001,N_28923);
xnor UO_1755 (O_1755,N_27550,N_28028);
xor UO_1756 (O_1756,N_27234,N_29652);
nor UO_1757 (O_1757,N_28402,N_29891);
xnor UO_1758 (O_1758,N_29118,N_29938);
nor UO_1759 (O_1759,N_28523,N_28190);
or UO_1760 (O_1760,N_27176,N_27073);
and UO_1761 (O_1761,N_29574,N_27791);
or UO_1762 (O_1762,N_28906,N_29471);
nor UO_1763 (O_1763,N_28823,N_27538);
or UO_1764 (O_1764,N_27068,N_28968);
nand UO_1765 (O_1765,N_29256,N_28846);
nor UO_1766 (O_1766,N_29748,N_29681);
nor UO_1767 (O_1767,N_29644,N_27729);
nor UO_1768 (O_1768,N_28028,N_27603);
or UO_1769 (O_1769,N_27728,N_28949);
xor UO_1770 (O_1770,N_29693,N_28947);
or UO_1771 (O_1771,N_29936,N_27232);
or UO_1772 (O_1772,N_28197,N_28611);
and UO_1773 (O_1773,N_28226,N_27378);
or UO_1774 (O_1774,N_29625,N_27954);
nand UO_1775 (O_1775,N_28229,N_27742);
and UO_1776 (O_1776,N_29103,N_27293);
nor UO_1777 (O_1777,N_27294,N_28599);
xnor UO_1778 (O_1778,N_28088,N_27866);
or UO_1779 (O_1779,N_27649,N_28906);
nand UO_1780 (O_1780,N_29328,N_27302);
nor UO_1781 (O_1781,N_27408,N_29687);
nor UO_1782 (O_1782,N_27697,N_28464);
nor UO_1783 (O_1783,N_29087,N_28142);
xor UO_1784 (O_1784,N_28852,N_28500);
nand UO_1785 (O_1785,N_29446,N_29652);
nand UO_1786 (O_1786,N_29980,N_27977);
nor UO_1787 (O_1787,N_29487,N_27208);
nor UO_1788 (O_1788,N_27992,N_29037);
xnor UO_1789 (O_1789,N_29177,N_27685);
nor UO_1790 (O_1790,N_27602,N_27392);
nand UO_1791 (O_1791,N_29451,N_28227);
nand UO_1792 (O_1792,N_27738,N_29068);
xor UO_1793 (O_1793,N_29274,N_29133);
or UO_1794 (O_1794,N_29550,N_29172);
nand UO_1795 (O_1795,N_29167,N_27591);
nor UO_1796 (O_1796,N_28670,N_29741);
and UO_1797 (O_1797,N_29041,N_29279);
nand UO_1798 (O_1798,N_27484,N_29342);
nor UO_1799 (O_1799,N_29342,N_27154);
nor UO_1800 (O_1800,N_29801,N_29673);
or UO_1801 (O_1801,N_27828,N_27240);
nand UO_1802 (O_1802,N_29428,N_29346);
nand UO_1803 (O_1803,N_29009,N_28157);
nor UO_1804 (O_1804,N_29325,N_29179);
or UO_1805 (O_1805,N_28992,N_29600);
nand UO_1806 (O_1806,N_28340,N_27822);
or UO_1807 (O_1807,N_27954,N_27443);
nor UO_1808 (O_1808,N_29121,N_29788);
or UO_1809 (O_1809,N_29461,N_28408);
nor UO_1810 (O_1810,N_29848,N_28509);
or UO_1811 (O_1811,N_27835,N_27970);
xnor UO_1812 (O_1812,N_29004,N_29884);
xor UO_1813 (O_1813,N_28884,N_29363);
or UO_1814 (O_1814,N_28510,N_29618);
xnor UO_1815 (O_1815,N_29747,N_27349);
nor UO_1816 (O_1816,N_27823,N_27548);
nor UO_1817 (O_1817,N_27103,N_27383);
xor UO_1818 (O_1818,N_28183,N_28639);
or UO_1819 (O_1819,N_29090,N_27127);
nand UO_1820 (O_1820,N_28363,N_29075);
nor UO_1821 (O_1821,N_27268,N_27122);
or UO_1822 (O_1822,N_29441,N_27019);
and UO_1823 (O_1823,N_28851,N_28374);
and UO_1824 (O_1824,N_27146,N_27607);
xor UO_1825 (O_1825,N_27583,N_29635);
nor UO_1826 (O_1826,N_27352,N_29003);
or UO_1827 (O_1827,N_27607,N_27891);
or UO_1828 (O_1828,N_27017,N_27870);
or UO_1829 (O_1829,N_29307,N_28054);
or UO_1830 (O_1830,N_28325,N_28420);
nor UO_1831 (O_1831,N_28235,N_28817);
or UO_1832 (O_1832,N_28530,N_27297);
nand UO_1833 (O_1833,N_28370,N_27490);
nor UO_1834 (O_1834,N_29524,N_28802);
xor UO_1835 (O_1835,N_27994,N_29259);
nor UO_1836 (O_1836,N_28375,N_29501);
or UO_1837 (O_1837,N_27496,N_27762);
nand UO_1838 (O_1838,N_28372,N_29225);
xor UO_1839 (O_1839,N_27925,N_29848);
and UO_1840 (O_1840,N_27383,N_27881);
xor UO_1841 (O_1841,N_29127,N_29384);
xnor UO_1842 (O_1842,N_27233,N_28901);
nor UO_1843 (O_1843,N_29153,N_28536);
nand UO_1844 (O_1844,N_28585,N_29765);
and UO_1845 (O_1845,N_27430,N_29635);
nor UO_1846 (O_1846,N_27077,N_27020);
and UO_1847 (O_1847,N_27264,N_27350);
and UO_1848 (O_1848,N_29843,N_27801);
and UO_1849 (O_1849,N_28810,N_28996);
xor UO_1850 (O_1850,N_28136,N_27287);
and UO_1851 (O_1851,N_28694,N_29030);
and UO_1852 (O_1852,N_28330,N_27902);
and UO_1853 (O_1853,N_29460,N_28051);
nor UO_1854 (O_1854,N_28139,N_28150);
nand UO_1855 (O_1855,N_27478,N_29794);
and UO_1856 (O_1856,N_29103,N_28232);
nor UO_1857 (O_1857,N_29726,N_28850);
xnor UO_1858 (O_1858,N_29056,N_27744);
nor UO_1859 (O_1859,N_27923,N_28862);
and UO_1860 (O_1860,N_28812,N_27834);
and UO_1861 (O_1861,N_29128,N_29567);
nor UO_1862 (O_1862,N_27859,N_29567);
xor UO_1863 (O_1863,N_29607,N_29321);
xor UO_1864 (O_1864,N_28874,N_29676);
or UO_1865 (O_1865,N_29158,N_29178);
xnor UO_1866 (O_1866,N_28250,N_29936);
xnor UO_1867 (O_1867,N_29884,N_28222);
or UO_1868 (O_1868,N_29046,N_27411);
xnor UO_1869 (O_1869,N_29986,N_28616);
xnor UO_1870 (O_1870,N_27103,N_27580);
and UO_1871 (O_1871,N_28060,N_29021);
nor UO_1872 (O_1872,N_29935,N_27644);
nand UO_1873 (O_1873,N_28831,N_28430);
or UO_1874 (O_1874,N_28874,N_29344);
nor UO_1875 (O_1875,N_27702,N_27400);
nor UO_1876 (O_1876,N_28139,N_29313);
nor UO_1877 (O_1877,N_29897,N_28224);
nand UO_1878 (O_1878,N_27935,N_28903);
and UO_1879 (O_1879,N_27876,N_27253);
xor UO_1880 (O_1880,N_29185,N_27252);
nor UO_1881 (O_1881,N_27266,N_29689);
xnor UO_1882 (O_1882,N_27015,N_29543);
or UO_1883 (O_1883,N_29549,N_27796);
nand UO_1884 (O_1884,N_29879,N_28354);
nor UO_1885 (O_1885,N_29238,N_28709);
nand UO_1886 (O_1886,N_29184,N_29191);
or UO_1887 (O_1887,N_27505,N_29872);
xnor UO_1888 (O_1888,N_27480,N_29579);
xor UO_1889 (O_1889,N_28666,N_27850);
nor UO_1890 (O_1890,N_28949,N_27799);
or UO_1891 (O_1891,N_28174,N_29783);
nor UO_1892 (O_1892,N_27155,N_29033);
xnor UO_1893 (O_1893,N_27025,N_28633);
nor UO_1894 (O_1894,N_29044,N_28374);
or UO_1895 (O_1895,N_29451,N_27985);
or UO_1896 (O_1896,N_29600,N_28477);
nor UO_1897 (O_1897,N_29517,N_28539);
nor UO_1898 (O_1898,N_29683,N_27394);
xnor UO_1899 (O_1899,N_29871,N_28343);
nor UO_1900 (O_1900,N_28799,N_27447);
or UO_1901 (O_1901,N_27395,N_29696);
or UO_1902 (O_1902,N_29612,N_29535);
xor UO_1903 (O_1903,N_28683,N_27144);
and UO_1904 (O_1904,N_28836,N_29483);
and UO_1905 (O_1905,N_29912,N_28606);
nor UO_1906 (O_1906,N_28776,N_29631);
nand UO_1907 (O_1907,N_27875,N_29844);
nor UO_1908 (O_1908,N_29795,N_27479);
xor UO_1909 (O_1909,N_29114,N_29326);
nand UO_1910 (O_1910,N_28756,N_29276);
nor UO_1911 (O_1911,N_29684,N_29495);
and UO_1912 (O_1912,N_29562,N_29956);
or UO_1913 (O_1913,N_27098,N_28278);
xnor UO_1914 (O_1914,N_29486,N_27024);
nor UO_1915 (O_1915,N_27368,N_27643);
nand UO_1916 (O_1916,N_29481,N_27273);
or UO_1917 (O_1917,N_28470,N_27942);
xnor UO_1918 (O_1918,N_28459,N_29291);
and UO_1919 (O_1919,N_29328,N_28799);
nand UO_1920 (O_1920,N_28126,N_27717);
nor UO_1921 (O_1921,N_27773,N_28652);
and UO_1922 (O_1922,N_28338,N_28436);
xnor UO_1923 (O_1923,N_27174,N_28980);
or UO_1924 (O_1924,N_29780,N_28701);
nor UO_1925 (O_1925,N_28432,N_27264);
xnor UO_1926 (O_1926,N_27212,N_27592);
nor UO_1927 (O_1927,N_29002,N_28266);
or UO_1928 (O_1928,N_28252,N_29961);
xor UO_1929 (O_1929,N_28735,N_28369);
and UO_1930 (O_1930,N_29959,N_29172);
or UO_1931 (O_1931,N_27902,N_27480);
nand UO_1932 (O_1932,N_27086,N_27346);
and UO_1933 (O_1933,N_27457,N_29087);
nand UO_1934 (O_1934,N_27609,N_27246);
nand UO_1935 (O_1935,N_27347,N_29788);
or UO_1936 (O_1936,N_29457,N_27029);
nor UO_1937 (O_1937,N_27106,N_29918);
and UO_1938 (O_1938,N_29218,N_29875);
nor UO_1939 (O_1939,N_29341,N_28406);
xnor UO_1940 (O_1940,N_29836,N_29480);
and UO_1941 (O_1941,N_29793,N_28089);
xnor UO_1942 (O_1942,N_28182,N_29630);
or UO_1943 (O_1943,N_28507,N_29946);
nor UO_1944 (O_1944,N_29104,N_29775);
nand UO_1945 (O_1945,N_29966,N_27503);
xor UO_1946 (O_1946,N_29438,N_28012);
nor UO_1947 (O_1947,N_28847,N_28241);
nand UO_1948 (O_1948,N_28431,N_27218);
or UO_1949 (O_1949,N_27018,N_27105);
nor UO_1950 (O_1950,N_27827,N_29449);
and UO_1951 (O_1951,N_27275,N_29241);
or UO_1952 (O_1952,N_28358,N_28773);
xor UO_1953 (O_1953,N_28788,N_28714);
and UO_1954 (O_1954,N_27732,N_28364);
nor UO_1955 (O_1955,N_27182,N_29413);
or UO_1956 (O_1956,N_28076,N_27532);
nand UO_1957 (O_1957,N_27716,N_28428);
nor UO_1958 (O_1958,N_27343,N_29642);
xnor UO_1959 (O_1959,N_29491,N_29790);
xor UO_1960 (O_1960,N_28562,N_29722);
and UO_1961 (O_1961,N_28905,N_29398);
nor UO_1962 (O_1962,N_28361,N_29261);
and UO_1963 (O_1963,N_28314,N_28136);
xor UO_1964 (O_1964,N_28097,N_28817);
or UO_1965 (O_1965,N_28708,N_28617);
or UO_1966 (O_1966,N_27187,N_27208);
or UO_1967 (O_1967,N_29607,N_28078);
or UO_1968 (O_1968,N_27683,N_28750);
nor UO_1969 (O_1969,N_29236,N_27362);
nand UO_1970 (O_1970,N_28643,N_28401);
xor UO_1971 (O_1971,N_28732,N_28960);
nor UO_1972 (O_1972,N_29051,N_29504);
nand UO_1973 (O_1973,N_28915,N_28742);
and UO_1974 (O_1974,N_28775,N_28708);
xor UO_1975 (O_1975,N_27048,N_27881);
nand UO_1976 (O_1976,N_27542,N_28027);
nor UO_1977 (O_1977,N_28370,N_28589);
and UO_1978 (O_1978,N_29706,N_28452);
xnor UO_1979 (O_1979,N_28576,N_27159);
xnor UO_1980 (O_1980,N_27709,N_29181);
xor UO_1981 (O_1981,N_29452,N_29310);
nor UO_1982 (O_1982,N_29475,N_27825);
xnor UO_1983 (O_1983,N_29351,N_28854);
nand UO_1984 (O_1984,N_27129,N_29984);
nor UO_1985 (O_1985,N_28807,N_27619);
nor UO_1986 (O_1986,N_27640,N_27779);
nand UO_1987 (O_1987,N_27472,N_27653);
or UO_1988 (O_1988,N_28112,N_27778);
nand UO_1989 (O_1989,N_28848,N_28571);
xnor UO_1990 (O_1990,N_27908,N_27098);
or UO_1991 (O_1991,N_27485,N_28627);
xor UO_1992 (O_1992,N_27223,N_28381);
nor UO_1993 (O_1993,N_27016,N_28147);
nor UO_1994 (O_1994,N_27754,N_27598);
and UO_1995 (O_1995,N_29048,N_28160);
or UO_1996 (O_1996,N_27728,N_29591);
and UO_1997 (O_1997,N_28730,N_27151);
nand UO_1998 (O_1998,N_27801,N_29752);
nand UO_1999 (O_1999,N_27961,N_27262);
nor UO_2000 (O_2000,N_29696,N_29885);
xor UO_2001 (O_2001,N_28858,N_28266);
nand UO_2002 (O_2002,N_28605,N_27675);
nor UO_2003 (O_2003,N_29596,N_29842);
or UO_2004 (O_2004,N_29826,N_28057);
and UO_2005 (O_2005,N_27080,N_28569);
and UO_2006 (O_2006,N_27572,N_28549);
and UO_2007 (O_2007,N_29844,N_27218);
xor UO_2008 (O_2008,N_27984,N_27054);
and UO_2009 (O_2009,N_29239,N_27704);
nor UO_2010 (O_2010,N_29635,N_27535);
and UO_2011 (O_2011,N_27095,N_27348);
nor UO_2012 (O_2012,N_29671,N_27557);
and UO_2013 (O_2013,N_29787,N_28422);
nand UO_2014 (O_2014,N_29063,N_27244);
xnor UO_2015 (O_2015,N_27541,N_29794);
or UO_2016 (O_2016,N_29161,N_29183);
nand UO_2017 (O_2017,N_29534,N_27437);
nor UO_2018 (O_2018,N_27748,N_29758);
nand UO_2019 (O_2019,N_27404,N_27558);
nand UO_2020 (O_2020,N_27732,N_29182);
nand UO_2021 (O_2021,N_29075,N_28578);
or UO_2022 (O_2022,N_27253,N_29048);
xnor UO_2023 (O_2023,N_28021,N_29057);
nor UO_2024 (O_2024,N_28187,N_27133);
or UO_2025 (O_2025,N_29667,N_28834);
and UO_2026 (O_2026,N_29059,N_27569);
nand UO_2027 (O_2027,N_29677,N_29243);
nor UO_2028 (O_2028,N_27131,N_27198);
or UO_2029 (O_2029,N_29883,N_28987);
xnor UO_2030 (O_2030,N_27389,N_27638);
nand UO_2031 (O_2031,N_27620,N_29710);
nand UO_2032 (O_2032,N_28617,N_27199);
and UO_2033 (O_2033,N_27185,N_29786);
or UO_2034 (O_2034,N_28450,N_29371);
or UO_2035 (O_2035,N_27865,N_28288);
nor UO_2036 (O_2036,N_29116,N_29563);
and UO_2037 (O_2037,N_29999,N_27376);
and UO_2038 (O_2038,N_27043,N_29799);
and UO_2039 (O_2039,N_29405,N_29941);
and UO_2040 (O_2040,N_28549,N_29793);
nor UO_2041 (O_2041,N_29415,N_29252);
nor UO_2042 (O_2042,N_28110,N_29606);
or UO_2043 (O_2043,N_29327,N_27880);
or UO_2044 (O_2044,N_27876,N_29289);
nor UO_2045 (O_2045,N_29209,N_28557);
xor UO_2046 (O_2046,N_27775,N_28518);
nand UO_2047 (O_2047,N_28610,N_27077);
nor UO_2048 (O_2048,N_28566,N_27823);
nand UO_2049 (O_2049,N_28096,N_29623);
or UO_2050 (O_2050,N_27532,N_27154);
and UO_2051 (O_2051,N_27765,N_27846);
and UO_2052 (O_2052,N_27627,N_29361);
and UO_2053 (O_2053,N_28443,N_28377);
nor UO_2054 (O_2054,N_27905,N_28366);
nor UO_2055 (O_2055,N_29982,N_27857);
nor UO_2056 (O_2056,N_27160,N_29696);
or UO_2057 (O_2057,N_28313,N_29667);
or UO_2058 (O_2058,N_28745,N_28990);
and UO_2059 (O_2059,N_29336,N_29782);
or UO_2060 (O_2060,N_28177,N_28278);
and UO_2061 (O_2061,N_28549,N_27310);
nor UO_2062 (O_2062,N_27032,N_29498);
and UO_2063 (O_2063,N_28592,N_28977);
or UO_2064 (O_2064,N_29606,N_27951);
xor UO_2065 (O_2065,N_29495,N_29574);
nor UO_2066 (O_2066,N_27811,N_29449);
and UO_2067 (O_2067,N_27323,N_29025);
nor UO_2068 (O_2068,N_28765,N_29843);
and UO_2069 (O_2069,N_28289,N_28735);
nor UO_2070 (O_2070,N_27227,N_28869);
nor UO_2071 (O_2071,N_29808,N_29829);
nand UO_2072 (O_2072,N_29284,N_28330);
or UO_2073 (O_2073,N_28461,N_27063);
and UO_2074 (O_2074,N_29549,N_28428);
and UO_2075 (O_2075,N_28766,N_28702);
and UO_2076 (O_2076,N_28371,N_29848);
or UO_2077 (O_2077,N_29566,N_29772);
xor UO_2078 (O_2078,N_27744,N_29452);
xor UO_2079 (O_2079,N_27461,N_28362);
or UO_2080 (O_2080,N_28155,N_29378);
and UO_2081 (O_2081,N_27881,N_28929);
xnor UO_2082 (O_2082,N_29526,N_29504);
and UO_2083 (O_2083,N_28460,N_28113);
or UO_2084 (O_2084,N_27046,N_27017);
and UO_2085 (O_2085,N_27430,N_28053);
nand UO_2086 (O_2086,N_28617,N_29428);
or UO_2087 (O_2087,N_27274,N_27486);
or UO_2088 (O_2088,N_27885,N_29674);
or UO_2089 (O_2089,N_29379,N_29482);
or UO_2090 (O_2090,N_27310,N_29607);
nor UO_2091 (O_2091,N_29507,N_28940);
xor UO_2092 (O_2092,N_29679,N_29689);
xnor UO_2093 (O_2093,N_29039,N_28887);
or UO_2094 (O_2094,N_29982,N_28789);
nand UO_2095 (O_2095,N_28691,N_29154);
nor UO_2096 (O_2096,N_28238,N_28315);
xor UO_2097 (O_2097,N_29556,N_28157);
or UO_2098 (O_2098,N_27388,N_29989);
xnor UO_2099 (O_2099,N_27947,N_27544);
or UO_2100 (O_2100,N_27789,N_27849);
nor UO_2101 (O_2101,N_27073,N_27501);
nand UO_2102 (O_2102,N_29710,N_28289);
nand UO_2103 (O_2103,N_28048,N_28724);
xnor UO_2104 (O_2104,N_29608,N_28997);
xnor UO_2105 (O_2105,N_28587,N_28219);
nand UO_2106 (O_2106,N_29077,N_28953);
xor UO_2107 (O_2107,N_28142,N_27844);
or UO_2108 (O_2108,N_27941,N_28970);
or UO_2109 (O_2109,N_28294,N_29498);
nor UO_2110 (O_2110,N_29455,N_29128);
and UO_2111 (O_2111,N_29325,N_27813);
or UO_2112 (O_2112,N_28390,N_29884);
or UO_2113 (O_2113,N_29979,N_27912);
or UO_2114 (O_2114,N_28878,N_29886);
xnor UO_2115 (O_2115,N_27283,N_29536);
or UO_2116 (O_2116,N_27892,N_29496);
xor UO_2117 (O_2117,N_29376,N_28002);
xor UO_2118 (O_2118,N_27717,N_27318);
or UO_2119 (O_2119,N_29313,N_29806);
xor UO_2120 (O_2120,N_27199,N_29140);
nor UO_2121 (O_2121,N_27403,N_29573);
nor UO_2122 (O_2122,N_28429,N_28851);
xor UO_2123 (O_2123,N_29749,N_29425);
nand UO_2124 (O_2124,N_29068,N_27029);
or UO_2125 (O_2125,N_29814,N_27328);
and UO_2126 (O_2126,N_27209,N_29062);
xor UO_2127 (O_2127,N_29906,N_28308);
and UO_2128 (O_2128,N_28770,N_27286);
and UO_2129 (O_2129,N_27173,N_27693);
and UO_2130 (O_2130,N_29770,N_27090);
and UO_2131 (O_2131,N_28845,N_28822);
nor UO_2132 (O_2132,N_28599,N_29996);
xnor UO_2133 (O_2133,N_28975,N_27413);
xor UO_2134 (O_2134,N_29628,N_28320);
nand UO_2135 (O_2135,N_28985,N_29683);
xor UO_2136 (O_2136,N_28521,N_27466);
or UO_2137 (O_2137,N_27930,N_27536);
and UO_2138 (O_2138,N_28217,N_29298);
nand UO_2139 (O_2139,N_29759,N_28213);
nor UO_2140 (O_2140,N_28961,N_28211);
nand UO_2141 (O_2141,N_28000,N_28707);
xor UO_2142 (O_2142,N_27576,N_27574);
nand UO_2143 (O_2143,N_29444,N_29552);
or UO_2144 (O_2144,N_27647,N_27978);
xnor UO_2145 (O_2145,N_29460,N_28856);
nor UO_2146 (O_2146,N_28805,N_28495);
nor UO_2147 (O_2147,N_28727,N_29633);
and UO_2148 (O_2148,N_28880,N_28173);
xor UO_2149 (O_2149,N_28539,N_29134);
xnor UO_2150 (O_2150,N_29446,N_29003);
nor UO_2151 (O_2151,N_27164,N_28074);
or UO_2152 (O_2152,N_27979,N_29783);
nor UO_2153 (O_2153,N_27562,N_29307);
xnor UO_2154 (O_2154,N_29918,N_29704);
or UO_2155 (O_2155,N_28721,N_27629);
nor UO_2156 (O_2156,N_28198,N_29955);
xnor UO_2157 (O_2157,N_29973,N_29888);
nor UO_2158 (O_2158,N_29024,N_29334);
or UO_2159 (O_2159,N_29269,N_27429);
and UO_2160 (O_2160,N_29162,N_29347);
nand UO_2161 (O_2161,N_27282,N_27693);
or UO_2162 (O_2162,N_28318,N_27477);
xnor UO_2163 (O_2163,N_28509,N_27006);
nor UO_2164 (O_2164,N_27079,N_29208);
nor UO_2165 (O_2165,N_28450,N_28676);
nor UO_2166 (O_2166,N_28307,N_28201);
nand UO_2167 (O_2167,N_29442,N_29112);
and UO_2168 (O_2168,N_27378,N_27889);
and UO_2169 (O_2169,N_27447,N_29270);
nand UO_2170 (O_2170,N_28619,N_27151);
or UO_2171 (O_2171,N_29705,N_29881);
and UO_2172 (O_2172,N_28338,N_27529);
and UO_2173 (O_2173,N_28075,N_28296);
xnor UO_2174 (O_2174,N_27451,N_28434);
or UO_2175 (O_2175,N_29013,N_28989);
nand UO_2176 (O_2176,N_27651,N_29696);
or UO_2177 (O_2177,N_28317,N_27860);
or UO_2178 (O_2178,N_28224,N_29365);
and UO_2179 (O_2179,N_27285,N_27360);
or UO_2180 (O_2180,N_27144,N_29229);
nor UO_2181 (O_2181,N_27878,N_29114);
and UO_2182 (O_2182,N_27621,N_27544);
or UO_2183 (O_2183,N_28721,N_29584);
and UO_2184 (O_2184,N_27324,N_28050);
and UO_2185 (O_2185,N_29272,N_29413);
xor UO_2186 (O_2186,N_28343,N_27348);
or UO_2187 (O_2187,N_29274,N_29458);
xnor UO_2188 (O_2188,N_27184,N_29103);
or UO_2189 (O_2189,N_27115,N_28719);
nor UO_2190 (O_2190,N_27895,N_27984);
nand UO_2191 (O_2191,N_28144,N_27590);
and UO_2192 (O_2192,N_27907,N_27417);
nand UO_2193 (O_2193,N_29061,N_28463);
or UO_2194 (O_2194,N_28085,N_29381);
nor UO_2195 (O_2195,N_28484,N_27571);
or UO_2196 (O_2196,N_28548,N_29867);
nor UO_2197 (O_2197,N_27383,N_28799);
and UO_2198 (O_2198,N_27056,N_29044);
xor UO_2199 (O_2199,N_29423,N_29847);
nor UO_2200 (O_2200,N_27442,N_27508);
and UO_2201 (O_2201,N_29184,N_29832);
xor UO_2202 (O_2202,N_28421,N_28447);
or UO_2203 (O_2203,N_29852,N_28119);
nand UO_2204 (O_2204,N_27283,N_27965);
nor UO_2205 (O_2205,N_29932,N_27928);
and UO_2206 (O_2206,N_27059,N_27101);
xnor UO_2207 (O_2207,N_28061,N_28523);
nor UO_2208 (O_2208,N_29807,N_29383);
or UO_2209 (O_2209,N_28316,N_29071);
nand UO_2210 (O_2210,N_28498,N_27875);
xor UO_2211 (O_2211,N_29010,N_27810);
nand UO_2212 (O_2212,N_28004,N_29915);
or UO_2213 (O_2213,N_28464,N_29564);
nand UO_2214 (O_2214,N_28366,N_27269);
nand UO_2215 (O_2215,N_27026,N_27768);
nand UO_2216 (O_2216,N_27107,N_28536);
nand UO_2217 (O_2217,N_29683,N_29328);
or UO_2218 (O_2218,N_29741,N_28462);
nand UO_2219 (O_2219,N_29552,N_28367);
xor UO_2220 (O_2220,N_28216,N_27948);
nor UO_2221 (O_2221,N_27764,N_27636);
or UO_2222 (O_2222,N_29201,N_28895);
nor UO_2223 (O_2223,N_27688,N_28013);
or UO_2224 (O_2224,N_27794,N_29639);
nand UO_2225 (O_2225,N_29789,N_29285);
or UO_2226 (O_2226,N_29211,N_28606);
nor UO_2227 (O_2227,N_28856,N_28310);
or UO_2228 (O_2228,N_28818,N_28465);
nor UO_2229 (O_2229,N_29453,N_27130);
nand UO_2230 (O_2230,N_29154,N_29723);
and UO_2231 (O_2231,N_28935,N_27675);
nand UO_2232 (O_2232,N_29476,N_27848);
and UO_2233 (O_2233,N_29824,N_29993);
or UO_2234 (O_2234,N_27641,N_29733);
nor UO_2235 (O_2235,N_29480,N_29238);
nand UO_2236 (O_2236,N_27040,N_28307);
and UO_2237 (O_2237,N_27125,N_29444);
nand UO_2238 (O_2238,N_27648,N_29168);
xor UO_2239 (O_2239,N_29607,N_27108);
nor UO_2240 (O_2240,N_28861,N_29757);
nor UO_2241 (O_2241,N_27946,N_28312);
nor UO_2242 (O_2242,N_28327,N_28524);
xnor UO_2243 (O_2243,N_29807,N_27700);
or UO_2244 (O_2244,N_28426,N_27644);
nor UO_2245 (O_2245,N_29025,N_27043);
and UO_2246 (O_2246,N_27298,N_28581);
nor UO_2247 (O_2247,N_29296,N_27904);
and UO_2248 (O_2248,N_28932,N_29571);
nor UO_2249 (O_2249,N_28925,N_27103);
nand UO_2250 (O_2250,N_27905,N_28725);
nand UO_2251 (O_2251,N_28303,N_27357);
and UO_2252 (O_2252,N_27453,N_29542);
or UO_2253 (O_2253,N_27787,N_28051);
or UO_2254 (O_2254,N_29919,N_28037);
nand UO_2255 (O_2255,N_28116,N_27926);
nor UO_2256 (O_2256,N_27003,N_28867);
nor UO_2257 (O_2257,N_27685,N_28283);
and UO_2258 (O_2258,N_29014,N_29646);
nand UO_2259 (O_2259,N_29216,N_28701);
nand UO_2260 (O_2260,N_27721,N_27655);
or UO_2261 (O_2261,N_29620,N_28355);
and UO_2262 (O_2262,N_29496,N_29142);
nand UO_2263 (O_2263,N_27152,N_27719);
and UO_2264 (O_2264,N_27024,N_28981);
and UO_2265 (O_2265,N_28213,N_28504);
or UO_2266 (O_2266,N_27877,N_28455);
and UO_2267 (O_2267,N_28455,N_28662);
xnor UO_2268 (O_2268,N_27162,N_29846);
nand UO_2269 (O_2269,N_28917,N_29830);
nor UO_2270 (O_2270,N_29515,N_29039);
nor UO_2271 (O_2271,N_29598,N_29691);
nand UO_2272 (O_2272,N_27612,N_29725);
or UO_2273 (O_2273,N_29900,N_29057);
nor UO_2274 (O_2274,N_29297,N_29811);
and UO_2275 (O_2275,N_27821,N_28432);
xnor UO_2276 (O_2276,N_27798,N_27759);
nand UO_2277 (O_2277,N_28245,N_29217);
or UO_2278 (O_2278,N_28308,N_27538);
or UO_2279 (O_2279,N_28955,N_28370);
xor UO_2280 (O_2280,N_28618,N_28693);
xor UO_2281 (O_2281,N_29202,N_27353);
nand UO_2282 (O_2282,N_27546,N_29252);
and UO_2283 (O_2283,N_27144,N_29311);
xor UO_2284 (O_2284,N_29606,N_27562);
and UO_2285 (O_2285,N_27407,N_28291);
xnor UO_2286 (O_2286,N_27494,N_27823);
nand UO_2287 (O_2287,N_28097,N_29411);
xnor UO_2288 (O_2288,N_29860,N_29055);
nor UO_2289 (O_2289,N_28053,N_28619);
and UO_2290 (O_2290,N_28759,N_27681);
nand UO_2291 (O_2291,N_28348,N_29537);
or UO_2292 (O_2292,N_27626,N_29421);
or UO_2293 (O_2293,N_28655,N_29507);
xnor UO_2294 (O_2294,N_27468,N_28504);
xnor UO_2295 (O_2295,N_28463,N_27210);
nand UO_2296 (O_2296,N_29762,N_29887);
nor UO_2297 (O_2297,N_29688,N_27771);
or UO_2298 (O_2298,N_29889,N_29978);
nand UO_2299 (O_2299,N_28342,N_28404);
and UO_2300 (O_2300,N_29066,N_29133);
or UO_2301 (O_2301,N_27107,N_28273);
nand UO_2302 (O_2302,N_29357,N_29982);
and UO_2303 (O_2303,N_29362,N_28612);
nand UO_2304 (O_2304,N_29360,N_27009);
or UO_2305 (O_2305,N_29866,N_29595);
or UO_2306 (O_2306,N_28642,N_28368);
and UO_2307 (O_2307,N_28702,N_27046);
nor UO_2308 (O_2308,N_28504,N_27327);
and UO_2309 (O_2309,N_28973,N_27889);
and UO_2310 (O_2310,N_28188,N_28929);
xor UO_2311 (O_2311,N_29814,N_28186);
and UO_2312 (O_2312,N_27776,N_28768);
nor UO_2313 (O_2313,N_27671,N_28769);
nand UO_2314 (O_2314,N_29205,N_27043);
nand UO_2315 (O_2315,N_29576,N_29396);
or UO_2316 (O_2316,N_27747,N_27560);
nand UO_2317 (O_2317,N_29839,N_29651);
nand UO_2318 (O_2318,N_27977,N_29060);
nor UO_2319 (O_2319,N_27341,N_27636);
nor UO_2320 (O_2320,N_29280,N_28969);
xnor UO_2321 (O_2321,N_27712,N_27356);
nor UO_2322 (O_2322,N_27946,N_29456);
nor UO_2323 (O_2323,N_28524,N_28683);
or UO_2324 (O_2324,N_28473,N_29117);
xnor UO_2325 (O_2325,N_28714,N_29695);
nor UO_2326 (O_2326,N_27326,N_27663);
or UO_2327 (O_2327,N_28369,N_29868);
nor UO_2328 (O_2328,N_27173,N_28682);
or UO_2329 (O_2329,N_27691,N_29297);
nand UO_2330 (O_2330,N_27578,N_28077);
and UO_2331 (O_2331,N_28146,N_28791);
nor UO_2332 (O_2332,N_29015,N_29206);
and UO_2333 (O_2333,N_27863,N_29509);
nand UO_2334 (O_2334,N_28639,N_27181);
nor UO_2335 (O_2335,N_28980,N_29271);
and UO_2336 (O_2336,N_27324,N_28719);
nand UO_2337 (O_2337,N_27364,N_28012);
and UO_2338 (O_2338,N_28223,N_28331);
xor UO_2339 (O_2339,N_29962,N_28366);
xor UO_2340 (O_2340,N_27781,N_27463);
nand UO_2341 (O_2341,N_28270,N_29486);
or UO_2342 (O_2342,N_29992,N_28650);
nand UO_2343 (O_2343,N_28138,N_28831);
or UO_2344 (O_2344,N_27196,N_29945);
and UO_2345 (O_2345,N_29553,N_28498);
nand UO_2346 (O_2346,N_27627,N_29285);
xor UO_2347 (O_2347,N_27245,N_28777);
xnor UO_2348 (O_2348,N_28007,N_27827);
and UO_2349 (O_2349,N_29954,N_27288);
nor UO_2350 (O_2350,N_27592,N_29211);
and UO_2351 (O_2351,N_27320,N_29461);
nor UO_2352 (O_2352,N_29779,N_28867);
xnor UO_2353 (O_2353,N_27033,N_29464);
or UO_2354 (O_2354,N_29558,N_29794);
nand UO_2355 (O_2355,N_28155,N_29467);
nand UO_2356 (O_2356,N_29015,N_28081);
nor UO_2357 (O_2357,N_27406,N_28083);
nand UO_2358 (O_2358,N_28039,N_27937);
nor UO_2359 (O_2359,N_28413,N_28988);
nand UO_2360 (O_2360,N_29612,N_27609);
xnor UO_2361 (O_2361,N_27630,N_29962);
nand UO_2362 (O_2362,N_27210,N_29978);
and UO_2363 (O_2363,N_29809,N_29189);
nor UO_2364 (O_2364,N_29009,N_29718);
xnor UO_2365 (O_2365,N_28022,N_28548);
and UO_2366 (O_2366,N_28492,N_28913);
and UO_2367 (O_2367,N_28867,N_28002);
nor UO_2368 (O_2368,N_27047,N_27874);
and UO_2369 (O_2369,N_27422,N_29690);
xor UO_2370 (O_2370,N_28851,N_27555);
nand UO_2371 (O_2371,N_27462,N_28529);
and UO_2372 (O_2372,N_28681,N_29796);
or UO_2373 (O_2373,N_28980,N_27891);
nand UO_2374 (O_2374,N_29417,N_29409);
nor UO_2375 (O_2375,N_28322,N_27733);
xor UO_2376 (O_2376,N_29834,N_28763);
xnor UO_2377 (O_2377,N_29167,N_27600);
nor UO_2378 (O_2378,N_27645,N_27922);
and UO_2379 (O_2379,N_29423,N_28776);
nand UO_2380 (O_2380,N_27045,N_28736);
or UO_2381 (O_2381,N_27954,N_28353);
nand UO_2382 (O_2382,N_27029,N_28353);
xor UO_2383 (O_2383,N_29325,N_27742);
or UO_2384 (O_2384,N_28142,N_27298);
xnor UO_2385 (O_2385,N_29348,N_28249);
nor UO_2386 (O_2386,N_27172,N_29940);
or UO_2387 (O_2387,N_29309,N_29622);
or UO_2388 (O_2388,N_28966,N_28605);
nor UO_2389 (O_2389,N_28853,N_28698);
nor UO_2390 (O_2390,N_27469,N_28853);
xor UO_2391 (O_2391,N_29960,N_28467);
nand UO_2392 (O_2392,N_29711,N_27556);
xnor UO_2393 (O_2393,N_29145,N_29409);
xor UO_2394 (O_2394,N_27582,N_28273);
xor UO_2395 (O_2395,N_28243,N_27625);
and UO_2396 (O_2396,N_29106,N_28709);
nor UO_2397 (O_2397,N_29691,N_27783);
or UO_2398 (O_2398,N_27431,N_29084);
nor UO_2399 (O_2399,N_28683,N_28937);
nor UO_2400 (O_2400,N_27999,N_28463);
xnor UO_2401 (O_2401,N_28594,N_29594);
nand UO_2402 (O_2402,N_29616,N_27710);
nor UO_2403 (O_2403,N_29776,N_27675);
nand UO_2404 (O_2404,N_28411,N_27583);
and UO_2405 (O_2405,N_28086,N_28483);
nand UO_2406 (O_2406,N_28526,N_27437);
nor UO_2407 (O_2407,N_29877,N_28278);
nand UO_2408 (O_2408,N_29485,N_27541);
nand UO_2409 (O_2409,N_29720,N_27064);
nand UO_2410 (O_2410,N_29965,N_28580);
or UO_2411 (O_2411,N_27560,N_27800);
xor UO_2412 (O_2412,N_29388,N_28574);
or UO_2413 (O_2413,N_27020,N_29080);
nor UO_2414 (O_2414,N_28417,N_27780);
xnor UO_2415 (O_2415,N_27267,N_28764);
xor UO_2416 (O_2416,N_29584,N_27519);
xnor UO_2417 (O_2417,N_28766,N_28360);
or UO_2418 (O_2418,N_28224,N_28701);
or UO_2419 (O_2419,N_29237,N_27373);
and UO_2420 (O_2420,N_27102,N_27114);
nor UO_2421 (O_2421,N_28741,N_27472);
or UO_2422 (O_2422,N_27072,N_29679);
nand UO_2423 (O_2423,N_28595,N_28524);
nor UO_2424 (O_2424,N_28018,N_28784);
nor UO_2425 (O_2425,N_27879,N_29714);
and UO_2426 (O_2426,N_28001,N_27293);
nor UO_2427 (O_2427,N_29506,N_27082);
or UO_2428 (O_2428,N_27066,N_29197);
xor UO_2429 (O_2429,N_28996,N_27327);
xnor UO_2430 (O_2430,N_28749,N_28166);
nor UO_2431 (O_2431,N_28274,N_29336);
nor UO_2432 (O_2432,N_28924,N_28051);
or UO_2433 (O_2433,N_28576,N_27767);
nor UO_2434 (O_2434,N_29197,N_27678);
xor UO_2435 (O_2435,N_27172,N_28261);
nor UO_2436 (O_2436,N_29729,N_28584);
xnor UO_2437 (O_2437,N_27494,N_27219);
xor UO_2438 (O_2438,N_28946,N_28275);
xor UO_2439 (O_2439,N_29574,N_28136);
nor UO_2440 (O_2440,N_28849,N_27569);
xnor UO_2441 (O_2441,N_27851,N_28787);
xor UO_2442 (O_2442,N_29276,N_27435);
or UO_2443 (O_2443,N_27062,N_28074);
or UO_2444 (O_2444,N_27893,N_27563);
nand UO_2445 (O_2445,N_28648,N_29879);
nand UO_2446 (O_2446,N_27179,N_28499);
nor UO_2447 (O_2447,N_28328,N_29704);
nand UO_2448 (O_2448,N_27483,N_29721);
or UO_2449 (O_2449,N_27779,N_28836);
or UO_2450 (O_2450,N_27402,N_27672);
and UO_2451 (O_2451,N_29968,N_29956);
xor UO_2452 (O_2452,N_29327,N_27610);
and UO_2453 (O_2453,N_29307,N_28212);
nor UO_2454 (O_2454,N_29258,N_29809);
nor UO_2455 (O_2455,N_29798,N_29873);
or UO_2456 (O_2456,N_29117,N_29103);
nand UO_2457 (O_2457,N_29547,N_29599);
nor UO_2458 (O_2458,N_28281,N_28384);
nor UO_2459 (O_2459,N_27534,N_28589);
nand UO_2460 (O_2460,N_29824,N_29839);
xnor UO_2461 (O_2461,N_29087,N_27741);
xor UO_2462 (O_2462,N_29808,N_28262);
nor UO_2463 (O_2463,N_29139,N_28889);
or UO_2464 (O_2464,N_27417,N_29864);
nor UO_2465 (O_2465,N_29036,N_27281);
xnor UO_2466 (O_2466,N_29175,N_29301);
nor UO_2467 (O_2467,N_27885,N_29841);
nor UO_2468 (O_2468,N_29057,N_28494);
xor UO_2469 (O_2469,N_27265,N_27671);
and UO_2470 (O_2470,N_29668,N_29135);
and UO_2471 (O_2471,N_27080,N_29380);
or UO_2472 (O_2472,N_29792,N_28351);
nor UO_2473 (O_2473,N_29223,N_29278);
and UO_2474 (O_2474,N_27553,N_29579);
and UO_2475 (O_2475,N_29998,N_27741);
nor UO_2476 (O_2476,N_28419,N_29706);
and UO_2477 (O_2477,N_28448,N_27875);
nand UO_2478 (O_2478,N_29106,N_29559);
nand UO_2479 (O_2479,N_27317,N_27772);
nand UO_2480 (O_2480,N_27183,N_29792);
nor UO_2481 (O_2481,N_29926,N_27182);
nor UO_2482 (O_2482,N_29129,N_29352);
nor UO_2483 (O_2483,N_29707,N_29480);
xnor UO_2484 (O_2484,N_29976,N_28904);
nor UO_2485 (O_2485,N_28771,N_28536);
nor UO_2486 (O_2486,N_29824,N_29246);
xor UO_2487 (O_2487,N_28395,N_29383);
or UO_2488 (O_2488,N_27398,N_29445);
nand UO_2489 (O_2489,N_27829,N_28593);
and UO_2490 (O_2490,N_27225,N_27478);
nand UO_2491 (O_2491,N_29060,N_28794);
nor UO_2492 (O_2492,N_28569,N_27488);
nor UO_2493 (O_2493,N_29382,N_27708);
and UO_2494 (O_2494,N_29434,N_28369);
xnor UO_2495 (O_2495,N_27495,N_29489);
xnor UO_2496 (O_2496,N_28087,N_27334);
nor UO_2497 (O_2497,N_27684,N_29204);
nand UO_2498 (O_2498,N_27968,N_27911);
nor UO_2499 (O_2499,N_27687,N_29369);
nand UO_2500 (O_2500,N_29110,N_29851);
and UO_2501 (O_2501,N_28623,N_29083);
nand UO_2502 (O_2502,N_29796,N_27374);
nor UO_2503 (O_2503,N_27171,N_28834);
nand UO_2504 (O_2504,N_27948,N_29362);
nand UO_2505 (O_2505,N_27898,N_27428);
xnor UO_2506 (O_2506,N_29282,N_28692);
nor UO_2507 (O_2507,N_27989,N_29343);
xnor UO_2508 (O_2508,N_27921,N_28820);
or UO_2509 (O_2509,N_27332,N_29306);
nor UO_2510 (O_2510,N_29034,N_28587);
and UO_2511 (O_2511,N_27519,N_27279);
or UO_2512 (O_2512,N_29537,N_28123);
or UO_2513 (O_2513,N_28819,N_29279);
or UO_2514 (O_2514,N_27123,N_28686);
or UO_2515 (O_2515,N_29750,N_28649);
nor UO_2516 (O_2516,N_29396,N_28522);
nand UO_2517 (O_2517,N_29019,N_27554);
xor UO_2518 (O_2518,N_28874,N_28135);
nand UO_2519 (O_2519,N_28004,N_28744);
and UO_2520 (O_2520,N_28082,N_28779);
and UO_2521 (O_2521,N_27462,N_27745);
and UO_2522 (O_2522,N_28214,N_28269);
xor UO_2523 (O_2523,N_28921,N_27062);
or UO_2524 (O_2524,N_29325,N_27610);
or UO_2525 (O_2525,N_27569,N_27380);
or UO_2526 (O_2526,N_27004,N_28287);
or UO_2527 (O_2527,N_29752,N_29713);
nor UO_2528 (O_2528,N_28108,N_29958);
nor UO_2529 (O_2529,N_29659,N_29466);
nand UO_2530 (O_2530,N_29662,N_28605);
nand UO_2531 (O_2531,N_28120,N_27990);
and UO_2532 (O_2532,N_28699,N_28420);
xor UO_2533 (O_2533,N_27114,N_28400);
or UO_2534 (O_2534,N_28160,N_27032);
xnor UO_2535 (O_2535,N_29232,N_28931);
nor UO_2536 (O_2536,N_29212,N_28973);
nand UO_2537 (O_2537,N_28674,N_28654);
or UO_2538 (O_2538,N_27569,N_28893);
xor UO_2539 (O_2539,N_29286,N_27273);
xor UO_2540 (O_2540,N_29514,N_27865);
nand UO_2541 (O_2541,N_29698,N_27866);
xnor UO_2542 (O_2542,N_28993,N_29173);
xor UO_2543 (O_2543,N_27987,N_28621);
or UO_2544 (O_2544,N_28138,N_27059);
nand UO_2545 (O_2545,N_28700,N_28562);
nor UO_2546 (O_2546,N_28713,N_27223);
nor UO_2547 (O_2547,N_27739,N_28365);
xnor UO_2548 (O_2548,N_27293,N_29407);
or UO_2549 (O_2549,N_29531,N_27345);
xnor UO_2550 (O_2550,N_28506,N_27827);
nor UO_2551 (O_2551,N_29320,N_27277);
nand UO_2552 (O_2552,N_29663,N_29256);
xor UO_2553 (O_2553,N_27493,N_29825);
and UO_2554 (O_2554,N_27847,N_28782);
and UO_2555 (O_2555,N_27688,N_29527);
and UO_2556 (O_2556,N_29467,N_28837);
xor UO_2557 (O_2557,N_27361,N_29119);
and UO_2558 (O_2558,N_28990,N_27351);
and UO_2559 (O_2559,N_28218,N_27742);
nand UO_2560 (O_2560,N_27046,N_29887);
or UO_2561 (O_2561,N_29421,N_27947);
or UO_2562 (O_2562,N_29568,N_29529);
nand UO_2563 (O_2563,N_28215,N_28769);
xor UO_2564 (O_2564,N_27372,N_28292);
or UO_2565 (O_2565,N_29604,N_28914);
nor UO_2566 (O_2566,N_28353,N_27194);
and UO_2567 (O_2567,N_29085,N_28386);
and UO_2568 (O_2568,N_29126,N_28299);
and UO_2569 (O_2569,N_28765,N_28048);
nand UO_2570 (O_2570,N_27000,N_29437);
and UO_2571 (O_2571,N_27720,N_27683);
nor UO_2572 (O_2572,N_28999,N_27185);
nor UO_2573 (O_2573,N_29022,N_28179);
xnor UO_2574 (O_2574,N_27431,N_29736);
xor UO_2575 (O_2575,N_28083,N_29139);
nor UO_2576 (O_2576,N_27731,N_29377);
and UO_2577 (O_2577,N_28440,N_27526);
nand UO_2578 (O_2578,N_28310,N_28831);
nand UO_2579 (O_2579,N_28421,N_29235);
or UO_2580 (O_2580,N_29143,N_29219);
xnor UO_2581 (O_2581,N_27897,N_28628);
and UO_2582 (O_2582,N_27439,N_28749);
or UO_2583 (O_2583,N_28743,N_28275);
xnor UO_2584 (O_2584,N_28171,N_28164);
nand UO_2585 (O_2585,N_27788,N_27389);
nand UO_2586 (O_2586,N_27334,N_29923);
and UO_2587 (O_2587,N_27090,N_27918);
nor UO_2588 (O_2588,N_28631,N_29613);
xnor UO_2589 (O_2589,N_28757,N_27190);
nand UO_2590 (O_2590,N_27921,N_29741);
xor UO_2591 (O_2591,N_29701,N_29062);
or UO_2592 (O_2592,N_27227,N_28426);
nor UO_2593 (O_2593,N_27374,N_29820);
nor UO_2594 (O_2594,N_28914,N_27124);
or UO_2595 (O_2595,N_28285,N_27687);
or UO_2596 (O_2596,N_28177,N_29133);
or UO_2597 (O_2597,N_28808,N_29360);
xnor UO_2598 (O_2598,N_27389,N_29168);
and UO_2599 (O_2599,N_29033,N_27100);
nand UO_2600 (O_2600,N_29010,N_28658);
or UO_2601 (O_2601,N_27036,N_29903);
or UO_2602 (O_2602,N_27821,N_29582);
nor UO_2603 (O_2603,N_28721,N_28706);
xnor UO_2604 (O_2604,N_27891,N_28730);
and UO_2605 (O_2605,N_29513,N_28827);
and UO_2606 (O_2606,N_28790,N_29946);
xnor UO_2607 (O_2607,N_28481,N_28589);
nor UO_2608 (O_2608,N_28319,N_27606);
xnor UO_2609 (O_2609,N_27743,N_29929);
or UO_2610 (O_2610,N_28570,N_27867);
nand UO_2611 (O_2611,N_27421,N_28231);
nor UO_2612 (O_2612,N_28716,N_29919);
and UO_2613 (O_2613,N_28793,N_28031);
nand UO_2614 (O_2614,N_29589,N_28733);
nor UO_2615 (O_2615,N_29359,N_28937);
xor UO_2616 (O_2616,N_29970,N_29698);
and UO_2617 (O_2617,N_27273,N_27561);
and UO_2618 (O_2618,N_29089,N_28356);
xor UO_2619 (O_2619,N_28203,N_27894);
nor UO_2620 (O_2620,N_28069,N_29408);
nor UO_2621 (O_2621,N_29858,N_29098);
nor UO_2622 (O_2622,N_28056,N_29444);
or UO_2623 (O_2623,N_27478,N_27130);
or UO_2624 (O_2624,N_29133,N_28172);
xnor UO_2625 (O_2625,N_28827,N_28760);
and UO_2626 (O_2626,N_27797,N_29151);
nor UO_2627 (O_2627,N_28911,N_29142);
nand UO_2628 (O_2628,N_28058,N_28356);
and UO_2629 (O_2629,N_29534,N_27362);
xor UO_2630 (O_2630,N_29388,N_27573);
and UO_2631 (O_2631,N_27822,N_27478);
nand UO_2632 (O_2632,N_28661,N_29718);
or UO_2633 (O_2633,N_28847,N_28917);
nand UO_2634 (O_2634,N_27445,N_27626);
nor UO_2635 (O_2635,N_29928,N_27591);
or UO_2636 (O_2636,N_27316,N_29501);
nand UO_2637 (O_2637,N_27778,N_27035);
nor UO_2638 (O_2638,N_27060,N_28098);
xor UO_2639 (O_2639,N_28813,N_27666);
nand UO_2640 (O_2640,N_27692,N_27627);
or UO_2641 (O_2641,N_28572,N_29804);
xnor UO_2642 (O_2642,N_27152,N_28262);
and UO_2643 (O_2643,N_28004,N_27437);
nor UO_2644 (O_2644,N_29121,N_27537);
xor UO_2645 (O_2645,N_29865,N_29489);
and UO_2646 (O_2646,N_29296,N_29692);
and UO_2647 (O_2647,N_28653,N_29294);
nor UO_2648 (O_2648,N_28203,N_27616);
xor UO_2649 (O_2649,N_27466,N_27752);
or UO_2650 (O_2650,N_27469,N_29946);
nor UO_2651 (O_2651,N_29727,N_27076);
nor UO_2652 (O_2652,N_28949,N_27134);
or UO_2653 (O_2653,N_27685,N_27849);
nor UO_2654 (O_2654,N_29422,N_27638);
and UO_2655 (O_2655,N_29801,N_27497);
nand UO_2656 (O_2656,N_28718,N_29457);
or UO_2657 (O_2657,N_27077,N_29999);
nor UO_2658 (O_2658,N_28449,N_28633);
or UO_2659 (O_2659,N_29549,N_27102);
nor UO_2660 (O_2660,N_28165,N_28046);
and UO_2661 (O_2661,N_27199,N_29985);
and UO_2662 (O_2662,N_28139,N_28928);
nor UO_2663 (O_2663,N_27318,N_29083);
or UO_2664 (O_2664,N_29340,N_29862);
and UO_2665 (O_2665,N_29218,N_28517);
xnor UO_2666 (O_2666,N_27687,N_29422);
nor UO_2667 (O_2667,N_29636,N_29039);
xnor UO_2668 (O_2668,N_29107,N_29357);
xnor UO_2669 (O_2669,N_27018,N_29377);
xnor UO_2670 (O_2670,N_29437,N_27073);
nand UO_2671 (O_2671,N_27876,N_27274);
xor UO_2672 (O_2672,N_28366,N_29003);
and UO_2673 (O_2673,N_27730,N_28981);
xor UO_2674 (O_2674,N_29860,N_28164);
nand UO_2675 (O_2675,N_29485,N_27469);
xnor UO_2676 (O_2676,N_29410,N_29997);
nor UO_2677 (O_2677,N_28086,N_27904);
xor UO_2678 (O_2678,N_28784,N_27307);
nor UO_2679 (O_2679,N_29299,N_29417);
nor UO_2680 (O_2680,N_27621,N_27699);
nand UO_2681 (O_2681,N_27048,N_28467);
nand UO_2682 (O_2682,N_29553,N_29338);
xnor UO_2683 (O_2683,N_29727,N_28840);
nand UO_2684 (O_2684,N_27857,N_27730);
and UO_2685 (O_2685,N_27001,N_27501);
nand UO_2686 (O_2686,N_28875,N_27026);
nor UO_2687 (O_2687,N_28959,N_29610);
nor UO_2688 (O_2688,N_29736,N_28221);
or UO_2689 (O_2689,N_27036,N_29787);
nand UO_2690 (O_2690,N_29293,N_27965);
nand UO_2691 (O_2691,N_28068,N_27924);
nand UO_2692 (O_2692,N_27083,N_27455);
nor UO_2693 (O_2693,N_28894,N_27505);
or UO_2694 (O_2694,N_29434,N_27529);
nand UO_2695 (O_2695,N_28906,N_28786);
xnor UO_2696 (O_2696,N_27949,N_28788);
xor UO_2697 (O_2697,N_29529,N_27868);
or UO_2698 (O_2698,N_29191,N_27877);
nor UO_2699 (O_2699,N_27266,N_27651);
nor UO_2700 (O_2700,N_29134,N_28004);
nor UO_2701 (O_2701,N_28417,N_29273);
nand UO_2702 (O_2702,N_27355,N_28441);
nor UO_2703 (O_2703,N_27317,N_27570);
xor UO_2704 (O_2704,N_27191,N_29995);
nor UO_2705 (O_2705,N_29763,N_29411);
nand UO_2706 (O_2706,N_27393,N_28829);
xnor UO_2707 (O_2707,N_27765,N_27604);
nor UO_2708 (O_2708,N_28103,N_28456);
and UO_2709 (O_2709,N_28174,N_28270);
nor UO_2710 (O_2710,N_29861,N_28496);
xor UO_2711 (O_2711,N_28588,N_28318);
nor UO_2712 (O_2712,N_29436,N_27589);
and UO_2713 (O_2713,N_28118,N_27103);
nor UO_2714 (O_2714,N_28753,N_28963);
nor UO_2715 (O_2715,N_28739,N_27176);
nor UO_2716 (O_2716,N_28383,N_28670);
or UO_2717 (O_2717,N_28461,N_27442);
or UO_2718 (O_2718,N_27075,N_29550);
xor UO_2719 (O_2719,N_28959,N_29611);
nor UO_2720 (O_2720,N_28070,N_28135);
xnor UO_2721 (O_2721,N_27175,N_29382);
and UO_2722 (O_2722,N_29916,N_27839);
nand UO_2723 (O_2723,N_27983,N_28001);
and UO_2724 (O_2724,N_27787,N_27347);
and UO_2725 (O_2725,N_28362,N_29271);
and UO_2726 (O_2726,N_29791,N_29093);
and UO_2727 (O_2727,N_27301,N_29285);
nand UO_2728 (O_2728,N_29718,N_27325);
or UO_2729 (O_2729,N_28913,N_27492);
nand UO_2730 (O_2730,N_27443,N_28680);
or UO_2731 (O_2731,N_28351,N_29557);
or UO_2732 (O_2732,N_27331,N_29630);
nand UO_2733 (O_2733,N_29988,N_27809);
and UO_2734 (O_2734,N_29388,N_29733);
and UO_2735 (O_2735,N_28440,N_29891);
or UO_2736 (O_2736,N_29563,N_27834);
nor UO_2737 (O_2737,N_28468,N_27858);
nand UO_2738 (O_2738,N_28254,N_29945);
or UO_2739 (O_2739,N_27179,N_28703);
xor UO_2740 (O_2740,N_28109,N_28398);
and UO_2741 (O_2741,N_29720,N_27768);
nor UO_2742 (O_2742,N_29267,N_27053);
or UO_2743 (O_2743,N_28023,N_27212);
or UO_2744 (O_2744,N_28555,N_29496);
or UO_2745 (O_2745,N_29415,N_28400);
and UO_2746 (O_2746,N_29797,N_27814);
nor UO_2747 (O_2747,N_28900,N_28164);
xor UO_2748 (O_2748,N_29553,N_27443);
xnor UO_2749 (O_2749,N_29772,N_28125);
nor UO_2750 (O_2750,N_28461,N_27334);
and UO_2751 (O_2751,N_29585,N_28360);
nor UO_2752 (O_2752,N_27638,N_27092);
nand UO_2753 (O_2753,N_29427,N_28207);
or UO_2754 (O_2754,N_28362,N_27044);
nor UO_2755 (O_2755,N_28316,N_28996);
or UO_2756 (O_2756,N_27249,N_29786);
nand UO_2757 (O_2757,N_29764,N_28940);
nand UO_2758 (O_2758,N_29185,N_29073);
nor UO_2759 (O_2759,N_28777,N_28904);
nor UO_2760 (O_2760,N_28797,N_27514);
and UO_2761 (O_2761,N_28190,N_28009);
xor UO_2762 (O_2762,N_28976,N_28453);
and UO_2763 (O_2763,N_27210,N_29796);
xor UO_2764 (O_2764,N_29455,N_29048);
xnor UO_2765 (O_2765,N_28418,N_28531);
and UO_2766 (O_2766,N_28154,N_27204);
and UO_2767 (O_2767,N_28253,N_29962);
or UO_2768 (O_2768,N_29923,N_27094);
and UO_2769 (O_2769,N_28556,N_29006);
nor UO_2770 (O_2770,N_27653,N_29770);
nand UO_2771 (O_2771,N_29464,N_29366);
or UO_2772 (O_2772,N_28602,N_28838);
or UO_2773 (O_2773,N_28973,N_28191);
or UO_2774 (O_2774,N_27214,N_28617);
or UO_2775 (O_2775,N_29514,N_29665);
xnor UO_2776 (O_2776,N_29569,N_28118);
and UO_2777 (O_2777,N_27556,N_28636);
nor UO_2778 (O_2778,N_27939,N_28425);
xnor UO_2779 (O_2779,N_27227,N_29075);
nand UO_2780 (O_2780,N_27284,N_27956);
nor UO_2781 (O_2781,N_29831,N_28725);
xor UO_2782 (O_2782,N_29327,N_28758);
or UO_2783 (O_2783,N_27583,N_28668);
and UO_2784 (O_2784,N_28795,N_29130);
or UO_2785 (O_2785,N_28567,N_28712);
and UO_2786 (O_2786,N_28344,N_27797);
and UO_2787 (O_2787,N_27646,N_28303);
xnor UO_2788 (O_2788,N_28466,N_29287);
nor UO_2789 (O_2789,N_27791,N_28439);
or UO_2790 (O_2790,N_29728,N_29924);
nand UO_2791 (O_2791,N_27887,N_28514);
or UO_2792 (O_2792,N_27188,N_27495);
xnor UO_2793 (O_2793,N_28417,N_29990);
nand UO_2794 (O_2794,N_27277,N_28827);
nand UO_2795 (O_2795,N_28857,N_29026);
or UO_2796 (O_2796,N_27059,N_28188);
nor UO_2797 (O_2797,N_27363,N_28793);
nor UO_2798 (O_2798,N_28871,N_28785);
xnor UO_2799 (O_2799,N_27940,N_27608);
and UO_2800 (O_2800,N_27985,N_27069);
nor UO_2801 (O_2801,N_28873,N_29719);
nor UO_2802 (O_2802,N_28102,N_28918);
nor UO_2803 (O_2803,N_29429,N_29447);
or UO_2804 (O_2804,N_28959,N_27388);
or UO_2805 (O_2805,N_27708,N_27372);
nand UO_2806 (O_2806,N_27417,N_27213);
or UO_2807 (O_2807,N_29547,N_27098);
nor UO_2808 (O_2808,N_29642,N_29934);
nand UO_2809 (O_2809,N_28960,N_27391);
and UO_2810 (O_2810,N_28802,N_28253);
nand UO_2811 (O_2811,N_28962,N_27486);
xnor UO_2812 (O_2812,N_27758,N_27409);
or UO_2813 (O_2813,N_28445,N_27997);
and UO_2814 (O_2814,N_29967,N_27655);
or UO_2815 (O_2815,N_28715,N_28568);
nor UO_2816 (O_2816,N_29192,N_27759);
and UO_2817 (O_2817,N_28523,N_29107);
and UO_2818 (O_2818,N_29041,N_28329);
or UO_2819 (O_2819,N_29156,N_27068);
nor UO_2820 (O_2820,N_27461,N_29011);
nand UO_2821 (O_2821,N_29924,N_28275);
nand UO_2822 (O_2822,N_28950,N_27587);
nand UO_2823 (O_2823,N_28305,N_27815);
and UO_2824 (O_2824,N_29819,N_27048);
nand UO_2825 (O_2825,N_29420,N_28840);
or UO_2826 (O_2826,N_28669,N_29764);
nand UO_2827 (O_2827,N_28076,N_29353);
xnor UO_2828 (O_2828,N_28710,N_29227);
or UO_2829 (O_2829,N_28650,N_27706);
nor UO_2830 (O_2830,N_29496,N_27456);
xnor UO_2831 (O_2831,N_27725,N_27994);
nand UO_2832 (O_2832,N_28871,N_29639);
xor UO_2833 (O_2833,N_29449,N_27453);
xor UO_2834 (O_2834,N_29279,N_29765);
nor UO_2835 (O_2835,N_28297,N_27030);
xnor UO_2836 (O_2836,N_28532,N_27166);
and UO_2837 (O_2837,N_27192,N_27646);
nor UO_2838 (O_2838,N_27046,N_29949);
nand UO_2839 (O_2839,N_27438,N_29176);
nor UO_2840 (O_2840,N_28757,N_28302);
nand UO_2841 (O_2841,N_29282,N_27851);
xor UO_2842 (O_2842,N_29778,N_27401);
or UO_2843 (O_2843,N_27189,N_29154);
nand UO_2844 (O_2844,N_27355,N_27320);
and UO_2845 (O_2845,N_29349,N_27756);
or UO_2846 (O_2846,N_29691,N_28518);
nor UO_2847 (O_2847,N_27695,N_29421);
nor UO_2848 (O_2848,N_27834,N_29349);
nor UO_2849 (O_2849,N_27275,N_29517);
xnor UO_2850 (O_2850,N_29543,N_28199);
xor UO_2851 (O_2851,N_27185,N_28071);
and UO_2852 (O_2852,N_29720,N_29495);
or UO_2853 (O_2853,N_27657,N_27700);
nand UO_2854 (O_2854,N_28335,N_29266);
or UO_2855 (O_2855,N_29043,N_28412);
and UO_2856 (O_2856,N_29933,N_28241);
or UO_2857 (O_2857,N_27158,N_27499);
nor UO_2858 (O_2858,N_29336,N_29969);
nor UO_2859 (O_2859,N_28539,N_27497);
nand UO_2860 (O_2860,N_29007,N_28413);
or UO_2861 (O_2861,N_27309,N_27751);
and UO_2862 (O_2862,N_28936,N_29322);
nor UO_2863 (O_2863,N_28079,N_28119);
nand UO_2864 (O_2864,N_28589,N_27554);
xor UO_2865 (O_2865,N_28077,N_28460);
xnor UO_2866 (O_2866,N_29626,N_27579);
and UO_2867 (O_2867,N_28262,N_29889);
or UO_2868 (O_2868,N_28412,N_28990);
nand UO_2869 (O_2869,N_29165,N_27179);
nor UO_2870 (O_2870,N_29721,N_29768);
xnor UO_2871 (O_2871,N_27022,N_29274);
or UO_2872 (O_2872,N_28898,N_27633);
and UO_2873 (O_2873,N_27837,N_28979);
and UO_2874 (O_2874,N_28261,N_27105);
nand UO_2875 (O_2875,N_27148,N_28779);
nor UO_2876 (O_2876,N_29160,N_28295);
or UO_2877 (O_2877,N_28724,N_28800);
nand UO_2878 (O_2878,N_29584,N_27291);
nand UO_2879 (O_2879,N_28107,N_27848);
or UO_2880 (O_2880,N_29569,N_27945);
nor UO_2881 (O_2881,N_28994,N_29095);
nand UO_2882 (O_2882,N_27480,N_27074);
xor UO_2883 (O_2883,N_28042,N_28678);
nand UO_2884 (O_2884,N_29634,N_28326);
nand UO_2885 (O_2885,N_28340,N_27268);
xor UO_2886 (O_2886,N_28949,N_27081);
xor UO_2887 (O_2887,N_29571,N_28659);
nor UO_2888 (O_2888,N_28315,N_28712);
nand UO_2889 (O_2889,N_27425,N_28131);
and UO_2890 (O_2890,N_28578,N_28505);
nand UO_2891 (O_2891,N_28083,N_27220);
and UO_2892 (O_2892,N_29313,N_29265);
nor UO_2893 (O_2893,N_27976,N_29291);
nor UO_2894 (O_2894,N_27943,N_27796);
nand UO_2895 (O_2895,N_28038,N_28505);
nor UO_2896 (O_2896,N_28349,N_27072);
nand UO_2897 (O_2897,N_29091,N_27343);
or UO_2898 (O_2898,N_28114,N_28484);
xnor UO_2899 (O_2899,N_28084,N_28595);
xnor UO_2900 (O_2900,N_28659,N_27664);
nand UO_2901 (O_2901,N_27975,N_29649);
and UO_2902 (O_2902,N_29269,N_27915);
nor UO_2903 (O_2903,N_27837,N_27902);
or UO_2904 (O_2904,N_28102,N_29961);
nand UO_2905 (O_2905,N_29310,N_27163);
or UO_2906 (O_2906,N_27521,N_29780);
and UO_2907 (O_2907,N_27385,N_29031);
nor UO_2908 (O_2908,N_28081,N_28534);
or UO_2909 (O_2909,N_28874,N_29259);
or UO_2910 (O_2910,N_29373,N_29846);
xnor UO_2911 (O_2911,N_28818,N_29462);
nor UO_2912 (O_2912,N_27106,N_29981);
nor UO_2913 (O_2913,N_27746,N_29425);
xnor UO_2914 (O_2914,N_27162,N_29787);
or UO_2915 (O_2915,N_27779,N_28061);
nand UO_2916 (O_2916,N_29116,N_29611);
or UO_2917 (O_2917,N_27105,N_28357);
or UO_2918 (O_2918,N_29645,N_28522);
nor UO_2919 (O_2919,N_27440,N_27242);
nand UO_2920 (O_2920,N_28206,N_28265);
or UO_2921 (O_2921,N_27897,N_27720);
nor UO_2922 (O_2922,N_27546,N_28105);
or UO_2923 (O_2923,N_27630,N_29396);
xor UO_2924 (O_2924,N_28051,N_28282);
xor UO_2925 (O_2925,N_28092,N_27958);
xnor UO_2926 (O_2926,N_28604,N_28531);
or UO_2927 (O_2927,N_29503,N_29784);
nand UO_2928 (O_2928,N_28196,N_29048);
xnor UO_2929 (O_2929,N_29138,N_27628);
or UO_2930 (O_2930,N_27070,N_29643);
nor UO_2931 (O_2931,N_27339,N_29343);
xor UO_2932 (O_2932,N_29887,N_27519);
or UO_2933 (O_2933,N_28934,N_28544);
or UO_2934 (O_2934,N_28797,N_28522);
or UO_2935 (O_2935,N_29393,N_28479);
xor UO_2936 (O_2936,N_29071,N_29173);
and UO_2937 (O_2937,N_27404,N_29101);
nand UO_2938 (O_2938,N_29453,N_27301);
xor UO_2939 (O_2939,N_29129,N_27384);
xor UO_2940 (O_2940,N_28436,N_27394);
nor UO_2941 (O_2941,N_27894,N_27563);
nand UO_2942 (O_2942,N_27869,N_27217);
xnor UO_2943 (O_2943,N_29150,N_27988);
or UO_2944 (O_2944,N_29940,N_27992);
nand UO_2945 (O_2945,N_28351,N_28760);
nor UO_2946 (O_2946,N_28038,N_29817);
and UO_2947 (O_2947,N_27270,N_28548);
nand UO_2948 (O_2948,N_27637,N_28321);
and UO_2949 (O_2949,N_29968,N_27177);
nand UO_2950 (O_2950,N_29514,N_28645);
nand UO_2951 (O_2951,N_27778,N_28236);
and UO_2952 (O_2952,N_27436,N_28089);
or UO_2953 (O_2953,N_28427,N_28804);
and UO_2954 (O_2954,N_27458,N_27454);
nand UO_2955 (O_2955,N_27850,N_29944);
and UO_2956 (O_2956,N_28542,N_28334);
xnor UO_2957 (O_2957,N_28387,N_29564);
nand UO_2958 (O_2958,N_28491,N_29791);
nand UO_2959 (O_2959,N_28075,N_29677);
or UO_2960 (O_2960,N_27625,N_29634);
nand UO_2961 (O_2961,N_28848,N_29220);
xor UO_2962 (O_2962,N_29598,N_27735);
and UO_2963 (O_2963,N_29556,N_29536);
nor UO_2964 (O_2964,N_27836,N_29272);
nor UO_2965 (O_2965,N_28848,N_29134);
nand UO_2966 (O_2966,N_29281,N_27557);
or UO_2967 (O_2967,N_29993,N_28937);
nor UO_2968 (O_2968,N_27474,N_29098);
xnor UO_2969 (O_2969,N_28426,N_27140);
nor UO_2970 (O_2970,N_27266,N_28377);
and UO_2971 (O_2971,N_27886,N_28092);
nor UO_2972 (O_2972,N_27092,N_29715);
nand UO_2973 (O_2973,N_28005,N_29107);
and UO_2974 (O_2974,N_29927,N_28317);
or UO_2975 (O_2975,N_27403,N_28366);
xor UO_2976 (O_2976,N_28161,N_27620);
nand UO_2977 (O_2977,N_27668,N_28930);
xor UO_2978 (O_2978,N_28752,N_28164);
or UO_2979 (O_2979,N_28916,N_28082);
nor UO_2980 (O_2980,N_28219,N_29679);
and UO_2981 (O_2981,N_29451,N_28475);
and UO_2982 (O_2982,N_28328,N_28722);
nor UO_2983 (O_2983,N_29329,N_29972);
nor UO_2984 (O_2984,N_27542,N_27485);
xor UO_2985 (O_2985,N_29197,N_29154);
or UO_2986 (O_2986,N_27717,N_27146);
and UO_2987 (O_2987,N_28860,N_29890);
nand UO_2988 (O_2988,N_27247,N_28123);
and UO_2989 (O_2989,N_29573,N_27022);
and UO_2990 (O_2990,N_27259,N_28712);
and UO_2991 (O_2991,N_28751,N_27221);
and UO_2992 (O_2992,N_27490,N_27198);
and UO_2993 (O_2993,N_29144,N_27045);
and UO_2994 (O_2994,N_27291,N_29401);
xor UO_2995 (O_2995,N_29372,N_29090);
and UO_2996 (O_2996,N_28795,N_29643);
xor UO_2997 (O_2997,N_29729,N_29638);
nand UO_2998 (O_2998,N_29153,N_29916);
and UO_2999 (O_2999,N_27339,N_27557);
and UO_3000 (O_3000,N_29269,N_27089);
or UO_3001 (O_3001,N_28542,N_28103);
and UO_3002 (O_3002,N_29087,N_28958);
and UO_3003 (O_3003,N_27099,N_27075);
or UO_3004 (O_3004,N_27336,N_27581);
nor UO_3005 (O_3005,N_28597,N_28407);
xor UO_3006 (O_3006,N_29305,N_27960);
nor UO_3007 (O_3007,N_29532,N_29174);
nor UO_3008 (O_3008,N_27679,N_29709);
nand UO_3009 (O_3009,N_27328,N_29153);
and UO_3010 (O_3010,N_28514,N_27533);
nand UO_3011 (O_3011,N_28798,N_28205);
nand UO_3012 (O_3012,N_28011,N_28128);
nand UO_3013 (O_3013,N_27971,N_28486);
xor UO_3014 (O_3014,N_29303,N_27455);
nor UO_3015 (O_3015,N_27420,N_27636);
nand UO_3016 (O_3016,N_28303,N_27895);
or UO_3017 (O_3017,N_27147,N_29143);
or UO_3018 (O_3018,N_28611,N_29091);
and UO_3019 (O_3019,N_29907,N_27418);
xor UO_3020 (O_3020,N_28746,N_28977);
or UO_3021 (O_3021,N_28670,N_29293);
nand UO_3022 (O_3022,N_28417,N_29536);
nand UO_3023 (O_3023,N_27635,N_28229);
nand UO_3024 (O_3024,N_29083,N_29147);
and UO_3025 (O_3025,N_28442,N_27311);
and UO_3026 (O_3026,N_28105,N_28804);
or UO_3027 (O_3027,N_27494,N_28379);
nand UO_3028 (O_3028,N_29206,N_29144);
nor UO_3029 (O_3029,N_27718,N_29562);
nor UO_3030 (O_3030,N_29658,N_27331);
xnor UO_3031 (O_3031,N_28490,N_27885);
nor UO_3032 (O_3032,N_27099,N_29612);
xnor UO_3033 (O_3033,N_29967,N_28390);
nor UO_3034 (O_3034,N_29790,N_29519);
xor UO_3035 (O_3035,N_29195,N_28835);
xor UO_3036 (O_3036,N_28647,N_28661);
xnor UO_3037 (O_3037,N_28679,N_29356);
xnor UO_3038 (O_3038,N_27379,N_29584);
and UO_3039 (O_3039,N_27363,N_29940);
nand UO_3040 (O_3040,N_28541,N_28414);
xor UO_3041 (O_3041,N_29650,N_29242);
nor UO_3042 (O_3042,N_29547,N_27638);
xor UO_3043 (O_3043,N_27474,N_29753);
nor UO_3044 (O_3044,N_27486,N_27798);
nor UO_3045 (O_3045,N_28229,N_28595);
nand UO_3046 (O_3046,N_29244,N_28547);
nand UO_3047 (O_3047,N_28284,N_27251);
and UO_3048 (O_3048,N_27577,N_28641);
or UO_3049 (O_3049,N_29901,N_27345);
or UO_3050 (O_3050,N_27628,N_28713);
nand UO_3051 (O_3051,N_27749,N_28117);
xnor UO_3052 (O_3052,N_27731,N_29037);
and UO_3053 (O_3053,N_28201,N_27768);
xnor UO_3054 (O_3054,N_27451,N_27411);
nand UO_3055 (O_3055,N_27545,N_27884);
nand UO_3056 (O_3056,N_28624,N_27984);
and UO_3057 (O_3057,N_28296,N_27289);
and UO_3058 (O_3058,N_29246,N_27583);
and UO_3059 (O_3059,N_29768,N_29041);
and UO_3060 (O_3060,N_28406,N_29333);
nor UO_3061 (O_3061,N_28677,N_27857);
nand UO_3062 (O_3062,N_27723,N_27071);
nand UO_3063 (O_3063,N_28047,N_27219);
xnor UO_3064 (O_3064,N_29164,N_29787);
and UO_3065 (O_3065,N_28583,N_28530);
xor UO_3066 (O_3066,N_27435,N_29515);
nor UO_3067 (O_3067,N_28404,N_29265);
or UO_3068 (O_3068,N_28282,N_29186);
xnor UO_3069 (O_3069,N_27259,N_27684);
or UO_3070 (O_3070,N_27468,N_27263);
xnor UO_3071 (O_3071,N_29533,N_29254);
xnor UO_3072 (O_3072,N_27100,N_28462);
and UO_3073 (O_3073,N_27989,N_27191);
xor UO_3074 (O_3074,N_29927,N_28655);
and UO_3075 (O_3075,N_29052,N_27398);
or UO_3076 (O_3076,N_28152,N_29716);
nor UO_3077 (O_3077,N_27007,N_27652);
or UO_3078 (O_3078,N_28846,N_29930);
nor UO_3079 (O_3079,N_29946,N_29016);
or UO_3080 (O_3080,N_28772,N_28395);
or UO_3081 (O_3081,N_29587,N_28222);
and UO_3082 (O_3082,N_28880,N_29777);
xnor UO_3083 (O_3083,N_28571,N_28171);
xnor UO_3084 (O_3084,N_29359,N_28388);
xor UO_3085 (O_3085,N_28988,N_28609);
and UO_3086 (O_3086,N_29156,N_29049);
and UO_3087 (O_3087,N_27550,N_27800);
or UO_3088 (O_3088,N_28278,N_27811);
nand UO_3089 (O_3089,N_29100,N_28734);
and UO_3090 (O_3090,N_29088,N_29584);
and UO_3091 (O_3091,N_28504,N_29561);
xor UO_3092 (O_3092,N_28052,N_29542);
xor UO_3093 (O_3093,N_27427,N_28260);
nor UO_3094 (O_3094,N_29556,N_29291);
xnor UO_3095 (O_3095,N_29382,N_29678);
or UO_3096 (O_3096,N_27988,N_29893);
nand UO_3097 (O_3097,N_28884,N_27807);
nor UO_3098 (O_3098,N_28548,N_28411);
and UO_3099 (O_3099,N_29173,N_27727);
nand UO_3100 (O_3100,N_29311,N_27599);
nor UO_3101 (O_3101,N_27520,N_29766);
and UO_3102 (O_3102,N_29559,N_29171);
nand UO_3103 (O_3103,N_28237,N_28607);
xor UO_3104 (O_3104,N_28714,N_29635);
or UO_3105 (O_3105,N_28156,N_28002);
nand UO_3106 (O_3106,N_28512,N_28184);
nor UO_3107 (O_3107,N_28082,N_28586);
xnor UO_3108 (O_3108,N_28083,N_28602);
nand UO_3109 (O_3109,N_28974,N_28124);
nand UO_3110 (O_3110,N_28296,N_27241);
nor UO_3111 (O_3111,N_29346,N_27830);
nand UO_3112 (O_3112,N_27880,N_28133);
or UO_3113 (O_3113,N_28791,N_28500);
nand UO_3114 (O_3114,N_27119,N_29251);
xor UO_3115 (O_3115,N_29352,N_29219);
xnor UO_3116 (O_3116,N_29817,N_27983);
nand UO_3117 (O_3117,N_28164,N_29423);
nand UO_3118 (O_3118,N_27932,N_28340);
nor UO_3119 (O_3119,N_29115,N_27497);
and UO_3120 (O_3120,N_29956,N_29603);
nand UO_3121 (O_3121,N_28216,N_29990);
nand UO_3122 (O_3122,N_28406,N_29345);
xor UO_3123 (O_3123,N_27436,N_29424);
and UO_3124 (O_3124,N_27976,N_28694);
nor UO_3125 (O_3125,N_28822,N_29953);
and UO_3126 (O_3126,N_29942,N_29189);
xnor UO_3127 (O_3127,N_29697,N_27828);
or UO_3128 (O_3128,N_27417,N_28135);
nand UO_3129 (O_3129,N_28810,N_29440);
and UO_3130 (O_3130,N_28772,N_27577);
nand UO_3131 (O_3131,N_29281,N_27243);
or UO_3132 (O_3132,N_29465,N_27309);
nand UO_3133 (O_3133,N_28209,N_27435);
nand UO_3134 (O_3134,N_27068,N_28492);
or UO_3135 (O_3135,N_27788,N_27132);
nor UO_3136 (O_3136,N_28210,N_28094);
nand UO_3137 (O_3137,N_29431,N_27554);
nand UO_3138 (O_3138,N_29781,N_29211);
or UO_3139 (O_3139,N_27687,N_28253);
and UO_3140 (O_3140,N_27274,N_29113);
nand UO_3141 (O_3141,N_29696,N_27912);
nor UO_3142 (O_3142,N_29202,N_28598);
or UO_3143 (O_3143,N_28840,N_29350);
xnor UO_3144 (O_3144,N_28671,N_27984);
or UO_3145 (O_3145,N_27467,N_29371);
nand UO_3146 (O_3146,N_28847,N_28464);
or UO_3147 (O_3147,N_29422,N_29461);
or UO_3148 (O_3148,N_28814,N_28177);
nor UO_3149 (O_3149,N_27620,N_27409);
xor UO_3150 (O_3150,N_27361,N_27792);
nand UO_3151 (O_3151,N_27606,N_28268);
xor UO_3152 (O_3152,N_29986,N_28202);
and UO_3153 (O_3153,N_27731,N_28233);
and UO_3154 (O_3154,N_29980,N_29835);
nand UO_3155 (O_3155,N_27807,N_27992);
xor UO_3156 (O_3156,N_28524,N_28571);
nand UO_3157 (O_3157,N_29328,N_27110);
xor UO_3158 (O_3158,N_27793,N_29912);
xnor UO_3159 (O_3159,N_29029,N_28271);
nor UO_3160 (O_3160,N_28653,N_29530);
nand UO_3161 (O_3161,N_29487,N_29013);
nand UO_3162 (O_3162,N_29657,N_28396);
nand UO_3163 (O_3163,N_28914,N_29810);
nor UO_3164 (O_3164,N_28361,N_27657);
xor UO_3165 (O_3165,N_27859,N_27749);
or UO_3166 (O_3166,N_29257,N_28216);
nor UO_3167 (O_3167,N_28832,N_29334);
nand UO_3168 (O_3168,N_27341,N_27309);
nor UO_3169 (O_3169,N_29948,N_29543);
and UO_3170 (O_3170,N_29546,N_29170);
or UO_3171 (O_3171,N_29685,N_27264);
and UO_3172 (O_3172,N_29702,N_29873);
nand UO_3173 (O_3173,N_28662,N_28854);
and UO_3174 (O_3174,N_29602,N_29309);
xnor UO_3175 (O_3175,N_27996,N_29311);
xor UO_3176 (O_3176,N_27303,N_28671);
xor UO_3177 (O_3177,N_29343,N_27013);
nand UO_3178 (O_3178,N_27717,N_27296);
and UO_3179 (O_3179,N_27069,N_28858);
nor UO_3180 (O_3180,N_27918,N_29572);
nand UO_3181 (O_3181,N_27185,N_29358);
xor UO_3182 (O_3182,N_27522,N_29247);
or UO_3183 (O_3183,N_29335,N_29741);
nand UO_3184 (O_3184,N_28491,N_27408);
xor UO_3185 (O_3185,N_27859,N_27389);
xnor UO_3186 (O_3186,N_28513,N_29018);
xnor UO_3187 (O_3187,N_29685,N_28401);
nor UO_3188 (O_3188,N_29817,N_27044);
and UO_3189 (O_3189,N_29728,N_27781);
xor UO_3190 (O_3190,N_27050,N_27120);
xor UO_3191 (O_3191,N_28345,N_27937);
nor UO_3192 (O_3192,N_27571,N_29627);
nand UO_3193 (O_3193,N_27864,N_27895);
xnor UO_3194 (O_3194,N_29796,N_27679);
and UO_3195 (O_3195,N_29358,N_29158);
and UO_3196 (O_3196,N_27395,N_28066);
nor UO_3197 (O_3197,N_27901,N_29253);
nor UO_3198 (O_3198,N_27602,N_27214);
xnor UO_3199 (O_3199,N_27389,N_28553);
and UO_3200 (O_3200,N_27944,N_28496);
nor UO_3201 (O_3201,N_29601,N_28284);
xnor UO_3202 (O_3202,N_29646,N_27722);
xor UO_3203 (O_3203,N_28071,N_27210);
xnor UO_3204 (O_3204,N_28921,N_28992);
and UO_3205 (O_3205,N_28079,N_27980);
and UO_3206 (O_3206,N_28217,N_27024);
nor UO_3207 (O_3207,N_28275,N_29369);
and UO_3208 (O_3208,N_27337,N_29128);
nand UO_3209 (O_3209,N_28267,N_28344);
xnor UO_3210 (O_3210,N_29585,N_28941);
nor UO_3211 (O_3211,N_28817,N_27386);
and UO_3212 (O_3212,N_29041,N_27540);
nand UO_3213 (O_3213,N_28601,N_28269);
nor UO_3214 (O_3214,N_27970,N_29684);
nor UO_3215 (O_3215,N_27181,N_27032);
xnor UO_3216 (O_3216,N_29180,N_29943);
nand UO_3217 (O_3217,N_27844,N_29041);
nor UO_3218 (O_3218,N_27923,N_28388);
or UO_3219 (O_3219,N_27007,N_27217);
nand UO_3220 (O_3220,N_28636,N_28003);
nor UO_3221 (O_3221,N_27464,N_27318);
and UO_3222 (O_3222,N_29532,N_28161);
nand UO_3223 (O_3223,N_29579,N_27524);
nor UO_3224 (O_3224,N_29496,N_27079);
nand UO_3225 (O_3225,N_29976,N_29710);
nor UO_3226 (O_3226,N_28639,N_27815);
nor UO_3227 (O_3227,N_27256,N_27818);
nor UO_3228 (O_3228,N_27955,N_27090);
xnor UO_3229 (O_3229,N_29971,N_29388);
nor UO_3230 (O_3230,N_29862,N_28702);
and UO_3231 (O_3231,N_27219,N_27373);
xor UO_3232 (O_3232,N_28141,N_28373);
nor UO_3233 (O_3233,N_28392,N_29928);
and UO_3234 (O_3234,N_27078,N_28057);
and UO_3235 (O_3235,N_27742,N_28496);
nand UO_3236 (O_3236,N_28384,N_29217);
xnor UO_3237 (O_3237,N_27022,N_28920);
nor UO_3238 (O_3238,N_29571,N_29268);
nor UO_3239 (O_3239,N_28027,N_28733);
or UO_3240 (O_3240,N_28325,N_28320);
nand UO_3241 (O_3241,N_28959,N_27458);
nand UO_3242 (O_3242,N_27540,N_27298);
nand UO_3243 (O_3243,N_29271,N_27430);
nand UO_3244 (O_3244,N_28457,N_29638);
xnor UO_3245 (O_3245,N_29346,N_27848);
xor UO_3246 (O_3246,N_27223,N_28771);
nor UO_3247 (O_3247,N_27578,N_29359);
and UO_3248 (O_3248,N_28014,N_27788);
xor UO_3249 (O_3249,N_29990,N_29000);
nand UO_3250 (O_3250,N_29588,N_28329);
or UO_3251 (O_3251,N_29179,N_28132);
nand UO_3252 (O_3252,N_29220,N_29069);
and UO_3253 (O_3253,N_27160,N_28048);
and UO_3254 (O_3254,N_27870,N_28873);
and UO_3255 (O_3255,N_29561,N_28973);
or UO_3256 (O_3256,N_27371,N_27704);
and UO_3257 (O_3257,N_27722,N_27715);
or UO_3258 (O_3258,N_27165,N_29399);
nor UO_3259 (O_3259,N_28067,N_27885);
or UO_3260 (O_3260,N_29249,N_28818);
and UO_3261 (O_3261,N_29583,N_29983);
nor UO_3262 (O_3262,N_27474,N_29786);
xnor UO_3263 (O_3263,N_29089,N_28552);
or UO_3264 (O_3264,N_27753,N_27530);
or UO_3265 (O_3265,N_29906,N_27688);
and UO_3266 (O_3266,N_27698,N_29485);
nor UO_3267 (O_3267,N_27361,N_27610);
and UO_3268 (O_3268,N_27546,N_27198);
nand UO_3269 (O_3269,N_29919,N_27532);
xnor UO_3270 (O_3270,N_29896,N_27209);
nand UO_3271 (O_3271,N_27760,N_29493);
nor UO_3272 (O_3272,N_29803,N_29420);
and UO_3273 (O_3273,N_29558,N_28831);
nand UO_3274 (O_3274,N_29662,N_28757);
xor UO_3275 (O_3275,N_28876,N_27573);
nand UO_3276 (O_3276,N_28103,N_29917);
nor UO_3277 (O_3277,N_27666,N_28123);
xor UO_3278 (O_3278,N_28840,N_29206);
and UO_3279 (O_3279,N_28634,N_29427);
xnor UO_3280 (O_3280,N_28517,N_28262);
and UO_3281 (O_3281,N_27930,N_29517);
or UO_3282 (O_3282,N_29794,N_28404);
xnor UO_3283 (O_3283,N_27576,N_29234);
or UO_3284 (O_3284,N_28799,N_29573);
nor UO_3285 (O_3285,N_29564,N_29498);
or UO_3286 (O_3286,N_28839,N_29972);
xnor UO_3287 (O_3287,N_29984,N_28415);
xor UO_3288 (O_3288,N_27619,N_27066);
and UO_3289 (O_3289,N_27937,N_27452);
nand UO_3290 (O_3290,N_28564,N_28306);
nor UO_3291 (O_3291,N_28375,N_28452);
nor UO_3292 (O_3292,N_29541,N_27431);
xnor UO_3293 (O_3293,N_27116,N_28432);
xor UO_3294 (O_3294,N_27968,N_28834);
xnor UO_3295 (O_3295,N_27239,N_29392);
xor UO_3296 (O_3296,N_27965,N_28285);
xnor UO_3297 (O_3297,N_28769,N_29305);
nor UO_3298 (O_3298,N_27131,N_27959);
xnor UO_3299 (O_3299,N_29089,N_27881);
and UO_3300 (O_3300,N_29231,N_28163);
or UO_3301 (O_3301,N_28007,N_28435);
and UO_3302 (O_3302,N_27339,N_28658);
and UO_3303 (O_3303,N_28312,N_27507);
nor UO_3304 (O_3304,N_27173,N_29400);
nand UO_3305 (O_3305,N_27603,N_29375);
nand UO_3306 (O_3306,N_28084,N_28793);
and UO_3307 (O_3307,N_28365,N_29058);
and UO_3308 (O_3308,N_28174,N_29139);
or UO_3309 (O_3309,N_27579,N_29299);
xnor UO_3310 (O_3310,N_29814,N_29872);
nand UO_3311 (O_3311,N_29933,N_29080);
xor UO_3312 (O_3312,N_29531,N_29791);
or UO_3313 (O_3313,N_28528,N_29216);
nor UO_3314 (O_3314,N_28343,N_27257);
xnor UO_3315 (O_3315,N_28409,N_27421);
or UO_3316 (O_3316,N_29114,N_29882);
xor UO_3317 (O_3317,N_28794,N_28749);
and UO_3318 (O_3318,N_28539,N_28668);
nor UO_3319 (O_3319,N_28020,N_27041);
and UO_3320 (O_3320,N_29985,N_28151);
xor UO_3321 (O_3321,N_27834,N_28207);
nand UO_3322 (O_3322,N_27952,N_29527);
xor UO_3323 (O_3323,N_28662,N_28708);
and UO_3324 (O_3324,N_29122,N_27907);
nor UO_3325 (O_3325,N_27028,N_27639);
nand UO_3326 (O_3326,N_29063,N_28979);
and UO_3327 (O_3327,N_28603,N_28681);
xnor UO_3328 (O_3328,N_27043,N_29515);
nand UO_3329 (O_3329,N_27784,N_28194);
xor UO_3330 (O_3330,N_28943,N_27790);
nor UO_3331 (O_3331,N_27326,N_27674);
or UO_3332 (O_3332,N_29038,N_28056);
nand UO_3333 (O_3333,N_28353,N_28981);
xor UO_3334 (O_3334,N_28089,N_28040);
or UO_3335 (O_3335,N_28930,N_29531);
and UO_3336 (O_3336,N_27774,N_27825);
nand UO_3337 (O_3337,N_29832,N_27984);
nor UO_3338 (O_3338,N_27994,N_27925);
or UO_3339 (O_3339,N_29128,N_27683);
and UO_3340 (O_3340,N_28740,N_27552);
or UO_3341 (O_3341,N_29301,N_27565);
and UO_3342 (O_3342,N_28029,N_29637);
nand UO_3343 (O_3343,N_29772,N_29257);
nor UO_3344 (O_3344,N_29880,N_28485);
nand UO_3345 (O_3345,N_27233,N_27699);
nor UO_3346 (O_3346,N_27815,N_29942);
xnor UO_3347 (O_3347,N_29459,N_29356);
nor UO_3348 (O_3348,N_29404,N_28796);
nand UO_3349 (O_3349,N_29568,N_27360);
and UO_3350 (O_3350,N_29682,N_29366);
or UO_3351 (O_3351,N_28269,N_28560);
xor UO_3352 (O_3352,N_29090,N_28756);
or UO_3353 (O_3353,N_29308,N_27716);
xor UO_3354 (O_3354,N_27969,N_28858);
nand UO_3355 (O_3355,N_29278,N_29948);
or UO_3356 (O_3356,N_27397,N_28855);
nand UO_3357 (O_3357,N_29402,N_28584);
or UO_3358 (O_3358,N_27091,N_29055);
xnor UO_3359 (O_3359,N_29014,N_28836);
nand UO_3360 (O_3360,N_27523,N_28567);
nor UO_3361 (O_3361,N_27181,N_27819);
and UO_3362 (O_3362,N_27488,N_29000);
or UO_3363 (O_3363,N_27784,N_28044);
nor UO_3364 (O_3364,N_29215,N_27556);
xnor UO_3365 (O_3365,N_28935,N_28664);
and UO_3366 (O_3366,N_28567,N_28463);
nand UO_3367 (O_3367,N_29364,N_28324);
or UO_3368 (O_3368,N_27997,N_29049);
nand UO_3369 (O_3369,N_28706,N_29582);
nand UO_3370 (O_3370,N_27480,N_28652);
nor UO_3371 (O_3371,N_28029,N_29419);
and UO_3372 (O_3372,N_29256,N_28962);
nand UO_3373 (O_3373,N_27025,N_27048);
or UO_3374 (O_3374,N_27328,N_29053);
or UO_3375 (O_3375,N_27625,N_27872);
nand UO_3376 (O_3376,N_29313,N_28501);
or UO_3377 (O_3377,N_28245,N_28436);
nand UO_3378 (O_3378,N_28311,N_28352);
nand UO_3379 (O_3379,N_28497,N_27560);
nor UO_3380 (O_3380,N_27592,N_27665);
xnor UO_3381 (O_3381,N_28772,N_29128);
nand UO_3382 (O_3382,N_29458,N_28035);
nand UO_3383 (O_3383,N_28605,N_29883);
and UO_3384 (O_3384,N_29009,N_29991);
nand UO_3385 (O_3385,N_28005,N_28173);
or UO_3386 (O_3386,N_29890,N_28488);
xnor UO_3387 (O_3387,N_27188,N_27835);
nand UO_3388 (O_3388,N_28808,N_28244);
nand UO_3389 (O_3389,N_29802,N_28250);
nand UO_3390 (O_3390,N_27031,N_29167);
nand UO_3391 (O_3391,N_27279,N_28727);
or UO_3392 (O_3392,N_28237,N_28446);
or UO_3393 (O_3393,N_27573,N_29921);
xor UO_3394 (O_3394,N_29662,N_29042);
xnor UO_3395 (O_3395,N_29104,N_29544);
nand UO_3396 (O_3396,N_28000,N_29591);
or UO_3397 (O_3397,N_27300,N_29640);
or UO_3398 (O_3398,N_29327,N_28348);
nand UO_3399 (O_3399,N_27247,N_28536);
nand UO_3400 (O_3400,N_29194,N_28938);
or UO_3401 (O_3401,N_27506,N_27476);
or UO_3402 (O_3402,N_27454,N_29324);
nor UO_3403 (O_3403,N_28684,N_27458);
xnor UO_3404 (O_3404,N_28279,N_28658);
xor UO_3405 (O_3405,N_28821,N_29270);
nor UO_3406 (O_3406,N_28582,N_27109);
xnor UO_3407 (O_3407,N_29215,N_28224);
and UO_3408 (O_3408,N_28971,N_29278);
xor UO_3409 (O_3409,N_27386,N_28951);
nand UO_3410 (O_3410,N_28323,N_29631);
nor UO_3411 (O_3411,N_29897,N_28070);
nor UO_3412 (O_3412,N_29302,N_27575);
nand UO_3413 (O_3413,N_28654,N_28394);
nand UO_3414 (O_3414,N_28638,N_28695);
or UO_3415 (O_3415,N_27430,N_27118);
and UO_3416 (O_3416,N_28041,N_28160);
or UO_3417 (O_3417,N_28982,N_29843);
or UO_3418 (O_3418,N_27761,N_28260);
nor UO_3419 (O_3419,N_28889,N_29277);
nor UO_3420 (O_3420,N_28704,N_28051);
xnor UO_3421 (O_3421,N_27663,N_29299);
and UO_3422 (O_3422,N_29690,N_28134);
or UO_3423 (O_3423,N_29133,N_27228);
xor UO_3424 (O_3424,N_28407,N_28255);
or UO_3425 (O_3425,N_28454,N_29607);
or UO_3426 (O_3426,N_27903,N_27150);
nor UO_3427 (O_3427,N_28934,N_29224);
nor UO_3428 (O_3428,N_28481,N_29474);
nand UO_3429 (O_3429,N_28339,N_27988);
nor UO_3430 (O_3430,N_29986,N_29286);
and UO_3431 (O_3431,N_29319,N_27427);
nand UO_3432 (O_3432,N_28865,N_29305);
nor UO_3433 (O_3433,N_27738,N_27165);
and UO_3434 (O_3434,N_29226,N_29285);
or UO_3435 (O_3435,N_28442,N_29000);
or UO_3436 (O_3436,N_28753,N_28676);
and UO_3437 (O_3437,N_27604,N_29710);
or UO_3438 (O_3438,N_27517,N_28470);
or UO_3439 (O_3439,N_29901,N_27486);
or UO_3440 (O_3440,N_29629,N_29225);
nor UO_3441 (O_3441,N_29100,N_28681);
or UO_3442 (O_3442,N_28322,N_28007);
or UO_3443 (O_3443,N_28288,N_29442);
or UO_3444 (O_3444,N_29462,N_28571);
nor UO_3445 (O_3445,N_29726,N_27242);
nand UO_3446 (O_3446,N_29763,N_27740);
nand UO_3447 (O_3447,N_29705,N_27218);
nand UO_3448 (O_3448,N_29915,N_27785);
or UO_3449 (O_3449,N_27554,N_28231);
nand UO_3450 (O_3450,N_29744,N_27610);
and UO_3451 (O_3451,N_27219,N_27666);
nor UO_3452 (O_3452,N_27970,N_28150);
nor UO_3453 (O_3453,N_28039,N_28467);
and UO_3454 (O_3454,N_29357,N_29106);
or UO_3455 (O_3455,N_29899,N_27900);
xor UO_3456 (O_3456,N_27424,N_27754);
xnor UO_3457 (O_3457,N_27679,N_29718);
xor UO_3458 (O_3458,N_28539,N_27099);
nand UO_3459 (O_3459,N_27083,N_27553);
nand UO_3460 (O_3460,N_29967,N_27740);
nand UO_3461 (O_3461,N_29692,N_28383);
and UO_3462 (O_3462,N_29023,N_28643);
and UO_3463 (O_3463,N_27986,N_29100);
and UO_3464 (O_3464,N_27029,N_27158);
or UO_3465 (O_3465,N_29522,N_29679);
xnor UO_3466 (O_3466,N_29138,N_28676);
and UO_3467 (O_3467,N_29698,N_29006);
and UO_3468 (O_3468,N_29367,N_29114);
or UO_3469 (O_3469,N_28309,N_28450);
and UO_3470 (O_3470,N_28682,N_29323);
and UO_3471 (O_3471,N_28381,N_28161);
xor UO_3472 (O_3472,N_28716,N_29846);
and UO_3473 (O_3473,N_29646,N_29197);
or UO_3474 (O_3474,N_28877,N_29895);
nand UO_3475 (O_3475,N_28110,N_27405);
nor UO_3476 (O_3476,N_27660,N_29933);
nor UO_3477 (O_3477,N_29906,N_29726);
or UO_3478 (O_3478,N_29454,N_29822);
nand UO_3479 (O_3479,N_29500,N_29125);
xor UO_3480 (O_3480,N_29170,N_27694);
nor UO_3481 (O_3481,N_27696,N_28852);
or UO_3482 (O_3482,N_28594,N_28859);
xnor UO_3483 (O_3483,N_27975,N_27925);
xor UO_3484 (O_3484,N_29916,N_29885);
xor UO_3485 (O_3485,N_29912,N_28379);
nor UO_3486 (O_3486,N_28161,N_29784);
nor UO_3487 (O_3487,N_28974,N_27053);
and UO_3488 (O_3488,N_28139,N_28961);
and UO_3489 (O_3489,N_27136,N_29838);
and UO_3490 (O_3490,N_28636,N_28774);
nor UO_3491 (O_3491,N_27342,N_29933);
or UO_3492 (O_3492,N_27460,N_29363);
and UO_3493 (O_3493,N_29306,N_28471);
nand UO_3494 (O_3494,N_27063,N_29262);
or UO_3495 (O_3495,N_29406,N_29590);
xnor UO_3496 (O_3496,N_29629,N_27085);
nand UO_3497 (O_3497,N_29242,N_29715);
xnor UO_3498 (O_3498,N_27448,N_28291);
or UO_3499 (O_3499,N_28785,N_29376);
endmodule