module basic_500_3000_500_3_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_259,In_112);
xor U1 (N_1,In_431,In_214);
nand U2 (N_2,In_458,In_359);
or U3 (N_3,In_292,In_143);
nor U4 (N_4,In_140,In_365);
and U5 (N_5,In_320,In_286);
and U6 (N_6,In_8,In_151);
nand U7 (N_7,In_170,In_402);
nor U8 (N_8,In_487,In_485);
nor U9 (N_9,In_194,In_148);
or U10 (N_10,In_264,In_212);
nor U11 (N_11,In_435,In_417);
and U12 (N_12,In_132,In_142);
nor U13 (N_13,In_375,In_316);
or U14 (N_14,In_12,In_276);
and U15 (N_15,In_237,In_413);
or U16 (N_16,In_342,In_400);
or U17 (N_17,In_309,In_275);
nand U18 (N_18,In_9,In_70);
and U19 (N_19,In_69,In_414);
and U20 (N_20,In_44,In_363);
or U21 (N_21,In_257,In_287);
or U22 (N_22,In_24,In_343);
nand U23 (N_23,In_36,In_465);
nand U24 (N_24,In_54,In_416);
or U25 (N_25,In_57,In_32);
nor U26 (N_26,In_354,In_131);
xor U27 (N_27,In_123,In_126);
xor U28 (N_28,In_238,In_491);
xnor U29 (N_29,In_436,In_93);
nand U30 (N_30,In_428,In_163);
or U31 (N_31,In_45,In_454);
and U32 (N_32,In_182,In_498);
and U33 (N_33,In_437,In_298);
and U34 (N_34,In_282,In_220);
and U35 (N_35,In_258,In_84);
or U36 (N_36,In_129,In_27);
or U37 (N_37,In_230,In_85);
and U38 (N_38,In_426,In_249);
nand U39 (N_39,In_154,In_392);
xnor U40 (N_40,In_105,In_33);
nor U41 (N_41,In_364,In_127);
nand U42 (N_42,In_216,In_450);
nor U43 (N_43,In_145,In_335);
or U44 (N_44,In_215,In_455);
xnor U45 (N_45,In_464,In_83);
nor U46 (N_46,In_373,In_334);
or U47 (N_47,In_441,In_374);
and U48 (N_48,In_94,In_56);
or U49 (N_49,In_284,In_277);
nor U50 (N_50,In_159,In_25);
xor U51 (N_51,In_13,In_442);
nand U52 (N_52,In_390,In_79);
nor U53 (N_53,In_474,In_100);
nand U54 (N_54,In_396,In_68);
and U55 (N_55,In_1,In_40);
nand U56 (N_56,In_256,In_62);
or U57 (N_57,In_307,In_80);
or U58 (N_58,In_19,In_87);
and U59 (N_59,In_421,In_3);
and U60 (N_60,In_95,In_248);
nand U61 (N_61,In_207,In_77);
and U62 (N_62,In_462,In_313);
nand U63 (N_63,In_218,In_326);
nor U64 (N_64,In_247,In_319);
nor U65 (N_65,In_254,In_378);
xnor U66 (N_66,In_469,In_337);
xnor U67 (N_67,In_231,In_39);
nand U68 (N_68,In_30,In_466);
xor U69 (N_69,In_196,In_0);
or U70 (N_70,In_353,In_299);
nand U71 (N_71,In_175,In_300);
nor U72 (N_72,In_324,In_246);
nor U73 (N_73,In_211,In_263);
and U74 (N_74,In_371,In_347);
nand U75 (N_75,In_481,In_162);
nor U76 (N_76,In_121,In_395);
and U77 (N_77,In_270,In_167);
xor U78 (N_78,In_409,In_340);
or U79 (N_79,In_47,In_76);
nor U80 (N_80,In_444,In_6);
or U81 (N_81,In_406,In_297);
or U82 (N_82,In_422,In_186);
nor U83 (N_83,In_141,In_133);
and U84 (N_84,In_329,In_296);
or U85 (N_85,In_72,In_43);
or U86 (N_86,In_89,In_193);
nor U87 (N_87,In_331,In_38);
and U88 (N_88,In_201,In_271);
and U89 (N_89,In_295,In_104);
nor U90 (N_90,In_244,In_323);
nor U91 (N_91,In_456,In_261);
xor U92 (N_92,In_479,In_16);
nor U93 (N_93,In_205,In_2);
and U94 (N_94,In_482,In_370);
nand U95 (N_95,In_478,In_403);
and U96 (N_96,In_438,In_302);
or U97 (N_97,In_191,In_433);
nand U98 (N_98,In_91,In_232);
xor U99 (N_99,In_368,In_117);
nor U100 (N_100,In_483,In_388);
nor U101 (N_101,In_168,In_171);
nand U102 (N_102,In_322,In_494);
or U103 (N_103,In_440,In_241);
nor U104 (N_104,In_497,In_475);
or U105 (N_105,In_7,In_360);
nor U106 (N_106,In_383,In_187);
nor U107 (N_107,In_155,In_495);
or U108 (N_108,In_172,In_147);
nor U109 (N_109,In_379,In_119);
nor U110 (N_110,In_273,In_108);
and U111 (N_111,In_17,In_22);
nand U112 (N_112,In_150,In_484);
or U113 (N_113,In_294,In_267);
nand U114 (N_114,In_389,In_423);
or U115 (N_115,In_219,In_46);
nand U116 (N_116,In_386,In_102);
and U117 (N_117,In_197,In_188);
and U118 (N_118,In_74,In_51);
or U119 (N_119,In_260,In_60);
or U120 (N_120,In_408,In_213);
or U121 (N_121,In_303,In_180);
xor U122 (N_122,In_425,In_137);
and U123 (N_123,In_285,In_125);
xnor U124 (N_124,In_21,In_149);
nor U125 (N_125,In_138,In_189);
nand U126 (N_126,In_120,In_449);
and U127 (N_127,In_208,In_473);
nor U128 (N_128,In_430,In_78);
nand U129 (N_129,In_177,In_198);
xor U130 (N_130,In_434,In_50);
and U131 (N_131,In_139,In_190);
or U132 (N_132,In_23,In_5);
nand U133 (N_133,In_288,In_445);
or U134 (N_134,In_245,In_448);
xnor U135 (N_135,In_181,In_461);
or U136 (N_136,In_136,In_317);
or U137 (N_137,In_361,In_34);
nor U138 (N_138,In_327,In_111);
or U139 (N_139,In_107,In_65);
nor U140 (N_140,In_10,In_471);
nand U141 (N_141,In_321,In_311);
and U142 (N_142,In_269,In_115);
nand U143 (N_143,In_217,In_199);
nor U144 (N_144,In_447,In_109);
nand U145 (N_145,In_352,In_28);
and U146 (N_146,In_58,In_463);
nor U147 (N_147,In_289,In_101);
nor U148 (N_148,In_63,In_439);
nor U149 (N_149,In_432,In_55);
or U150 (N_150,In_18,In_429);
nor U151 (N_151,In_266,In_411);
nor U152 (N_152,In_357,In_274);
or U153 (N_153,In_156,In_135);
nor U154 (N_154,In_86,In_272);
and U155 (N_155,In_235,In_15);
nand U156 (N_156,In_233,In_96);
nor U157 (N_157,In_480,In_452);
or U158 (N_158,In_176,In_377);
nor U159 (N_159,In_81,In_407);
nor U160 (N_160,In_476,In_158);
xnor U161 (N_161,In_164,In_418);
or U162 (N_162,In_489,In_173);
or U163 (N_163,In_226,In_397);
and U164 (N_164,In_460,In_355);
nand U165 (N_165,In_486,In_410);
nand U166 (N_166,In_467,In_468);
nand U167 (N_167,In_268,In_399);
nand U168 (N_168,In_92,In_174);
nand U169 (N_169,In_443,In_384);
and U170 (N_170,In_393,In_160);
or U171 (N_171,In_252,In_376);
nor U172 (N_172,In_203,In_349);
nand U173 (N_173,In_255,In_310);
nor U174 (N_174,In_446,In_496);
and U175 (N_175,In_262,In_48);
and U176 (N_176,In_103,In_493);
nand U177 (N_177,In_380,In_308);
or U178 (N_178,In_293,In_183);
nand U179 (N_179,In_225,In_283);
or U180 (N_180,In_52,In_451);
and U181 (N_181,In_394,In_169);
or U182 (N_182,In_239,In_346);
and U183 (N_183,In_49,In_339);
and U184 (N_184,In_37,In_66);
or U185 (N_185,In_457,In_291);
and U186 (N_186,In_195,In_348);
nor U187 (N_187,In_166,In_41);
nand U188 (N_188,In_116,In_209);
and U189 (N_189,In_26,In_35);
and U190 (N_190,In_387,In_114);
and U191 (N_191,In_401,In_382);
or U192 (N_192,In_250,In_315);
and U193 (N_193,In_332,In_229);
nand U194 (N_194,In_279,In_124);
and U195 (N_195,In_67,In_192);
nand U196 (N_196,In_234,In_318);
nor U197 (N_197,In_253,In_152);
nor U198 (N_198,In_351,In_64);
or U199 (N_199,In_369,In_71);
xor U200 (N_200,In_356,In_31);
nor U201 (N_201,In_73,In_204);
or U202 (N_202,In_345,In_398);
xnor U203 (N_203,In_330,In_14);
nand U204 (N_204,In_146,In_210);
nor U205 (N_205,In_122,In_98);
or U206 (N_206,In_75,In_490);
and U207 (N_207,In_381,In_366);
nor U208 (N_208,In_341,In_202);
xnor U209 (N_209,In_222,In_367);
or U210 (N_210,In_42,In_420);
or U211 (N_211,In_224,In_470);
nor U212 (N_212,In_492,In_499);
nand U213 (N_213,In_290,In_82);
and U214 (N_214,In_4,In_328);
nor U215 (N_215,In_336,In_228);
nand U216 (N_216,In_280,In_178);
nand U217 (N_217,In_240,In_206);
xor U218 (N_218,In_236,In_61);
and U219 (N_219,In_11,In_372);
and U220 (N_220,In_165,In_184);
nor U221 (N_221,In_391,In_312);
xor U222 (N_222,In_242,In_53);
nand U223 (N_223,In_325,In_179);
nor U224 (N_224,In_333,In_128);
xnor U225 (N_225,In_453,In_412);
nand U226 (N_226,In_130,In_278);
nand U227 (N_227,In_424,In_110);
xor U228 (N_228,In_243,In_144);
nand U229 (N_229,In_305,In_419);
nand U230 (N_230,In_459,In_134);
nor U231 (N_231,In_118,In_20);
nand U232 (N_232,In_227,In_488);
or U233 (N_233,In_99,In_415);
nor U234 (N_234,In_344,In_221);
nand U235 (N_235,In_161,In_90);
nor U236 (N_236,In_59,In_301);
or U237 (N_237,In_157,In_223);
and U238 (N_238,In_265,In_97);
or U239 (N_239,In_185,In_200);
and U240 (N_240,In_314,In_477);
or U241 (N_241,In_350,In_88);
nand U242 (N_242,In_281,In_29);
and U243 (N_243,In_472,In_405);
xor U244 (N_244,In_427,In_113);
nor U245 (N_245,In_362,In_153);
or U246 (N_246,In_304,In_385);
or U247 (N_247,In_338,In_306);
or U248 (N_248,In_358,In_404);
nor U249 (N_249,In_251,In_106);
nor U250 (N_250,In_183,In_405);
nand U251 (N_251,In_130,In_431);
or U252 (N_252,In_433,In_311);
nand U253 (N_253,In_79,In_473);
xor U254 (N_254,In_258,In_250);
and U255 (N_255,In_240,In_310);
and U256 (N_256,In_328,In_357);
xor U257 (N_257,In_132,In_355);
or U258 (N_258,In_487,In_214);
and U259 (N_259,In_243,In_434);
nand U260 (N_260,In_480,In_308);
or U261 (N_261,In_291,In_169);
nand U262 (N_262,In_187,In_116);
nand U263 (N_263,In_398,In_228);
nor U264 (N_264,In_390,In_186);
nand U265 (N_265,In_153,In_111);
or U266 (N_266,In_428,In_76);
nand U267 (N_267,In_406,In_36);
and U268 (N_268,In_148,In_168);
nor U269 (N_269,In_374,In_48);
nor U270 (N_270,In_265,In_217);
nand U271 (N_271,In_288,In_188);
nor U272 (N_272,In_488,In_295);
nor U273 (N_273,In_248,In_57);
and U274 (N_274,In_288,In_387);
nor U275 (N_275,In_397,In_2);
nand U276 (N_276,In_323,In_352);
nand U277 (N_277,In_75,In_384);
nand U278 (N_278,In_220,In_157);
xnor U279 (N_279,In_17,In_183);
nand U280 (N_280,In_245,In_246);
xnor U281 (N_281,In_298,In_384);
or U282 (N_282,In_483,In_482);
or U283 (N_283,In_17,In_234);
and U284 (N_284,In_401,In_367);
nand U285 (N_285,In_333,In_411);
nand U286 (N_286,In_472,In_395);
nand U287 (N_287,In_203,In_297);
nand U288 (N_288,In_464,In_339);
and U289 (N_289,In_81,In_28);
nand U290 (N_290,In_12,In_302);
nor U291 (N_291,In_92,In_416);
and U292 (N_292,In_347,In_485);
and U293 (N_293,In_134,In_231);
and U294 (N_294,In_330,In_12);
xor U295 (N_295,In_111,In_336);
xor U296 (N_296,In_114,In_432);
or U297 (N_297,In_148,In_421);
nor U298 (N_298,In_368,In_362);
and U299 (N_299,In_34,In_415);
or U300 (N_300,In_92,In_85);
and U301 (N_301,In_122,In_398);
nand U302 (N_302,In_23,In_210);
nand U303 (N_303,In_459,In_82);
nor U304 (N_304,In_457,In_272);
nand U305 (N_305,In_355,In_346);
nor U306 (N_306,In_159,In_329);
or U307 (N_307,In_410,In_499);
or U308 (N_308,In_170,In_367);
nand U309 (N_309,In_117,In_50);
and U310 (N_310,In_246,In_456);
or U311 (N_311,In_90,In_152);
and U312 (N_312,In_327,In_331);
nand U313 (N_313,In_464,In_352);
or U314 (N_314,In_187,In_314);
nor U315 (N_315,In_360,In_490);
and U316 (N_316,In_160,In_443);
or U317 (N_317,In_228,In_213);
nand U318 (N_318,In_101,In_355);
and U319 (N_319,In_259,In_4);
and U320 (N_320,In_173,In_34);
and U321 (N_321,In_2,In_312);
nand U322 (N_322,In_268,In_30);
nand U323 (N_323,In_306,In_420);
nand U324 (N_324,In_151,In_13);
nor U325 (N_325,In_140,In_271);
xnor U326 (N_326,In_40,In_364);
or U327 (N_327,In_315,In_171);
nand U328 (N_328,In_113,In_13);
nor U329 (N_329,In_401,In_275);
nand U330 (N_330,In_313,In_328);
nand U331 (N_331,In_323,In_106);
nor U332 (N_332,In_443,In_63);
and U333 (N_333,In_324,In_494);
xor U334 (N_334,In_295,In_415);
and U335 (N_335,In_58,In_405);
or U336 (N_336,In_470,In_133);
nand U337 (N_337,In_292,In_78);
and U338 (N_338,In_53,In_387);
and U339 (N_339,In_42,In_419);
and U340 (N_340,In_118,In_221);
xnor U341 (N_341,In_188,In_391);
and U342 (N_342,In_20,In_55);
or U343 (N_343,In_325,In_25);
or U344 (N_344,In_104,In_462);
nor U345 (N_345,In_325,In_452);
nand U346 (N_346,In_213,In_91);
nor U347 (N_347,In_150,In_464);
nand U348 (N_348,In_97,In_171);
xnor U349 (N_349,In_217,In_435);
nand U350 (N_350,In_242,In_286);
nand U351 (N_351,In_16,In_349);
xnor U352 (N_352,In_31,In_419);
nor U353 (N_353,In_418,In_49);
nor U354 (N_354,In_388,In_253);
and U355 (N_355,In_456,In_275);
nor U356 (N_356,In_307,In_384);
and U357 (N_357,In_39,In_189);
nand U358 (N_358,In_348,In_409);
or U359 (N_359,In_330,In_162);
nor U360 (N_360,In_21,In_280);
nand U361 (N_361,In_280,In_10);
or U362 (N_362,In_101,In_353);
or U363 (N_363,In_125,In_154);
or U364 (N_364,In_452,In_113);
or U365 (N_365,In_35,In_436);
and U366 (N_366,In_340,In_106);
and U367 (N_367,In_427,In_439);
xnor U368 (N_368,In_196,In_348);
or U369 (N_369,In_421,In_35);
or U370 (N_370,In_352,In_441);
or U371 (N_371,In_375,In_366);
nor U372 (N_372,In_357,In_279);
nand U373 (N_373,In_163,In_487);
nor U374 (N_374,In_248,In_489);
nand U375 (N_375,In_44,In_367);
and U376 (N_376,In_393,In_304);
nor U377 (N_377,In_147,In_2);
nor U378 (N_378,In_166,In_321);
nand U379 (N_379,In_9,In_253);
nor U380 (N_380,In_454,In_50);
nor U381 (N_381,In_250,In_81);
and U382 (N_382,In_353,In_188);
nor U383 (N_383,In_223,In_260);
nor U384 (N_384,In_330,In_305);
and U385 (N_385,In_217,In_132);
nand U386 (N_386,In_334,In_115);
and U387 (N_387,In_318,In_482);
nor U388 (N_388,In_128,In_106);
and U389 (N_389,In_42,In_8);
and U390 (N_390,In_301,In_2);
nand U391 (N_391,In_488,In_421);
or U392 (N_392,In_140,In_182);
nand U393 (N_393,In_301,In_449);
nor U394 (N_394,In_104,In_105);
nand U395 (N_395,In_269,In_268);
nand U396 (N_396,In_358,In_48);
and U397 (N_397,In_475,In_460);
nor U398 (N_398,In_29,In_367);
nor U399 (N_399,In_249,In_342);
and U400 (N_400,In_149,In_252);
or U401 (N_401,In_232,In_421);
xor U402 (N_402,In_178,In_98);
nand U403 (N_403,In_102,In_390);
and U404 (N_404,In_346,In_307);
nand U405 (N_405,In_255,In_400);
nor U406 (N_406,In_408,In_199);
nor U407 (N_407,In_333,In_124);
or U408 (N_408,In_352,In_495);
xnor U409 (N_409,In_484,In_257);
nand U410 (N_410,In_325,In_352);
or U411 (N_411,In_59,In_309);
nor U412 (N_412,In_208,In_170);
or U413 (N_413,In_266,In_362);
nor U414 (N_414,In_448,In_317);
or U415 (N_415,In_58,In_86);
or U416 (N_416,In_428,In_44);
nor U417 (N_417,In_156,In_490);
nand U418 (N_418,In_165,In_454);
nand U419 (N_419,In_77,In_232);
or U420 (N_420,In_137,In_255);
or U421 (N_421,In_137,In_13);
nand U422 (N_422,In_189,In_339);
nand U423 (N_423,In_64,In_359);
and U424 (N_424,In_27,In_361);
or U425 (N_425,In_229,In_2);
nand U426 (N_426,In_267,In_468);
nand U427 (N_427,In_54,In_272);
or U428 (N_428,In_72,In_476);
and U429 (N_429,In_18,In_27);
nor U430 (N_430,In_234,In_280);
or U431 (N_431,In_465,In_485);
nand U432 (N_432,In_144,In_323);
nand U433 (N_433,In_360,In_279);
and U434 (N_434,In_86,In_26);
or U435 (N_435,In_320,In_71);
and U436 (N_436,In_140,In_137);
or U437 (N_437,In_272,In_100);
nor U438 (N_438,In_244,In_246);
nor U439 (N_439,In_481,In_384);
nor U440 (N_440,In_43,In_149);
and U441 (N_441,In_359,In_190);
nor U442 (N_442,In_164,In_436);
and U443 (N_443,In_146,In_414);
nand U444 (N_444,In_388,In_180);
nor U445 (N_445,In_39,In_0);
or U446 (N_446,In_316,In_280);
and U447 (N_447,In_403,In_483);
and U448 (N_448,In_185,In_160);
nor U449 (N_449,In_479,In_149);
xnor U450 (N_450,In_171,In_328);
or U451 (N_451,In_225,In_154);
and U452 (N_452,In_66,In_403);
or U453 (N_453,In_454,In_412);
and U454 (N_454,In_433,In_356);
and U455 (N_455,In_377,In_368);
nand U456 (N_456,In_445,In_203);
or U457 (N_457,In_234,In_421);
nor U458 (N_458,In_309,In_348);
nand U459 (N_459,In_413,In_202);
and U460 (N_460,In_445,In_499);
nor U461 (N_461,In_342,In_322);
nand U462 (N_462,In_388,In_277);
xor U463 (N_463,In_438,In_482);
and U464 (N_464,In_161,In_212);
nand U465 (N_465,In_235,In_398);
nor U466 (N_466,In_462,In_260);
nor U467 (N_467,In_362,In_175);
and U468 (N_468,In_396,In_314);
nor U469 (N_469,In_362,In_182);
or U470 (N_470,In_275,In_101);
nor U471 (N_471,In_182,In_64);
and U472 (N_472,In_97,In_268);
or U473 (N_473,In_168,In_115);
nand U474 (N_474,In_166,In_480);
xnor U475 (N_475,In_475,In_113);
nand U476 (N_476,In_167,In_110);
or U477 (N_477,In_417,In_414);
nor U478 (N_478,In_419,In_405);
nand U479 (N_479,In_95,In_329);
and U480 (N_480,In_382,In_141);
nand U481 (N_481,In_110,In_334);
nand U482 (N_482,In_71,In_108);
nand U483 (N_483,In_0,In_341);
and U484 (N_484,In_114,In_34);
nor U485 (N_485,In_132,In_171);
xor U486 (N_486,In_44,In_119);
nor U487 (N_487,In_251,In_259);
nor U488 (N_488,In_490,In_298);
nand U489 (N_489,In_48,In_429);
nand U490 (N_490,In_244,In_222);
nor U491 (N_491,In_28,In_482);
nand U492 (N_492,In_402,In_347);
or U493 (N_493,In_426,In_67);
or U494 (N_494,In_130,In_464);
and U495 (N_495,In_244,In_162);
and U496 (N_496,In_492,In_405);
nand U497 (N_497,In_115,In_498);
and U498 (N_498,In_487,In_279);
nor U499 (N_499,In_405,In_312);
or U500 (N_500,In_318,In_29);
and U501 (N_501,In_373,In_240);
or U502 (N_502,In_6,In_316);
nor U503 (N_503,In_347,In_257);
or U504 (N_504,In_404,In_328);
nor U505 (N_505,In_163,In_118);
nor U506 (N_506,In_215,In_85);
and U507 (N_507,In_4,In_281);
nor U508 (N_508,In_99,In_277);
xnor U509 (N_509,In_273,In_292);
and U510 (N_510,In_231,In_213);
nand U511 (N_511,In_444,In_259);
or U512 (N_512,In_434,In_399);
nor U513 (N_513,In_17,In_431);
nor U514 (N_514,In_252,In_495);
nor U515 (N_515,In_166,In_308);
and U516 (N_516,In_124,In_344);
or U517 (N_517,In_31,In_401);
nor U518 (N_518,In_156,In_247);
nand U519 (N_519,In_361,In_150);
and U520 (N_520,In_95,In_173);
or U521 (N_521,In_50,In_76);
nand U522 (N_522,In_226,In_389);
or U523 (N_523,In_118,In_465);
and U524 (N_524,In_100,In_321);
and U525 (N_525,In_78,In_405);
or U526 (N_526,In_107,In_216);
or U527 (N_527,In_72,In_15);
and U528 (N_528,In_195,In_406);
nand U529 (N_529,In_143,In_211);
or U530 (N_530,In_332,In_365);
or U531 (N_531,In_284,In_370);
and U532 (N_532,In_88,In_362);
nor U533 (N_533,In_119,In_444);
nand U534 (N_534,In_437,In_422);
xnor U535 (N_535,In_129,In_435);
nand U536 (N_536,In_175,In_94);
nand U537 (N_537,In_176,In_66);
nor U538 (N_538,In_126,In_323);
or U539 (N_539,In_106,In_289);
nor U540 (N_540,In_418,In_415);
nor U541 (N_541,In_309,In_431);
and U542 (N_542,In_228,In_455);
nand U543 (N_543,In_120,In_208);
xnor U544 (N_544,In_454,In_247);
or U545 (N_545,In_226,In_127);
nor U546 (N_546,In_383,In_27);
or U547 (N_547,In_12,In_171);
and U548 (N_548,In_93,In_129);
nor U549 (N_549,In_339,In_29);
nand U550 (N_550,In_441,In_346);
and U551 (N_551,In_367,In_397);
nor U552 (N_552,In_3,In_401);
and U553 (N_553,In_426,In_86);
and U554 (N_554,In_366,In_451);
or U555 (N_555,In_322,In_260);
nor U556 (N_556,In_259,In_208);
nand U557 (N_557,In_204,In_182);
nor U558 (N_558,In_234,In_38);
and U559 (N_559,In_337,In_268);
nor U560 (N_560,In_255,In_53);
and U561 (N_561,In_433,In_264);
or U562 (N_562,In_174,In_357);
nor U563 (N_563,In_264,In_403);
or U564 (N_564,In_73,In_372);
nand U565 (N_565,In_16,In_51);
xnor U566 (N_566,In_235,In_489);
or U567 (N_567,In_27,In_181);
or U568 (N_568,In_298,In_250);
and U569 (N_569,In_189,In_440);
nand U570 (N_570,In_224,In_19);
or U571 (N_571,In_106,In_195);
xor U572 (N_572,In_320,In_307);
or U573 (N_573,In_136,In_413);
nand U574 (N_574,In_46,In_209);
or U575 (N_575,In_16,In_216);
or U576 (N_576,In_425,In_27);
nand U577 (N_577,In_129,In_252);
xnor U578 (N_578,In_255,In_233);
or U579 (N_579,In_14,In_90);
nor U580 (N_580,In_198,In_355);
nor U581 (N_581,In_235,In_332);
nand U582 (N_582,In_412,In_466);
nor U583 (N_583,In_322,In_281);
or U584 (N_584,In_303,In_81);
nor U585 (N_585,In_250,In_413);
or U586 (N_586,In_157,In_282);
and U587 (N_587,In_354,In_468);
or U588 (N_588,In_434,In_395);
and U589 (N_589,In_132,In_246);
and U590 (N_590,In_153,In_141);
nor U591 (N_591,In_250,In_56);
and U592 (N_592,In_396,In_230);
and U593 (N_593,In_223,In_141);
nor U594 (N_594,In_487,In_60);
nor U595 (N_595,In_377,In_175);
and U596 (N_596,In_38,In_337);
nor U597 (N_597,In_147,In_382);
and U598 (N_598,In_473,In_47);
and U599 (N_599,In_173,In_428);
or U600 (N_600,In_461,In_389);
nor U601 (N_601,In_25,In_346);
nand U602 (N_602,In_443,In_272);
and U603 (N_603,In_152,In_150);
and U604 (N_604,In_85,In_248);
nor U605 (N_605,In_492,In_265);
nand U606 (N_606,In_304,In_285);
xnor U607 (N_607,In_180,In_416);
nor U608 (N_608,In_409,In_175);
nor U609 (N_609,In_328,In_469);
nor U610 (N_610,In_446,In_454);
nor U611 (N_611,In_308,In_230);
and U612 (N_612,In_308,In_136);
or U613 (N_613,In_12,In_156);
or U614 (N_614,In_326,In_398);
or U615 (N_615,In_164,In_440);
or U616 (N_616,In_245,In_325);
and U617 (N_617,In_231,In_162);
or U618 (N_618,In_483,In_448);
xnor U619 (N_619,In_280,In_247);
and U620 (N_620,In_176,In_103);
nor U621 (N_621,In_351,In_432);
or U622 (N_622,In_455,In_12);
nand U623 (N_623,In_205,In_369);
nor U624 (N_624,In_382,In_345);
nand U625 (N_625,In_158,In_421);
or U626 (N_626,In_398,In_29);
or U627 (N_627,In_301,In_389);
and U628 (N_628,In_389,In_267);
nand U629 (N_629,In_496,In_263);
nor U630 (N_630,In_212,In_210);
nand U631 (N_631,In_440,In_79);
xnor U632 (N_632,In_330,In_452);
nand U633 (N_633,In_310,In_225);
nand U634 (N_634,In_200,In_469);
and U635 (N_635,In_273,In_306);
and U636 (N_636,In_70,In_334);
nand U637 (N_637,In_416,In_408);
or U638 (N_638,In_327,In_141);
and U639 (N_639,In_354,In_343);
nand U640 (N_640,In_266,In_25);
or U641 (N_641,In_37,In_339);
nor U642 (N_642,In_214,In_249);
xnor U643 (N_643,In_244,In_395);
nor U644 (N_644,In_353,In_42);
and U645 (N_645,In_302,In_340);
nand U646 (N_646,In_319,In_493);
nand U647 (N_647,In_146,In_346);
and U648 (N_648,In_472,In_361);
or U649 (N_649,In_350,In_141);
or U650 (N_650,In_321,In_372);
or U651 (N_651,In_83,In_321);
nor U652 (N_652,In_197,In_491);
and U653 (N_653,In_61,In_444);
or U654 (N_654,In_479,In_207);
nor U655 (N_655,In_369,In_164);
or U656 (N_656,In_130,In_427);
nand U657 (N_657,In_323,In_39);
and U658 (N_658,In_21,In_414);
and U659 (N_659,In_379,In_86);
nor U660 (N_660,In_484,In_184);
or U661 (N_661,In_486,In_485);
nand U662 (N_662,In_31,In_191);
or U663 (N_663,In_165,In_176);
and U664 (N_664,In_485,In_125);
or U665 (N_665,In_83,In_343);
and U666 (N_666,In_225,In_315);
nor U667 (N_667,In_279,In_168);
nor U668 (N_668,In_121,In_147);
nand U669 (N_669,In_192,In_59);
and U670 (N_670,In_143,In_188);
nor U671 (N_671,In_93,In_109);
nor U672 (N_672,In_167,In_6);
xor U673 (N_673,In_221,In_430);
nand U674 (N_674,In_431,In_73);
nor U675 (N_675,In_79,In_215);
nand U676 (N_676,In_389,In_183);
xor U677 (N_677,In_12,In_77);
nor U678 (N_678,In_454,In_283);
nor U679 (N_679,In_186,In_424);
or U680 (N_680,In_469,In_52);
and U681 (N_681,In_237,In_25);
xnor U682 (N_682,In_295,In_348);
nor U683 (N_683,In_45,In_444);
or U684 (N_684,In_425,In_441);
nor U685 (N_685,In_88,In_201);
and U686 (N_686,In_33,In_276);
xor U687 (N_687,In_371,In_365);
nand U688 (N_688,In_334,In_226);
nor U689 (N_689,In_454,In_292);
nand U690 (N_690,In_389,In_62);
and U691 (N_691,In_100,In_260);
or U692 (N_692,In_402,In_234);
and U693 (N_693,In_436,In_499);
nand U694 (N_694,In_293,In_24);
or U695 (N_695,In_361,In_220);
nand U696 (N_696,In_187,In_472);
or U697 (N_697,In_35,In_278);
nand U698 (N_698,In_258,In_63);
xnor U699 (N_699,In_436,In_196);
and U700 (N_700,In_172,In_296);
or U701 (N_701,In_376,In_25);
or U702 (N_702,In_57,In_373);
nand U703 (N_703,In_332,In_63);
or U704 (N_704,In_418,In_110);
or U705 (N_705,In_172,In_233);
or U706 (N_706,In_310,In_300);
xnor U707 (N_707,In_414,In_425);
nand U708 (N_708,In_325,In_101);
nor U709 (N_709,In_120,In_53);
nor U710 (N_710,In_36,In_322);
and U711 (N_711,In_75,In_210);
xor U712 (N_712,In_402,In_380);
or U713 (N_713,In_255,In_50);
nand U714 (N_714,In_50,In_71);
nand U715 (N_715,In_50,In_275);
nand U716 (N_716,In_334,In_431);
and U717 (N_717,In_291,In_410);
nor U718 (N_718,In_211,In_177);
nand U719 (N_719,In_137,In_87);
and U720 (N_720,In_18,In_79);
nand U721 (N_721,In_273,In_395);
nand U722 (N_722,In_121,In_324);
nand U723 (N_723,In_250,In_452);
nor U724 (N_724,In_416,In_31);
or U725 (N_725,In_147,In_324);
xnor U726 (N_726,In_391,In_137);
nor U727 (N_727,In_145,In_124);
nor U728 (N_728,In_330,In_180);
or U729 (N_729,In_215,In_490);
and U730 (N_730,In_416,In_480);
nor U731 (N_731,In_314,In_319);
xor U732 (N_732,In_202,In_404);
nor U733 (N_733,In_399,In_69);
nand U734 (N_734,In_122,In_475);
nor U735 (N_735,In_111,In_176);
and U736 (N_736,In_108,In_88);
nor U737 (N_737,In_208,In_10);
nand U738 (N_738,In_86,In_411);
nand U739 (N_739,In_167,In_20);
or U740 (N_740,In_145,In_192);
xor U741 (N_741,In_84,In_146);
and U742 (N_742,In_216,In_192);
or U743 (N_743,In_195,In_367);
xnor U744 (N_744,In_115,In_240);
or U745 (N_745,In_170,In_12);
or U746 (N_746,In_361,In_19);
nor U747 (N_747,In_131,In_182);
xnor U748 (N_748,In_77,In_277);
or U749 (N_749,In_479,In_391);
or U750 (N_750,In_178,In_151);
nand U751 (N_751,In_411,In_149);
and U752 (N_752,In_27,In_256);
or U753 (N_753,In_494,In_94);
and U754 (N_754,In_388,In_467);
or U755 (N_755,In_289,In_388);
xnor U756 (N_756,In_225,In_172);
nor U757 (N_757,In_18,In_114);
or U758 (N_758,In_68,In_231);
and U759 (N_759,In_165,In_142);
nor U760 (N_760,In_368,In_123);
or U761 (N_761,In_477,In_42);
and U762 (N_762,In_5,In_124);
xor U763 (N_763,In_271,In_49);
or U764 (N_764,In_354,In_48);
and U765 (N_765,In_285,In_300);
or U766 (N_766,In_273,In_389);
nand U767 (N_767,In_434,In_187);
and U768 (N_768,In_65,In_459);
and U769 (N_769,In_200,In_44);
and U770 (N_770,In_442,In_210);
and U771 (N_771,In_298,In_31);
or U772 (N_772,In_181,In_424);
nor U773 (N_773,In_110,In_344);
nand U774 (N_774,In_284,In_138);
nor U775 (N_775,In_78,In_134);
and U776 (N_776,In_100,In_38);
nand U777 (N_777,In_108,In_23);
nand U778 (N_778,In_144,In_33);
and U779 (N_779,In_456,In_116);
or U780 (N_780,In_370,In_394);
xnor U781 (N_781,In_117,In_445);
nor U782 (N_782,In_240,In_132);
nand U783 (N_783,In_109,In_385);
or U784 (N_784,In_348,In_66);
or U785 (N_785,In_202,In_299);
nor U786 (N_786,In_440,In_265);
nor U787 (N_787,In_207,In_377);
nand U788 (N_788,In_450,In_407);
nand U789 (N_789,In_292,In_246);
nand U790 (N_790,In_284,In_116);
nand U791 (N_791,In_135,In_354);
or U792 (N_792,In_297,In_235);
nor U793 (N_793,In_440,In_107);
nor U794 (N_794,In_392,In_119);
nor U795 (N_795,In_437,In_17);
or U796 (N_796,In_50,In_102);
or U797 (N_797,In_366,In_329);
nand U798 (N_798,In_165,In_146);
xor U799 (N_799,In_390,In_477);
xor U800 (N_800,In_254,In_459);
and U801 (N_801,In_284,In_243);
and U802 (N_802,In_331,In_499);
nand U803 (N_803,In_478,In_301);
xor U804 (N_804,In_473,In_130);
and U805 (N_805,In_324,In_32);
nand U806 (N_806,In_162,In_28);
or U807 (N_807,In_425,In_316);
xnor U808 (N_808,In_408,In_437);
and U809 (N_809,In_110,In_239);
and U810 (N_810,In_146,In_171);
xnor U811 (N_811,In_215,In_400);
and U812 (N_812,In_481,In_230);
and U813 (N_813,In_263,In_164);
nand U814 (N_814,In_138,In_261);
nor U815 (N_815,In_484,In_417);
and U816 (N_816,In_60,In_445);
nor U817 (N_817,In_10,In_73);
and U818 (N_818,In_433,In_210);
or U819 (N_819,In_212,In_479);
nand U820 (N_820,In_249,In_72);
nor U821 (N_821,In_456,In_495);
nor U822 (N_822,In_325,In_471);
nand U823 (N_823,In_420,In_421);
and U824 (N_824,In_63,In_268);
and U825 (N_825,In_335,In_170);
or U826 (N_826,In_327,In_170);
and U827 (N_827,In_240,In_154);
or U828 (N_828,In_69,In_298);
xor U829 (N_829,In_460,In_332);
nand U830 (N_830,In_38,In_355);
xor U831 (N_831,In_150,In_305);
nand U832 (N_832,In_127,In_439);
nand U833 (N_833,In_48,In_140);
or U834 (N_834,In_127,In_278);
nor U835 (N_835,In_13,In_454);
xor U836 (N_836,In_429,In_335);
and U837 (N_837,In_207,In_320);
nor U838 (N_838,In_48,In_153);
nor U839 (N_839,In_405,In_394);
nand U840 (N_840,In_32,In_122);
and U841 (N_841,In_72,In_46);
nor U842 (N_842,In_373,In_255);
nor U843 (N_843,In_380,In_356);
and U844 (N_844,In_221,In_156);
nand U845 (N_845,In_430,In_433);
and U846 (N_846,In_285,In_180);
and U847 (N_847,In_7,In_218);
and U848 (N_848,In_197,In_108);
nand U849 (N_849,In_319,In_183);
nor U850 (N_850,In_286,In_494);
or U851 (N_851,In_161,In_148);
xnor U852 (N_852,In_438,In_64);
nor U853 (N_853,In_403,In_430);
nand U854 (N_854,In_105,In_218);
or U855 (N_855,In_409,In_456);
nor U856 (N_856,In_187,In_124);
and U857 (N_857,In_311,In_262);
or U858 (N_858,In_143,In_244);
nand U859 (N_859,In_225,In_390);
and U860 (N_860,In_458,In_445);
or U861 (N_861,In_169,In_448);
or U862 (N_862,In_263,In_424);
or U863 (N_863,In_199,In_354);
nand U864 (N_864,In_372,In_382);
and U865 (N_865,In_348,In_294);
or U866 (N_866,In_77,In_476);
nand U867 (N_867,In_189,In_93);
nor U868 (N_868,In_15,In_125);
nor U869 (N_869,In_397,In_378);
or U870 (N_870,In_291,In_353);
or U871 (N_871,In_338,In_339);
nand U872 (N_872,In_434,In_39);
and U873 (N_873,In_252,In_71);
nor U874 (N_874,In_316,In_333);
nor U875 (N_875,In_259,In_65);
nand U876 (N_876,In_470,In_418);
or U877 (N_877,In_303,In_176);
xnor U878 (N_878,In_172,In_496);
nor U879 (N_879,In_6,In_163);
nor U880 (N_880,In_377,In_268);
and U881 (N_881,In_432,In_77);
or U882 (N_882,In_122,In_135);
or U883 (N_883,In_300,In_416);
nor U884 (N_884,In_352,In_97);
nand U885 (N_885,In_248,In_197);
and U886 (N_886,In_115,In_51);
and U887 (N_887,In_347,In_316);
nand U888 (N_888,In_436,In_344);
xnor U889 (N_889,In_485,In_116);
and U890 (N_890,In_47,In_327);
nand U891 (N_891,In_181,In_140);
nor U892 (N_892,In_201,In_340);
or U893 (N_893,In_417,In_496);
xor U894 (N_894,In_228,In_297);
nand U895 (N_895,In_261,In_1);
nor U896 (N_896,In_375,In_235);
and U897 (N_897,In_134,In_436);
nand U898 (N_898,In_351,In_422);
nor U899 (N_899,In_143,In_267);
and U900 (N_900,In_269,In_65);
and U901 (N_901,In_28,In_255);
and U902 (N_902,In_305,In_456);
xnor U903 (N_903,In_439,In_476);
nand U904 (N_904,In_224,In_9);
nand U905 (N_905,In_311,In_476);
nor U906 (N_906,In_127,In_173);
nand U907 (N_907,In_495,In_363);
nand U908 (N_908,In_136,In_429);
xnor U909 (N_909,In_375,In_97);
nor U910 (N_910,In_310,In_53);
nor U911 (N_911,In_139,In_351);
nand U912 (N_912,In_338,In_385);
nor U913 (N_913,In_410,In_294);
nor U914 (N_914,In_383,In_298);
or U915 (N_915,In_116,In_447);
nand U916 (N_916,In_303,In_100);
nor U917 (N_917,In_459,In_135);
and U918 (N_918,In_441,In_418);
nand U919 (N_919,In_315,In_179);
xnor U920 (N_920,In_409,In_279);
nand U921 (N_921,In_13,In_256);
and U922 (N_922,In_283,In_497);
nand U923 (N_923,In_376,In_493);
and U924 (N_924,In_120,In_224);
nor U925 (N_925,In_309,In_44);
nor U926 (N_926,In_471,In_182);
and U927 (N_927,In_343,In_184);
or U928 (N_928,In_446,In_220);
nand U929 (N_929,In_213,In_444);
or U930 (N_930,In_52,In_65);
nand U931 (N_931,In_332,In_396);
nor U932 (N_932,In_14,In_220);
nor U933 (N_933,In_26,In_114);
or U934 (N_934,In_372,In_298);
nand U935 (N_935,In_352,In_360);
and U936 (N_936,In_315,In_381);
or U937 (N_937,In_268,In_279);
nand U938 (N_938,In_468,In_87);
xor U939 (N_939,In_366,In_32);
nand U940 (N_940,In_135,In_304);
nand U941 (N_941,In_385,In_262);
xnor U942 (N_942,In_314,In_84);
nand U943 (N_943,In_21,In_224);
xnor U944 (N_944,In_66,In_350);
nand U945 (N_945,In_42,In_407);
and U946 (N_946,In_66,In_21);
and U947 (N_947,In_102,In_279);
nand U948 (N_948,In_419,In_287);
nor U949 (N_949,In_449,In_143);
nor U950 (N_950,In_450,In_145);
or U951 (N_951,In_77,In_441);
nand U952 (N_952,In_64,In_71);
nor U953 (N_953,In_325,In_348);
nor U954 (N_954,In_40,In_407);
nor U955 (N_955,In_198,In_202);
and U956 (N_956,In_190,In_331);
nor U957 (N_957,In_344,In_155);
nand U958 (N_958,In_389,In_99);
and U959 (N_959,In_307,In_485);
nand U960 (N_960,In_258,In_16);
nand U961 (N_961,In_412,In_75);
and U962 (N_962,In_166,In_174);
nor U963 (N_963,In_147,In_99);
xor U964 (N_964,In_298,In_287);
and U965 (N_965,In_24,In_218);
or U966 (N_966,In_235,In_152);
or U967 (N_967,In_311,In_434);
nand U968 (N_968,In_60,In_281);
or U969 (N_969,In_265,In_143);
or U970 (N_970,In_168,In_426);
or U971 (N_971,In_2,In_236);
nor U972 (N_972,In_280,In_112);
nand U973 (N_973,In_292,In_465);
xnor U974 (N_974,In_93,In_403);
nand U975 (N_975,In_293,In_424);
or U976 (N_976,In_307,In_222);
or U977 (N_977,In_35,In_141);
nand U978 (N_978,In_59,In_139);
nand U979 (N_979,In_22,In_452);
and U980 (N_980,In_363,In_199);
and U981 (N_981,In_480,In_486);
xnor U982 (N_982,In_380,In_413);
xnor U983 (N_983,In_347,In_9);
nor U984 (N_984,In_121,In_379);
nor U985 (N_985,In_136,In_491);
and U986 (N_986,In_61,In_120);
and U987 (N_987,In_10,In_480);
or U988 (N_988,In_328,In_87);
nor U989 (N_989,In_338,In_204);
nor U990 (N_990,In_282,In_38);
or U991 (N_991,In_470,In_407);
and U992 (N_992,In_130,In_304);
or U993 (N_993,In_28,In_498);
and U994 (N_994,In_418,In_48);
nor U995 (N_995,In_96,In_322);
nand U996 (N_996,In_482,In_66);
nand U997 (N_997,In_484,In_451);
nor U998 (N_998,In_396,In_152);
or U999 (N_999,In_203,In_202);
nor U1000 (N_1000,N_201,N_632);
xor U1001 (N_1001,N_797,N_572);
and U1002 (N_1002,N_492,N_153);
nand U1003 (N_1003,N_991,N_329);
xor U1004 (N_1004,N_152,N_868);
and U1005 (N_1005,N_178,N_699);
or U1006 (N_1006,N_247,N_530);
xor U1007 (N_1007,N_902,N_437);
and U1008 (N_1008,N_385,N_396);
xor U1009 (N_1009,N_583,N_562);
nor U1010 (N_1010,N_244,N_468);
nand U1011 (N_1011,N_367,N_341);
nand U1012 (N_1012,N_159,N_491);
or U1013 (N_1013,N_208,N_581);
xnor U1014 (N_1014,N_865,N_218);
xnor U1015 (N_1015,N_554,N_604);
nor U1016 (N_1016,N_227,N_771);
nand U1017 (N_1017,N_648,N_23);
xnor U1018 (N_1018,N_597,N_843);
xor U1019 (N_1019,N_977,N_4);
nor U1020 (N_1020,N_747,N_743);
xnor U1021 (N_1021,N_140,N_413);
or U1022 (N_1022,N_296,N_688);
nand U1023 (N_1023,N_525,N_904);
and U1024 (N_1024,N_948,N_175);
or U1025 (N_1025,N_284,N_974);
nor U1026 (N_1026,N_123,N_461);
xnor U1027 (N_1027,N_307,N_231);
xor U1028 (N_1028,N_476,N_148);
nand U1029 (N_1029,N_186,N_196);
xor U1030 (N_1030,N_533,N_886);
nor U1031 (N_1031,N_466,N_749);
nor U1032 (N_1032,N_858,N_852);
or U1033 (N_1033,N_363,N_757);
nor U1034 (N_1034,N_862,N_481);
nor U1035 (N_1035,N_933,N_680);
and U1036 (N_1036,N_518,N_839);
and U1037 (N_1037,N_378,N_42);
or U1038 (N_1038,N_573,N_734);
nor U1039 (N_1039,N_718,N_350);
nand U1040 (N_1040,N_596,N_156);
xor U1041 (N_1041,N_469,N_428);
nand U1042 (N_1042,N_854,N_857);
nor U1043 (N_1043,N_311,N_15);
and U1044 (N_1044,N_789,N_48);
and U1045 (N_1045,N_549,N_76);
and U1046 (N_1046,N_65,N_470);
nand U1047 (N_1047,N_220,N_906);
xnor U1048 (N_1048,N_932,N_464);
or U1049 (N_1049,N_801,N_912);
or U1050 (N_1050,N_856,N_911);
nand U1051 (N_1051,N_520,N_927);
and U1052 (N_1052,N_373,N_321);
nor U1053 (N_1053,N_835,N_986);
or U1054 (N_1054,N_303,N_937);
xnor U1055 (N_1055,N_391,N_769);
nor U1056 (N_1056,N_668,N_931);
or U1057 (N_1057,N_57,N_582);
nand U1058 (N_1058,N_654,N_869);
nand U1059 (N_1059,N_664,N_47);
nand U1060 (N_1060,N_5,N_655);
or U1061 (N_1061,N_358,N_364);
or U1062 (N_1062,N_269,N_340);
nor U1063 (N_1063,N_593,N_704);
or U1064 (N_1064,N_922,N_901);
nor U1065 (N_1065,N_696,N_760);
and U1066 (N_1066,N_71,N_320);
nand U1067 (N_1067,N_864,N_874);
and U1068 (N_1068,N_619,N_56);
nor U1069 (N_1069,N_756,N_193);
or U1070 (N_1070,N_427,N_762);
nand U1071 (N_1071,N_863,N_434);
nand U1072 (N_1072,N_878,N_891);
nand U1073 (N_1073,N_577,N_3);
nor U1074 (N_1074,N_216,N_452);
nor U1075 (N_1075,N_449,N_925);
nand U1076 (N_1076,N_641,N_450);
xnor U1077 (N_1077,N_149,N_333);
nand U1078 (N_1078,N_982,N_81);
or U1079 (N_1079,N_954,N_649);
nor U1080 (N_1080,N_214,N_314);
or U1081 (N_1081,N_574,N_431);
nand U1082 (N_1082,N_77,N_997);
or U1083 (N_1083,N_895,N_945);
and U1084 (N_1084,N_523,N_197);
nand U1085 (N_1085,N_145,N_844);
or U1086 (N_1086,N_213,N_657);
or U1087 (N_1087,N_758,N_325);
or U1088 (N_1088,N_827,N_104);
and U1089 (N_1089,N_976,N_301);
or U1090 (N_1090,N_16,N_894);
nor U1091 (N_1091,N_989,N_105);
nand U1092 (N_1092,N_184,N_690);
nand U1093 (N_1093,N_800,N_158);
or U1094 (N_1094,N_753,N_386);
and U1095 (N_1095,N_570,N_488);
and U1096 (N_1096,N_403,N_274);
and U1097 (N_1097,N_354,N_271);
xor U1098 (N_1098,N_224,N_280);
xnor U1099 (N_1099,N_84,N_513);
or U1100 (N_1100,N_971,N_832);
nor U1101 (N_1101,N_348,N_448);
and U1102 (N_1102,N_88,N_887);
xnor U1103 (N_1103,N_144,N_293);
nor U1104 (N_1104,N_667,N_262);
or U1105 (N_1105,N_546,N_605);
or U1106 (N_1106,N_748,N_475);
or U1107 (N_1107,N_251,N_795);
or U1108 (N_1108,N_265,N_405);
and U1109 (N_1109,N_783,N_478);
or U1110 (N_1110,N_558,N_327);
nand U1111 (N_1111,N_205,N_623);
nand U1112 (N_1112,N_509,N_560);
and U1113 (N_1113,N_728,N_715);
and U1114 (N_1114,N_836,N_256);
nand U1115 (N_1115,N_259,N_199);
or U1116 (N_1116,N_831,N_459);
nand U1117 (N_1117,N_228,N_133);
or U1118 (N_1118,N_91,N_784);
nand U1119 (N_1119,N_489,N_312);
nor U1120 (N_1120,N_684,N_441);
or U1121 (N_1121,N_99,N_647);
and U1122 (N_1122,N_221,N_585);
xor U1123 (N_1123,N_686,N_618);
and U1124 (N_1124,N_870,N_44);
xnor U1125 (N_1125,N_967,N_75);
and U1126 (N_1126,N_820,N_162);
and U1127 (N_1127,N_38,N_399);
nand U1128 (N_1128,N_934,N_115);
nand U1129 (N_1129,N_495,N_642);
and U1130 (N_1130,N_750,N_659);
or U1131 (N_1131,N_181,N_745);
and U1132 (N_1132,N_682,N_248);
or U1133 (N_1133,N_818,N_643);
and U1134 (N_1134,N_936,N_479);
nor U1135 (N_1135,N_587,N_418);
nor U1136 (N_1136,N_374,N_317);
and U1137 (N_1137,N_805,N_826);
nand U1138 (N_1138,N_442,N_74);
xnor U1139 (N_1139,N_482,N_200);
nand U1140 (N_1140,N_598,N_683);
and U1141 (N_1141,N_187,N_432);
nand U1142 (N_1142,N_167,N_362);
or U1143 (N_1143,N_407,N_236);
nor U1144 (N_1144,N_444,N_923);
nor U1145 (N_1145,N_130,N_781);
and U1146 (N_1146,N_589,N_798);
nor U1147 (N_1147,N_480,N_792);
xor U1148 (N_1148,N_628,N_959);
or U1149 (N_1149,N_599,N_981);
nor U1150 (N_1150,N_13,N_310);
nor U1151 (N_1151,N_487,N_393);
nor U1152 (N_1152,N_714,N_810);
and U1153 (N_1153,N_634,N_903);
nor U1154 (N_1154,N_171,N_86);
xnor U1155 (N_1155,N_586,N_440);
nor U1156 (N_1156,N_796,N_166);
and U1157 (N_1157,N_861,N_9);
or U1158 (N_1158,N_723,N_420);
and U1159 (N_1159,N_414,N_567);
or U1160 (N_1160,N_866,N_292);
or U1161 (N_1161,N_304,N_794);
and U1162 (N_1162,N_892,N_421);
or U1163 (N_1163,N_701,N_661);
or U1164 (N_1164,N_339,N_819);
nor U1165 (N_1165,N_958,N_551);
or U1166 (N_1166,N_893,N_838);
xor U1167 (N_1167,N_534,N_477);
or U1168 (N_1168,N_561,N_283);
nor U1169 (N_1169,N_883,N_559);
or U1170 (N_1170,N_608,N_964);
nor U1171 (N_1171,N_51,N_368);
nor U1172 (N_1172,N_451,N_834);
nand U1173 (N_1173,N_910,N_250);
or U1174 (N_1174,N_744,N_535);
nand U1175 (N_1175,N_650,N_968);
or U1176 (N_1176,N_300,N_527);
or U1177 (N_1177,N_31,N_966);
or U1178 (N_1178,N_621,N_277);
xnor U1179 (N_1179,N_95,N_316);
nand U1180 (N_1180,N_384,N_829);
and U1181 (N_1181,N_693,N_369);
and U1182 (N_1182,N_571,N_729);
or U1183 (N_1183,N_397,N_359);
nor U1184 (N_1184,N_89,N_849);
xnor U1185 (N_1185,N_249,N_241);
or U1186 (N_1186,N_299,N_266);
nand U1187 (N_1187,N_603,N_806);
nor U1188 (N_1188,N_970,N_962);
and U1189 (N_1189,N_500,N_370);
and U1190 (N_1190,N_49,N_980);
or U1191 (N_1191,N_322,N_681);
or U1192 (N_1192,N_467,N_692);
xor U1193 (N_1193,N_871,N_833);
xnor U1194 (N_1194,N_334,N_25);
and U1195 (N_1195,N_78,N_987);
nor U1196 (N_1196,N_411,N_889);
and U1197 (N_1197,N_978,N_345);
xnor U1198 (N_1198,N_872,N_935);
nand U1199 (N_1199,N_360,N_335);
or U1200 (N_1200,N_388,N_463);
and U1201 (N_1201,N_484,N_22);
or U1202 (N_1202,N_626,N_899);
or U1203 (N_1203,N_302,N_409);
and U1204 (N_1204,N_436,N_174);
or U1205 (N_1205,N_636,N_644);
nand U1206 (N_1206,N_999,N_281);
nand U1207 (N_1207,N_157,N_486);
nand U1208 (N_1208,N_782,N_267);
nor U1209 (N_1209,N_417,N_506);
nand U1210 (N_1210,N_183,N_288);
nand U1211 (N_1211,N_557,N_730);
and U1212 (N_1212,N_37,N_924);
xor U1213 (N_1213,N_263,N_32);
xnor U1214 (N_1214,N_122,N_136);
or U1215 (N_1215,N_888,N_775);
nand U1216 (N_1216,N_1,N_401);
or U1217 (N_1217,N_698,N_60);
nand U1218 (N_1218,N_627,N_20);
or U1219 (N_1219,N_677,N_629);
and U1220 (N_1220,N_791,N_652);
and U1221 (N_1221,N_483,N_2);
nand U1222 (N_1222,N_27,N_568);
nor U1223 (N_1223,N_639,N_947);
and U1224 (N_1224,N_779,N_995);
and U1225 (N_1225,N_656,N_415);
or U1226 (N_1226,N_64,N_100);
or U1227 (N_1227,N_702,N_837);
and U1228 (N_1228,N_988,N_939);
or U1229 (N_1229,N_209,N_344);
and U1230 (N_1230,N_768,N_717);
and U1231 (N_1231,N_103,N_875);
and U1232 (N_1232,N_705,N_96);
nand U1233 (N_1233,N_678,N_41);
and U1234 (N_1234,N_92,N_809);
and U1235 (N_1235,N_382,N_462);
and U1236 (N_1236,N_703,N_860);
nor U1237 (N_1237,N_445,N_965);
and U1238 (N_1238,N_98,N_788);
nand U1239 (N_1239,N_548,N_337);
nor U1240 (N_1240,N_46,N_419);
or U1241 (N_1241,N_324,N_503);
or U1242 (N_1242,N_859,N_944);
nor U1243 (N_1243,N_80,N_816);
or U1244 (N_1244,N_458,N_297);
nand U1245 (N_1245,N_349,N_108);
and U1246 (N_1246,N_102,N_55);
and U1247 (N_1247,N_54,N_777);
or U1248 (N_1248,N_165,N_700);
or U1249 (N_1249,N_106,N_447);
or U1250 (N_1250,N_261,N_135);
nand U1251 (N_1251,N_607,N_660);
or U1252 (N_1252,N_695,N_517);
nand U1253 (N_1253,N_828,N_710);
nor U1254 (N_1254,N_614,N_356);
nand U1255 (N_1255,N_217,N_630);
nor U1256 (N_1256,N_516,N_651);
nand U1257 (N_1257,N_996,N_438);
nand U1258 (N_1258,N_640,N_510);
or U1259 (N_1259,N_433,N_291);
xnor U1260 (N_1260,N_815,N_169);
nand U1261 (N_1261,N_953,N_776);
and U1262 (N_1262,N_381,N_59);
and U1263 (N_1263,N_613,N_260);
nand U1264 (N_1264,N_882,N_232);
and U1265 (N_1265,N_876,N_772);
nor U1266 (N_1266,N_515,N_867);
nor U1267 (N_1267,N_87,N_514);
and U1268 (N_1268,N_594,N_375);
and U1269 (N_1269,N_52,N_817);
or U1270 (N_1270,N_270,N_624);
nor U1271 (N_1271,N_62,N_134);
or U1272 (N_1272,N_770,N_202);
and U1273 (N_1273,N_993,N_917);
and U1274 (N_1274,N_675,N_313);
xnor U1275 (N_1275,N_823,N_138);
nand U1276 (N_1276,N_785,N_215);
and U1277 (N_1277,N_40,N_410);
nor U1278 (N_1278,N_600,N_556);
nor U1279 (N_1279,N_132,N_58);
nor U1280 (N_1280,N_851,N_120);
nand U1281 (N_1281,N_207,N_955);
or U1282 (N_1282,N_204,N_473);
or U1283 (N_1283,N_740,N_595);
and U1284 (N_1284,N_383,N_279);
and U1285 (N_1285,N_620,N_82);
or U1286 (N_1286,N_246,N_918);
nand U1287 (N_1287,N_637,N_28);
nand U1288 (N_1288,N_786,N_371);
nor U1289 (N_1289,N_323,N_879);
and U1290 (N_1290,N_763,N_191);
and U1291 (N_1291,N_471,N_168);
nand U1292 (N_1292,N_505,N_143);
or U1293 (N_1293,N_332,N_720);
and U1294 (N_1294,N_315,N_956);
nand U1295 (N_1295,N_584,N_840);
nand U1296 (N_1296,N_422,N_146);
nand U1297 (N_1297,N_460,N_164);
or U1298 (N_1298,N_240,N_242);
and U1299 (N_1299,N_726,N_230);
and U1300 (N_1300,N_767,N_907);
nor U1301 (N_1301,N_180,N_873);
and U1302 (N_1302,N_545,N_353);
nand U1303 (N_1303,N_670,N_490);
nand U1304 (N_1304,N_137,N_497);
or U1305 (N_1305,N_716,N_646);
or U1306 (N_1306,N_243,N_550);
nor U1307 (N_1307,N_346,N_131);
nand U1308 (N_1308,N_493,N_252);
nand U1309 (N_1309,N_177,N_914);
or U1310 (N_1310,N_790,N_443);
and U1311 (N_1311,N_124,N_496);
nor U1312 (N_1312,N_128,N_163);
and U1313 (N_1313,N_524,N_521);
nor U1314 (N_1314,N_210,N_848);
nor U1315 (N_1315,N_0,N_590);
or U1316 (N_1316,N_119,N_273);
nand U1317 (N_1317,N_685,N_824);
and U1318 (N_1318,N_93,N_669);
or U1319 (N_1319,N_24,N_66);
xnor U1320 (N_1320,N_663,N_121);
nor U1321 (N_1321,N_983,N_116);
nand U1322 (N_1322,N_127,N_569);
nor U1323 (N_1323,N_766,N_635);
or U1324 (N_1324,N_107,N_541);
nor U1325 (N_1325,N_219,N_278);
and U1326 (N_1326,N_921,N_542);
nor U1327 (N_1327,N_812,N_814);
and U1328 (N_1328,N_674,N_564);
nor U1329 (N_1329,N_606,N_926);
or U1330 (N_1330,N_7,N_176);
nand U1331 (N_1331,N_532,N_6);
nand U1332 (N_1332,N_206,N_161);
and U1333 (N_1333,N_531,N_426);
nand U1334 (N_1334,N_402,N_969);
or U1335 (N_1335,N_203,N_408);
and U1336 (N_1336,N_170,N_578);
and U1337 (N_1337,N_793,N_537);
or U1338 (N_1338,N_712,N_807);
and U1339 (N_1339,N_960,N_735);
or U1340 (N_1340,N_973,N_616);
nor U1341 (N_1341,N_755,N_539);
nand U1342 (N_1342,N_985,N_845);
or U1343 (N_1343,N_658,N_631);
xor U1344 (N_1344,N_237,N_342);
or U1345 (N_1345,N_392,N_97);
nor U1346 (N_1346,N_689,N_366);
or U1347 (N_1347,N_276,N_881);
and U1348 (N_1348,N_679,N_282);
xnor U1349 (N_1349,N_275,N_190);
nor U1350 (N_1350,N_225,N_14);
or U1351 (N_1351,N_326,N_129);
and U1352 (N_1352,N_540,N_802);
nor U1353 (N_1353,N_406,N_429);
and U1354 (N_1354,N_672,N_709);
nor U1355 (N_1355,N_526,N_940);
nor U1356 (N_1356,N_351,N_258);
nand U1357 (N_1357,N_11,N_994);
or U1358 (N_1358,N_439,N_555);
nand U1359 (N_1359,N_395,N_900);
and U1360 (N_1360,N_853,N_938);
nand U1361 (N_1361,N_151,N_253);
nand U1362 (N_1362,N_697,N_719);
nor U1363 (N_1363,N_830,N_61);
nand U1364 (N_1364,N_736,N_376);
xnor U1365 (N_1365,N_591,N_412);
nand U1366 (N_1366,N_12,N_821);
nor U1367 (N_1367,N_622,N_17);
nand U1368 (N_1368,N_264,N_69);
xnor U1369 (N_1369,N_233,N_125);
or U1370 (N_1370,N_453,N_528);
nand U1371 (N_1371,N_379,N_19);
xnor U1372 (N_1372,N_502,N_942);
and U1373 (N_1373,N_909,N_754);
or U1374 (N_1374,N_160,N_880);
or U1375 (N_1375,N_961,N_485);
or U1376 (N_1376,N_179,N_239);
nand U1377 (N_1377,N_309,N_285);
nand U1378 (N_1378,N_673,N_741);
and U1379 (N_1379,N_50,N_972);
and U1380 (N_1380,N_943,N_331);
nand U1381 (N_1381,N_272,N_941);
nand U1382 (N_1382,N_126,N_26);
nand U1383 (N_1383,N_885,N_67);
and U1384 (N_1384,N_380,N_355);
nand U1385 (N_1385,N_289,N_377);
nor U1386 (N_1386,N_446,N_36);
and U1387 (N_1387,N_111,N_72);
nand U1388 (N_1388,N_198,N_457);
nand U1389 (N_1389,N_498,N_665);
and U1390 (N_1390,N_662,N_565);
and U1391 (N_1391,N_841,N_761);
or U1392 (N_1392,N_150,N_949);
or U1393 (N_1393,N_588,N_154);
and U1394 (N_1394,N_739,N_727);
and U1395 (N_1395,N_890,N_724);
nor U1396 (N_1396,N_139,N_294);
nand U1397 (N_1397,N_306,N_538);
nand U1398 (N_1398,N_601,N_390);
or U1399 (N_1399,N_950,N_638);
or U1400 (N_1400,N_387,N_575);
xnor U1401 (N_1401,N_235,N_822);
nor U1402 (N_1402,N_211,N_913);
and U1403 (N_1403,N_773,N_94);
nor U1404 (N_1404,N_617,N_430);
and U1405 (N_1405,N_552,N_255);
nor U1406 (N_1406,N_147,N_751);
nor U1407 (N_1407,N_666,N_915);
and U1408 (N_1408,N_963,N_990);
and U1409 (N_1409,N_508,N_268);
and U1410 (N_1410,N_29,N_361);
xnor U1411 (N_1411,N_691,N_511);
nand U1412 (N_1412,N_30,N_234);
nand U1413 (N_1413,N_298,N_21);
or U1414 (N_1414,N_855,N_499);
nand U1415 (N_1415,N_117,N_929);
nor U1416 (N_1416,N_172,N_615);
nor U1417 (N_1417,N_110,N_687);
nand U1418 (N_1418,N_877,N_580);
nand U1419 (N_1419,N_738,N_811);
or U1420 (N_1420,N_404,N_10);
or U1421 (N_1421,N_957,N_504);
and U1422 (N_1422,N_713,N_522);
or U1423 (N_1423,N_394,N_916);
nor U1424 (N_1424,N_33,N_547);
or U1425 (N_1425,N_286,N_529);
and U1426 (N_1426,N_998,N_774);
nor U1427 (N_1427,N_155,N_194);
nand U1428 (N_1428,N_984,N_804);
nand U1429 (N_1429,N_79,N_287);
nor U1430 (N_1430,N_223,N_722);
nor U1431 (N_1431,N_842,N_290);
xnor U1432 (N_1432,N_389,N_212);
or U1433 (N_1433,N_141,N_787);
and U1434 (N_1434,N_456,N_778);
nor U1435 (N_1435,N_90,N_455);
and U1436 (N_1436,N_592,N_34);
nor U1437 (N_1437,N_711,N_229);
nand U1438 (N_1438,N_930,N_425);
or U1439 (N_1439,N_192,N_653);
nand U1440 (N_1440,N_63,N_733);
nand U1441 (N_1441,N_238,N_18);
or U1442 (N_1442,N_73,N_759);
xor U1443 (N_1443,N_318,N_611);
nor U1444 (N_1444,N_919,N_319);
and U1445 (N_1445,N_70,N_112);
or U1446 (N_1446,N_897,N_946);
nor U1447 (N_1447,N_563,N_898);
and U1448 (N_1448,N_928,N_905);
nand U1449 (N_1449,N_609,N_645);
and U1450 (N_1450,N_847,N_610);
and U1451 (N_1451,N_952,N_519);
or U1452 (N_1452,N_737,N_254);
xor U1453 (N_1453,N_908,N_707);
and U1454 (N_1454,N_109,N_222);
and U1455 (N_1455,N_780,N_39);
or U1456 (N_1456,N_764,N_708);
and U1457 (N_1457,N_896,N_752);
xor U1458 (N_1458,N_400,N_765);
xnor U1459 (N_1459,N_305,N_474);
and U1460 (N_1460,N_465,N_732);
and U1461 (N_1461,N_951,N_357);
or U1462 (N_1462,N_536,N_226);
nand U1463 (N_1463,N_189,N_694);
or U1464 (N_1464,N_182,N_343);
or U1465 (N_1465,N_338,N_336);
or U1466 (N_1466,N_35,N_633);
and U1467 (N_1467,N_566,N_101);
nor U1468 (N_1468,N_416,N_731);
nand U1469 (N_1469,N_543,N_113);
nand U1470 (N_1470,N_721,N_676);
and U1471 (N_1471,N_553,N_424);
xor U1472 (N_1472,N_142,N_706);
nand U1473 (N_1473,N_884,N_423);
nand U1474 (N_1474,N_602,N_53);
nor U1475 (N_1475,N_920,N_799);
and U1476 (N_1476,N_195,N_579);
xnor U1477 (N_1477,N_625,N_494);
xor U1478 (N_1478,N_257,N_671);
and U1479 (N_1479,N_114,N_813);
nor U1480 (N_1480,N_118,N_825);
nand U1481 (N_1481,N_85,N_83);
or U1482 (N_1482,N_328,N_742);
and U1483 (N_1483,N_472,N_846);
or U1484 (N_1484,N_512,N_746);
nor U1485 (N_1485,N_975,N_245);
nor U1486 (N_1486,N_372,N_576);
nor U1487 (N_1487,N_365,N_347);
or U1488 (N_1488,N_185,N_43);
or U1489 (N_1489,N_435,N_398);
nand U1490 (N_1490,N_308,N_352);
nor U1491 (N_1491,N_979,N_173);
nor U1492 (N_1492,N_454,N_501);
or U1493 (N_1493,N_188,N_612);
and U1494 (N_1494,N_330,N_803);
nor U1495 (N_1495,N_808,N_544);
nand U1496 (N_1496,N_295,N_68);
and U1497 (N_1497,N_8,N_725);
nand U1498 (N_1498,N_992,N_507);
nor U1499 (N_1499,N_45,N_850);
or U1500 (N_1500,N_943,N_993);
or U1501 (N_1501,N_989,N_970);
or U1502 (N_1502,N_856,N_186);
or U1503 (N_1503,N_928,N_532);
and U1504 (N_1504,N_189,N_973);
nor U1505 (N_1505,N_7,N_99);
and U1506 (N_1506,N_383,N_834);
nor U1507 (N_1507,N_613,N_540);
and U1508 (N_1508,N_375,N_977);
and U1509 (N_1509,N_355,N_206);
or U1510 (N_1510,N_855,N_750);
and U1511 (N_1511,N_466,N_790);
nand U1512 (N_1512,N_979,N_989);
or U1513 (N_1513,N_853,N_708);
nor U1514 (N_1514,N_434,N_502);
and U1515 (N_1515,N_879,N_468);
nor U1516 (N_1516,N_195,N_585);
and U1517 (N_1517,N_813,N_485);
nor U1518 (N_1518,N_138,N_462);
or U1519 (N_1519,N_32,N_852);
or U1520 (N_1520,N_658,N_780);
xnor U1521 (N_1521,N_297,N_521);
or U1522 (N_1522,N_361,N_264);
or U1523 (N_1523,N_749,N_776);
nor U1524 (N_1524,N_677,N_544);
and U1525 (N_1525,N_743,N_1);
and U1526 (N_1526,N_237,N_791);
nor U1527 (N_1527,N_483,N_92);
xnor U1528 (N_1528,N_913,N_173);
nand U1529 (N_1529,N_541,N_80);
or U1530 (N_1530,N_912,N_812);
or U1531 (N_1531,N_941,N_82);
and U1532 (N_1532,N_358,N_143);
or U1533 (N_1533,N_597,N_697);
nand U1534 (N_1534,N_726,N_466);
or U1535 (N_1535,N_177,N_54);
or U1536 (N_1536,N_290,N_503);
or U1537 (N_1537,N_347,N_669);
and U1538 (N_1538,N_319,N_17);
nand U1539 (N_1539,N_8,N_307);
or U1540 (N_1540,N_103,N_576);
and U1541 (N_1541,N_110,N_307);
and U1542 (N_1542,N_429,N_203);
nor U1543 (N_1543,N_797,N_528);
nor U1544 (N_1544,N_782,N_606);
and U1545 (N_1545,N_937,N_754);
nor U1546 (N_1546,N_389,N_136);
xor U1547 (N_1547,N_677,N_61);
xor U1548 (N_1548,N_543,N_438);
nand U1549 (N_1549,N_389,N_978);
nor U1550 (N_1550,N_926,N_388);
nor U1551 (N_1551,N_670,N_841);
or U1552 (N_1552,N_225,N_201);
nor U1553 (N_1553,N_80,N_469);
and U1554 (N_1554,N_987,N_492);
or U1555 (N_1555,N_188,N_20);
nand U1556 (N_1556,N_597,N_161);
or U1557 (N_1557,N_738,N_762);
and U1558 (N_1558,N_586,N_788);
xor U1559 (N_1559,N_979,N_604);
xor U1560 (N_1560,N_115,N_471);
xor U1561 (N_1561,N_444,N_942);
nand U1562 (N_1562,N_74,N_127);
nor U1563 (N_1563,N_113,N_261);
and U1564 (N_1564,N_144,N_214);
nand U1565 (N_1565,N_684,N_103);
nand U1566 (N_1566,N_962,N_248);
and U1567 (N_1567,N_254,N_849);
nand U1568 (N_1568,N_349,N_757);
xor U1569 (N_1569,N_147,N_151);
nand U1570 (N_1570,N_64,N_362);
nor U1571 (N_1571,N_970,N_263);
or U1572 (N_1572,N_927,N_820);
nor U1573 (N_1573,N_909,N_874);
and U1574 (N_1574,N_138,N_157);
nand U1575 (N_1575,N_535,N_465);
xnor U1576 (N_1576,N_166,N_189);
and U1577 (N_1577,N_190,N_289);
nor U1578 (N_1578,N_377,N_624);
nand U1579 (N_1579,N_945,N_909);
nor U1580 (N_1580,N_367,N_600);
or U1581 (N_1581,N_115,N_323);
nand U1582 (N_1582,N_925,N_300);
and U1583 (N_1583,N_19,N_848);
and U1584 (N_1584,N_483,N_343);
nand U1585 (N_1585,N_204,N_881);
nor U1586 (N_1586,N_184,N_818);
nand U1587 (N_1587,N_324,N_435);
or U1588 (N_1588,N_773,N_44);
or U1589 (N_1589,N_159,N_817);
nor U1590 (N_1590,N_366,N_487);
or U1591 (N_1591,N_220,N_216);
and U1592 (N_1592,N_663,N_72);
or U1593 (N_1593,N_358,N_195);
nor U1594 (N_1594,N_910,N_995);
nand U1595 (N_1595,N_666,N_876);
and U1596 (N_1596,N_9,N_160);
or U1597 (N_1597,N_762,N_977);
or U1598 (N_1598,N_493,N_621);
and U1599 (N_1599,N_328,N_262);
and U1600 (N_1600,N_992,N_572);
nor U1601 (N_1601,N_338,N_240);
or U1602 (N_1602,N_310,N_717);
or U1603 (N_1603,N_872,N_781);
nand U1604 (N_1604,N_521,N_652);
nor U1605 (N_1605,N_39,N_429);
and U1606 (N_1606,N_552,N_753);
nand U1607 (N_1607,N_600,N_526);
or U1608 (N_1608,N_597,N_333);
nor U1609 (N_1609,N_816,N_786);
xnor U1610 (N_1610,N_906,N_573);
or U1611 (N_1611,N_232,N_66);
and U1612 (N_1612,N_251,N_712);
nand U1613 (N_1613,N_768,N_329);
xor U1614 (N_1614,N_615,N_144);
and U1615 (N_1615,N_918,N_421);
and U1616 (N_1616,N_571,N_315);
nor U1617 (N_1617,N_837,N_902);
nor U1618 (N_1618,N_274,N_141);
xnor U1619 (N_1619,N_105,N_824);
nand U1620 (N_1620,N_879,N_118);
nand U1621 (N_1621,N_636,N_102);
nor U1622 (N_1622,N_437,N_777);
nor U1623 (N_1623,N_811,N_597);
and U1624 (N_1624,N_183,N_917);
and U1625 (N_1625,N_230,N_562);
nor U1626 (N_1626,N_235,N_352);
nand U1627 (N_1627,N_231,N_928);
and U1628 (N_1628,N_184,N_24);
nand U1629 (N_1629,N_687,N_618);
and U1630 (N_1630,N_296,N_911);
and U1631 (N_1631,N_672,N_840);
nor U1632 (N_1632,N_165,N_827);
nand U1633 (N_1633,N_223,N_262);
and U1634 (N_1634,N_236,N_617);
nor U1635 (N_1635,N_184,N_761);
or U1636 (N_1636,N_697,N_299);
nor U1637 (N_1637,N_325,N_289);
nor U1638 (N_1638,N_301,N_363);
nand U1639 (N_1639,N_18,N_391);
or U1640 (N_1640,N_429,N_658);
xor U1641 (N_1641,N_554,N_371);
or U1642 (N_1642,N_171,N_143);
nor U1643 (N_1643,N_63,N_257);
and U1644 (N_1644,N_299,N_7);
and U1645 (N_1645,N_391,N_875);
nand U1646 (N_1646,N_448,N_20);
xnor U1647 (N_1647,N_377,N_850);
or U1648 (N_1648,N_339,N_382);
nand U1649 (N_1649,N_690,N_170);
nor U1650 (N_1650,N_977,N_943);
or U1651 (N_1651,N_738,N_554);
nand U1652 (N_1652,N_229,N_237);
nor U1653 (N_1653,N_203,N_571);
or U1654 (N_1654,N_748,N_432);
or U1655 (N_1655,N_189,N_316);
or U1656 (N_1656,N_498,N_912);
and U1657 (N_1657,N_596,N_273);
nand U1658 (N_1658,N_369,N_595);
or U1659 (N_1659,N_345,N_395);
nand U1660 (N_1660,N_104,N_962);
or U1661 (N_1661,N_886,N_937);
and U1662 (N_1662,N_585,N_147);
or U1663 (N_1663,N_964,N_641);
or U1664 (N_1664,N_722,N_517);
and U1665 (N_1665,N_859,N_529);
and U1666 (N_1666,N_591,N_79);
and U1667 (N_1667,N_669,N_700);
and U1668 (N_1668,N_736,N_456);
nand U1669 (N_1669,N_252,N_791);
nor U1670 (N_1670,N_297,N_264);
xor U1671 (N_1671,N_878,N_184);
and U1672 (N_1672,N_245,N_940);
nor U1673 (N_1673,N_124,N_398);
and U1674 (N_1674,N_191,N_834);
nor U1675 (N_1675,N_748,N_375);
nor U1676 (N_1676,N_80,N_158);
nor U1677 (N_1677,N_675,N_797);
nand U1678 (N_1678,N_701,N_953);
nand U1679 (N_1679,N_906,N_726);
nand U1680 (N_1680,N_897,N_176);
nor U1681 (N_1681,N_131,N_488);
nand U1682 (N_1682,N_304,N_725);
nand U1683 (N_1683,N_576,N_512);
nand U1684 (N_1684,N_819,N_203);
nor U1685 (N_1685,N_626,N_615);
nand U1686 (N_1686,N_450,N_766);
or U1687 (N_1687,N_76,N_523);
nand U1688 (N_1688,N_334,N_257);
nand U1689 (N_1689,N_937,N_340);
nor U1690 (N_1690,N_297,N_454);
nand U1691 (N_1691,N_314,N_824);
nor U1692 (N_1692,N_463,N_293);
or U1693 (N_1693,N_370,N_566);
nor U1694 (N_1694,N_669,N_216);
nor U1695 (N_1695,N_380,N_162);
nor U1696 (N_1696,N_746,N_445);
and U1697 (N_1697,N_267,N_167);
and U1698 (N_1698,N_692,N_802);
nor U1699 (N_1699,N_40,N_259);
nand U1700 (N_1700,N_905,N_678);
and U1701 (N_1701,N_921,N_403);
nor U1702 (N_1702,N_63,N_159);
and U1703 (N_1703,N_43,N_464);
and U1704 (N_1704,N_911,N_849);
nand U1705 (N_1705,N_227,N_523);
or U1706 (N_1706,N_492,N_497);
and U1707 (N_1707,N_639,N_511);
nor U1708 (N_1708,N_161,N_704);
nor U1709 (N_1709,N_835,N_710);
or U1710 (N_1710,N_540,N_628);
nand U1711 (N_1711,N_520,N_157);
nand U1712 (N_1712,N_134,N_563);
nand U1713 (N_1713,N_217,N_188);
nand U1714 (N_1714,N_786,N_895);
nand U1715 (N_1715,N_322,N_116);
nor U1716 (N_1716,N_641,N_730);
or U1717 (N_1717,N_855,N_808);
nor U1718 (N_1718,N_820,N_12);
nand U1719 (N_1719,N_651,N_262);
and U1720 (N_1720,N_730,N_426);
and U1721 (N_1721,N_398,N_167);
nand U1722 (N_1722,N_806,N_751);
xor U1723 (N_1723,N_245,N_126);
and U1724 (N_1724,N_499,N_444);
xor U1725 (N_1725,N_815,N_554);
and U1726 (N_1726,N_741,N_492);
nand U1727 (N_1727,N_264,N_564);
nor U1728 (N_1728,N_508,N_984);
nand U1729 (N_1729,N_669,N_729);
nor U1730 (N_1730,N_225,N_614);
nor U1731 (N_1731,N_551,N_859);
nand U1732 (N_1732,N_668,N_459);
nor U1733 (N_1733,N_568,N_704);
and U1734 (N_1734,N_588,N_197);
nand U1735 (N_1735,N_96,N_240);
nor U1736 (N_1736,N_113,N_459);
xor U1737 (N_1737,N_851,N_511);
and U1738 (N_1738,N_887,N_253);
nor U1739 (N_1739,N_745,N_635);
xnor U1740 (N_1740,N_230,N_543);
xor U1741 (N_1741,N_929,N_49);
or U1742 (N_1742,N_414,N_63);
nor U1743 (N_1743,N_326,N_20);
and U1744 (N_1744,N_391,N_81);
nor U1745 (N_1745,N_876,N_644);
or U1746 (N_1746,N_389,N_429);
nor U1747 (N_1747,N_843,N_613);
or U1748 (N_1748,N_874,N_359);
and U1749 (N_1749,N_213,N_980);
xor U1750 (N_1750,N_616,N_169);
nor U1751 (N_1751,N_918,N_53);
nand U1752 (N_1752,N_424,N_8);
or U1753 (N_1753,N_363,N_455);
nor U1754 (N_1754,N_806,N_905);
or U1755 (N_1755,N_539,N_807);
or U1756 (N_1756,N_605,N_355);
nor U1757 (N_1757,N_772,N_950);
or U1758 (N_1758,N_979,N_397);
xor U1759 (N_1759,N_957,N_146);
or U1760 (N_1760,N_985,N_910);
nor U1761 (N_1761,N_883,N_614);
nand U1762 (N_1762,N_220,N_936);
nand U1763 (N_1763,N_901,N_939);
nor U1764 (N_1764,N_937,N_805);
and U1765 (N_1765,N_630,N_848);
nand U1766 (N_1766,N_613,N_179);
xor U1767 (N_1767,N_174,N_954);
nor U1768 (N_1768,N_392,N_877);
nor U1769 (N_1769,N_581,N_570);
and U1770 (N_1770,N_327,N_716);
nor U1771 (N_1771,N_387,N_253);
or U1772 (N_1772,N_332,N_683);
nor U1773 (N_1773,N_54,N_482);
or U1774 (N_1774,N_480,N_872);
nor U1775 (N_1775,N_92,N_341);
or U1776 (N_1776,N_126,N_268);
or U1777 (N_1777,N_678,N_752);
nor U1778 (N_1778,N_27,N_635);
nand U1779 (N_1779,N_389,N_525);
and U1780 (N_1780,N_843,N_326);
nand U1781 (N_1781,N_858,N_576);
or U1782 (N_1782,N_218,N_618);
nor U1783 (N_1783,N_182,N_753);
nor U1784 (N_1784,N_26,N_623);
nor U1785 (N_1785,N_680,N_148);
nand U1786 (N_1786,N_569,N_214);
nand U1787 (N_1787,N_209,N_874);
nor U1788 (N_1788,N_819,N_451);
and U1789 (N_1789,N_59,N_614);
nor U1790 (N_1790,N_678,N_994);
nor U1791 (N_1791,N_970,N_260);
nor U1792 (N_1792,N_131,N_336);
nor U1793 (N_1793,N_770,N_302);
or U1794 (N_1794,N_193,N_508);
nor U1795 (N_1795,N_87,N_829);
and U1796 (N_1796,N_916,N_424);
xnor U1797 (N_1797,N_400,N_978);
nor U1798 (N_1798,N_648,N_721);
or U1799 (N_1799,N_224,N_430);
nor U1800 (N_1800,N_276,N_972);
and U1801 (N_1801,N_496,N_662);
xor U1802 (N_1802,N_768,N_554);
and U1803 (N_1803,N_294,N_114);
or U1804 (N_1804,N_670,N_510);
nand U1805 (N_1805,N_26,N_227);
xor U1806 (N_1806,N_98,N_960);
xnor U1807 (N_1807,N_811,N_235);
xnor U1808 (N_1808,N_528,N_145);
nand U1809 (N_1809,N_601,N_629);
or U1810 (N_1810,N_727,N_960);
nand U1811 (N_1811,N_137,N_452);
nor U1812 (N_1812,N_279,N_714);
nand U1813 (N_1813,N_5,N_888);
and U1814 (N_1814,N_582,N_496);
or U1815 (N_1815,N_917,N_405);
and U1816 (N_1816,N_15,N_23);
nor U1817 (N_1817,N_190,N_728);
or U1818 (N_1818,N_457,N_847);
and U1819 (N_1819,N_532,N_373);
xor U1820 (N_1820,N_534,N_306);
or U1821 (N_1821,N_167,N_450);
nor U1822 (N_1822,N_819,N_895);
and U1823 (N_1823,N_233,N_993);
and U1824 (N_1824,N_830,N_574);
and U1825 (N_1825,N_515,N_562);
or U1826 (N_1826,N_641,N_260);
nor U1827 (N_1827,N_501,N_209);
nand U1828 (N_1828,N_818,N_984);
nand U1829 (N_1829,N_414,N_914);
or U1830 (N_1830,N_461,N_526);
nor U1831 (N_1831,N_765,N_47);
nand U1832 (N_1832,N_949,N_943);
and U1833 (N_1833,N_520,N_24);
nand U1834 (N_1834,N_852,N_959);
and U1835 (N_1835,N_507,N_420);
or U1836 (N_1836,N_989,N_336);
nor U1837 (N_1837,N_228,N_58);
and U1838 (N_1838,N_864,N_735);
xnor U1839 (N_1839,N_413,N_993);
and U1840 (N_1840,N_481,N_110);
and U1841 (N_1841,N_949,N_472);
nor U1842 (N_1842,N_876,N_824);
and U1843 (N_1843,N_616,N_40);
nand U1844 (N_1844,N_346,N_912);
and U1845 (N_1845,N_550,N_737);
and U1846 (N_1846,N_921,N_238);
nor U1847 (N_1847,N_105,N_355);
and U1848 (N_1848,N_824,N_539);
and U1849 (N_1849,N_951,N_858);
nor U1850 (N_1850,N_654,N_919);
or U1851 (N_1851,N_510,N_239);
or U1852 (N_1852,N_740,N_313);
or U1853 (N_1853,N_295,N_281);
nand U1854 (N_1854,N_133,N_376);
and U1855 (N_1855,N_172,N_255);
and U1856 (N_1856,N_141,N_618);
or U1857 (N_1857,N_748,N_275);
nor U1858 (N_1858,N_464,N_550);
nand U1859 (N_1859,N_911,N_764);
or U1860 (N_1860,N_95,N_913);
xor U1861 (N_1861,N_272,N_51);
or U1862 (N_1862,N_826,N_173);
or U1863 (N_1863,N_46,N_751);
nand U1864 (N_1864,N_34,N_978);
nor U1865 (N_1865,N_796,N_697);
and U1866 (N_1866,N_339,N_289);
or U1867 (N_1867,N_443,N_372);
and U1868 (N_1868,N_467,N_984);
or U1869 (N_1869,N_40,N_628);
and U1870 (N_1870,N_353,N_1);
or U1871 (N_1871,N_820,N_166);
nor U1872 (N_1872,N_832,N_786);
or U1873 (N_1873,N_32,N_227);
nor U1874 (N_1874,N_869,N_630);
or U1875 (N_1875,N_639,N_907);
or U1876 (N_1876,N_460,N_121);
nor U1877 (N_1877,N_32,N_64);
nor U1878 (N_1878,N_126,N_510);
and U1879 (N_1879,N_615,N_256);
or U1880 (N_1880,N_629,N_46);
nor U1881 (N_1881,N_647,N_64);
nor U1882 (N_1882,N_592,N_725);
and U1883 (N_1883,N_293,N_698);
and U1884 (N_1884,N_995,N_553);
nand U1885 (N_1885,N_99,N_442);
nor U1886 (N_1886,N_851,N_705);
nor U1887 (N_1887,N_972,N_827);
or U1888 (N_1888,N_429,N_830);
and U1889 (N_1889,N_222,N_296);
nand U1890 (N_1890,N_731,N_280);
nor U1891 (N_1891,N_510,N_411);
nand U1892 (N_1892,N_241,N_849);
nor U1893 (N_1893,N_563,N_769);
nand U1894 (N_1894,N_709,N_413);
nor U1895 (N_1895,N_355,N_640);
or U1896 (N_1896,N_419,N_898);
and U1897 (N_1897,N_790,N_782);
or U1898 (N_1898,N_721,N_347);
and U1899 (N_1899,N_47,N_276);
or U1900 (N_1900,N_155,N_405);
or U1901 (N_1901,N_504,N_862);
or U1902 (N_1902,N_808,N_0);
nand U1903 (N_1903,N_581,N_602);
and U1904 (N_1904,N_20,N_753);
nand U1905 (N_1905,N_747,N_6);
nand U1906 (N_1906,N_148,N_580);
or U1907 (N_1907,N_672,N_750);
or U1908 (N_1908,N_139,N_99);
nor U1909 (N_1909,N_490,N_663);
or U1910 (N_1910,N_529,N_785);
and U1911 (N_1911,N_164,N_990);
nor U1912 (N_1912,N_644,N_45);
and U1913 (N_1913,N_677,N_120);
and U1914 (N_1914,N_183,N_19);
and U1915 (N_1915,N_130,N_528);
and U1916 (N_1916,N_121,N_495);
and U1917 (N_1917,N_862,N_801);
nor U1918 (N_1918,N_848,N_701);
nor U1919 (N_1919,N_49,N_873);
nor U1920 (N_1920,N_898,N_76);
nand U1921 (N_1921,N_131,N_490);
nor U1922 (N_1922,N_460,N_399);
nand U1923 (N_1923,N_195,N_858);
and U1924 (N_1924,N_518,N_140);
nor U1925 (N_1925,N_146,N_547);
nor U1926 (N_1926,N_37,N_573);
nor U1927 (N_1927,N_228,N_476);
and U1928 (N_1928,N_274,N_426);
nand U1929 (N_1929,N_619,N_55);
or U1930 (N_1930,N_628,N_436);
or U1931 (N_1931,N_419,N_402);
nand U1932 (N_1932,N_377,N_460);
nor U1933 (N_1933,N_996,N_175);
and U1934 (N_1934,N_105,N_773);
and U1935 (N_1935,N_542,N_421);
nor U1936 (N_1936,N_461,N_43);
or U1937 (N_1937,N_371,N_47);
and U1938 (N_1938,N_658,N_550);
and U1939 (N_1939,N_404,N_196);
nor U1940 (N_1940,N_522,N_404);
nor U1941 (N_1941,N_479,N_174);
and U1942 (N_1942,N_52,N_839);
and U1943 (N_1943,N_650,N_335);
or U1944 (N_1944,N_449,N_83);
and U1945 (N_1945,N_45,N_499);
or U1946 (N_1946,N_728,N_835);
nor U1947 (N_1947,N_444,N_743);
and U1948 (N_1948,N_38,N_996);
nor U1949 (N_1949,N_163,N_538);
or U1950 (N_1950,N_287,N_149);
and U1951 (N_1951,N_668,N_427);
or U1952 (N_1952,N_805,N_134);
or U1953 (N_1953,N_517,N_172);
xnor U1954 (N_1954,N_675,N_780);
xor U1955 (N_1955,N_73,N_925);
or U1956 (N_1956,N_594,N_87);
nor U1957 (N_1957,N_983,N_618);
or U1958 (N_1958,N_583,N_636);
nand U1959 (N_1959,N_319,N_526);
nor U1960 (N_1960,N_652,N_380);
nand U1961 (N_1961,N_927,N_410);
xor U1962 (N_1962,N_501,N_392);
nor U1963 (N_1963,N_735,N_694);
and U1964 (N_1964,N_647,N_888);
and U1965 (N_1965,N_538,N_979);
nor U1966 (N_1966,N_792,N_518);
xnor U1967 (N_1967,N_25,N_267);
and U1968 (N_1968,N_581,N_390);
nor U1969 (N_1969,N_784,N_390);
and U1970 (N_1970,N_332,N_112);
xor U1971 (N_1971,N_18,N_432);
or U1972 (N_1972,N_729,N_719);
and U1973 (N_1973,N_128,N_235);
nor U1974 (N_1974,N_790,N_522);
nor U1975 (N_1975,N_674,N_986);
nor U1976 (N_1976,N_349,N_890);
xor U1977 (N_1977,N_813,N_272);
xor U1978 (N_1978,N_858,N_893);
and U1979 (N_1979,N_662,N_299);
nand U1980 (N_1980,N_485,N_814);
xnor U1981 (N_1981,N_823,N_371);
nand U1982 (N_1982,N_748,N_53);
nor U1983 (N_1983,N_286,N_940);
or U1984 (N_1984,N_340,N_399);
or U1985 (N_1985,N_58,N_467);
nor U1986 (N_1986,N_922,N_882);
nand U1987 (N_1987,N_209,N_84);
or U1988 (N_1988,N_623,N_955);
and U1989 (N_1989,N_130,N_934);
nor U1990 (N_1990,N_14,N_932);
xnor U1991 (N_1991,N_165,N_0);
or U1992 (N_1992,N_802,N_327);
xor U1993 (N_1993,N_182,N_659);
nor U1994 (N_1994,N_917,N_579);
and U1995 (N_1995,N_487,N_499);
or U1996 (N_1996,N_953,N_207);
xnor U1997 (N_1997,N_474,N_819);
and U1998 (N_1998,N_988,N_349);
nand U1999 (N_1999,N_227,N_350);
nand U2000 (N_2000,N_1295,N_1030);
or U2001 (N_2001,N_1644,N_1163);
or U2002 (N_2002,N_1015,N_1941);
nor U2003 (N_2003,N_1390,N_1619);
nor U2004 (N_2004,N_1288,N_1009);
nand U2005 (N_2005,N_1817,N_1429);
nand U2006 (N_2006,N_1379,N_1061);
or U2007 (N_2007,N_1326,N_1764);
nor U2008 (N_2008,N_1417,N_1242);
nand U2009 (N_2009,N_1062,N_1026);
nor U2010 (N_2010,N_1317,N_1907);
or U2011 (N_2011,N_1477,N_1999);
or U2012 (N_2012,N_1141,N_1189);
or U2013 (N_2013,N_1557,N_1331);
or U2014 (N_2014,N_1554,N_1636);
or U2015 (N_2015,N_1630,N_1475);
and U2016 (N_2016,N_1919,N_1432);
nor U2017 (N_2017,N_1830,N_1401);
or U2018 (N_2018,N_1212,N_1466);
or U2019 (N_2019,N_1013,N_1053);
xnor U2020 (N_2020,N_1089,N_1542);
and U2021 (N_2021,N_1765,N_1543);
and U2022 (N_2022,N_1454,N_1057);
xor U2023 (N_2023,N_1760,N_1665);
or U2024 (N_2024,N_1544,N_1837);
and U2025 (N_2025,N_1244,N_1794);
xnor U2026 (N_2026,N_1786,N_1305);
and U2027 (N_2027,N_1458,N_1949);
and U2028 (N_2028,N_1133,N_1670);
nand U2029 (N_2029,N_1376,N_1103);
or U2030 (N_2030,N_1097,N_1289);
or U2031 (N_2031,N_1732,N_1952);
xor U2032 (N_2032,N_1444,N_1783);
and U2033 (N_2033,N_1253,N_1613);
or U2034 (N_2034,N_1398,N_1781);
and U2035 (N_2035,N_1622,N_1523);
xnor U2036 (N_2036,N_1079,N_1286);
nor U2037 (N_2037,N_1790,N_1927);
nand U2038 (N_2038,N_1032,N_1007);
or U2039 (N_2039,N_1124,N_1671);
or U2040 (N_2040,N_1093,N_1452);
and U2041 (N_2041,N_1056,N_1277);
and U2042 (N_2042,N_1074,N_1058);
nand U2043 (N_2043,N_1176,N_1433);
nor U2044 (N_2044,N_1945,N_1535);
and U2045 (N_2045,N_1712,N_1036);
nand U2046 (N_2046,N_1096,N_1998);
nor U2047 (N_2047,N_1421,N_1939);
and U2048 (N_2048,N_1227,N_1263);
or U2049 (N_2049,N_1327,N_1348);
or U2050 (N_2050,N_1791,N_1268);
nor U2051 (N_2051,N_1855,N_1083);
or U2052 (N_2052,N_1947,N_1406);
xnor U2053 (N_2053,N_1891,N_1371);
nand U2054 (N_2054,N_1487,N_1434);
nand U2055 (N_2055,N_1601,N_1785);
and U2056 (N_2056,N_1462,N_1898);
nor U2057 (N_2057,N_1142,N_1967);
and U2058 (N_2058,N_1003,N_1109);
and U2059 (N_2059,N_1116,N_1873);
nor U2060 (N_2060,N_1615,N_1533);
nand U2061 (N_2061,N_1235,N_1372);
or U2062 (N_2062,N_1981,N_1121);
nand U2063 (N_2063,N_1568,N_1384);
nand U2064 (N_2064,N_1735,N_1408);
xor U2065 (N_2065,N_1006,N_1337);
and U2066 (N_2066,N_1809,N_1382);
nor U2067 (N_2067,N_1257,N_1662);
nand U2068 (N_2068,N_1208,N_1834);
and U2069 (N_2069,N_1004,N_1190);
nand U2070 (N_2070,N_1739,N_1342);
nand U2071 (N_2071,N_1883,N_1717);
nand U2072 (N_2072,N_1367,N_1266);
xor U2073 (N_2073,N_1740,N_1146);
or U2074 (N_2074,N_1890,N_1493);
and U2075 (N_2075,N_1234,N_1490);
and U2076 (N_2076,N_1815,N_1117);
nand U2077 (N_2077,N_1660,N_1343);
nand U2078 (N_2078,N_1931,N_1860);
or U2079 (N_2079,N_1932,N_1411);
or U2080 (N_2080,N_1370,N_1674);
nand U2081 (N_2081,N_1605,N_1221);
nor U2082 (N_2082,N_1249,N_1374);
and U2083 (N_2083,N_1726,N_1409);
or U2084 (N_2084,N_1905,N_1933);
and U2085 (N_2085,N_1233,N_1831);
and U2086 (N_2086,N_1736,N_1574);
or U2087 (N_2087,N_1780,N_1361);
xor U2088 (N_2088,N_1494,N_1778);
nand U2089 (N_2089,N_1969,N_1037);
and U2090 (N_2090,N_1697,N_1914);
or U2091 (N_2091,N_1561,N_1756);
and U2092 (N_2092,N_1196,N_1521);
or U2093 (N_2093,N_1456,N_1629);
or U2094 (N_2094,N_1415,N_1140);
or U2095 (N_2095,N_1170,N_1090);
nor U2096 (N_2096,N_1708,N_1526);
xnor U2097 (N_2097,N_1642,N_1306);
nor U2098 (N_2098,N_1298,N_1530);
nor U2099 (N_2099,N_1446,N_1813);
nand U2100 (N_2100,N_1795,N_1394);
nor U2101 (N_2101,N_1168,N_1645);
nand U2102 (N_2102,N_1843,N_1748);
nor U2103 (N_2103,N_1839,N_1151);
and U2104 (N_2104,N_1852,N_1256);
nand U2105 (N_2105,N_1631,N_1934);
and U2106 (N_2106,N_1112,N_1745);
and U2107 (N_2107,N_1024,N_1471);
and U2108 (N_2108,N_1937,N_1548);
or U2109 (N_2109,N_1144,N_1733);
or U2110 (N_2110,N_1159,N_1826);
or U2111 (N_2111,N_1413,N_1846);
and U2112 (N_2112,N_1049,N_1127);
and U2113 (N_2113,N_1495,N_1857);
and U2114 (N_2114,N_1624,N_1206);
and U2115 (N_2115,N_1796,N_1874);
nor U2116 (N_2116,N_1359,N_1237);
nor U2117 (N_2117,N_1023,N_1270);
nand U2118 (N_2118,N_1640,N_1747);
or U2119 (N_2119,N_1593,N_1333);
or U2120 (N_2120,N_1546,N_1005);
and U2121 (N_2121,N_1767,N_1822);
nand U2122 (N_2122,N_1279,N_1885);
nor U2123 (N_2123,N_1008,N_1910);
or U2124 (N_2124,N_1152,N_1291);
or U2125 (N_2125,N_1000,N_1325);
nor U2126 (N_2126,N_1391,N_1908);
nand U2127 (N_2127,N_1847,N_1243);
nor U2128 (N_2128,N_1590,N_1556);
nand U2129 (N_2129,N_1179,N_1913);
and U2130 (N_2130,N_1186,N_1070);
xnor U2131 (N_2131,N_1115,N_1858);
nor U2132 (N_2132,N_1532,N_1819);
nand U2133 (N_2133,N_1854,N_1978);
or U2134 (N_2134,N_1431,N_1191);
xnor U2135 (N_2135,N_1862,N_1218);
nor U2136 (N_2136,N_1380,N_1692);
and U2137 (N_2137,N_1650,N_1600);
xor U2138 (N_2138,N_1872,N_1626);
or U2139 (N_2139,N_1255,N_1617);
and U2140 (N_2140,N_1531,N_1924);
nor U2141 (N_2141,N_1805,N_1352);
or U2142 (N_2142,N_1609,N_1893);
nand U2143 (N_2143,N_1219,N_1559);
xor U2144 (N_2144,N_1536,N_1264);
nor U2145 (N_2145,N_1480,N_1051);
nor U2146 (N_2146,N_1287,N_1994);
and U2147 (N_2147,N_1293,N_1727);
nand U2148 (N_2148,N_1982,N_1566);
and U2149 (N_2149,N_1766,N_1016);
nand U2150 (N_2150,N_1020,N_1110);
or U2151 (N_2151,N_1679,N_1746);
nor U2152 (N_2152,N_1555,N_1154);
or U2153 (N_2153,N_1840,N_1467);
nand U2154 (N_2154,N_1938,N_1001);
nand U2155 (N_2155,N_1503,N_1158);
nor U2156 (N_2156,N_1285,N_1461);
or U2157 (N_2157,N_1699,N_1749);
and U2158 (N_2158,N_1841,N_1358);
nor U2159 (N_2159,N_1602,N_1684);
nor U2160 (N_2160,N_1131,N_1029);
or U2161 (N_2161,N_1076,N_1311);
nor U2162 (N_2162,N_1041,N_1492);
nand U2163 (N_2163,N_1845,N_1483);
or U2164 (N_2164,N_1213,N_1788);
or U2165 (N_2165,N_1563,N_1031);
nand U2166 (N_2166,N_1971,N_1060);
nand U2167 (N_2167,N_1887,N_1988);
nand U2168 (N_2168,N_1484,N_1018);
nand U2169 (N_2169,N_1725,N_1129);
and U2170 (N_2170,N_1851,N_1420);
nand U2171 (N_2171,N_1039,N_1412);
and U2172 (N_2172,N_1918,N_1375);
xnor U2173 (N_2173,N_1299,N_1976);
nor U2174 (N_2174,N_1632,N_1324);
nand U2175 (N_2175,N_1260,N_1996);
nand U2176 (N_2176,N_1405,N_1126);
nand U2177 (N_2177,N_1538,N_1486);
and U2178 (N_2178,N_1661,N_1312);
or U2179 (N_2179,N_1050,N_1455);
nand U2180 (N_2180,N_1332,N_1681);
nand U2181 (N_2181,N_1956,N_1214);
nor U2182 (N_2182,N_1201,N_1386);
nor U2183 (N_2183,N_1625,N_1782);
and U2184 (N_2184,N_1621,N_1957);
xnor U2185 (N_2185,N_1321,N_1125);
nand U2186 (N_2186,N_1750,N_1876);
nor U2187 (N_2187,N_1950,N_1596);
or U2188 (N_2188,N_1025,N_1118);
nand U2189 (N_2189,N_1022,N_1534);
or U2190 (N_2190,N_1868,N_1866);
and U2191 (N_2191,N_1155,N_1247);
and U2192 (N_2192,N_1936,N_1239);
nand U2193 (N_2193,N_1620,N_1067);
and U2194 (N_2194,N_1635,N_1842);
xor U2195 (N_2195,N_1357,N_1094);
or U2196 (N_2196,N_1687,N_1637);
nand U2197 (N_2197,N_1741,N_1071);
nand U2198 (N_2198,N_1985,N_1719);
nand U2199 (N_2199,N_1106,N_1187);
or U2200 (N_2200,N_1519,N_1731);
or U2201 (N_2201,N_1423,N_1283);
xnor U2202 (N_2202,N_1202,N_1280);
or U2203 (N_2203,N_1643,N_1803);
xor U2204 (N_2204,N_1442,N_1604);
nor U2205 (N_2205,N_1181,N_1368);
or U2206 (N_2206,N_1571,N_1930);
nand U2207 (N_2207,N_1792,N_1450);
and U2208 (N_2208,N_1870,N_1838);
nor U2209 (N_2209,N_1504,N_1236);
nor U2210 (N_2210,N_1799,N_1821);
and U2211 (N_2211,N_1459,N_1677);
or U2212 (N_2212,N_1111,N_1698);
nor U2213 (N_2213,N_1192,N_1329);
and U2214 (N_2214,N_1909,N_1722);
and U2215 (N_2215,N_1120,N_1652);
or U2216 (N_2216,N_1054,N_1364);
xor U2217 (N_2217,N_1979,N_1033);
nor U2218 (N_2218,N_1867,N_1658);
nand U2219 (N_2219,N_1258,N_1162);
nand U2220 (N_2220,N_1537,N_1232);
nor U2221 (N_2221,N_1506,N_1606);
or U2222 (N_2222,N_1246,N_1425);
or U2223 (N_2223,N_1577,N_1254);
nand U2224 (N_2224,N_1498,N_1438);
nor U2225 (N_2225,N_1355,N_1922);
or U2226 (N_2226,N_1528,N_1775);
nor U2227 (N_2227,N_1128,N_1203);
or U2228 (N_2228,N_1171,N_1638);
and U2229 (N_2229,N_1585,N_1426);
and U2230 (N_2230,N_1292,N_1850);
nor U2231 (N_2231,N_1964,N_1558);
nor U2232 (N_2232,N_1871,N_1634);
nor U2233 (N_2233,N_1685,N_1771);
nor U2234 (N_2234,N_1592,N_1248);
nand U2235 (N_2235,N_1511,N_1776);
or U2236 (N_2236,N_1073,N_1449);
and U2237 (N_2237,N_1149,N_1951);
and U2238 (N_2238,N_1586,N_1319);
and U2239 (N_2239,N_1104,N_1308);
and U2240 (N_2240,N_1579,N_1849);
nor U2241 (N_2241,N_1238,N_1385);
xor U2242 (N_2242,N_1896,N_1944);
nand U2243 (N_2243,N_1188,N_1989);
nand U2244 (N_2244,N_1307,N_1017);
nor U2245 (N_2245,N_1578,N_1935);
and U2246 (N_2246,N_1465,N_1844);
or U2247 (N_2247,N_1360,N_1728);
nor U2248 (N_2248,N_1512,N_1588);
nand U2249 (N_2249,N_1345,N_1993);
nor U2250 (N_2250,N_1430,N_1177);
nand U2251 (N_2251,N_1216,N_1628);
nor U2252 (N_2252,N_1474,N_1276);
or U2253 (N_2253,N_1925,N_1055);
nand U2254 (N_2254,N_1567,N_1565);
and U2255 (N_2255,N_1804,N_1770);
nor U2256 (N_2256,N_1199,N_1589);
nor U2257 (N_2257,N_1928,N_1545);
nand U2258 (N_2258,N_1403,N_1655);
nand U2259 (N_2259,N_1410,N_1920);
and U2260 (N_2260,N_1524,N_1965);
xor U2261 (N_2261,N_1829,N_1211);
nor U2262 (N_2262,N_1422,N_1877);
or U2263 (N_2263,N_1691,N_1863);
nand U2264 (N_2264,N_1614,N_1878);
nor U2265 (N_2265,N_1014,N_1737);
xor U2266 (N_2266,N_1427,N_1836);
xnor U2267 (N_2267,N_1608,N_1448);
xor U2268 (N_2268,N_1711,N_1833);
nor U2269 (N_2269,N_1975,N_1706);
nor U2270 (N_2270,N_1653,N_1469);
or U2271 (N_2271,N_1942,N_1916);
nand U2272 (N_2272,N_1646,N_1575);
and U2273 (N_2273,N_1397,N_1986);
nand U2274 (N_2274,N_1100,N_1439);
xnor U2275 (N_2275,N_1482,N_1353);
nand U2276 (N_2276,N_1603,N_1987);
and U2277 (N_2277,N_1716,N_1564);
or U2278 (N_2278,N_1570,N_1085);
and U2279 (N_2279,N_1832,N_1540);
and U2280 (N_2280,N_1225,N_1378);
or U2281 (N_2281,N_1940,N_1095);
nor U2282 (N_2282,N_1848,N_1294);
nor U2283 (N_2283,N_1946,N_1798);
or U2284 (N_2284,N_1065,N_1241);
nand U2285 (N_2285,N_1599,N_1172);
or U2286 (N_2286,N_1997,N_1668);
nor U2287 (N_2287,N_1086,N_1729);
xnor U2288 (N_2288,N_1879,N_1262);
nor U2289 (N_2289,N_1088,N_1441);
and U2290 (N_2290,N_1539,N_1572);
nand U2291 (N_2291,N_1806,N_1991);
or U2292 (N_2292,N_1198,N_1515);
nand U2293 (N_2293,N_1346,N_1954);
and U2294 (N_2294,N_1688,N_1028);
nor U2295 (N_2295,N_1560,N_1464);
nor U2296 (N_2296,N_1335,N_1436);
xor U2297 (N_2297,N_1700,N_1451);
and U2298 (N_2298,N_1251,N_1812);
nand U2299 (N_2299,N_1396,N_1105);
and U2300 (N_2300,N_1087,N_1864);
xor U2301 (N_2301,N_1911,N_1948);
nor U2302 (N_2302,N_1267,N_1774);
or U2303 (N_2303,N_1281,N_1800);
nor U2304 (N_2304,N_1414,N_1044);
nor U2305 (N_2305,N_1443,N_1607);
or U2306 (N_2306,N_1892,N_1479);
xnor U2307 (N_2307,N_1906,N_1362);
and U2308 (N_2308,N_1943,N_1808);
nand U2309 (N_2309,N_1481,N_1721);
nor U2310 (N_2310,N_1310,N_1145);
or U2311 (N_2311,N_1713,N_1252);
nor U2312 (N_2312,N_1974,N_1921);
nor U2313 (N_2313,N_1389,N_1334);
and U2314 (N_2314,N_1753,N_1673);
nor U2315 (N_2315,N_1040,N_1823);
nor U2316 (N_2316,N_1816,N_1797);
nor U2317 (N_2317,N_1064,N_1897);
or U2318 (N_2318,N_1156,N_1597);
or U2319 (N_2319,N_1047,N_1224);
nand U2320 (N_2320,N_1768,N_1350);
and U2321 (N_2321,N_1875,N_1761);
nor U2322 (N_2322,N_1404,N_1099);
nand U2323 (N_2323,N_1138,N_1365);
nand U2324 (N_2324,N_1340,N_1549);
xor U2325 (N_2325,N_1820,N_1669);
nand U2326 (N_2326,N_1314,N_1101);
nor U2327 (N_2327,N_1166,N_1595);
nand U2328 (N_2328,N_1884,N_1393);
and U2329 (N_2329,N_1447,N_1207);
nor U2330 (N_2330,N_1139,N_1656);
nand U2331 (N_2331,N_1730,N_1010);
nand U2332 (N_2332,N_1265,N_1338);
nand U2333 (N_2333,N_1894,N_1983);
or U2334 (N_2334,N_1197,N_1366);
and U2335 (N_2335,N_1966,N_1758);
or U2336 (N_2336,N_1869,N_1261);
nand U2337 (N_2337,N_1541,N_1777);
or U2338 (N_2338,N_1807,N_1284);
and U2339 (N_2339,N_1694,N_1082);
xor U2340 (N_2340,N_1108,N_1363);
and U2341 (N_2341,N_1977,N_1463);
or U2342 (N_2342,N_1175,N_1183);
nor U2343 (N_2343,N_1381,N_1714);
xor U2344 (N_2344,N_1701,N_1742);
nand U2345 (N_2345,N_1369,N_1383);
nor U2346 (N_2346,N_1724,N_1297);
and U2347 (N_2347,N_1980,N_1702);
or U2348 (N_2348,N_1553,N_1787);
nor U2349 (N_2349,N_1217,N_1328);
and U2350 (N_2350,N_1814,N_1686);
nand U2351 (N_2351,N_1098,N_1339);
or U2352 (N_2352,N_1901,N_1587);
nor U2353 (N_2353,N_1437,N_1923);
and U2354 (N_2354,N_1160,N_1757);
xor U2355 (N_2355,N_1204,N_1984);
nand U2356 (N_2356,N_1042,N_1223);
nor U2357 (N_2357,N_1195,N_1752);
nor U2358 (N_2358,N_1762,N_1066);
and U2359 (N_2359,N_1418,N_1580);
xnor U2360 (N_2360,N_1229,N_1509);
and U2361 (N_2361,N_1323,N_1550);
or U2362 (N_2362,N_1205,N_1759);
nor U2363 (N_2363,N_1419,N_1853);
or U2364 (N_2364,N_1081,N_1672);
or U2365 (N_2365,N_1667,N_1402);
nand U2366 (N_2366,N_1573,N_1865);
nor U2367 (N_2367,N_1802,N_1569);
nor U2368 (N_2368,N_1959,N_1773);
and U2369 (N_2369,N_1835,N_1228);
xor U2370 (N_2370,N_1072,N_1598);
or U2371 (N_2371,N_1926,N_1178);
or U2372 (N_2372,N_1510,N_1610);
or U2373 (N_2373,N_1710,N_1581);
or U2374 (N_2374,N_1522,N_1990);
nor U2375 (N_2375,N_1027,N_1651);
nand U2376 (N_2376,N_1755,N_1676);
nand U2377 (N_2377,N_1612,N_1882);
or U2378 (N_2378,N_1972,N_1904);
nand U2379 (N_2379,N_1069,N_1903);
nor U2380 (N_2380,N_1659,N_1738);
nand U2381 (N_2381,N_1290,N_1516);
nand U2382 (N_2382,N_1473,N_1084);
xor U2383 (N_2383,N_1157,N_1301);
nand U2384 (N_2384,N_1318,N_1011);
nand U2385 (N_2385,N_1518,N_1859);
xnor U2386 (N_2386,N_1664,N_1052);
and U2387 (N_2387,N_1351,N_1502);
nand U2388 (N_2388,N_1395,N_1165);
or U2389 (N_2389,N_1185,N_1038);
nand U2390 (N_2390,N_1703,N_1616);
nand U2391 (N_2391,N_1784,N_1690);
or U2392 (N_2392,N_1618,N_1696);
nand U2393 (N_2393,N_1330,N_1682);
and U2394 (N_2394,N_1693,N_1271);
nor U2395 (N_2395,N_1012,N_1476);
nor U2396 (N_2396,N_1824,N_1445);
or U2397 (N_2397,N_1961,N_1496);
and U2398 (N_2398,N_1886,N_1046);
or U2399 (N_2399,N_1460,N_1734);
or U2400 (N_2400,N_1272,N_1695);
or U2401 (N_2401,N_1303,N_1316);
xor U2402 (N_2402,N_1387,N_1043);
xor U2403 (N_2403,N_1440,N_1880);
nor U2404 (N_2404,N_1917,N_1705);
xor U2405 (N_2405,N_1153,N_1527);
nand U2406 (N_2406,N_1763,N_1407);
or U2407 (N_2407,N_1611,N_1416);
or U2408 (N_2408,N_1130,N_1551);
nor U2409 (N_2409,N_1889,N_1173);
xnor U2410 (N_2410,N_1349,N_1341);
or U2411 (N_2411,N_1274,N_1915);
nor U2412 (N_2412,N_1769,N_1373);
and U2413 (N_2413,N_1507,N_1594);
and U2414 (N_2414,N_1059,N_1754);
nor U2415 (N_2415,N_1226,N_1513);
and U2416 (N_2416,N_1275,N_1900);
or U2417 (N_2417,N_1282,N_1304);
xnor U2418 (N_2418,N_1744,N_1075);
and U2419 (N_2419,N_1184,N_1514);
xor U2420 (N_2420,N_1743,N_1751);
nand U2421 (N_2421,N_1488,N_1584);
nor U2422 (N_2422,N_1347,N_1167);
nor U2423 (N_2423,N_1666,N_1478);
and U2424 (N_2424,N_1718,N_1623);
nand U2425 (N_2425,N_1973,N_1472);
and U2426 (N_2426,N_1428,N_1517);
nor U2427 (N_2427,N_1077,N_1647);
nand U2428 (N_2428,N_1035,N_1680);
and U2429 (N_2429,N_1215,N_1278);
or U2430 (N_2430,N_1136,N_1639);
nor U2431 (N_2431,N_1720,N_1723);
nand U2432 (N_2432,N_1772,N_1960);
nor U2433 (N_2433,N_1861,N_1457);
nand U2434 (N_2434,N_1470,N_1648);
xnor U2435 (N_2435,N_1547,N_1525);
and U2436 (N_2436,N_1633,N_1180);
and U2437 (N_2437,N_1995,N_1148);
or U2438 (N_2438,N_1194,N_1309);
nor U2439 (N_2439,N_1888,N_1649);
or U2440 (N_2440,N_1302,N_1955);
nand U2441 (N_2441,N_1529,N_1881);
nand U2442 (N_2442,N_1508,N_1675);
nand U2443 (N_2443,N_1811,N_1827);
nand U2444 (N_2444,N_1825,N_1063);
nand U2445 (N_2445,N_1678,N_1068);
nor U2446 (N_2446,N_1552,N_1895);
and U2447 (N_2447,N_1134,N_1968);
and U2448 (N_2448,N_1657,N_1641);
nor U2449 (N_2449,N_1135,N_1322);
and U2450 (N_2450,N_1501,N_1091);
nand U2451 (N_2451,N_1929,N_1002);
or U2452 (N_2452,N_1222,N_1627);
or U2453 (N_2453,N_1200,N_1245);
and U2454 (N_2454,N_1182,N_1045);
nor U2455 (N_2455,N_1856,N_1582);
xnor U2456 (N_2456,N_1107,N_1021);
nor U2457 (N_2457,N_1992,N_1259);
and U2458 (N_2458,N_1715,N_1576);
and U2459 (N_2459,N_1210,N_1828);
and U2460 (N_2460,N_1485,N_1810);
or U2461 (N_2461,N_1174,N_1500);
nand U2462 (N_2462,N_1132,N_1269);
and U2463 (N_2463,N_1663,N_1080);
nor U2464 (N_2464,N_1497,N_1399);
nand U2465 (N_2465,N_1654,N_1970);
nor U2466 (N_2466,N_1161,N_1801);
nor U2467 (N_2467,N_1520,N_1143);
and U2468 (N_2468,N_1344,N_1250);
nor U2469 (N_2469,N_1779,N_1707);
and U2470 (N_2470,N_1123,N_1562);
and U2471 (N_2471,N_1435,N_1377);
or U2472 (N_2472,N_1113,N_1209);
and U2473 (N_2473,N_1899,N_1953);
and U2474 (N_2474,N_1356,N_1468);
and U2475 (N_2475,N_1392,N_1963);
nor U2476 (N_2476,N_1793,N_1499);
nand U2477 (N_2477,N_1704,N_1147);
nor U2478 (N_2478,N_1150,N_1231);
and U2479 (N_2479,N_1709,N_1102);
xor U2480 (N_2480,N_1034,N_1689);
xor U2481 (N_2481,N_1119,N_1583);
and U2482 (N_2482,N_1240,N_1313);
and U2483 (N_2483,N_1491,N_1424);
xnor U2484 (N_2484,N_1164,N_1818);
or U2485 (N_2485,N_1019,N_1354);
or U2486 (N_2486,N_1169,N_1300);
nor U2487 (N_2487,N_1273,N_1114);
or U2488 (N_2488,N_1092,N_1505);
and U2489 (N_2489,N_1320,N_1315);
nand U2490 (N_2490,N_1137,N_1962);
or U2491 (N_2491,N_1296,N_1789);
nor U2492 (N_2492,N_1388,N_1902);
and U2493 (N_2493,N_1193,N_1489);
nor U2494 (N_2494,N_1683,N_1591);
or U2495 (N_2495,N_1958,N_1912);
and U2496 (N_2496,N_1220,N_1453);
and U2497 (N_2497,N_1336,N_1230);
or U2498 (N_2498,N_1078,N_1048);
or U2499 (N_2499,N_1400,N_1122);
nand U2500 (N_2500,N_1374,N_1884);
or U2501 (N_2501,N_1207,N_1056);
nand U2502 (N_2502,N_1648,N_1143);
xor U2503 (N_2503,N_1551,N_1422);
and U2504 (N_2504,N_1289,N_1678);
nor U2505 (N_2505,N_1296,N_1220);
nand U2506 (N_2506,N_1880,N_1229);
xnor U2507 (N_2507,N_1266,N_1053);
and U2508 (N_2508,N_1083,N_1301);
and U2509 (N_2509,N_1244,N_1396);
xnor U2510 (N_2510,N_1254,N_1903);
nand U2511 (N_2511,N_1469,N_1772);
nor U2512 (N_2512,N_1355,N_1819);
nand U2513 (N_2513,N_1926,N_1731);
or U2514 (N_2514,N_1337,N_1644);
nor U2515 (N_2515,N_1144,N_1245);
or U2516 (N_2516,N_1771,N_1478);
and U2517 (N_2517,N_1640,N_1943);
xnor U2518 (N_2518,N_1819,N_1513);
nand U2519 (N_2519,N_1286,N_1321);
nor U2520 (N_2520,N_1423,N_1425);
or U2521 (N_2521,N_1923,N_1909);
nor U2522 (N_2522,N_1957,N_1520);
and U2523 (N_2523,N_1956,N_1736);
and U2524 (N_2524,N_1370,N_1918);
nand U2525 (N_2525,N_1035,N_1076);
nand U2526 (N_2526,N_1754,N_1367);
and U2527 (N_2527,N_1174,N_1981);
or U2528 (N_2528,N_1147,N_1863);
or U2529 (N_2529,N_1485,N_1835);
or U2530 (N_2530,N_1760,N_1086);
and U2531 (N_2531,N_1406,N_1228);
and U2532 (N_2532,N_1898,N_1224);
xor U2533 (N_2533,N_1326,N_1598);
and U2534 (N_2534,N_1615,N_1481);
and U2535 (N_2535,N_1767,N_1037);
nor U2536 (N_2536,N_1156,N_1813);
or U2537 (N_2537,N_1923,N_1106);
nor U2538 (N_2538,N_1820,N_1918);
and U2539 (N_2539,N_1311,N_1684);
nor U2540 (N_2540,N_1373,N_1121);
xor U2541 (N_2541,N_1870,N_1218);
and U2542 (N_2542,N_1057,N_1486);
nor U2543 (N_2543,N_1310,N_1760);
nor U2544 (N_2544,N_1311,N_1160);
nor U2545 (N_2545,N_1336,N_1612);
nor U2546 (N_2546,N_1488,N_1209);
xor U2547 (N_2547,N_1468,N_1195);
and U2548 (N_2548,N_1335,N_1958);
and U2549 (N_2549,N_1518,N_1675);
and U2550 (N_2550,N_1208,N_1405);
nor U2551 (N_2551,N_1585,N_1736);
or U2552 (N_2552,N_1236,N_1654);
or U2553 (N_2553,N_1844,N_1635);
nand U2554 (N_2554,N_1567,N_1595);
nor U2555 (N_2555,N_1170,N_1065);
nor U2556 (N_2556,N_1863,N_1067);
and U2557 (N_2557,N_1576,N_1312);
xor U2558 (N_2558,N_1796,N_1156);
nor U2559 (N_2559,N_1179,N_1733);
xnor U2560 (N_2560,N_1600,N_1615);
and U2561 (N_2561,N_1594,N_1949);
nand U2562 (N_2562,N_1863,N_1286);
nor U2563 (N_2563,N_1675,N_1973);
or U2564 (N_2564,N_1675,N_1222);
nand U2565 (N_2565,N_1964,N_1089);
xnor U2566 (N_2566,N_1947,N_1364);
nor U2567 (N_2567,N_1114,N_1778);
or U2568 (N_2568,N_1097,N_1702);
or U2569 (N_2569,N_1258,N_1979);
and U2570 (N_2570,N_1874,N_1787);
nand U2571 (N_2571,N_1256,N_1379);
nor U2572 (N_2572,N_1098,N_1363);
xnor U2573 (N_2573,N_1959,N_1611);
nand U2574 (N_2574,N_1132,N_1464);
nand U2575 (N_2575,N_1666,N_1250);
nand U2576 (N_2576,N_1813,N_1454);
and U2577 (N_2577,N_1952,N_1703);
and U2578 (N_2578,N_1320,N_1579);
nor U2579 (N_2579,N_1378,N_1900);
nand U2580 (N_2580,N_1997,N_1360);
or U2581 (N_2581,N_1159,N_1652);
nand U2582 (N_2582,N_1621,N_1536);
nand U2583 (N_2583,N_1183,N_1561);
or U2584 (N_2584,N_1950,N_1576);
and U2585 (N_2585,N_1296,N_1534);
nor U2586 (N_2586,N_1259,N_1545);
nand U2587 (N_2587,N_1492,N_1317);
and U2588 (N_2588,N_1731,N_1161);
nand U2589 (N_2589,N_1518,N_1363);
nor U2590 (N_2590,N_1872,N_1848);
and U2591 (N_2591,N_1572,N_1892);
nor U2592 (N_2592,N_1482,N_1662);
nor U2593 (N_2593,N_1378,N_1927);
nor U2594 (N_2594,N_1606,N_1661);
nand U2595 (N_2595,N_1585,N_1616);
nand U2596 (N_2596,N_1117,N_1699);
xor U2597 (N_2597,N_1410,N_1924);
or U2598 (N_2598,N_1276,N_1847);
and U2599 (N_2599,N_1534,N_1879);
or U2600 (N_2600,N_1057,N_1851);
or U2601 (N_2601,N_1513,N_1411);
or U2602 (N_2602,N_1227,N_1601);
or U2603 (N_2603,N_1637,N_1001);
or U2604 (N_2604,N_1507,N_1606);
xor U2605 (N_2605,N_1325,N_1594);
and U2606 (N_2606,N_1530,N_1823);
xnor U2607 (N_2607,N_1907,N_1616);
nor U2608 (N_2608,N_1477,N_1879);
nand U2609 (N_2609,N_1116,N_1658);
nor U2610 (N_2610,N_1308,N_1522);
and U2611 (N_2611,N_1171,N_1535);
xnor U2612 (N_2612,N_1523,N_1764);
or U2613 (N_2613,N_1866,N_1302);
nand U2614 (N_2614,N_1604,N_1504);
nor U2615 (N_2615,N_1123,N_1721);
xnor U2616 (N_2616,N_1236,N_1680);
nand U2617 (N_2617,N_1373,N_1061);
xor U2618 (N_2618,N_1104,N_1351);
and U2619 (N_2619,N_1706,N_1919);
and U2620 (N_2620,N_1409,N_1092);
xnor U2621 (N_2621,N_1166,N_1254);
xnor U2622 (N_2622,N_1500,N_1898);
nor U2623 (N_2623,N_1835,N_1339);
nor U2624 (N_2624,N_1368,N_1946);
nor U2625 (N_2625,N_1523,N_1856);
nand U2626 (N_2626,N_1727,N_1981);
nor U2627 (N_2627,N_1002,N_1665);
nor U2628 (N_2628,N_1808,N_1999);
nor U2629 (N_2629,N_1819,N_1267);
or U2630 (N_2630,N_1161,N_1391);
xnor U2631 (N_2631,N_1091,N_1834);
or U2632 (N_2632,N_1448,N_1711);
nand U2633 (N_2633,N_1929,N_1992);
nand U2634 (N_2634,N_1555,N_1562);
xnor U2635 (N_2635,N_1852,N_1278);
nor U2636 (N_2636,N_1382,N_1886);
nor U2637 (N_2637,N_1820,N_1392);
or U2638 (N_2638,N_1878,N_1567);
nand U2639 (N_2639,N_1981,N_1436);
nor U2640 (N_2640,N_1077,N_1221);
nor U2641 (N_2641,N_1089,N_1842);
nor U2642 (N_2642,N_1310,N_1496);
nor U2643 (N_2643,N_1109,N_1936);
and U2644 (N_2644,N_1524,N_1579);
and U2645 (N_2645,N_1461,N_1636);
nor U2646 (N_2646,N_1919,N_1481);
nand U2647 (N_2647,N_1015,N_1604);
or U2648 (N_2648,N_1703,N_1937);
or U2649 (N_2649,N_1577,N_1461);
nand U2650 (N_2650,N_1352,N_1497);
nor U2651 (N_2651,N_1639,N_1931);
and U2652 (N_2652,N_1017,N_1104);
nand U2653 (N_2653,N_1976,N_1977);
or U2654 (N_2654,N_1343,N_1507);
nand U2655 (N_2655,N_1640,N_1940);
or U2656 (N_2656,N_1107,N_1501);
nor U2657 (N_2657,N_1477,N_1914);
nand U2658 (N_2658,N_1267,N_1202);
and U2659 (N_2659,N_1416,N_1332);
or U2660 (N_2660,N_1059,N_1904);
or U2661 (N_2661,N_1599,N_1251);
xor U2662 (N_2662,N_1362,N_1552);
xor U2663 (N_2663,N_1538,N_1794);
and U2664 (N_2664,N_1094,N_1342);
or U2665 (N_2665,N_1859,N_1223);
or U2666 (N_2666,N_1380,N_1746);
nand U2667 (N_2667,N_1426,N_1323);
nand U2668 (N_2668,N_1001,N_1599);
nand U2669 (N_2669,N_1720,N_1979);
nand U2670 (N_2670,N_1706,N_1750);
nand U2671 (N_2671,N_1296,N_1086);
or U2672 (N_2672,N_1357,N_1717);
nand U2673 (N_2673,N_1558,N_1836);
or U2674 (N_2674,N_1572,N_1102);
and U2675 (N_2675,N_1555,N_1210);
or U2676 (N_2676,N_1043,N_1415);
nand U2677 (N_2677,N_1458,N_1819);
and U2678 (N_2678,N_1242,N_1280);
xnor U2679 (N_2679,N_1900,N_1983);
xnor U2680 (N_2680,N_1306,N_1536);
and U2681 (N_2681,N_1366,N_1096);
nand U2682 (N_2682,N_1894,N_1140);
or U2683 (N_2683,N_1928,N_1964);
nor U2684 (N_2684,N_1584,N_1256);
nor U2685 (N_2685,N_1990,N_1702);
nor U2686 (N_2686,N_1545,N_1663);
or U2687 (N_2687,N_1184,N_1033);
and U2688 (N_2688,N_1106,N_1713);
nand U2689 (N_2689,N_1818,N_1473);
nor U2690 (N_2690,N_1150,N_1097);
xnor U2691 (N_2691,N_1855,N_1767);
nor U2692 (N_2692,N_1439,N_1319);
nor U2693 (N_2693,N_1365,N_1731);
nor U2694 (N_2694,N_1070,N_1905);
nand U2695 (N_2695,N_1001,N_1351);
nand U2696 (N_2696,N_1303,N_1402);
nand U2697 (N_2697,N_1426,N_1108);
and U2698 (N_2698,N_1867,N_1636);
or U2699 (N_2699,N_1839,N_1245);
nand U2700 (N_2700,N_1780,N_1486);
or U2701 (N_2701,N_1544,N_1471);
or U2702 (N_2702,N_1486,N_1709);
nand U2703 (N_2703,N_1098,N_1028);
nor U2704 (N_2704,N_1897,N_1490);
or U2705 (N_2705,N_1611,N_1712);
xnor U2706 (N_2706,N_1780,N_1035);
nor U2707 (N_2707,N_1519,N_1609);
nor U2708 (N_2708,N_1333,N_1379);
nor U2709 (N_2709,N_1720,N_1525);
and U2710 (N_2710,N_1801,N_1861);
nor U2711 (N_2711,N_1533,N_1387);
nor U2712 (N_2712,N_1415,N_1446);
nand U2713 (N_2713,N_1927,N_1516);
or U2714 (N_2714,N_1667,N_1476);
and U2715 (N_2715,N_1258,N_1200);
or U2716 (N_2716,N_1980,N_1204);
and U2717 (N_2717,N_1535,N_1898);
or U2718 (N_2718,N_1342,N_1469);
or U2719 (N_2719,N_1075,N_1323);
nand U2720 (N_2720,N_1534,N_1237);
xnor U2721 (N_2721,N_1060,N_1667);
nor U2722 (N_2722,N_1238,N_1120);
nor U2723 (N_2723,N_1963,N_1805);
or U2724 (N_2724,N_1895,N_1688);
nand U2725 (N_2725,N_1465,N_1726);
nor U2726 (N_2726,N_1421,N_1718);
or U2727 (N_2727,N_1095,N_1081);
and U2728 (N_2728,N_1696,N_1815);
nand U2729 (N_2729,N_1172,N_1068);
nor U2730 (N_2730,N_1360,N_1188);
or U2731 (N_2731,N_1435,N_1151);
nor U2732 (N_2732,N_1597,N_1345);
and U2733 (N_2733,N_1792,N_1861);
and U2734 (N_2734,N_1233,N_1030);
nand U2735 (N_2735,N_1056,N_1297);
xor U2736 (N_2736,N_1854,N_1531);
nor U2737 (N_2737,N_1925,N_1857);
nand U2738 (N_2738,N_1885,N_1766);
and U2739 (N_2739,N_1038,N_1900);
nand U2740 (N_2740,N_1363,N_1505);
xnor U2741 (N_2741,N_1053,N_1527);
nand U2742 (N_2742,N_1843,N_1004);
nor U2743 (N_2743,N_1160,N_1776);
nor U2744 (N_2744,N_1335,N_1561);
or U2745 (N_2745,N_1986,N_1853);
nor U2746 (N_2746,N_1055,N_1964);
nor U2747 (N_2747,N_1027,N_1128);
nand U2748 (N_2748,N_1490,N_1268);
or U2749 (N_2749,N_1858,N_1381);
nand U2750 (N_2750,N_1517,N_1114);
and U2751 (N_2751,N_1240,N_1033);
nand U2752 (N_2752,N_1157,N_1276);
and U2753 (N_2753,N_1964,N_1530);
and U2754 (N_2754,N_1449,N_1229);
nand U2755 (N_2755,N_1497,N_1588);
nand U2756 (N_2756,N_1919,N_1247);
nor U2757 (N_2757,N_1216,N_1152);
nand U2758 (N_2758,N_1591,N_1111);
nor U2759 (N_2759,N_1946,N_1590);
or U2760 (N_2760,N_1953,N_1361);
nand U2761 (N_2761,N_1288,N_1552);
nor U2762 (N_2762,N_1448,N_1475);
xor U2763 (N_2763,N_1143,N_1863);
nand U2764 (N_2764,N_1305,N_1303);
and U2765 (N_2765,N_1996,N_1029);
and U2766 (N_2766,N_1323,N_1237);
nor U2767 (N_2767,N_1549,N_1723);
nand U2768 (N_2768,N_1629,N_1720);
or U2769 (N_2769,N_1274,N_1684);
and U2770 (N_2770,N_1672,N_1745);
and U2771 (N_2771,N_1434,N_1008);
or U2772 (N_2772,N_1833,N_1385);
or U2773 (N_2773,N_1304,N_1968);
nor U2774 (N_2774,N_1795,N_1664);
and U2775 (N_2775,N_1307,N_1169);
and U2776 (N_2776,N_1421,N_1984);
nand U2777 (N_2777,N_1441,N_1062);
nor U2778 (N_2778,N_1171,N_1109);
and U2779 (N_2779,N_1542,N_1999);
and U2780 (N_2780,N_1549,N_1429);
or U2781 (N_2781,N_1503,N_1917);
or U2782 (N_2782,N_1789,N_1573);
or U2783 (N_2783,N_1952,N_1698);
and U2784 (N_2784,N_1635,N_1146);
nor U2785 (N_2785,N_1760,N_1472);
nand U2786 (N_2786,N_1426,N_1969);
nor U2787 (N_2787,N_1797,N_1361);
nor U2788 (N_2788,N_1625,N_1244);
and U2789 (N_2789,N_1642,N_1842);
nor U2790 (N_2790,N_1769,N_1831);
nand U2791 (N_2791,N_1623,N_1183);
and U2792 (N_2792,N_1038,N_1042);
or U2793 (N_2793,N_1240,N_1530);
or U2794 (N_2794,N_1135,N_1989);
and U2795 (N_2795,N_1625,N_1669);
nand U2796 (N_2796,N_1879,N_1238);
and U2797 (N_2797,N_1436,N_1748);
nor U2798 (N_2798,N_1373,N_1058);
nor U2799 (N_2799,N_1695,N_1427);
nand U2800 (N_2800,N_1036,N_1637);
nand U2801 (N_2801,N_1932,N_1360);
xnor U2802 (N_2802,N_1314,N_1953);
and U2803 (N_2803,N_1171,N_1921);
or U2804 (N_2804,N_1652,N_1438);
or U2805 (N_2805,N_1931,N_1984);
nand U2806 (N_2806,N_1442,N_1319);
or U2807 (N_2807,N_1021,N_1373);
nand U2808 (N_2808,N_1373,N_1867);
nor U2809 (N_2809,N_1163,N_1035);
nand U2810 (N_2810,N_1827,N_1894);
nor U2811 (N_2811,N_1367,N_1383);
nor U2812 (N_2812,N_1493,N_1182);
nor U2813 (N_2813,N_1773,N_1780);
and U2814 (N_2814,N_1962,N_1026);
or U2815 (N_2815,N_1422,N_1150);
and U2816 (N_2816,N_1842,N_1040);
or U2817 (N_2817,N_1691,N_1789);
or U2818 (N_2818,N_1902,N_1176);
nor U2819 (N_2819,N_1550,N_1088);
or U2820 (N_2820,N_1911,N_1507);
or U2821 (N_2821,N_1382,N_1272);
or U2822 (N_2822,N_1984,N_1679);
and U2823 (N_2823,N_1255,N_1388);
and U2824 (N_2824,N_1399,N_1495);
xnor U2825 (N_2825,N_1289,N_1611);
xor U2826 (N_2826,N_1433,N_1941);
and U2827 (N_2827,N_1359,N_1771);
nor U2828 (N_2828,N_1055,N_1365);
nand U2829 (N_2829,N_1279,N_1540);
and U2830 (N_2830,N_1000,N_1985);
and U2831 (N_2831,N_1104,N_1503);
nor U2832 (N_2832,N_1887,N_1294);
or U2833 (N_2833,N_1052,N_1206);
nor U2834 (N_2834,N_1934,N_1613);
nor U2835 (N_2835,N_1783,N_1612);
nor U2836 (N_2836,N_1876,N_1840);
or U2837 (N_2837,N_1254,N_1227);
nor U2838 (N_2838,N_1564,N_1430);
nor U2839 (N_2839,N_1098,N_1044);
nor U2840 (N_2840,N_1679,N_1407);
nand U2841 (N_2841,N_1862,N_1271);
xor U2842 (N_2842,N_1464,N_1386);
nor U2843 (N_2843,N_1695,N_1028);
and U2844 (N_2844,N_1278,N_1532);
xor U2845 (N_2845,N_1196,N_1114);
nor U2846 (N_2846,N_1078,N_1894);
nand U2847 (N_2847,N_1008,N_1159);
or U2848 (N_2848,N_1214,N_1731);
xor U2849 (N_2849,N_1601,N_1180);
or U2850 (N_2850,N_1179,N_1268);
nand U2851 (N_2851,N_1951,N_1836);
nor U2852 (N_2852,N_1170,N_1401);
nor U2853 (N_2853,N_1215,N_1495);
and U2854 (N_2854,N_1784,N_1224);
nor U2855 (N_2855,N_1500,N_1932);
nor U2856 (N_2856,N_1519,N_1668);
and U2857 (N_2857,N_1737,N_1732);
and U2858 (N_2858,N_1509,N_1149);
nand U2859 (N_2859,N_1679,N_1663);
nor U2860 (N_2860,N_1620,N_1628);
and U2861 (N_2861,N_1200,N_1704);
nand U2862 (N_2862,N_1057,N_1012);
xnor U2863 (N_2863,N_1539,N_1307);
nor U2864 (N_2864,N_1148,N_1285);
xnor U2865 (N_2865,N_1614,N_1676);
or U2866 (N_2866,N_1294,N_1250);
or U2867 (N_2867,N_1271,N_1450);
nor U2868 (N_2868,N_1652,N_1516);
nand U2869 (N_2869,N_1697,N_1841);
nor U2870 (N_2870,N_1868,N_1023);
or U2871 (N_2871,N_1017,N_1326);
or U2872 (N_2872,N_1412,N_1184);
or U2873 (N_2873,N_1970,N_1139);
nor U2874 (N_2874,N_1507,N_1092);
nor U2875 (N_2875,N_1509,N_1299);
or U2876 (N_2876,N_1913,N_1233);
nand U2877 (N_2877,N_1028,N_1856);
and U2878 (N_2878,N_1885,N_1870);
and U2879 (N_2879,N_1602,N_1367);
and U2880 (N_2880,N_1039,N_1368);
or U2881 (N_2881,N_1525,N_1772);
nor U2882 (N_2882,N_1692,N_1531);
or U2883 (N_2883,N_1243,N_1121);
or U2884 (N_2884,N_1256,N_1141);
or U2885 (N_2885,N_1166,N_1876);
nand U2886 (N_2886,N_1157,N_1910);
or U2887 (N_2887,N_1049,N_1308);
xor U2888 (N_2888,N_1624,N_1636);
nand U2889 (N_2889,N_1506,N_1537);
nand U2890 (N_2890,N_1931,N_1886);
nand U2891 (N_2891,N_1245,N_1595);
xnor U2892 (N_2892,N_1300,N_1805);
or U2893 (N_2893,N_1704,N_1479);
nor U2894 (N_2894,N_1754,N_1585);
or U2895 (N_2895,N_1728,N_1784);
and U2896 (N_2896,N_1591,N_1130);
nand U2897 (N_2897,N_1094,N_1221);
nand U2898 (N_2898,N_1556,N_1878);
and U2899 (N_2899,N_1770,N_1342);
and U2900 (N_2900,N_1769,N_1401);
xnor U2901 (N_2901,N_1279,N_1471);
xnor U2902 (N_2902,N_1793,N_1518);
or U2903 (N_2903,N_1147,N_1028);
nor U2904 (N_2904,N_1801,N_1335);
nand U2905 (N_2905,N_1332,N_1430);
xnor U2906 (N_2906,N_1137,N_1033);
or U2907 (N_2907,N_1387,N_1322);
and U2908 (N_2908,N_1758,N_1312);
or U2909 (N_2909,N_1477,N_1648);
nor U2910 (N_2910,N_1054,N_1573);
and U2911 (N_2911,N_1819,N_1419);
xnor U2912 (N_2912,N_1355,N_1101);
and U2913 (N_2913,N_1741,N_1416);
nor U2914 (N_2914,N_1574,N_1635);
nand U2915 (N_2915,N_1888,N_1632);
nand U2916 (N_2916,N_1371,N_1545);
nor U2917 (N_2917,N_1498,N_1366);
or U2918 (N_2918,N_1451,N_1083);
or U2919 (N_2919,N_1636,N_1448);
and U2920 (N_2920,N_1599,N_1132);
or U2921 (N_2921,N_1867,N_1405);
and U2922 (N_2922,N_1012,N_1976);
and U2923 (N_2923,N_1787,N_1944);
and U2924 (N_2924,N_1130,N_1267);
or U2925 (N_2925,N_1708,N_1188);
and U2926 (N_2926,N_1189,N_1691);
and U2927 (N_2927,N_1652,N_1402);
and U2928 (N_2928,N_1942,N_1906);
nand U2929 (N_2929,N_1963,N_1134);
nand U2930 (N_2930,N_1408,N_1064);
and U2931 (N_2931,N_1238,N_1361);
xnor U2932 (N_2932,N_1399,N_1027);
nor U2933 (N_2933,N_1994,N_1752);
and U2934 (N_2934,N_1904,N_1296);
nand U2935 (N_2935,N_1597,N_1402);
nand U2936 (N_2936,N_1534,N_1880);
nand U2937 (N_2937,N_1243,N_1604);
nand U2938 (N_2938,N_1179,N_1008);
nor U2939 (N_2939,N_1054,N_1350);
nor U2940 (N_2940,N_1456,N_1663);
and U2941 (N_2941,N_1093,N_1275);
and U2942 (N_2942,N_1485,N_1111);
and U2943 (N_2943,N_1433,N_1801);
nand U2944 (N_2944,N_1848,N_1483);
nor U2945 (N_2945,N_1004,N_1659);
nand U2946 (N_2946,N_1889,N_1142);
or U2947 (N_2947,N_1520,N_1724);
nand U2948 (N_2948,N_1825,N_1540);
and U2949 (N_2949,N_1278,N_1007);
or U2950 (N_2950,N_1449,N_1118);
or U2951 (N_2951,N_1115,N_1391);
or U2952 (N_2952,N_1290,N_1612);
and U2953 (N_2953,N_1060,N_1508);
xnor U2954 (N_2954,N_1966,N_1424);
or U2955 (N_2955,N_1916,N_1508);
nand U2956 (N_2956,N_1910,N_1246);
and U2957 (N_2957,N_1145,N_1488);
nor U2958 (N_2958,N_1234,N_1371);
nand U2959 (N_2959,N_1408,N_1872);
xor U2960 (N_2960,N_1801,N_1121);
xor U2961 (N_2961,N_1974,N_1121);
nor U2962 (N_2962,N_1837,N_1004);
nand U2963 (N_2963,N_1201,N_1089);
nand U2964 (N_2964,N_1275,N_1482);
nand U2965 (N_2965,N_1998,N_1987);
or U2966 (N_2966,N_1346,N_1778);
nor U2967 (N_2967,N_1482,N_1134);
and U2968 (N_2968,N_1508,N_1914);
or U2969 (N_2969,N_1925,N_1105);
nor U2970 (N_2970,N_1381,N_1009);
nand U2971 (N_2971,N_1176,N_1879);
xor U2972 (N_2972,N_1253,N_1974);
or U2973 (N_2973,N_1914,N_1619);
or U2974 (N_2974,N_1488,N_1364);
or U2975 (N_2975,N_1053,N_1936);
or U2976 (N_2976,N_1202,N_1805);
nor U2977 (N_2977,N_1362,N_1731);
or U2978 (N_2978,N_1169,N_1051);
and U2979 (N_2979,N_1444,N_1238);
nor U2980 (N_2980,N_1838,N_1037);
nand U2981 (N_2981,N_1415,N_1789);
xnor U2982 (N_2982,N_1685,N_1262);
nor U2983 (N_2983,N_1515,N_1246);
nor U2984 (N_2984,N_1081,N_1833);
nand U2985 (N_2985,N_1637,N_1339);
and U2986 (N_2986,N_1642,N_1163);
xor U2987 (N_2987,N_1760,N_1153);
and U2988 (N_2988,N_1367,N_1196);
nand U2989 (N_2989,N_1099,N_1012);
nand U2990 (N_2990,N_1538,N_1878);
or U2991 (N_2991,N_1969,N_1029);
xnor U2992 (N_2992,N_1050,N_1316);
or U2993 (N_2993,N_1579,N_1288);
nand U2994 (N_2994,N_1565,N_1009);
xor U2995 (N_2995,N_1418,N_1181);
or U2996 (N_2996,N_1017,N_1345);
or U2997 (N_2997,N_1508,N_1076);
and U2998 (N_2998,N_1536,N_1963);
or U2999 (N_2999,N_1190,N_1517);
nand UO_0 (O_0,N_2940,N_2269);
xnor UO_1 (O_1,N_2572,N_2726);
and UO_2 (O_2,N_2605,N_2597);
nand UO_3 (O_3,N_2689,N_2471);
nand UO_4 (O_4,N_2228,N_2058);
nor UO_5 (O_5,N_2032,N_2417);
nand UO_6 (O_6,N_2793,N_2264);
nand UO_7 (O_7,N_2346,N_2511);
or UO_8 (O_8,N_2991,N_2255);
nor UO_9 (O_9,N_2443,N_2157);
nand UO_10 (O_10,N_2720,N_2507);
nand UO_11 (O_11,N_2132,N_2618);
nor UO_12 (O_12,N_2513,N_2355);
and UO_13 (O_13,N_2257,N_2781);
and UO_14 (O_14,N_2531,N_2743);
and UO_15 (O_15,N_2460,N_2772);
or UO_16 (O_16,N_2634,N_2410);
and UO_17 (O_17,N_2037,N_2093);
nand UO_18 (O_18,N_2150,N_2935);
nand UO_19 (O_19,N_2898,N_2801);
nand UO_20 (O_20,N_2496,N_2843);
nand UO_21 (O_21,N_2331,N_2756);
or UO_22 (O_22,N_2595,N_2985);
and UO_23 (O_23,N_2375,N_2939);
or UO_24 (O_24,N_2796,N_2553);
nand UO_25 (O_25,N_2860,N_2609);
or UO_26 (O_26,N_2842,N_2327);
nor UO_27 (O_27,N_2428,N_2524);
xnor UO_28 (O_28,N_2998,N_2626);
and UO_29 (O_29,N_2418,N_2266);
nand UO_30 (O_30,N_2035,N_2329);
nor UO_31 (O_31,N_2218,N_2321);
or UO_32 (O_32,N_2240,N_2876);
nand UO_33 (O_33,N_2527,N_2112);
nor UO_34 (O_34,N_2232,N_2712);
xor UO_35 (O_35,N_2462,N_2281);
nor UO_36 (O_36,N_2302,N_2859);
or UO_37 (O_37,N_2092,N_2352);
nand UO_38 (O_38,N_2691,N_2052);
and UO_39 (O_39,N_2326,N_2811);
nor UO_40 (O_40,N_2825,N_2676);
and UO_41 (O_41,N_2661,N_2474);
nand UO_42 (O_42,N_2668,N_2891);
and UO_43 (O_43,N_2837,N_2763);
nor UO_44 (O_44,N_2630,N_2555);
and UO_45 (O_45,N_2742,N_2459);
xnor UO_46 (O_46,N_2751,N_2980);
nor UO_47 (O_47,N_2386,N_2768);
nand UO_48 (O_48,N_2739,N_2650);
and UO_49 (O_49,N_2340,N_2581);
and UO_50 (O_50,N_2864,N_2614);
or UO_51 (O_51,N_2397,N_2186);
xnor UO_52 (O_52,N_2065,N_2688);
nor UO_53 (O_53,N_2493,N_2006);
nor UO_54 (O_54,N_2559,N_2197);
nor UO_55 (O_55,N_2760,N_2078);
nor UO_56 (O_56,N_2219,N_2530);
and UO_57 (O_57,N_2239,N_2425);
nor UO_58 (O_58,N_2131,N_2335);
and UO_59 (O_59,N_2512,N_2012);
or UO_60 (O_60,N_2631,N_2115);
nand UO_61 (O_61,N_2855,N_2441);
and UO_62 (O_62,N_2976,N_2633);
and UO_63 (O_63,N_2705,N_2299);
nor UO_64 (O_64,N_2519,N_2127);
nor UO_65 (O_65,N_2722,N_2996);
nor UO_66 (O_66,N_2217,N_2072);
and UO_67 (O_67,N_2350,N_2806);
or UO_68 (O_68,N_2666,N_2292);
and UO_69 (O_69,N_2000,N_2649);
and UO_70 (O_70,N_2967,N_2448);
nand UO_71 (O_71,N_2194,N_2371);
and UO_72 (O_72,N_2883,N_2258);
or UO_73 (O_73,N_2180,N_2869);
and UO_74 (O_74,N_2695,N_2918);
nor UO_75 (O_75,N_2674,N_2522);
and UO_76 (O_76,N_2309,N_2424);
nor UO_77 (O_77,N_2393,N_2546);
xnor UO_78 (O_78,N_2048,N_2728);
nand UO_79 (O_79,N_2889,N_2771);
nor UO_80 (O_80,N_2933,N_2733);
nand UO_81 (O_81,N_2243,N_2044);
nand UO_82 (O_82,N_2685,N_2830);
nand UO_83 (O_83,N_2794,N_2323);
and UO_84 (O_84,N_2066,N_2617);
nand UO_85 (O_85,N_2042,N_2168);
nand UO_86 (O_86,N_2322,N_2560);
and UO_87 (O_87,N_2364,N_2149);
or UO_88 (O_88,N_2382,N_2420);
and UO_89 (O_89,N_2916,N_2995);
nor UO_90 (O_90,N_2325,N_2818);
nand UO_91 (O_91,N_2815,N_2189);
and UO_92 (O_92,N_2455,N_2971);
xnor UO_93 (O_93,N_2039,N_2023);
or UO_94 (O_94,N_2964,N_2170);
nor UO_95 (O_95,N_2759,N_2658);
or UO_96 (O_96,N_2261,N_2449);
nor UO_97 (O_97,N_2308,N_2200);
nand UO_98 (O_98,N_2749,N_2025);
xor UO_99 (O_99,N_2556,N_2736);
nand UO_100 (O_100,N_2061,N_2005);
nor UO_101 (O_101,N_2354,N_2670);
or UO_102 (O_102,N_2268,N_2171);
xnor UO_103 (O_103,N_2704,N_2063);
nor UO_104 (O_104,N_2642,N_2349);
nand UO_105 (O_105,N_2604,N_2205);
or UO_106 (O_106,N_2653,N_2900);
or UO_107 (O_107,N_2176,N_2946);
nor UO_108 (O_108,N_2782,N_2886);
nand UO_109 (O_109,N_2358,N_2646);
nand UO_110 (O_110,N_2136,N_2094);
nor UO_111 (O_111,N_2706,N_2026);
or UO_112 (O_112,N_2224,N_2682);
nand UO_113 (O_113,N_2922,N_2960);
nand UO_114 (O_114,N_2125,N_2095);
nand UO_115 (O_115,N_2117,N_2036);
xor UO_116 (O_116,N_2421,N_2096);
xnor UO_117 (O_117,N_2056,N_2100);
nand UO_118 (O_118,N_2901,N_2550);
and UO_119 (O_119,N_2993,N_2831);
or UO_120 (O_120,N_2001,N_2896);
or UO_121 (O_121,N_2684,N_2403);
and UO_122 (O_122,N_2923,N_2506);
xnor UO_123 (O_123,N_2129,N_2526);
and UO_124 (O_124,N_2988,N_2019);
xor UO_125 (O_125,N_2256,N_2948);
nand UO_126 (O_126,N_2997,N_2810);
and UO_127 (O_127,N_2865,N_2592);
nor UO_128 (O_128,N_2235,N_2033);
and UO_129 (O_129,N_2499,N_2687);
nor UO_130 (O_130,N_2483,N_2582);
nand UO_131 (O_131,N_2740,N_2930);
xor UO_132 (O_132,N_2637,N_2043);
or UO_133 (O_133,N_2868,N_2612);
nand UO_134 (O_134,N_2181,N_2450);
xnor UO_135 (O_135,N_2076,N_2490);
nand UO_136 (O_136,N_2639,N_2333);
and UO_137 (O_137,N_2757,N_2857);
nand UO_138 (O_138,N_2416,N_2401);
nor UO_139 (O_139,N_2298,N_2412);
and UO_140 (O_140,N_2353,N_2015);
and UO_141 (O_141,N_2681,N_2284);
or UO_142 (O_142,N_2011,N_2797);
nand UO_143 (O_143,N_2594,N_2301);
and UO_144 (O_144,N_2716,N_2476);
nor UO_145 (O_145,N_2725,N_2764);
nor UO_146 (O_146,N_2404,N_2558);
or UO_147 (O_147,N_2521,N_2500);
nand UO_148 (O_148,N_2178,N_2209);
nor UO_149 (O_149,N_2941,N_2854);
nor UO_150 (O_150,N_2481,N_2529);
or UO_151 (O_151,N_2698,N_2040);
or UO_152 (O_152,N_2858,N_2847);
nor UO_153 (O_153,N_2875,N_2746);
nor UO_154 (O_154,N_2737,N_2138);
nor UO_155 (O_155,N_2657,N_2366);
nor UO_156 (O_156,N_2315,N_2505);
and UO_157 (O_157,N_2169,N_2177);
nor UO_158 (O_158,N_2850,N_2575);
and UO_159 (O_159,N_2250,N_2047);
or UO_160 (O_160,N_2758,N_2342);
nor UO_161 (O_161,N_2908,N_2028);
nor UO_162 (O_162,N_2562,N_2151);
nand UO_163 (O_163,N_2709,N_2290);
nor UO_164 (O_164,N_2973,N_2091);
nand UO_165 (O_165,N_2910,N_2950);
and UO_166 (O_166,N_2641,N_2718);
or UO_167 (O_167,N_2405,N_2565);
nand UO_168 (O_168,N_2338,N_2834);
nor UO_169 (O_169,N_2584,N_2753);
or UO_170 (O_170,N_2271,N_2598);
nand UO_171 (O_171,N_2934,N_2599);
or UO_172 (O_172,N_2501,N_2602);
nand UO_173 (O_173,N_2369,N_2291);
or UO_174 (O_174,N_2692,N_2391);
nand UO_175 (O_175,N_2162,N_2396);
or UO_176 (O_176,N_2557,N_2356);
and UO_177 (O_177,N_2894,N_2016);
nand UO_178 (O_178,N_2947,N_2153);
and UO_179 (O_179,N_2683,N_2172);
and UO_180 (O_180,N_2206,N_2114);
nor UO_181 (O_181,N_2696,N_2220);
nand UO_182 (O_182,N_2300,N_2738);
nor UO_183 (O_183,N_2080,N_2254);
nor UO_184 (O_184,N_2729,N_2362);
nor UO_185 (O_185,N_2824,N_2148);
nor UO_186 (O_186,N_2427,N_2635);
nand UO_187 (O_187,N_2880,N_2345);
and UO_188 (O_188,N_2183,N_2943);
nor UO_189 (O_189,N_2547,N_2890);
xor UO_190 (O_190,N_2456,N_2365);
nor UO_191 (O_191,N_2675,N_2415);
or UO_192 (O_192,N_2789,N_2344);
xnor UO_193 (O_193,N_2663,N_2139);
or UO_194 (O_194,N_2222,N_2051);
nand UO_195 (O_195,N_2246,N_2179);
nand UO_196 (O_196,N_2379,N_2786);
xor UO_197 (O_197,N_2569,N_2014);
or UO_198 (O_198,N_2199,N_2402);
nor UO_199 (O_199,N_2770,N_2775);
nand UO_200 (O_200,N_2422,N_2102);
nor UO_201 (O_201,N_2343,N_2929);
nand UO_202 (O_202,N_2158,N_2510);
and UO_203 (O_203,N_2981,N_2542);
and UO_204 (O_204,N_2750,N_2237);
nor UO_205 (O_205,N_2370,N_2808);
xnor UO_206 (O_206,N_2748,N_2226);
or UO_207 (O_207,N_2881,N_2103);
and UO_208 (O_208,N_2377,N_2866);
and UO_209 (O_209,N_2776,N_2593);
or UO_210 (O_210,N_2374,N_2059);
and UO_211 (O_211,N_2468,N_2089);
and UO_212 (O_212,N_2204,N_2230);
nor UO_213 (O_213,N_2304,N_2931);
nor UO_214 (O_214,N_2699,N_2234);
nor UO_215 (O_215,N_2451,N_2777);
xor UO_216 (O_216,N_2965,N_2260);
nor UO_217 (O_217,N_2549,N_2090);
or UO_218 (O_218,N_2765,N_2068);
or UO_219 (O_219,N_2975,N_2434);
nand UO_220 (O_220,N_2472,N_2307);
nor UO_221 (O_221,N_2174,N_2487);
nor UO_222 (O_222,N_2970,N_2816);
nand UO_223 (O_223,N_2086,N_2134);
nand UO_224 (O_224,N_2719,N_2341);
and UO_225 (O_225,N_2400,N_2892);
nand UO_226 (O_226,N_2795,N_2537);
and UO_227 (O_227,N_2045,N_2805);
nor UO_228 (O_228,N_2485,N_2312);
nor UO_229 (O_229,N_2671,N_2735);
or UO_230 (O_230,N_2785,N_2587);
or UO_231 (O_231,N_2282,N_2407);
nand UO_232 (O_232,N_2479,N_2055);
and UO_233 (O_233,N_2579,N_2924);
or UO_234 (O_234,N_2192,N_2867);
nand UO_235 (O_235,N_2648,N_2060);
or UO_236 (O_236,N_2589,N_2050);
nor UO_237 (O_237,N_2762,N_2724);
nor UO_238 (O_238,N_2741,N_2440);
nor UO_239 (O_239,N_2439,N_2606);
or UO_240 (O_240,N_2885,N_2084);
nand UO_241 (O_241,N_2478,N_2141);
nand UO_242 (O_242,N_2914,N_2018);
nor UO_243 (O_243,N_2774,N_2387);
xor UO_244 (O_244,N_2638,N_2295);
nor UO_245 (O_245,N_2314,N_2798);
nand UO_246 (O_246,N_2380,N_2423);
xnor UO_247 (O_247,N_2809,N_2913);
nand UO_248 (O_248,N_2128,N_2098);
or UO_249 (O_249,N_2899,N_2730);
nand UO_250 (O_250,N_2987,N_2853);
nand UO_251 (O_251,N_2679,N_2160);
nor UO_252 (O_252,N_2215,N_2389);
nor UO_253 (O_253,N_2544,N_2624);
nor UO_254 (O_254,N_2070,N_2419);
or UO_255 (O_255,N_2273,N_2755);
and UO_256 (O_256,N_2673,N_2182);
nor UO_257 (O_257,N_2841,N_2074);
nor UO_258 (O_258,N_2385,N_2664);
and UO_259 (O_259,N_2953,N_2475);
nor UO_260 (O_260,N_2390,N_2357);
nand UO_261 (O_261,N_2373,N_2442);
or UO_262 (O_262,N_2120,N_2836);
nor UO_263 (O_263,N_2911,N_2662);
or UO_264 (O_264,N_2937,N_2305);
and UO_265 (O_265,N_2840,N_2458);
or UO_266 (O_266,N_2878,N_2586);
xor UO_267 (O_267,N_2164,N_2887);
or UO_268 (O_268,N_2804,N_2163);
or UO_269 (O_269,N_2942,N_2888);
nor UO_270 (O_270,N_2381,N_2064);
nor UO_271 (O_271,N_2480,N_2278);
nor UO_272 (O_272,N_2852,N_2191);
nor UO_273 (O_273,N_2022,N_2118);
xnor UO_274 (O_274,N_2792,N_2293);
nand UO_275 (O_275,N_2715,N_2613);
and UO_276 (O_276,N_2821,N_2140);
nand UO_277 (O_277,N_2503,N_2528);
nor UO_278 (O_278,N_2359,N_2956);
nand UO_279 (O_279,N_2137,N_2938);
and UO_280 (O_280,N_2539,N_2372);
xor UO_281 (O_281,N_2625,N_2360);
xnor UO_282 (O_282,N_2202,N_2190);
nor UO_283 (O_283,N_2660,N_2807);
nand UO_284 (O_284,N_2915,N_2651);
nand UO_285 (O_285,N_2893,N_2665);
nor UO_286 (O_286,N_2655,N_2540);
nor UO_287 (O_287,N_2464,N_2551);
nor UO_288 (O_288,N_2436,N_2925);
or UO_289 (O_289,N_2536,N_2603);
nor UO_290 (O_290,N_2520,N_2962);
nand UO_291 (O_291,N_2337,N_2591);
nand UO_292 (O_292,N_2251,N_2465);
nor UO_293 (O_293,N_2285,N_2645);
and UO_294 (O_294,N_2632,N_2690);
or UO_295 (O_295,N_2989,N_2969);
nand UO_296 (O_296,N_2780,N_2640);
nor UO_297 (O_297,N_2723,N_2152);
or UO_298 (O_298,N_2124,N_2361);
xor UO_299 (O_299,N_2242,N_2870);
or UO_300 (O_300,N_2259,N_2504);
and UO_301 (O_301,N_2761,N_2498);
or UO_302 (O_302,N_2701,N_2784);
nor UO_303 (O_303,N_2802,N_2435);
or UO_304 (O_304,N_2845,N_2009);
nand UO_305 (O_305,N_2588,N_2561);
nand UO_306 (O_306,N_2057,N_2656);
nor UO_307 (O_307,N_2570,N_2945);
and UO_308 (O_308,N_2453,N_2654);
nand UO_309 (O_309,N_2972,N_2438);
and UO_310 (O_310,N_2992,N_2351);
xnor UO_311 (O_311,N_2534,N_2488);
nor UO_312 (O_312,N_2144,N_2067);
or UO_313 (O_313,N_2769,N_2306);
and UO_314 (O_314,N_2328,N_2311);
nand UO_315 (O_315,N_2707,N_2253);
nor UO_316 (O_316,N_2245,N_2029);
or UO_317 (O_317,N_2819,N_2848);
nand UO_318 (O_318,N_2585,N_2431);
and UO_319 (O_319,N_2932,N_2007);
xor UO_320 (O_320,N_2610,N_2324);
or UO_321 (O_321,N_2823,N_2813);
and UO_322 (O_322,N_2210,N_2517);
nand UO_323 (O_323,N_2754,N_2779);
and UO_324 (O_324,N_2203,N_2686);
nand UO_325 (O_325,N_2008,N_2252);
or UO_326 (O_326,N_2188,N_2999);
xor UO_327 (O_327,N_2608,N_2708);
and UO_328 (O_328,N_2949,N_2954);
and UO_329 (O_329,N_2013,N_2574);
or UO_330 (O_330,N_2142,N_2541);
and UO_331 (O_331,N_2073,N_2905);
or UO_332 (O_332,N_2467,N_2263);
or UO_333 (O_333,N_2790,N_2231);
nor UO_334 (O_334,N_2473,N_2238);
nand UO_335 (O_335,N_2079,N_2062);
and UO_336 (O_336,N_2334,N_2053);
or UO_337 (O_337,N_2452,N_2123);
and UO_338 (O_338,N_2835,N_2430);
nor UO_339 (O_339,N_2814,N_2249);
or UO_340 (O_340,N_2484,N_2839);
and UO_341 (O_341,N_2482,N_2270);
xor UO_342 (O_342,N_2196,N_2702);
nor UO_343 (O_343,N_2310,N_2677);
nor UO_344 (O_344,N_2316,N_2897);
or UO_345 (O_345,N_2554,N_2088);
nor UO_346 (O_346,N_2703,N_2629);
or UO_347 (O_347,N_2447,N_2580);
nor UO_348 (O_348,N_2108,N_2611);
nor UO_349 (O_349,N_2248,N_2126);
nand UO_350 (O_350,N_2038,N_2236);
and UO_351 (O_351,N_2184,N_2083);
xnor UO_352 (O_352,N_2395,N_2336);
xor UO_353 (O_353,N_2669,N_2514);
or UO_354 (O_354,N_2982,N_2966);
nand UO_355 (O_355,N_2844,N_2783);
or UO_356 (O_356,N_2958,N_2223);
xnor UO_357 (O_357,N_2207,N_2116);
and UO_358 (O_358,N_2347,N_2659);
nor UO_359 (O_359,N_2921,N_2318);
and UO_360 (O_360,N_2021,N_2732);
and UO_361 (O_361,N_2213,N_2647);
nand UO_362 (O_362,N_2607,N_2272);
or UO_363 (O_363,N_2927,N_2030);
or UO_364 (O_364,N_2974,N_2099);
nand UO_365 (O_365,N_2984,N_2919);
and UO_366 (O_366,N_2577,N_2445);
nor UO_367 (O_367,N_2486,N_2075);
xnor UO_368 (O_368,N_2829,N_2983);
and UO_369 (O_369,N_2154,N_2216);
or UO_370 (O_370,N_2429,N_2461);
or UO_371 (O_371,N_2902,N_2077);
and UO_372 (O_372,N_2004,N_2071);
or UO_373 (O_373,N_2294,N_2469);
and UO_374 (O_374,N_2145,N_2296);
nand UO_375 (O_375,N_2225,N_2024);
nor UO_376 (O_376,N_2135,N_2874);
nand UO_377 (O_377,N_2087,N_2247);
nand UO_378 (O_378,N_2986,N_2313);
nor UO_379 (O_379,N_2515,N_2838);
and UO_380 (O_380,N_2041,N_2884);
nand UO_381 (O_381,N_2622,N_2319);
nand UO_382 (O_382,N_2494,N_2143);
nor UO_383 (O_383,N_2863,N_2773);
nand UO_384 (O_384,N_2265,N_2167);
and UO_385 (O_385,N_2409,N_2408);
or UO_386 (O_386,N_2563,N_2297);
nand UO_387 (O_387,N_2470,N_2107);
xor UO_388 (O_388,N_2856,N_2959);
nor UO_389 (O_389,N_2615,N_2745);
nand UO_390 (O_390,N_2303,N_2895);
or UO_391 (O_391,N_2846,N_2851);
and UO_392 (O_392,N_2525,N_2627);
xnor UO_393 (O_393,N_2928,N_2332);
nand UO_394 (O_394,N_2110,N_2714);
nor UO_395 (O_395,N_2518,N_2491);
nor UO_396 (O_396,N_2376,N_2523);
xnor UO_397 (O_397,N_2713,N_2165);
and UO_398 (O_398,N_2968,N_2276);
nor UO_399 (O_399,N_2803,N_2229);
xor UO_400 (O_400,N_2185,N_2616);
nand UO_401 (O_401,N_2680,N_2198);
and UO_402 (O_402,N_2046,N_2262);
and UO_403 (O_403,N_2552,N_2717);
or UO_404 (O_404,N_2398,N_2017);
nand UO_405 (O_405,N_2119,N_2466);
nand UO_406 (O_406,N_2951,N_2978);
and UO_407 (O_407,N_2944,N_2787);
nor UO_408 (O_408,N_2620,N_2567);
nand UO_409 (O_409,N_2516,N_2414);
xnor UO_410 (O_410,N_2643,N_2275);
and UO_411 (O_411,N_2054,N_2214);
and UO_412 (O_412,N_2105,N_2623);
nor UO_413 (O_413,N_2492,N_2384);
xnor UO_414 (O_414,N_2600,N_2367);
or UO_415 (O_415,N_2903,N_2121);
xnor UO_416 (O_416,N_2437,N_2678);
nand UO_417 (O_417,N_2446,N_2081);
and UO_418 (O_418,N_2721,N_2672);
nand UO_419 (O_419,N_2287,N_2509);
xnor UO_420 (O_420,N_2233,N_2828);
and UO_421 (O_421,N_2952,N_2211);
nor UO_422 (O_422,N_2882,N_2788);
nor UO_423 (O_423,N_2477,N_2936);
nor UO_424 (O_424,N_2454,N_2871);
and UO_425 (O_425,N_2538,N_2432);
and UO_426 (O_426,N_2161,N_2832);
and UO_427 (O_427,N_2003,N_2977);
and UO_428 (O_428,N_2700,N_2990);
nor UO_429 (O_429,N_2020,N_2113);
nor UO_430 (O_430,N_2621,N_2862);
and UO_431 (O_431,N_2731,N_2727);
nor UO_432 (O_432,N_2348,N_2752);
or UO_433 (O_433,N_2636,N_2106);
or UO_434 (O_434,N_2155,N_2861);
nor UO_435 (O_435,N_2535,N_2800);
nor UO_436 (O_436,N_2693,N_2566);
nor UO_437 (O_437,N_2010,N_2027);
nand UO_438 (O_438,N_2320,N_2049);
and UO_439 (O_439,N_2279,N_2069);
or UO_440 (O_440,N_2280,N_2920);
xor UO_441 (O_441,N_2583,N_2533);
nor UO_442 (O_442,N_2159,N_2175);
or UO_443 (O_443,N_2545,N_2747);
xnor UO_444 (O_444,N_2963,N_2208);
and UO_445 (O_445,N_2244,N_2957);
nand UO_446 (O_446,N_2394,N_2444);
or UO_447 (O_447,N_2433,N_2388);
or UO_448 (O_448,N_2212,N_2339);
and UO_449 (O_449,N_2791,N_2590);
and UO_450 (O_450,N_2564,N_2392);
nor UO_451 (O_451,N_2457,N_2286);
and UO_452 (O_452,N_2917,N_2601);
or UO_453 (O_453,N_2368,N_2697);
nand UO_454 (O_454,N_2101,N_2097);
nand UO_455 (O_455,N_2873,N_2744);
nor UO_456 (O_456,N_2822,N_2111);
nor UO_457 (O_457,N_2833,N_2495);
xnor UO_458 (O_458,N_2694,N_2193);
nor UO_459 (O_459,N_2667,N_2330);
nor UO_460 (O_460,N_2879,N_2104);
or UO_461 (O_461,N_2082,N_2543);
nor UO_462 (O_462,N_2912,N_2767);
or UO_463 (O_463,N_2926,N_2872);
and UO_464 (O_464,N_2573,N_2133);
nor UO_465 (O_465,N_2778,N_2644);
nor UO_466 (O_466,N_2317,N_2532);
nor UO_467 (O_467,N_2508,N_2267);
or UO_468 (O_468,N_2241,N_2994);
or UO_469 (O_469,N_2277,N_2195);
or UO_470 (O_470,N_2288,N_2274);
or UO_471 (O_471,N_2399,N_2378);
or UO_472 (O_472,N_2961,N_2799);
or UO_473 (O_473,N_2221,N_2817);
or UO_474 (O_474,N_2187,N_2578);
or UO_475 (O_475,N_2571,N_2147);
nor UO_476 (O_476,N_2826,N_2652);
nand UO_477 (O_477,N_2122,N_2734);
xnor UO_478 (O_478,N_2201,N_2909);
and UO_479 (O_479,N_2031,N_2548);
nand UO_480 (O_480,N_2426,N_2130);
and UO_481 (O_481,N_2146,N_2812);
nor UO_482 (O_482,N_2576,N_2411);
and UO_483 (O_483,N_2227,N_2827);
or UO_484 (O_484,N_2166,N_2955);
xnor UO_485 (O_485,N_2489,N_2109);
nand UO_486 (O_486,N_2173,N_2766);
and UO_487 (O_487,N_2979,N_2413);
or UO_488 (O_488,N_2283,N_2710);
nand UO_489 (O_489,N_2463,N_2849);
nor UO_490 (O_490,N_2596,N_2711);
nand UO_491 (O_491,N_2002,N_2383);
xor UO_492 (O_492,N_2363,N_2502);
nand UO_493 (O_493,N_2820,N_2497);
and UO_494 (O_494,N_2406,N_2289);
and UO_495 (O_495,N_2877,N_2085);
nor UO_496 (O_496,N_2628,N_2907);
and UO_497 (O_497,N_2906,N_2619);
xor UO_498 (O_498,N_2904,N_2034);
and UO_499 (O_499,N_2568,N_2156);
endmodule