module basic_2000_20000_2500_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_157,In_300);
xor U1 (N_1,In_52,In_1635);
nor U2 (N_2,In_1995,In_586);
or U3 (N_3,In_521,In_140);
and U4 (N_4,In_516,In_1082);
nor U5 (N_5,In_874,In_1420);
or U6 (N_6,In_1352,In_1592);
nand U7 (N_7,In_452,In_1699);
or U8 (N_8,In_371,In_348);
nor U9 (N_9,In_724,In_1717);
nor U10 (N_10,In_396,In_1353);
or U11 (N_11,In_70,In_1528);
nand U12 (N_12,In_962,In_675);
and U13 (N_13,In_109,In_1093);
and U14 (N_14,In_957,In_856);
nor U15 (N_15,In_1524,In_1697);
xnor U16 (N_16,In_1614,In_1870);
and U17 (N_17,In_1947,In_459);
nor U18 (N_18,In_1006,In_1398);
xor U19 (N_19,In_794,In_1465);
nand U20 (N_20,In_15,In_1990);
and U21 (N_21,In_583,In_1944);
xnor U22 (N_22,In_515,In_935);
nand U23 (N_23,In_1847,In_118);
nand U24 (N_24,In_872,In_863);
nand U25 (N_25,In_661,In_295);
and U26 (N_26,In_1732,In_1129);
or U27 (N_27,In_1103,In_1652);
nor U28 (N_28,In_1919,In_1740);
or U29 (N_29,In_1039,In_1135);
nor U30 (N_30,In_153,In_254);
or U31 (N_31,In_1337,In_623);
and U32 (N_32,In_1473,In_734);
or U33 (N_33,In_106,In_400);
xnor U34 (N_34,In_1609,In_1536);
or U35 (N_35,In_1974,In_242);
or U36 (N_36,In_479,In_1704);
nand U37 (N_37,In_1326,In_318);
nand U38 (N_38,In_87,In_1969);
nand U39 (N_39,In_1375,In_510);
or U40 (N_40,In_1387,In_1959);
xor U41 (N_41,In_893,In_575);
nor U42 (N_42,In_1727,In_1053);
and U43 (N_43,In_548,In_1810);
and U44 (N_44,In_1767,In_220);
nor U45 (N_45,In_1071,In_223);
xor U46 (N_46,In_1057,In_438);
and U47 (N_47,In_1126,In_1456);
nand U48 (N_48,In_1687,In_1922);
and U49 (N_49,In_687,In_145);
nand U50 (N_50,In_264,In_782);
nor U51 (N_51,In_1920,In_85);
xor U52 (N_52,In_977,In_889);
nor U53 (N_53,In_232,In_78);
or U54 (N_54,In_466,In_1940);
nand U55 (N_55,In_244,In_1662);
nor U56 (N_56,In_1745,In_439);
or U57 (N_57,In_156,In_595);
or U58 (N_58,In_308,In_776);
and U59 (N_59,In_1871,In_394);
or U60 (N_60,In_1065,In_382);
xnor U61 (N_61,In_21,In_1038);
nor U62 (N_62,In_1162,In_1855);
nand U63 (N_63,In_1265,In_1440);
or U64 (N_64,In_370,In_130);
nor U65 (N_65,In_1287,In_317);
nand U66 (N_66,In_1088,In_1030);
nor U67 (N_67,In_496,In_128);
nand U68 (N_68,In_1410,In_557);
and U69 (N_69,In_955,In_1522);
xnor U70 (N_70,In_1333,In_1453);
and U71 (N_71,In_76,In_1862);
nor U72 (N_72,In_1642,In_1820);
and U73 (N_73,In_1497,In_1393);
xnor U74 (N_74,In_816,In_1963);
or U75 (N_75,In_1016,In_1324);
and U76 (N_76,In_468,In_288);
nor U77 (N_77,In_1476,In_947);
or U78 (N_78,In_77,In_1683);
nor U79 (N_79,In_1489,In_1252);
and U80 (N_80,In_658,In_450);
and U81 (N_81,In_34,In_455);
nand U82 (N_82,In_171,In_427);
nand U83 (N_83,In_1828,In_1939);
nand U84 (N_84,In_1112,In_234);
xor U85 (N_85,In_1827,In_179);
nor U86 (N_86,In_1094,In_218);
xor U87 (N_87,In_255,In_596);
nand U88 (N_88,In_131,In_174);
and U89 (N_89,In_1396,In_1421);
xnor U90 (N_90,In_1452,In_885);
xnor U91 (N_91,In_1728,In_1354);
nor U92 (N_92,In_123,In_1208);
and U93 (N_93,In_1150,In_1293);
and U94 (N_94,In_1183,In_347);
nand U95 (N_95,In_344,In_941);
and U96 (N_96,In_1599,In_1160);
nand U97 (N_97,In_667,In_1863);
nor U98 (N_98,In_748,In_681);
xor U99 (N_99,In_670,In_587);
xnor U100 (N_100,In_1673,In_1931);
or U101 (N_101,In_895,In_1665);
nand U102 (N_102,In_192,In_737);
or U103 (N_103,In_1374,In_97);
and U104 (N_104,In_48,In_1807);
and U105 (N_105,In_1554,In_789);
and U106 (N_106,In_1432,In_208);
nor U107 (N_107,In_688,In_1679);
xnor U108 (N_108,In_1917,In_1362);
nand U109 (N_109,In_1022,In_907);
nor U110 (N_110,In_1884,In_716);
nor U111 (N_111,In_936,In_475);
xnor U112 (N_112,In_3,In_1641);
or U113 (N_113,In_451,In_817);
or U114 (N_114,In_473,In_1534);
nand U115 (N_115,In_804,In_840);
nor U116 (N_116,In_1175,In_1461);
nand U117 (N_117,In_1838,In_1546);
nand U118 (N_118,In_119,In_1466);
xor U119 (N_119,In_531,In_1230);
nor U120 (N_120,In_666,In_321);
and U121 (N_121,In_188,In_126);
xnor U122 (N_122,In_1986,In_1760);
or U123 (N_123,In_1334,In_1253);
xor U124 (N_124,In_701,In_1753);
nand U125 (N_125,In_1806,In_1189);
nand U126 (N_126,In_1771,In_559);
xor U127 (N_127,In_967,In_960);
or U128 (N_128,In_1493,In_1992);
and U129 (N_129,In_1226,In_704);
nor U130 (N_130,In_1236,In_1729);
nand U131 (N_131,In_80,In_1779);
nand U132 (N_132,In_1224,In_378);
xor U133 (N_133,In_1074,In_831);
and U134 (N_134,In_942,In_10);
nand U135 (N_135,In_913,In_229);
and U136 (N_136,In_779,In_1267);
and U137 (N_137,In_993,In_1164);
or U138 (N_138,In_1763,In_855);
and U139 (N_139,In_1765,In_1243);
xor U140 (N_140,In_1210,In_965);
and U141 (N_141,In_564,In_1594);
nand U142 (N_142,In_454,In_339);
nand U143 (N_143,In_1975,In_26);
and U144 (N_144,In_115,In_671);
xor U145 (N_145,In_1613,In_607);
or U146 (N_146,In_983,In_576);
or U147 (N_147,In_1902,In_281);
and U148 (N_148,In_602,In_1297);
xnor U149 (N_149,In_1882,In_1171);
nor U150 (N_150,In_968,In_1589);
or U151 (N_151,In_1711,In_4);
nor U152 (N_152,In_530,In_245);
xnor U153 (N_153,In_110,In_1842);
xor U154 (N_154,In_1789,In_383);
and U155 (N_155,In_1218,In_1706);
and U156 (N_156,In_618,In_273);
nor U157 (N_157,In_1597,In_922);
or U158 (N_158,In_762,In_642);
nand U159 (N_159,In_702,In_172);
nand U160 (N_160,In_1301,In_517);
or U161 (N_161,In_127,In_1887);
nand U162 (N_162,In_1626,In_1719);
xnor U163 (N_163,In_163,In_1621);
xnor U164 (N_164,In_1978,In_198);
nor U165 (N_165,In_176,In_235);
nand U166 (N_166,In_1379,In_37);
xor U167 (N_167,In_945,In_1743);
nand U168 (N_168,In_937,In_1075);
nand U169 (N_169,In_205,In_259);
or U170 (N_170,In_1068,In_1303);
and U171 (N_171,In_565,In_1705);
xnor U172 (N_172,In_1795,In_1272);
nor U173 (N_173,In_1018,In_1754);
nor U174 (N_174,In_134,In_1904);
nor U175 (N_175,In_801,In_1143);
nand U176 (N_176,In_1369,In_585);
xnor U177 (N_177,In_665,In_1217);
nor U178 (N_178,In_1013,In_566);
and U179 (N_179,In_89,In_1624);
and U180 (N_180,In_1105,In_1858);
nand U181 (N_181,In_703,In_851);
or U182 (N_182,In_1578,In_270);
or U183 (N_183,In_1158,In_16);
or U184 (N_184,In_543,In_66);
or U185 (N_185,In_1487,In_1535);
and U186 (N_186,In_59,In_1181);
nor U187 (N_187,In_1390,In_1401);
or U188 (N_188,In_1012,In_714);
and U189 (N_189,In_546,In_750);
nand U190 (N_190,In_568,In_946);
nor U191 (N_191,In_1099,In_1320);
and U192 (N_192,In_726,In_1304);
or U193 (N_193,In_64,In_1223);
nand U194 (N_194,In_973,In_753);
nand U195 (N_195,In_732,In_833);
or U196 (N_196,In_1721,In_307);
or U197 (N_197,In_1238,In_470);
or U198 (N_198,In_843,In_1394);
or U199 (N_199,In_940,In_492);
or U200 (N_200,In_1259,In_1197);
nand U201 (N_201,In_165,In_303);
nor U202 (N_202,In_579,In_1734);
or U203 (N_203,In_1331,In_1671);
and U204 (N_204,In_465,In_1824);
and U205 (N_205,In_249,In_177);
or U206 (N_206,In_1176,In_1058);
nand U207 (N_207,In_1319,In_323);
nand U208 (N_208,In_1428,In_1967);
nor U209 (N_209,In_857,In_1108);
and U210 (N_210,In_436,In_1646);
or U211 (N_211,In_33,In_632);
or U212 (N_212,In_98,In_1868);
or U213 (N_213,In_1182,In_1214);
nand U214 (N_214,In_1669,In_99);
nor U215 (N_215,In_201,In_1172);
or U216 (N_216,In_1233,In_1101);
xor U217 (N_217,In_1275,In_739);
xor U218 (N_218,In_1072,In_1141);
and U219 (N_219,In_669,In_1376);
xor U220 (N_220,In_614,In_1908);
xor U221 (N_221,In_1231,In_409);
nor U222 (N_222,In_482,In_590);
nand U223 (N_223,In_164,In_1332);
and U224 (N_224,In_353,In_1933);
and U225 (N_225,In_1104,In_1695);
nand U226 (N_226,In_100,In_1981);
and U227 (N_227,In_214,In_886);
nand U228 (N_228,In_637,In_181);
xor U229 (N_229,In_712,In_1268);
nand U230 (N_230,In_194,In_810);
nor U231 (N_231,In_803,In_1564);
and U232 (N_232,In_1895,In_340);
nor U233 (N_233,In_178,In_1366);
nor U234 (N_234,In_631,In_1349);
nand U235 (N_235,In_562,In_368);
nor U236 (N_236,In_221,In_360);
and U237 (N_237,In_1288,In_1144);
xnor U238 (N_238,In_293,In_639);
nor U239 (N_239,In_297,In_1755);
and U240 (N_240,In_1344,In_711);
nand U241 (N_241,In_437,In_897);
nor U242 (N_242,In_1764,In_1644);
nand U243 (N_243,In_662,In_375);
nor U244 (N_244,In_320,In_1980);
and U245 (N_245,In_1741,In_729);
nor U246 (N_246,In_1970,In_1608);
xnor U247 (N_247,In_584,In_1212);
xor U248 (N_248,In_1571,In_1124);
nor U249 (N_249,In_733,In_1431);
xor U250 (N_250,In_362,In_916);
nand U251 (N_251,In_679,In_1911);
xnor U252 (N_252,In_1336,In_755);
xnor U253 (N_253,In_182,In_1234);
or U254 (N_254,In_1888,In_1549);
nand U255 (N_255,In_556,In_812);
nor U256 (N_256,In_405,In_393);
nor U257 (N_257,In_20,In_747);
nand U258 (N_258,In_133,In_351);
and U259 (N_259,In_1110,In_1941);
or U260 (N_260,In_180,In_341);
nand U261 (N_261,In_1423,In_685);
and U262 (N_262,In_535,In_1270);
nor U263 (N_263,In_1508,In_744);
nand U264 (N_264,In_891,In_786);
nand U265 (N_265,In_630,In_1748);
and U266 (N_266,In_219,In_286);
nand U267 (N_267,In_1961,In_252);
or U268 (N_268,In_1467,In_1060);
nand U269 (N_269,In_974,In_979);
or U270 (N_270,In_668,In_1836);
or U271 (N_271,In_1418,In_1165);
xnor U272 (N_272,In_1501,In_1221);
and U273 (N_273,In_1232,In_291);
and U274 (N_274,In_1616,In_1298);
and U275 (N_275,In_1837,In_1);
nand U276 (N_276,In_1693,In_868);
nand U277 (N_277,In_431,In_1523);
and U278 (N_278,In_1503,In_1269);
nor U279 (N_279,In_1676,In_1346);
or U280 (N_280,In_796,In_1159);
xor U281 (N_281,In_1260,In_1627);
or U282 (N_282,In_1169,In_534);
or U283 (N_283,In_1170,In_558);
nand U284 (N_284,In_1985,In_480);
or U285 (N_285,In_1185,In_689);
nand U286 (N_286,In_1296,In_1382);
or U287 (N_287,In_952,In_1485);
and U288 (N_288,In_1548,In_1762);
and U289 (N_289,In_1115,In_1010);
xnor U290 (N_290,In_691,In_283);
and U291 (N_291,In_1347,In_1808);
nor U292 (N_292,In_1912,In_1496);
and U293 (N_293,In_1800,In_1802);
nor U294 (N_294,In_19,In_251);
nor U295 (N_295,In_767,In_1651);
xor U296 (N_296,In_545,In_384);
xor U297 (N_297,In_992,In_1356);
or U298 (N_298,In_832,In_1723);
nor U299 (N_299,In_1483,In_346);
xnor U300 (N_300,In_1591,In_333);
or U301 (N_301,In_659,In_250);
xor U302 (N_302,In_1861,In_299);
and U303 (N_303,In_1562,In_877);
xnor U304 (N_304,In_683,In_800);
nor U305 (N_305,In_92,In_463);
nand U306 (N_306,In_55,In_1315);
xor U307 (N_307,In_1064,In_481);
and U308 (N_308,In_419,In_1814);
or U309 (N_309,In_1604,In_329);
nor U310 (N_310,In_1688,In_1584);
and U311 (N_311,In_700,In_484);
or U312 (N_312,In_445,In_905);
xnor U313 (N_313,In_1419,In_1195);
xnor U314 (N_314,In_1161,In_1459);
and U315 (N_315,In_1874,In_961);
and U316 (N_316,In_723,In_386);
nor U317 (N_317,In_1752,In_908);
xor U318 (N_318,In_483,In_90);
or U319 (N_319,In_412,In_1803);
nand U320 (N_320,In_598,In_1063);
nand U321 (N_321,In_1738,In_862);
xor U322 (N_322,In_61,In_67);
and U323 (N_323,In_1282,In_1610);
nand U324 (N_324,In_939,In_697);
nor U325 (N_325,In_190,In_1650);
or U326 (N_326,In_988,In_1632);
or U327 (N_327,In_969,In_1623);
nor U328 (N_328,In_253,In_376);
or U329 (N_329,In_207,In_1775);
xnor U330 (N_330,In_985,In_1736);
or U331 (N_331,In_1994,In_1251);
xor U332 (N_332,In_603,In_1574);
nand U333 (N_333,In_883,In_1425);
or U334 (N_334,In_1345,In_1935);
nor U335 (N_335,In_853,In_1817);
nand U336 (N_336,In_953,In_1527);
or U337 (N_337,In_336,In_11);
and U338 (N_338,In_674,In_1015);
and U339 (N_339,In_616,In_417);
or U340 (N_340,In_1153,In_316);
nor U341 (N_341,In_1426,In_1950);
nor U342 (N_342,In_1749,In_1516);
nand U343 (N_343,In_997,In_1097);
nor U344 (N_344,In_1383,In_1271);
and U345 (N_345,In_95,In_1844);
nand U346 (N_346,In_1948,In_228);
nand U347 (N_347,In_276,In_1629);
xor U348 (N_348,In_696,In_1102);
xnor U349 (N_349,In_1184,In_440);
nand U350 (N_350,In_1377,In_783);
or U351 (N_351,In_1831,In_301);
and U352 (N_352,In_1913,In_442);
nand U353 (N_353,In_772,In_699);
xnor U354 (N_354,In_655,In_571);
xnor U355 (N_355,In_151,In_1849);
xor U356 (N_356,In_1696,In_1631);
or U357 (N_357,In_124,In_1883);
and U358 (N_358,In_5,In_524);
or U359 (N_359,In_121,In_1330);
and U360 (N_360,In_673,In_934);
and U361 (N_361,In_1596,In_764);
nor U362 (N_362,In_995,In_1403);
xnor U363 (N_363,In_1569,In_589);
xor U364 (N_364,In_1285,In_1113);
nor U365 (N_365,In_1953,In_1540);
xor U366 (N_366,In_322,In_453);
nand U367 (N_367,In_196,In_1017);
nand U368 (N_368,In_1859,In_1077);
nor U369 (N_369,In_1323,In_765);
or U370 (N_370,In_1742,In_1885);
and U371 (N_371,In_1648,In_41);
and U372 (N_372,In_1279,In_391);
xor U373 (N_373,In_1019,In_330);
or U374 (N_374,In_240,In_788);
nand U375 (N_375,In_415,In_197);
and U376 (N_376,In_651,In_1843);
and U377 (N_377,In_785,In_1951);
xnor U378 (N_378,In_808,In_821);
nor U379 (N_379,In_1921,In_797);
nor U380 (N_380,In_1056,In_1167);
nor U381 (N_381,In_806,In_1095);
xor U382 (N_382,In_918,In_469);
nand U383 (N_383,In_1388,In_1694);
xor U384 (N_384,In_1890,In_628);
xor U385 (N_385,In_111,In_108);
nand U386 (N_386,In_1580,In_925);
or U387 (N_387,In_313,In_433);
nor U388 (N_388,In_101,In_924);
xnor U389 (N_389,In_870,In_1000);
or U390 (N_390,In_1875,In_999);
nand U391 (N_391,In_63,In_1080);
nor U392 (N_392,In_476,In_512);
nor U393 (N_393,In_1768,In_741);
and U394 (N_394,In_1772,In_1338);
nand U395 (N_395,In_514,In_1001);
nand U396 (N_396,In_1027,In_643);
xnor U397 (N_397,In_650,In_1850);
and U398 (N_398,In_1114,In_1905);
and U399 (N_399,In_331,In_1942);
nand U400 (N_400,In_22,In_1313);
xnor U401 (N_401,In_1261,In_1916);
xnor U402 (N_402,In_1712,In_1051);
nand U403 (N_403,In_1138,In_1965);
nand U404 (N_404,In_305,In_200);
and U405 (N_405,In_392,In_1906);
xor U406 (N_406,In_1145,In_1826);
nand U407 (N_407,In_1494,In_791);
or U408 (N_408,In_413,In_1096);
or U409 (N_409,In_170,In_257);
or U410 (N_410,In_46,In_1537);
nor U411 (N_411,In_1146,In_756);
nor U412 (N_412,In_1405,In_1718);
or U413 (N_413,In_1305,In_763);
xor U414 (N_414,In_267,In_599);
xor U415 (N_415,In_1896,In_69);
xnor U416 (N_416,In_1770,In_68);
or U417 (N_417,In_1543,In_1774);
nand U418 (N_418,In_792,In_807);
and U419 (N_419,In_1378,In_1823);
or U420 (N_420,In_1500,In_148);
nand U421 (N_421,In_1668,In_1923);
and U422 (N_422,In_943,In_1555);
nand U423 (N_423,In_1188,In_422);
or U424 (N_424,In_577,In_1934);
or U425 (N_425,In_719,In_93);
or U426 (N_426,In_1989,In_625);
nor U427 (N_427,In_7,In_1449);
nor U428 (N_428,In_1321,In_1825);
or U429 (N_429,In_1411,In_781);
or U430 (N_430,In_1131,In_608);
xor U431 (N_431,In_1776,In_715);
nor U432 (N_432,In_1044,In_1550);
or U433 (N_433,In_406,In_407);
or U434 (N_434,In_1299,In_410);
xor U435 (N_435,In_29,In_835);
nand U436 (N_436,In_1120,In_1525);
or U437 (N_437,In_561,In_211);
nor U438 (N_438,In_154,In_441);
nor U439 (N_439,In_206,In_162);
or U440 (N_440,In_397,In_224);
nand U441 (N_441,In_636,In_275);
nor U442 (N_442,In_1155,In_1028);
and U443 (N_443,In_284,In_1385);
and U444 (N_444,In_1661,In_705);
xnor U445 (N_445,In_1792,In_745);
or U446 (N_446,In_1083,In_1869);
or U447 (N_447,In_828,In_256);
or U448 (N_448,In_660,In_1539);
and U449 (N_449,In_1227,In_1892);
and U450 (N_450,In_1470,In_1572);
or U451 (N_451,In_1193,In_51);
nand U452 (N_452,In_146,In_1122);
or U453 (N_453,In_1241,In_981);
and U454 (N_454,In_1225,In_1482);
xor U455 (N_455,In_58,In_186);
xor U456 (N_456,In_1907,In_1515);
nor U457 (N_457,In_1180,In_225);
nor U458 (N_458,In_758,In_271);
nand U459 (N_459,In_513,In_457);
or U460 (N_460,In_837,In_147);
and U461 (N_461,In_1045,In_1703);
and U462 (N_462,In_1142,In_1085);
and U463 (N_463,In_462,In_1451);
nor U464 (N_464,In_735,In_903);
and U465 (N_465,In_1373,In_1481);
xnor U466 (N_466,In_1499,In_1450);
nand U467 (N_467,In_1791,In_1702);
or U468 (N_468,In_1972,In_695);
nand U469 (N_469,In_263,In_421);
or U470 (N_470,In_1520,In_1943);
and U471 (N_471,In_954,In_597);
or U472 (N_472,In_91,In_1833);
nand U473 (N_473,In_248,In_495);
xor U474 (N_474,In_418,In_1035);
nor U475 (N_475,In_277,In_1340);
or U476 (N_476,In_629,In_1812);
nor U477 (N_477,In_1049,In_648);
nand U478 (N_478,In_949,In_357);
nand U479 (N_479,In_1603,In_617);
and U480 (N_480,In_1203,In_921);
or U481 (N_481,In_841,In_527);
nand U482 (N_482,In_28,In_551);
or U483 (N_483,In_1945,In_1198);
nand U484 (N_484,In_434,In_580);
nor U485 (N_485,In_149,In_1325);
and U486 (N_486,In_1707,In_487);
nor U487 (N_487,In_202,In_47);
nor U488 (N_488,In_1878,In_1292);
nand U489 (N_489,In_1168,In_1590);
and U490 (N_490,In_1645,In_1316);
nand U491 (N_491,In_570,In_1794);
or U492 (N_492,In_672,In_743);
nand U493 (N_493,In_302,In_60);
xor U494 (N_494,In_994,In_1746);
or U495 (N_495,In_644,In_1544);
or U496 (N_496,In_1698,In_166);
or U497 (N_497,In_1048,In_216);
nand U498 (N_498,In_823,In_167);
nor U499 (N_499,In_1200,In_1587);
xnor U500 (N_500,In_1041,In_1686);
xor U501 (N_501,In_1462,In_1491);
nor U502 (N_502,In_1036,In_1134);
and U503 (N_503,In_829,In_1533);
or U504 (N_504,In_1722,In_183);
nor U505 (N_505,In_38,In_1936);
or U506 (N_506,In_1342,In_1486);
or U507 (N_507,In_88,In_1713);
nand U508 (N_508,In_1894,In_1506);
or U509 (N_509,In_1715,In_1607);
nand U510 (N_510,In_1778,In_1598);
nand U511 (N_511,In_1443,In_731);
nor U512 (N_512,In_1435,In_444);
or U513 (N_513,In_1274,In_1682);
nand U514 (N_514,In_1903,In_79);
and U515 (N_515,In_1365,In_1938);
and U516 (N_516,In_684,In_1512);
or U517 (N_517,In_464,In_1620);
xnor U518 (N_518,In_1625,In_1518);
or U519 (N_519,In_775,In_1918);
xnor U520 (N_520,In_81,In_613);
nand U521 (N_521,In_1979,In_1005);
and U522 (N_522,In_1372,In_555);
xor U523 (N_523,In_847,In_826);
and U524 (N_524,In_621,In_900);
nand U525 (N_525,In_342,In_114);
nor U526 (N_526,In_1566,In_1196);
nor U527 (N_527,In_365,In_845);
nor U528 (N_528,In_591,In_1242);
xor U529 (N_529,In_986,In_1593);
xor U530 (N_530,In_1343,In_290);
nand U531 (N_531,In_1192,In_1612);
xor U532 (N_532,In_1628,In_1585);
nand U533 (N_533,In_1222,In_1559);
xor U534 (N_534,In_718,In_1829);
and U535 (N_535,In_710,In_243);
or U536 (N_536,In_1899,In_74);
or U537 (N_537,In_1781,In_324);
nor U538 (N_538,In_1993,In_72);
nor U539 (N_539,In_282,In_1561);
or U540 (N_540,In_1577,In_815);
xor U541 (N_541,In_814,In_203);
or U542 (N_542,In_1886,In_266);
nor U543 (N_543,In_1983,In_83);
xnor U544 (N_544,In_367,In_1438);
nand U545 (N_545,In_472,In_1283);
xor U546 (N_546,In_1790,In_1851);
xor U547 (N_547,In_1684,In_884);
nand U548 (N_548,In_882,In_594);
nor U549 (N_549,In_790,In_998);
and U550 (N_550,In_633,In_873);
and U551 (N_551,In_606,In_1202);
or U552 (N_552,In_1997,In_887);
nor U553 (N_553,In_1355,In_1846);
xor U554 (N_554,In_1955,In_1194);
xnor U555 (N_555,In_560,In_1505);
nand U556 (N_556,In_552,In_722);
or U557 (N_557,In_938,In_125);
or U558 (N_558,In_507,In_611);
and U559 (N_559,In_1551,In_395);
xnor U560 (N_560,In_811,In_377);
nor U561 (N_561,In_519,In_1002);
nand U562 (N_562,In_909,In_1029);
xor U563 (N_563,In_888,In_1724);
or U564 (N_564,In_930,In_113);
nand U565 (N_565,In_498,In_1581);
nand U566 (N_566,In_1307,In_1123);
and U567 (N_567,In_1220,In_1675);
and U568 (N_568,In_1444,In_30);
nor U569 (N_569,In_1893,In_494);
xnor U570 (N_570,In_1530,In_1777);
or U571 (N_571,In_1973,In_1091);
nand U572 (N_572,In_1381,In_420);
xor U573 (N_573,In_1408,In_1249);
nand U574 (N_574,In_31,In_1949);
nor U575 (N_575,In_388,In_296);
nor U576 (N_576,In_261,In_774);
xnor U577 (N_577,In_1617,In_1880);
nor U578 (N_578,In_1284,In_866);
nor U579 (N_579,In_1787,In_1341);
xor U580 (N_580,In_1720,In_1186);
nand U581 (N_581,In_1084,In_1174);
and U582 (N_582,In_1925,In_1213);
xor U583 (N_583,In_898,In_1689);
nand U584 (N_584,In_1132,In_1455);
or U585 (N_585,In_760,In_708);
and U586 (N_586,In_653,In_485);
or U587 (N_587,In_865,In_359);
and U588 (N_588,In_12,In_861);
xnor U589 (N_589,In_757,In_1128);
nor U590 (N_590,In_1678,In_1576);
nor U591 (N_591,In_1239,In_859);
and U592 (N_592,In_1025,In_1910);
or U593 (N_593,In_553,In_759);
or U594 (N_594,In_210,In_1240);
nor U595 (N_595,In_541,In_522);
or U596 (N_596,In_447,In_1228);
xor U597 (N_597,In_443,In_1109);
nor U598 (N_598,In_1758,In_75);
nor U599 (N_599,In_1475,In_610);
or U600 (N_600,In_57,In_740);
and U601 (N_601,In_1424,In_1111);
nand U602 (N_602,In_285,In_247);
or U603 (N_603,In_1206,In_448);
nor U604 (N_604,In_24,In_1579);
and U605 (N_605,In_1414,In_361);
nor U606 (N_606,In_1988,In_802);
nor U607 (N_607,In_899,In_1266);
nor U608 (N_608,In_523,In_902);
and U609 (N_609,In_1464,In_634);
nand U610 (N_610,In_104,In_429);
nand U611 (N_611,In_1647,In_25);
nor U612 (N_612,In_168,In_1291);
or U613 (N_613,In_1602,In_96);
nand U614 (N_614,In_686,In_1670);
xor U615 (N_615,In_1783,In_1448);
and U616 (N_616,In_1964,In_780);
or U617 (N_617,In_1046,In_73);
or U618 (N_618,In_195,In_71);
or U619 (N_619,In_825,In_278);
nor U620 (N_620,In_1956,In_915);
or U621 (N_621,In_1976,In_1649);
nand U622 (N_622,In_720,In_1107);
xnor U623 (N_623,In_17,In_272);
xor U624 (N_624,In_944,In_1009);
xor U625 (N_625,In_236,In_1835);
nor U626 (N_626,In_1773,In_191);
xor U627 (N_627,In_1509,In_500);
xor U628 (N_628,In_1469,In_1066);
nor U629 (N_629,In_622,In_1857);
xor U630 (N_630,In_1119,In_1630);
nand U631 (N_631,In_1205,In_1553);
xnor U632 (N_632,In_350,In_1422);
xor U633 (N_633,In_518,In_528);
nor U634 (N_634,In_638,In_227);
nand U635 (N_635,In_948,In_1092);
and U636 (N_636,In_1657,In_503);
xnor U637 (N_637,In_635,In_260);
and U638 (N_638,In_1034,In_645);
or U639 (N_639,In_1457,In_1690);
nor U640 (N_640,In_49,In_1257);
xor U641 (N_641,In_1417,In_526);
or U642 (N_642,In_707,In_499);
xor U643 (N_643,In_477,In_795);
nor U644 (N_644,In_1759,In_1805);
and U645 (N_645,In_423,In_1519);
nand U646 (N_646,In_910,In_1042);
xnor U647 (N_647,In_1788,In_1127);
and U648 (N_648,In_1701,In_1380);
nand U649 (N_649,In_36,In_403);
nor U650 (N_650,In_920,In_919);
xnor U651 (N_651,In_1477,In_567);
and U652 (N_652,In_1560,In_1819);
nand U653 (N_653,In_975,In_1557);
nand U654 (N_654,In_231,In_23);
nor U655 (N_655,In_1659,In_1492);
nor U656 (N_656,In_1666,In_1757);
nor U657 (N_657,In_850,In_1575);
nor U658 (N_658,In_1570,In_258);
nor U659 (N_659,In_1258,In_1937);
and U660 (N_660,In_1306,In_1327);
xor U661 (N_661,In_694,In_1495);
or U662 (N_662,In_1932,In_1078);
nand U663 (N_663,In_615,In_1310);
and U664 (N_664,In_1490,In_1600);
nand U665 (N_665,In_1339,In_860);
and U666 (N_666,In_1619,In_1430);
nor U667 (N_667,In_1139,In_294);
or U668 (N_668,In_458,In_1809);
and U669 (N_669,In_972,In_959);
xor U670 (N_670,In_1709,In_770);
nand U671 (N_671,In_489,In_355);
xor U672 (N_672,In_328,In_1395);
and U673 (N_673,In_1219,In_1137);
nand U674 (N_674,In_1361,In_1840);
nor U675 (N_675,In_325,In_1052);
xnor U676 (N_676,In_354,In_1839);
nand U677 (N_677,In_572,In_917);
nor U678 (N_678,In_601,In_1478);
nor U679 (N_679,In_573,In_337);
nand U680 (N_680,In_369,In_150);
or U681 (N_681,In_996,In_416);
nand U682 (N_682,In_45,In_1914);
and U683 (N_683,In_1502,In_1348);
xnor U684 (N_684,In_509,In_193);
nand U685 (N_685,In_1148,In_117);
and U686 (N_686,In_213,In_1363);
or U687 (N_687,In_1402,In_1853);
xor U688 (N_688,In_582,In_1416);
nor U689 (N_689,In_1474,In_1007);
xor U690 (N_690,In_1924,In_749);
xnor U691 (N_691,In_1930,In_612);
nand U692 (N_692,In_204,In_746);
and U693 (N_693,In_1215,In_1601);
and U694 (N_694,In_239,In_1565);
nand U695 (N_695,In_1639,In_1636);
nand U696 (N_696,In_1680,In_677);
nand U697 (N_697,In_1946,In_460);
or U698 (N_698,In_736,In_554);
nand U699 (N_699,In_1308,In_950);
xor U700 (N_700,In_399,In_690);
and U701 (N_701,In_1011,In_1458);
nor U702 (N_702,In_1484,In_1998);
xnor U703 (N_703,In_449,In_1247);
nor U704 (N_704,In_752,In_2);
or U705 (N_705,In_1076,In_1716);
and U706 (N_706,In_262,In_141);
or U707 (N_707,In_1118,In_1881);
and U708 (N_708,In_890,In_1877);
or U709 (N_709,In_1664,In_1412);
xnor U710 (N_710,In_1061,In_1656);
xnor U711 (N_711,In_827,In_1404);
nand U712 (N_712,In_425,In_1538);
nor U713 (N_713,In_1653,In_1441);
and U714 (N_714,In_467,In_1798);
nor U715 (N_715,In_246,In_1116);
nor U716 (N_716,In_1898,In_1351);
nand U717 (N_717,In_1434,In_692);
or U718 (N_718,In_1179,In_604);
and U719 (N_719,In_768,In_120);
or U720 (N_720,In_1317,In_289);
xor U721 (N_721,In_1087,In_1460);
or U722 (N_722,In_838,In_1860);
xnor U723 (N_723,In_408,In_238);
nand U724 (N_724,In_678,In_505);
xnor U725 (N_725,In_846,In_1360);
or U726 (N_726,In_1573,In_310);
and U727 (N_727,In_1386,In_569);
nor U728 (N_728,In_1731,In_1856);
nand U729 (N_729,In_199,In_706);
nand U730 (N_730,In_1445,In_144);
and U731 (N_731,In_1400,In_43);
nand U732 (N_732,In_1987,In_1479);
nand U733 (N_733,In_547,In_878);
and U734 (N_734,In_1250,In_32);
and U735 (N_735,In_542,In_830);
or U736 (N_736,In_18,In_1816);
and U737 (N_737,In_1685,In_1446);
nor U738 (N_738,In_881,In_1531);
nand U739 (N_739,In_1278,In_769);
xor U740 (N_740,In_1517,In_414);
and U741 (N_741,In_646,In_1154);
and U742 (N_742,In_327,In_138);
nor U743 (N_743,In_1468,In_1872);
xnor U744 (N_744,In_401,In_544);
and U745 (N_745,In_1854,In_923);
xor U746 (N_746,In_834,In_682);
nand U747 (N_747,In_1793,In_929);
or U748 (N_748,In_536,In_230);
or U749 (N_749,In_1329,In_1003);
nand U750 (N_750,In_173,In_1915);
nor U751 (N_751,In_338,In_132);
nand U752 (N_752,In_1954,In_620);
nor U753 (N_753,In_493,In_461);
nor U754 (N_754,In_1971,In_928);
and U755 (N_755,In_904,In_849);
and U756 (N_756,In_1098,In_428);
xnor U757 (N_757,In_1818,In_1674);
and U758 (N_758,In_1618,In_550);
and U759 (N_759,In_1384,In_1055);
nand U760 (N_760,In_1229,In_1804);
xor U761 (N_761,In_1737,In_1900);
xor U762 (N_762,In_839,In_1615);
nand U763 (N_763,In_848,In_1480);
nor U764 (N_764,In_1929,In_605);
nand U765 (N_765,In_1957,In_298);
and U766 (N_766,In_1047,In_381);
and U767 (N_767,In_1996,In_1409);
or U768 (N_768,In_488,In_292);
xor U769 (N_769,In_279,In_1472);
and U770 (N_770,In_1873,In_1677);
nor U771 (N_771,In_27,In_1568);
nand U772 (N_772,In_432,In_1140);
xnor U773 (N_773,In_269,In_784);
nand U774 (N_774,In_364,In_1436);
xor U775 (N_775,In_486,In_1542);
xor U776 (N_776,In_1442,In_619);
xnor U777 (N_777,In_1514,In_980);
and U778 (N_778,In_1050,In_366);
or U779 (N_779,In_1309,In_1962);
and U780 (N_780,In_892,In_1427);
nand U781 (N_781,In_189,In_549);
nand U782 (N_782,In_738,In_1605);
or U783 (N_783,In_693,In_426);
and U784 (N_784,In_649,In_0);
or U785 (N_785,In_1672,In_1314);
xor U786 (N_786,In_1216,In_1583);
and U787 (N_787,In_158,In_1244);
and U788 (N_788,In_1811,In_717);
nand U789 (N_789,In_1359,In_1952);
or U790 (N_790,In_9,In_155);
nor U791 (N_791,In_754,In_1595);
and U792 (N_792,In_446,In_824);
and U793 (N_793,In_1062,In_540);
and U794 (N_794,In_1190,In_1834);
and U795 (N_795,In_1876,In_1173);
or U796 (N_796,In_987,In_896);
and U797 (N_797,In_869,In_1782);
or U798 (N_798,In_1813,In_1389);
nor U799 (N_799,In_656,In_1879);
and U800 (N_800,In_1177,In_1927);
or U801 (N_801,In_184,In_1841);
xnor U802 (N_802,In_1691,In_112);
nor U803 (N_803,In_1801,In_578);
or U804 (N_804,In_508,In_1660);
xor U805 (N_805,In_217,In_1471);
nand U806 (N_806,In_778,In_520);
xnor U807 (N_807,In_506,In_389);
nor U808 (N_808,In_13,In_1264);
and U809 (N_809,In_588,In_1246);
or U810 (N_810,In_1407,In_1130);
or U811 (N_811,In_1909,In_627);
nor U812 (N_812,In_529,In_1785);
xor U813 (N_813,In_1611,In_1991);
xnor U814 (N_814,In_1552,In_894);
xnor U815 (N_815,In_1033,In_185);
nor U816 (N_816,In_581,In_1406);
nand U817 (N_817,In_713,In_363);
xnor U818 (N_818,In_1867,In_1498);
or U819 (N_819,In_39,In_809);
and U820 (N_820,In_82,In_1008);
and U821 (N_821,In_725,In_1769);
xnor U822 (N_822,In_511,In_349);
and U823 (N_823,In_1799,In_1796);
and U824 (N_824,In_1586,In_777);
nand U825 (N_825,In_1147,In_139);
nand U826 (N_826,In_1043,In_373);
nor U827 (N_827,In_1504,In_761);
and U828 (N_828,In_1311,In_982);
nor U829 (N_829,In_8,In_1290);
or U830 (N_830,In_1822,In_730);
nor U831 (N_831,In_1558,In_574);
and U832 (N_832,In_268,In_1368);
nand U833 (N_833,In_122,In_352);
or U834 (N_834,In_497,In_241);
nor U835 (N_835,In_44,In_129);
nand U836 (N_836,In_116,In_1488);
or U837 (N_837,In_306,In_390);
xnor U838 (N_838,In_1563,In_136);
nor U839 (N_839,In_107,In_1784);
and U840 (N_840,In_435,In_343);
nand U841 (N_841,In_1655,In_50);
and U842 (N_842,In_728,In_1852);
and U843 (N_843,In_663,In_42);
and U844 (N_844,In_1541,In_626);
and U845 (N_845,In_1152,In_1014);
and U846 (N_846,In_35,In_1780);
and U847 (N_847,In_345,In_1766);
nand U848 (N_848,In_742,In_1744);
nand U849 (N_849,In_1897,In_1437);
or U850 (N_850,In_818,In_842);
nand U851 (N_851,In_309,In_358);
nor U852 (N_852,In_1532,In_1606);
nor U853 (N_853,In_319,In_1245);
nand U854 (N_854,In_152,In_1026);
nor U855 (N_855,In_385,In_727);
nor U856 (N_856,In_533,In_914);
xor U857 (N_857,In_1926,In_1207);
xnor U858 (N_858,In_1622,In_1199);
xnor U859 (N_859,In_926,In_1023);
and U860 (N_860,In_525,In_1255);
xor U861 (N_861,In_1725,In_1281);
and U862 (N_862,In_86,In_640);
and U863 (N_863,In_991,In_1262);
nor U864 (N_864,In_1367,In_978);
nor U865 (N_865,In_1507,In_94);
and U866 (N_866,In_1658,In_1889);
or U867 (N_867,In_1276,In_334);
xnor U868 (N_868,In_820,In_398);
or U869 (N_869,In_356,In_1067);
nor U870 (N_870,In_1582,In_374);
nand U871 (N_871,In_1037,In_504);
xnor U872 (N_872,In_402,In_901);
nand U873 (N_873,In_1237,In_1335);
nor U874 (N_874,In_1747,In_1588);
nand U875 (N_875,In_1663,In_1714);
nor U876 (N_876,In_876,In_1370);
nand U877 (N_877,In_1751,In_1726);
nor U878 (N_878,In_430,In_647);
and U879 (N_879,In_805,In_592);
and U880 (N_880,In_532,In_1235);
and U881 (N_881,In_539,In_1090);
or U882 (N_882,In_1739,In_858);
and U883 (N_883,In_1821,In_641);
nand U884 (N_884,In_864,In_1848);
xnor U885 (N_885,In_1106,In_1070);
or U886 (N_886,In_813,In_54);
or U887 (N_887,In_1786,In_490);
and U888 (N_888,In_1750,In_280);
nand U889 (N_889,In_799,In_159);
and U890 (N_890,In_1526,In_1358);
nor U891 (N_891,In_867,In_1521);
nor U892 (N_892,In_215,In_1121);
nand U893 (N_893,In_1392,In_1510);
nor U894 (N_894,In_1413,In_1735);
nor U895 (N_895,In_142,In_287);
nand U896 (N_896,In_880,In_1069);
and U897 (N_897,In_1248,In_135);
nand U898 (N_898,In_1032,In_1364);
nand U899 (N_899,In_222,In_1511);
nor U900 (N_900,In_844,In_1209);
and U901 (N_901,In_1371,In_664);
or U902 (N_902,In_1204,In_1263);
nor U903 (N_903,In_1634,In_879);
and U904 (N_904,In_471,In_53);
xnor U905 (N_905,In_933,In_600);
nand U906 (N_906,In_456,In_474);
xnor U907 (N_907,In_1157,In_65);
nand U908 (N_908,In_1031,In_1254);
or U909 (N_909,In_335,In_676);
nand U910 (N_910,In_563,In_1454);
or U911 (N_911,In_1865,In_609);
nor U912 (N_912,In_766,In_1866);
xnor U913 (N_913,In_1958,In_1891);
nor U914 (N_914,In_1125,In_1201);
nand U915 (N_915,In_971,In_721);
nand U916 (N_916,In_1567,In_1982);
nand U917 (N_917,In_1117,In_1156);
or U918 (N_918,In_1977,In_326);
or U919 (N_919,In_956,In_1312);
nand U920 (N_920,In_1643,In_911);
or U921 (N_921,In_1667,In_233);
or U922 (N_922,In_964,In_990);
and U923 (N_923,In_1681,In_709);
xnor U924 (N_924,In_1322,In_1020);
nor U925 (N_925,In_1756,In_1513);
nor U926 (N_926,In_62,In_927);
nand U927 (N_927,In_14,In_984);
nand U928 (N_928,In_1054,In_912);
xor U929 (N_929,In_274,In_237);
or U930 (N_930,In_1399,In_372);
nor U931 (N_931,In_424,In_1832);
nor U932 (N_932,In_1187,In_906);
nor U933 (N_933,In_1463,In_1700);
and U934 (N_934,In_1638,In_854);
or U935 (N_935,In_963,In_951);
nand U936 (N_936,In_332,In_1984);
nand U937 (N_937,In_1086,In_698);
nor U938 (N_938,In_1295,In_1640);
or U939 (N_939,In_105,In_1191);
and U940 (N_940,In_1300,In_1024);
and U941 (N_941,In_478,In_187);
nor U942 (N_942,In_304,In_1273);
xor U943 (N_943,In_143,In_793);
or U944 (N_944,In_315,In_1692);
xnor U945 (N_945,In_1529,In_209);
or U946 (N_946,In_593,In_538);
or U947 (N_947,In_1136,In_137);
nor U948 (N_948,In_1178,In_1059);
and U949 (N_949,In_836,In_1040);
and U950 (N_950,In_1901,In_1429);
xor U951 (N_951,In_1968,In_1081);
and U952 (N_952,In_1864,In_102);
xnor U953 (N_953,In_932,In_314);
and U954 (N_954,In_1289,In_1830);
nand U955 (N_955,In_379,In_1733);
or U956 (N_956,In_380,In_40);
xnor U957 (N_957,In_1928,In_1633);
xor U958 (N_958,In_265,In_1277);
nor U959 (N_959,In_103,In_1761);
nor U960 (N_960,In_875,In_226);
and U961 (N_961,In_169,In_311);
nand U962 (N_962,In_871,In_819);
nor U963 (N_963,In_411,In_787);
nand U964 (N_964,In_1079,In_654);
nand U965 (N_965,In_1100,In_1999);
nor U966 (N_966,In_1637,In_1654);
and U967 (N_967,In_56,In_652);
xor U968 (N_968,In_161,In_537);
xnor U969 (N_969,In_751,In_624);
and U970 (N_970,In_1286,In_1710);
or U971 (N_971,In_491,In_1280);
or U972 (N_972,In_1328,In_958);
and U973 (N_973,In_771,In_1302);
or U974 (N_974,In_84,In_1966);
nor U975 (N_975,In_502,In_1133);
and U976 (N_976,In_1797,In_1845);
and U977 (N_977,In_1960,In_1073);
nor U978 (N_978,In_1815,In_175);
nor U979 (N_979,In_6,In_1547);
xor U980 (N_980,In_1256,In_1166);
nor U981 (N_981,In_1357,In_312);
nand U982 (N_982,In_1211,In_773);
xnor U983 (N_983,In_501,In_657);
and U984 (N_984,In_1151,In_680);
nor U985 (N_985,In_1350,In_852);
nand U986 (N_986,In_1397,In_970);
and U987 (N_987,In_798,In_160);
and U988 (N_988,In_1163,In_989);
nor U989 (N_989,In_1439,In_1556);
nand U990 (N_990,In_822,In_966);
nor U991 (N_991,In_1294,In_931);
and U992 (N_992,In_387,In_1149);
nand U993 (N_993,In_404,In_212);
nand U994 (N_994,In_1021,In_1415);
xnor U995 (N_995,In_1089,In_1447);
xor U996 (N_996,In_1545,In_1708);
xnor U997 (N_997,In_1433,In_1730);
xnor U998 (N_998,In_1391,In_1004);
or U999 (N_999,In_1318,In_976);
nand U1000 (N_1000,In_552,In_1128);
nor U1001 (N_1001,In_1494,In_1637);
and U1002 (N_1002,In_1739,In_1848);
or U1003 (N_1003,In_6,In_1957);
or U1004 (N_1004,In_640,In_954);
nor U1005 (N_1005,In_381,In_0);
nand U1006 (N_1006,In_1177,In_1532);
or U1007 (N_1007,In_507,In_962);
xor U1008 (N_1008,In_584,In_1314);
xnor U1009 (N_1009,In_436,In_797);
nor U1010 (N_1010,In_1516,In_602);
nand U1011 (N_1011,In_1882,In_21);
nand U1012 (N_1012,In_523,In_641);
nand U1013 (N_1013,In_1607,In_1166);
or U1014 (N_1014,In_923,In_536);
or U1015 (N_1015,In_1450,In_628);
or U1016 (N_1016,In_400,In_1904);
or U1017 (N_1017,In_1337,In_1071);
nand U1018 (N_1018,In_1326,In_1721);
and U1019 (N_1019,In_1868,In_1079);
nand U1020 (N_1020,In_69,In_1890);
or U1021 (N_1021,In_1889,In_414);
or U1022 (N_1022,In_1765,In_421);
xnor U1023 (N_1023,In_111,In_79);
or U1024 (N_1024,In_1496,In_1209);
and U1025 (N_1025,In_1136,In_503);
and U1026 (N_1026,In_430,In_1113);
and U1027 (N_1027,In_1941,In_1506);
nor U1028 (N_1028,In_270,In_1128);
or U1029 (N_1029,In_1559,In_422);
and U1030 (N_1030,In_1318,In_1678);
nand U1031 (N_1031,In_1004,In_1783);
or U1032 (N_1032,In_1369,In_664);
nor U1033 (N_1033,In_858,In_1614);
nor U1034 (N_1034,In_1262,In_1782);
xnor U1035 (N_1035,In_1568,In_1110);
xor U1036 (N_1036,In_1582,In_537);
and U1037 (N_1037,In_1780,In_764);
or U1038 (N_1038,In_498,In_923);
nor U1039 (N_1039,In_544,In_1702);
xor U1040 (N_1040,In_190,In_963);
nor U1041 (N_1041,In_1679,In_765);
xor U1042 (N_1042,In_1665,In_1837);
or U1043 (N_1043,In_637,In_697);
nand U1044 (N_1044,In_12,In_1531);
nor U1045 (N_1045,In_1833,In_1699);
nand U1046 (N_1046,In_1683,In_103);
nand U1047 (N_1047,In_907,In_1379);
or U1048 (N_1048,In_747,In_341);
or U1049 (N_1049,In_719,In_670);
or U1050 (N_1050,In_1320,In_65);
and U1051 (N_1051,In_17,In_1830);
and U1052 (N_1052,In_1282,In_191);
nand U1053 (N_1053,In_168,In_415);
and U1054 (N_1054,In_1511,In_1448);
nor U1055 (N_1055,In_1689,In_1667);
or U1056 (N_1056,In_1157,In_1381);
nor U1057 (N_1057,In_268,In_1624);
and U1058 (N_1058,In_1162,In_678);
nand U1059 (N_1059,In_931,In_1724);
or U1060 (N_1060,In_767,In_962);
nor U1061 (N_1061,In_1446,In_706);
xor U1062 (N_1062,In_1234,In_1652);
nor U1063 (N_1063,In_488,In_1782);
xor U1064 (N_1064,In_1469,In_655);
nor U1065 (N_1065,In_965,In_736);
nand U1066 (N_1066,In_534,In_1022);
and U1067 (N_1067,In_226,In_1797);
or U1068 (N_1068,In_29,In_1330);
xnor U1069 (N_1069,In_668,In_864);
xnor U1070 (N_1070,In_531,In_1625);
xor U1071 (N_1071,In_521,In_27);
nand U1072 (N_1072,In_1179,In_907);
or U1073 (N_1073,In_362,In_1276);
nor U1074 (N_1074,In_220,In_374);
nor U1075 (N_1075,In_1325,In_1975);
nand U1076 (N_1076,In_769,In_198);
nor U1077 (N_1077,In_1344,In_1210);
xor U1078 (N_1078,In_1932,In_1701);
xnor U1079 (N_1079,In_0,In_355);
or U1080 (N_1080,In_1196,In_1481);
xor U1081 (N_1081,In_872,In_1529);
or U1082 (N_1082,In_980,In_702);
xor U1083 (N_1083,In_170,In_745);
and U1084 (N_1084,In_306,In_1206);
nor U1085 (N_1085,In_1939,In_1975);
or U1086 (N_1086,In_1019,In_1590);
and U1087 (N_1087,In_342,In_1791);
nor U1088 (N_1088,In_365,In_849);
nand U1089 (N_1089,In_1973,In_392);
or U1090 (N_1090,In_1521,In_1952);
and U1091 (N_1091,In_1697,In_1449);
xnor U1092 (N_1092,In_1434,In_1240);
and U1093 (N_1093,In_839,In_1878);
nor U1094 (N_1094,In_672,In_227);
nor U1095 (N_1095,In_865,In_1247);
xnor U1096 (N_1096,In_423,In_1361);
and U1097 (N_1097,In_910,In_1614);
or U1098 (N_1098,In_172,In_792);
xnor U1099 (N_1099,In_1878,In_1248);
xnor U1100 (N_1100,In_512,In_670);
or U1101 (N_1101,In_1544,In_1769);
nand U1102 (N_1102,In_1282,In_1481);
and U1103 (N_1103,In_664,In_1412);
nor U1104 (N_1104,In_29,In_548);
nand U1105 (N_1105,In_1699,In_1641);
or U1106 (N_1106,In_1203,In_1432);
or U1107 (N_1107,In_1785,In_447);
nand U1108 (N_1108,In_61,In_730);
and U1109 (N_1109,In_760,In_1193);
or U1110 (N_1110,In_1404,In_1820);
xor U1111 (N_1111,In_1355,In_179);
nand U1112 (N_1112,In_950,In_796);
or U1113 (N_1113,In_983,In_892);
nand U1114 (N_1114,In_332,In_868);
or U1115 (N_1115,In_760,In_1020);
nand U1116 (N_1116,In_1462,In_729);
xor U1117 (N_1117,In_1883,In_557);
or U1118 (N_1118,In_263,In_1568);
and U1119 (N_1119,In_1457,In_734);
xor U1120 (N_1120,In_754,In_350);
and U1121 (N_1121,In_152,In_399);
and U1122 (N_1122,In_1076,In_1255);
nor U1123 (N_1123,In_473,In_973);
and U1124 (N_1124,In_358,In_764);
or U1125 (N_1125,In_828,In_494);
nand U1126 (N_1126,In_1685,In_1545);
xor U1127 (N_1127,In_472,In_1133);
or U1128 (N_1128,In_90,In_903);
or U1129 (N_1129,In_709,In_41);
nor U1130 (N_1130,In_1501,In_1125);
or U1131 (N_1131,In_887,In_1371);
xor U1132 (N_1132,In_1421,In_691);
or U1133 (N_1133,In_164,In_1297);
and U1134 (N_1134,In_1630,In_1362);
xor U1135 (N_1135,In_640,In_946);
and U1136 (N_1136,In_1882,In_694);
or U1137 (N_1137,In_1811,In_815);
nor U1138 (N_1138,In_1434,In_926);
nor U1139 (N_1139,In_116,In_150);
or U1140 (N_1140,In_1785,In_1061);
nor U1141 (N_1141,In_1327,In_731);
xnor U1142 (N_1142,In_1510,In_594);
nand U1143 (N_1143,In_1850,In_1445);
nand U1144 (N_1144,In_1094,In_1061);
or U1145 (N_1145,In_1456,In_934);
nand U1146 (N_1146,In_398,In_1878);
nand U1147 (N_1147,In_1523,In_1771);
nand U1148 (N_1148,In_1327,In_907);
or U1149 (N_1149,In_1239,In_263);
nand U1150 (N_1150,In_1433,In_117);
and U1151 (N_1151,In_232,In_1480);
nand U1152 (N_1152,In_530,In_1425);
nor U1153 (N_1153,In_1402,In_1662);
nand U1154 (N_1154,In_1949,In_1151);
nor U1155 (N_1155,In_1246,In_73);
xnor U1156 (N_1156,In_757,In_465);
and U1157 (N_1157,In_1788,In_467);
xnor U1158 (N_1158,In_1661,In_1956);
nand U1159 (N_1159,In_258,In_1497);
nor U1160 (N_1160,In_1533,In_581);
nor U1161 (N_1161,In_1641,In_396);
xor U1162 (N_1162,In_725,In_407);
nor U1163 (N_1163,In_1166,In_1424);
nor U1164 (N_1164,In_1881,In_855);
and U1165 (N_1165,In_1980,In_1320);
nand U1166 (N_1166,In_113,In_491);
or U1167 (N_1167,In_871,In_990);
nor U1168 (N_1168,In_175,In_215);
or U1169 (N_1169,In_1564,In_1286);
xor U1170 (N_1170,In_436,In_865);
nor U1171 (N_1171,In_829,In_1085);
nand U1172 (N_1172,In_693,In_1292);
and U1173 (N_1173,In_1802,In_74);
xor U1174 (N_1174,In_1093,In_1421);
nor U1175 (N_1175,In_1719,In_1154);
and U1176 (N_1176,In_1566,In_970);
nor U1177 (N_1177,In_629,In_1979);
nand U1178 (N_1178,In_1628,In_206);
nand U1179 (N_1179,In_1853,In_412);
nor U1180 (N_1180,In_866,In_238);
nor U1181 (N_1181,In_123,In_1657);
and U1182 (N_1182,In_682,In_212);
nor U1183 (N_1183,In_374,In_812);
and U1184 (N_1184,In_513,In_1032);
nor U1185 (N_1185,In_53,In_373);
or U1186 (N_1186,In_635,In_367);
nand U1187 (N_1187,In_1430,In_1346);
nor U1188 (N_1188,In_1593,In_1148);
xnor U1189 (N_1189,In_1384,In_1179);
nor U1190 (N_1190,In_1529,In_198);
nand U1191 (N_1191,In_1962,In_408);
nor U1192 (N_1192,In_186,In_565);
xnor U1193 (N_1193,In_1800,In_1469);
nor U1194 (N_1194,In_1982,In_1437);
xor U1195 (N_1195,In_1058,In_443);
or U1196 (N_1196,In_991,In_1613);
and U1197 (N_1197,In_437,In_1422);
xnor U1198 (N_1198,In_477,In_502);
nor U1199 (N_1199,In_1118,In_1029);
nor U1200 (N_1200,In_95,In_928);
nand U1201 (N_1201,In_468,In_1013);
and U1202 (N_1202,In_1603,In_1471);
xor U1203 (N_1203,In_1279,In_1579);
or U1204 (N_1204,In_1738,In_1364);
and U1205 (N_1205,In_1034,In_1893);
nand U1206 (N_1206,In_531,In_533);
or U1207 (N_1207,In_1620,In_1467);
or U1208 (N_1208,In_30,In_1457);
or U1209 (N_1209,In_1504,In_1194);
and U1210 (N_1210,In_942,In_1438);
xor U1211 (N_1211,In_1397,In_378);
xnor U1212 (N_1212,In_1914,In_436);
nand U1213 (N_1213,In_1446,In_1136);
or U1214 (N_1214,In_1917,In_1133);
or U1215 (N_1215,In_700,In_1826);
xor U1216 (N_1216,In_191,In_1478);
nor U1217 (N_1217,In_746,In_811);
or U1218 (N_1218,In_367,In_1627);
xor U1219 (N_1219,In_1289,In_1775);
and U1220 (N_1220,In_1115,In_1162);
xor U1221 (N_1221,In_971,In_881);
nand U1222 (N_1222,In_1487,In_460);
and U1223 (N_1223,In_1602,In_581);
xnor U1224 (N_1224,In_1352,In_317);
or U1225 (N_1225,In_680,In_906);
nor U1226 (N_1226,In_513,In_279);
nor U1227 (N_1227,In_1315,In_1284);
xnor U1228 (N_1228,In_1121,In_1028);
or U1229 (N_1229,In_93,In_1105);
and U1230 (N_1230,In_544,In_1492);
nor U1231 (N_1231,In_1413,In_1820);
or U1232 (N_1232,In_340,In_497);
xnor U1233 (N_1233,In_248,In_1312);
or U1234 (N_1234,In_10,In_113);
and U1235 (N_1235,In_778,In_317);
nand U1236 (N_1236,In_221,In_1606);
or U1237 (N_1237,In_1811,In_1257);
and U1238 (N_1238,In_150,In_1042);
nand U1239 (N_1239,In_514,In_133);
nand U1240 (N_1240,In_1680,In_913);
nand U1241 (N_1241,In_539,In_1129);
xnor U1242 (N_1242,In_853,In_880);
nand U1243 (N_1243,In_1288,In_1933);
and U1244 (N_1244,In_1418,In_1125);
nand U1245 (N_1245,In_1674,In_672);
nand U1246 (N_1246,In_598,In_780);
nor U1247 (N_1247,In_238,In_1035);
or U1248 (N_1248,In_106,In_192);
or U1249 (N_1249,In_1101,In_1121);
or U1250 (N_1250,In_210,In_1457);
and U1251 (N_1251,In_876,In_1587);
and U1252 (N_1252,In_567,In_1555);
and U1253 (N_1253,In_1543,In_932);
or U1254 (N_1254,In_964,In_1915);
or U1255 (N_1255,In_1408,In_1052);
or U1256 (N_1256,In_494,In_764);
xor U1257 (N_1257,In_915,In_261);
and U1258 (N_1258,In_1124,In_315);
nor U1259 (N_1259,In_1155,In_1214);
xor U1260 (N_1260,In_100,In_1693);
or U1261 (N_1261,In_522,In_825);
or U1262 (N_1262,In_87,In_1720);
and U1263 (N_1263,In_305,In_866);
nand U1264 (N_1264,In_1474,In_1887);
and U1265 (N_1265,In_18,In_391);
nand U1266 (N_1266,In_1127,In_1835);
or U1267 (N_1267,In_691,In_1960);
xor U1268 (N_1268,In_1148,In_377);
and U1269 (N_1269,In_315,In_391);
nand U1270 (N_1270,In_1010,In_1131);
and U1271 (N_1271,In_1059,In_149);
and U1272 (N_1272,In_826,In_626);
nand U1273 (N_1273,In_782,In_1073);
or U1274 (N_1274,In_374,In_1632);
nor U1275 (N_1275,In_1464,In_274);
nor U1276 (N_1276,In_1513,In_1061);
or U1277 (N_1277,In_1347,In_123);
xor U1278 (N_1278,In_1974,In_61);
xnor U1279 (N_1279,In_1965,In_1872);
xnor U1280 (N_1280,In_98,In_1936);
nand U1281 (N_1281,In_473,In_606);
xor U1282 (N_1282,In_1617,In_1277);
xor U1283 (N_1283,In_729,In_1049);
or U1284 (N_1284,In_970,In_1166);
nand U1285 (N_1285,In_626,In_718);
nor U1286 (N_1286,In_606,In_1623);
nor U1287 (N_1287,In_289,In_1730);
nand U1288 (N_1288,In_1578,In_269);
xor U1289 (N_1289,In_104,In_177);
and U1290 (N_1290,In_611,In_399);
and U1291 (N_1291,In_349,In_561);
nor U1292 (N_1292,In_45,In_1466);
nand U1293 (N_1293,In_1133,In_496);
xor U1294 (N_1294,In_698,In_1178);
nand U1295 (N_1295,In_1405,In_463);
or U1296 (N_1296,In_332,In_1692);
nor U1297 (N_1297,In_1718,In_1651);
xor U1298 (N_1298,In_820,In_998);
nor U1299 (N_1299,In_751,In_99);
and U1300 (N_1300,In_815,In_813);
or U1301 (N_1301,In_444,In_1693);
xnor U1302 (N_1302,In_1120,In_1640);
nand U1303 (N_1303,In_1274,In_162);
and U1304 (N_1304,In_1874,In_1774);
or U1305 (N_1305,In_1302,In_1023);
nand U1306 (N_1306,In_783,In_1638);
nand U1307 (N_1307,In_144,In_1182);
xnor U1308 (N_1308,In_1400,In_1576);
nor U1309 (N_1309,In_1380,In_1410);
nand U1310 (N_1310,In_796,In_1366);
nand U1311 (N_1311,In_1135,In_1914);
and U1312 (N_1312,In_1386,In_1502);
nor U1313 (N_1313,In_1065,In_1410);
nand U1314 (N_1314,In_1734,In_1864);
nor U1315 (N_1315,In_971,In_543);
nor U1316 (N_1316,In_597,In_1303);
xnor U1317 (N_1317,In_1194,In_587);
nor U1318 (N_1318,In_232,In_1758);
or U1319 (N_1319,In_351,In_1916);
and U1320 (N_1320,In_253,In_1347);
xor U1321 (N_1321,In_1585,In_1235);
or U1322 (N_1322,In_472,In_1655);
xnor U1323 (N_1323,In_851,In_1930);
nand U1324 (N_1324,In_830,In_1676);
and U1325 (N_1325,In_1747,In_224);
or U1326 (N_1326,In_473,In_882);
or U1327 (N_1327,In_447,In_1638);
nand U1328 (N_1328,In_776,In_1207);
nor U1329 (N_1329,In_973,In_1477);
nand U1330 (N_1330,In_429,In_499);
or U1331 (N_1331,In_678,In_112);
and U1332 (N_1332,In_1388,In_622);
nor U1333 (N_1333,In_1581,In_928);
nor U1334 (N_1334,In_1476,In_705);
or U1335 (N_1335,In_244,In_1312);
nor U1336 (N_1336,In_1590,In_1346);
or U1337 (N_1337,In_1363,In_57);
nor U1338 (N_1338,In_1371,In_44);
nand U1339 (N_1339,In_1977,In_760);
and U1340 (N_1340,In_344,In_1409);
nor U1341 (N_1341,In_1708,In_777);
xnor U1342 (N_1342,In_1756,In_1119);
nand U1343 (N_1343,In_1106,In_145);
and U1344 (N_1344,In_1968,In_840);
nand U1345 (N_1345,In_1922,In_482);
or U1346 (N_1346,In_557,In_1008);
nor U1347 (N_1347,In_925,In_804);
or U1348 (N_1348,In_1053,In_395);
nand U1349 (N_1349,In_1462,In_699);
or U1350 (N_1350,In_168,In_44);
and U1351 (N_1351,In_270,In_715);
nand U1352 (N_1352,In_1787,In_884);
nor U1353 (N_1353,In_963,In_1104);
nand U1354 (N_1354,In_1417,In_426);
nor U1355 (N_1355,In_995,In_1976);
nand U1356 (N_1356,In_1207,In_498);
or U1357 (N_1357,In_322,In_1955);
nand U1358 (N_1358,In_1385,In_238);
and U1359 (N_1359,In_1492,In_423);
and U1360 (N_1360,In_533,In_1193);
and U1361 (N_1361,In_683,In_1505);
nand U1362 (N_1362,In_1215,In_1304);
xor U1363 (N_1363,In_249,In_1551);
nand U1364 (N_1364,In_1185,In_1564);
nor U1365 (N_1365,In_1545,In_1019);
and U1366 (N_1366,In_1846,In_1594);
nand U1367 (N_1367,In_1000,In_1012);
nor U1368 (N_1368,In_182,In_70);
and U1369 (N_1369,In_355,In_1161);
and U1370 (N_1370,In_1825,In_1110);
and U1371 (N_1371,In_1093,In_1558);
and U1372 (N_1372,In_424,In_750);
xor U1373 (N_1373,In_1694,In_579);
nand U1374 (N_1374,In_349,In_799);
nor U1375 (N_1375,In_504,In_747);
nor U1376 (N_1376,In_364,In_1307);
xnor U1377 (N_1377,In_512,In_828);
xnor U1378 (N_1378,In_137,In_558);
xnor U1379 (N_1379,In_179,In_65);
or U1380 (N_1380,In_1549,In_1590);
and U1381 (N_1381,In_427,In_1133);
and U1382 (N_1382,In_703,In_1754);
nand U1383 (N_1383,In_1201,In_814);
nand U1384 (N_1384,In_435,In_1001);
nand U1385 (N_1385,In_417,In_688);
xnor U1386 (N_1386,In_1326,In_1692);
and U1387 (N_1387,In_1755,In_1665);
nor U1388 (N_1388,In_323,In_614);
nor U1389 (N_1389,In_1547,In_1005);
xnor U1390 (N_1390,In_361,In_255);
or U1391 (N_1391,In_922,In_1097);
and U1392 (N_1392,In_112,In_1249);
nor U1393 (N_1393,In_199,In_571);
nand U1394 (N_1394,In_1559,In_1731);
and U1395 (N_1395,In_1903,In_573);
xor U1396 (N_1396,In_199,In_906);
nand U1397 (N_1397,In_1803,In_1977);
xor U1398 (N_1398,In_5,In_1226);
xnor U1399 (N_1399,In_737,In_1313);
nand U1400 (N_1400,In_1468,In_1953);
xor U1401 (N_1401,In_319,In_212);
nor U1402 (N_1402,In_1210,In_1594);
xnor U1403 (N_1403,In_1545,In_1580);
and U1404 (N_1404,In_1541,In_231);
nor U1405 (N_1405,In_1263,In_1008);
nand U1406 (N_1406,In_926,In_550);
nand U1407 (N_1407,In_1013,In_1129);
nand U1408 (N_1408,In_1886,In_1890);
and U1409 (N_1409,In_1614,In_1633);
and U1410 (N_1410,In_1933,In_1611);
nand U1411 (N_1411,In_351,In_1381);
nor U1412 (N_1412,In_1158,In_525);
xnor U1413 (N_1413,In_38,In_1052);
or U1414 (N_1414,In_450,In_242);
nand U1415 (N_1415,In_866,In_198);
or U1416 (N_1416,In_1896,In_1959);
nand U1417 (N_1417,In_1901,In_989);
nand U1418 (N_1418,In_521,In_1767);
nor U1419 (N_1419,In_1925,In_1513);
or U1420 (N_1420,In_1120,In_985);
nor U1421 (N_1421,In_569,In_270);
nand U1422 (N_1422,In_1437,In_1505);
nor U1423 (N_1423,In_257,In_1958);
nand U1424 (N_1424,In_1397,In_1271);
xor U1425 (N_1425,In_1328,In_1928);
xor U1426 (N_1426,In_1124,In_1804);
or U1427 (N_1427,In_1172,In_1623);
or U1428 (N_1428,In_756,In_1550);
and U1429 (N_1429,In_1895,In_701);
xor U1430 (N_1430,In_1804,In_1850);
and U1431 (N_1431,In_538,In_177);
nor U1432 (N_1432,In_953,In_1659);
xor U1433 (N_1433,In_1794,In_227);
and U1434 (N_1434,In_1296,In_1258);
nor U1435 (N_1435,In_1572,In_521);
or U1436 (N_1436,In_733,In_1152);
and U1437 (N_1437,In_1055,In_1046);
xor U1438 (N_1438,In_1579,In_1821);
nor U1439 (N_1439,In_1379,In_1771);
nor U1440 (N_1440,In_900,In_484);
nand U1441 (N_1441,In_427,In_769);
or U1442 (N_1442,In_157,In_148);
xor U1443 (N_1443,In_1910,In_405);
or U1444 (N_1444,In_291,In_721);
nor U1445 (N_1445,In_1346,In_94);
nand U1446 (N_1446,In_676,In_640);
nand U1447 (N_1447,In_770,In_1356);
xor U1448 (N_1448,In_1661,In_600);
or U1449 (N_1449,In_71,In_536);
nand U1450 (N_1450,In_813,In_471);
nand U1451 (N_1451,In_1309,In_1917);
nand U1452 (N_1452,In_1179,In_1615);
or U1453 (N_1453,In_390,In_836);
nor U1454 (N_1454,In_1106,In_1247);
nor U1455 (N_1455,In_998,In_1558);
nand U1456 (N_1456,In_473,In_407);
nand U1457 (N_1457,In_1218,In_177);
nand U1458 (N_1458,In_915,In_1764);
nand U1459 (N_1459,In_1135,In_1206);
xnor U1460 (N_1460,In_1942,In_77);
nand U1461 (N_1461,In_885,In_71);
and U1462 (N_1462,In_168,In_24);
nand U1463 (N_1463,In_825,In_542);
and U1464 (N_1464,In_294,In_1638);
or U1465 (N_1465,In_1117,In_940);
xor U1466 (N_1466,In_935,In_353);
nand U1467 (N_1467,In_941,In_1245);
and U1468 (N_1468,In_1122,In_711);
or U1469 (N_1469,In_1750,In_1353);
xnor U1470 (N_1470,In_1426,In_1240);
or U1471 (N_1471,In_1680,In_134);
or U1472 (N_1472,In_1952,In_860);
xor U1473 (N_1473,In_893,In_1304);
nand U1474 (N_1474,In_1104,In_1176);
or U1475 (N_1475,In_593,In_1190);
xnor U1476 (N_1476,In_372,In_1367);
nand U1477 (N_1477,In_1557,In_1469);
nor U1478 (N_1478,In_1337,In_1784);
xnor U1479 (N_1479,In_661,In_667);
xor U1480 (N_1480,In_1491,In_200);
and U1481 (N_1481,In_899,In_1223);
and U1482 (N_1482,In_924,In_1394);
and U1483 (N_1483,In_243,In_413);
xnor U1484 (N_1484,In_43,In_1115);
or U1485 (N_1485,In_691,In_11);
nand U1486 (N_1486,In_1887,In_1053);
xnor U1487 (N_1487,In_349,In_737);
or U1488 (N_1488,In_644,In_1708);
xnor U1489 (N_1489,In_471,In_639);
or U1490 (N_1490,In_750,In_1755);
nor U1491 (N_1491,In_87,In_1184);
or U1492 (N_1492,In_1376,In_123);
xor U1493 (N_1493,In_266,In_593);
nor U1494 (N_1494,In_633,In_1189);
or U1495 (N_1495,In_190,In_1458);
or U1496 (N_1496,In_1860,In_1711);
nand U1497 (N_1497,In_989,In_1155);
and U1498 (N_1498,In_922,In_639);
or U1499 (N_1499,In_461,In_164);
nor U1500 (N_1500,In_829,In_1078);
and U1501 (N_1501,In_1637,In_812);
xor U1502 (N_1502,In_899,In_1976);
xnor U1503 (N_1503,In_747,In_870);
or U1504 (N_1504,In_1472,In_384);
and U1505 (N_1505,In_1839,In_776);
and U1506 (N_1506,In_157,In_1664);
nand U1507 (N_1507,In_224,In_1766);
nand U1508 (N_1508,In_938,In_1632);
xor U1509 (N_1509,In_909,In_889);
and U1510 (N_1510,In_663,In_289);
or U1511 (N_1511,In_289,In_1852);
or U1512 (N_1512,In_1126,In_767);
and U1513 (N_1513,In_1679,In_94);
and U1514 (N_1514,In_15,In_1189);
xor U1515 (N_1515,In_1380,In_208);
xor U1516 (N_1516,In_1263,In_1741);
and U1517 (N_1517,In_1939,In_1218);
nor U1518 (N_1518,In_25,In_108);
nor U1519 (N_1519,In_922,In_1231);
or U1520 (N_1520,In_1587,In_742);
or U1521 (N_1521,In_1023,In_280);
or U1522 (N_1522,In_387,In_265);
nor U1523 (N_1523,In_609,In_840);
nor U1524 (N_1524,In_1406,In_247);
nor U1525 (N_1525,In_1163,In_1265);
or U1526 (N_1526,In_1803,In_7);
and U1527 (N_1527,In_1575,In_1187);
xnor U1528 (N_1528,In_1438,In_1582);
xor U1529 (N_1529,In_1022,In_1521);
and U1530 (N_1530,In_399,In_257);
or U1531 (N_1531,In_1739,In_1510);
nor U1532 (N_1532,In_80,In_756);
or U1533 (N_1533,In_221,In_825);
xor U1534 (N_1534,In_1243,In_1760);
and U1535 (N_1535,In_848,In_1921);
nand U1536 (N_1536,In_750,In_1793);
xor U1537 (N_1537,In_759,In_690);
nand U1538 (N_1538,In_919,In_1797);
xor U1539 (N_1539,In_1167,In_1640);
or U1540 (N_1540,In_1575,In_180);
or U1541 (N_1541,In_1624,In_712);
or U1542 (N_1542,In_1697,In_500);
nor U1543 (N_1543,In_273,In_1978);
xnor U1544 (N_1544,In_269,In_775);
and U1545 (N_1545,In_576,In_213);
xor U1546 (N_1546,In_987,In_869);
xor U1547 (N_1547,In_1585,In_376);
nor U1548 (N_1548,In_152,In_110);
xor U1549 (N_1549,In_1020,In_1886);
or U1550 (N_1550,In_1691,In_1685);
and U1551 (N_1551,In_1499,In_1435);
xnor U1552 (N_1552,In_424,In_1814);
and U1553 (N_1553,In_593,In_591);
nand U1554 (N_1554,In_282,In_1037);
nor U1555 (N_1555,In_1138,In_1820);
or U1556 (N_1556,In_1843,In_1658);
or U1557 (N_1557,In_1041,In_204);
and U1558 (N_1558,In_827,In_172);
and U1559 (N_1559,In_925,In_1097);
or U1560 (N_1560,In_100,In_1345);
or U1561 (N_1561,In_1689,In_416);
and U1562 (N_1562,In_1110,In_469);
and U1563 (N_1563,In_1901,In_210);
nor U1564 (N_1564,In_705,In_17);
and U1565 (N_1565,In_787,In_502);
or U1566 (N_1566,In_204,In_236);
nor U1567 (N_1567,In_403,In_1143);
or U1568 (N_1568,In_260,In_907);
nor U1569 (N_1569,In_1588,In_1700);
nor U1570 (N_1570,In_1938,In_967);
nand U1571 (N_1571,In_1787,In_1286);
and U1572 (N_1572,In_762,In_1707);
and U1573 (N_1573,In_1668,In_845);
or U1574 (N_1574,In_1083,In_375);
nor U1575 (N_1575,In_505,In_1715);
xor U1576 (N_1576,In_888,In_1474);
nand U1577 (N_1577,In_1741,In_1039);
nor U1578 (N_1578,In_1094,In_1867);
nor U1579 (N_1579,In_489,In_231);
nand U1580 (N_1580,In_1343,In_1544);
or U1581 (N_1581,In_840,In_520);
nand U1582 (N_1582,In_622,In_589);
nor U1583 (N_1583,In_1473,In_264);
and U1584 (N_1584,In_1594,In_45);
nand U1585 (N_1585,In_410,In_797);
nand U1586 (N_1586,In_810,In_374);
and U1587 (N_1587,In_1780,In_1519);
nor U1588 (N_1588,In_1053,In_798);
nand U1589 (N_1589,In_185,In_1561);
xnor U1590 (N_1590,In_508,In_991);
nand U1591 (N_1591,In_335,In_1210);
nor U1592 (N_1592,In_1212,In_1211);
nand U1593 (N_1593,In_597,In_655);
nor U1594 (N_1594,In_1282,In_576);
or U1595 (N_1595,In_908,In_1924);
or U1596 (N_1596,In_1653,In_144);
and U1597 (N_1597,In_557,In_978);
or U1598 (N_1598,In_1534,In_275);
nand U1599 (N_1599,In_1256,In_819);
nand U1600 (N_1600,In_660,In_850);
nor U1601 (N_1601,In_1418,In_774);
nor U1602 (N_1602,In_163,In_1480);
and U1603 (N_1603,In_808,In_134);
and U1604 (N_1604,In_1195,In_69);
xor U1605 (N_1605,In_225,In_1457);
xor U1606 (N_1606,In_373,In_1765);
or U1607 (N_1607,In_293,In_676);
nand U1608 (N_1608,In_84,In_1027);
nor U1609 (N_1609,In_1524,In_1356);
nor U1610 (N_1610,In_409,In_1216);
nor U1611 (N_1611,In_1207,In_1147);
and U1612 (N_1612,In_1129,In_1574);
nor U1613 (N_1613,In_137,In_1305);
or U1614 (N_1614,In_358,In_1931);
nor U1615 (N_1615,In_1150,In_367);
nand U1616 (N_1616,In_1623,In_34);
or U1617 (N_1617,In_1556,In_73);
nand U1618 (N_1618,In_747,In_561);
or U1619 (N_1619,In_1781,In_874);
and U1620 (N_1620,In_320,In_1374);
xnor U1621 (N_1621,In_1772,In_1798);
and U1622 (N_1622,In_941,In_1369);
xnor U1623 (N_1623,In_1355,In_1790);
and U1624 (N_1624,In_234,In_1128);
nand U1625 (N_1625,In_1954,In_125);
nand U1626 (N_1626,In_1138,In_882);
and U1627 (N_1627,In_707,In_1069);
nor U1628 (N_1628,In_38,In_169);
xor U1629 (N_1629,In_1594,In_76);
xnor U1630 (N_1630,In_1456,In_1946);
or U1631 (N_1631,In_871,In_445);
or U1632 (N_1632,In_1291,In_1213);
nor U1633 (N_1633,In_102,In_1840);
nand U1634 (N_1634,In_86,In_449);
xor U1635 (N_1635,In_592,In_917);
xor U1636 (N_1636,In_388,In_723);
and U1637 (N_1637,In_870,In_724);
and U1638 (N_1638,In_1158,In_577);
or U1639 (N_1639,In_1606,In_1917);
or U1640 (N_1640,In_410,In_1353);
nand U1641 (N_1641,In_1934,In_1145);
nor U1642 (N_1642,In_1263,In_606);
xor U1643 (N_1643,In_1103,In_1333);
nand U1644 (N_1644,In_1991,In_389);
or U1645 (N_1645,In_1584,In_1681);
nand U1646 (N_1646,In_1458,In_920);
nor U1647 (N_1647,In_1890,In_259);
xnor U1648 (N_1648,In_484,In_1623);
nor U1649 (N_1649,In_190,In_1740);
and U1650 (N_1650,In_31,In_1348);
nor U1651 (N_1651,In_1606,In_1701);
nor U1652 (N_1652,In_193,In_970);
or U1653 (N_1653,In_1080,In_1642);
nor U1654 (N_1654,In_867,In_1776);
nand U1655 (N_1655,In_245,In_319);
xnor U1656 (N_1656,In_1556,In_1977);
nand U1657 (N_1657,In_1223,In_970);
nand U1658 (N_1658,In_1373,In_995);
and U1659 (N_1659,In_1032,In_1201);
xor U1660 (N_1660,In_676,In_1103);
nor U1661 (N_1661,In_1567,In_394);
or U1662 (N_1662,In_310,In_32);
xnor U1663 (N_1663,In_427,In_1544);
and U1664 (N_1664,In_437,In_1137);
and U1665 (N_1665,In_1445,In_165);
nand U1666 (N_1666,In_1841,In_1233);
nand U1667 (N_1667,In_1207,In_1349);
nor U1668 (N_1668,In_261,In_1150);
and U1669 (N_1669,In_68,In_1076);
or U1670 (N_1670,In_411,In_1569);
nor U1671 (N_1671,In_989,In_1002);
and U1672 (N_1672,In_377,In_1308);
nor U1673 (N_1673,In_188,In_989);
or U1674 (N_1674,In_947,In_332);
xor U1675 (N_1675,In_1930,In_1215);
xor U1676 (N_1676,In_339,In_238);
xor U1677 (N_1677,In_558,In_1364);
nand U1678 (N_1678,In_768,In_648);
xnor U1679 (N_1679,In_1801,In_1302);
nand U1680 (N_1680,In_231,In_764);
or U1681 (N_1681,In_341,In_1683);
and U1682 (N_1682,In_1028,In_1344);
or U1683 (N_1683,In_681,In_1588);
or U1684 (N_1684,In_178,In_720);
and U1685 (N_1685,In_754,In_1941);
or U1686 (N_1686,In_1578,In_287);
or U1687 (N_1687,In_1268,In_1475);
nor U1688 (N_1688,In_722,In_1106);
xnor U1689 (N_1689,In_787,In_477);
and U1690 (N_1690,In_361,In_1328);
nor U1691 (N_1691,In_1214,In_57);
and U1692 (N_1692,In_1480,In_929);
nor U1693 (N_1693,In_1823,In_1110);
nor U1694 (N_1694,In_233,In_145);
nor U1695 (N_1695,In_392,In_987);
xor U1696 (N_1696,In_1536,In_758);
and U1697 (N_1697,In_1384,In_751);
nor U1698 (N_1698,In_392,In_1149);
nor U1699 (N_1699,In_1618,In_1508);
nand U1700 (N_1700,In_860,In_414);
nor U1701 (N_1701,In_965,In_279);
nor U1702 (N_1702,In_1202,In_195);
or U1703 (N_1703,In_179,In_1086);
nand U1704 (N_1704,In_155,In_1747);
nand U1705 (N_1705,In_851,In_547);
and U1706 (N_1706,In_33,In_1113);
and U1707 (N_1707,In_435,In_671);
xor U1708 (N_1708,In_1332,In_546);
xor U1709 (N_1709,In_589,In_1876);
xor U1710 (N_1710,In_1345,In_1775);
nand U1711 (N_1711,In_921,In_76);
or U1712 (N_1712,In_1155,In_257);
xnor U1713 (N_1713,In_1272,In_1390);
and U1714 (N_1714,In_1664,In_316);
nand U1715 (N_1715,In_1108,In_601);
and U1716 (N_1716,In_1806,In_516);
nor U1717 (N_1717,In_1601,In_1248);
nand U1718 (N_1718,In_92,In_733);
or U1719 (N_1719,In_1914,In_1465);
xnor U1720 (N_1720,In_1646,In_595);
nand U1721 (N_1721,In_912,In_1327);
xnor U1722 (N_1722,In_356,In_1586);
nand U1723 (N_1723,In_1906,In_1303);
nand U1724 (N_1724,In_1855,In_110);
nand U1725 (N_1725,In_1469,In_1423);
nor U1726 (N_1726,In_1888,In_753);
xnor U1727 (N_1727,In_252,In_26);
or U1728 (N_1728,In_415,In_1834);
nand U1729 (N_1729,In_1978,In_773);
or U1730 (N_1730,In_1931,In_1667);
or U1731 (N_1731,In_1052,In_1692);
nor U1732 (N_1732,In_1698,In_1343);
xnor U1733 (N_1733,In_580,In_298);
and U1734 (N_1734,In_1281,In_11);
and U1735 (N_1735,In_1316,In_1344);
or U1736 (N_1736,In_752,In_393);
nor U1737 (N_1737,In_416,In_629);
or U1738 (N_1738,In_1878,In_507);
or U1739 (N_1739,In_539,In_1314);
nand U1740 (N_1740,In_315,In_1521);
xor U1741 (N_1741,In_1199,In_1689);
or U1742 (N_1742,In_1150,In_1187);
nand U1743 (N_1743,In_1390,In_179);
and U1744 (N_1744,In_1341,In_192);
or U1745 (N_1745,In_1318,In_752);
nor U1746 (N_1746,In_1683,In_721);
nor U1747 (N_1747,In_41,In_1425);
nor U1748 (N_1748,In_1689,In_1048);
or U1749 (N_1749,In_796,In_1411);
xor U1750 (N_1750,In_1833,In_1082);
or U1751 (N_1751,In_1421,In_1525);
nand U1752 (N_1752,In_917,In_1380);
nor U1753 (N_1753,In_1671,In_1729);
nand U1754 (N_1754,In_1360,In_714);
and U1755 (N_1755,In_1003,In_1701);
or U1756 (N_1756,In_446,In_1667);
xor U1757 (N_1757,In_1345,In_1346);
nor U1758 (N_1758,In_484,In_28);
or U1759 (N_1759,In_1469,In_1426);
xor U1760 (N_1760,In_1875,In_917);
xnor U1761 (N_1761,In_989,In_73);
nand U1762 (N_1762,In_11,In_1662);
and U1763 (N_1763,In_757,In_572);
and U1764 (N_1764,In_1183,In_1649);
nor U1765 (N_1765,In_1778,In_1621);
nor U1766 (N_1766,In_986,In_452);
nand U1767 (N_1767,In_635,In_303);
nand U1768 (N_1768,In_1015,In_259);
nor U1769 (N_1769,In_224,In_1009);
or U1770 (N_1770,In_1178,In_1211);
xor U1771 (N_1771,In_781,In_234);
nor U1772 (N_1772,In_149,In_889);
or U1773 (N_1773,In_1584,In_189);
xor U1774 (N_1774,In_993,In_213);
nand U1775 (N_1775,In_108,In_1540);
or U1776 (N_1776,In_1594,In_534);
and U1777 (N_1777,In_596,In_1266);
xor U1778 (N_1778,In_1204,In_1247);
nor U1779 (N_1779,In_1700,In_387);
nand U1780 (N_1780,In_134,In_47);
and U1781 (N_1781,In_1560,In_1818);
nand U1782 (N_1782,In_853,In_1228);
or U1783 (N_1783,In_1092,In_1808);
and U1784 (N_1784,In_1807,In_626);
or U1785 (N_1785,In_1584,In_273);
or U1786 (N_1786,In_1172,In_2);
and U1787 (N_1787,In_1351,In_1011);
nand U1788 (N_1788,In_1906,In_1214);
xor U1789 (N_1789,In_1957,In_1398);
nor U1790 (N_1790,In_412,In_295);
or U1791 (N_1791,In_1368,In_504);
or U1792 (N_1792,In_39,In_1069);
xor U1793 (N_1793,In_1353,In_332);
nor U1794 (N_1794,In_308,In_1591);
nor U1795 (N_1795,In_811,In_228);
nand U1796 (N_1796,In_165,In_513);
or U1797 (N_1797,In_1844,In_266);
nor U1798 (N_1798,In_124,In_237);
and U1799 (N_1799,In_1354,In_713);
and U1800 (N_1800,In_1831,In_1793);
nor U1801 (N_1801,In_1699,In_1200);
xnor U1802 (N_1802,In_1803,In_266);
xor U1803 (N_1803,In_1079,In_1145);
nand U1804 (N_1804,In_49,In_1042);
nand U1805 (N_1805,In_1535,In_106);
nor U1806 (N_1806,In_347,In_1997);
nor U1807 (N_1807,In_352,In_850);
and U1808 (N_1808,In_1952,In_908);
xnor U1809 (N_1809,In_1259,In_1484);
and U1810 (N_1810,In_364,In_1449);
and U1811 (N_1811,In_26,In_49);
nand U1812 (N_1812,In_1651,In_893);
and U1813 (N_1813,In_138,In_1031);
nand U1814 (N_1814,In_1177,In_973);
or U1815 (N_1815,In_1383,In_1952);
xor U1816 (N_1816,In_1732,In_661);
and U1817 (N_1817,In_1651,In_1352);
nor U1818 (N_1818,In_760,In_1825);
nor U1819 (N_1819,In_97,In_1247);
nand U1820 (N_1820,In_404,In_218);
nand U1821 (N_1821,In_1461,In_819);
or U1822 (N_1822,In_1446,In_1908);
and U1823 (N_1823,In_1388,In_1474);
xor U1824 (N_1824,In_1957,In_1605);
nand U1825 (N_1825,In_275,In_1585);
xnor U1826 (N_1826,In_1517,In_796);
and U1827 (N_1827,In_1526,In_1773);
and U1828 (N_1828,In_974,In_267);
nor U1829 (N_1829,In_1048,In_129);
xor U1830 (N_1830,In_143,In_1123);
nand U1831 (N_1831,In_498,In_981);
nor U1832 (N_1832,In_904,In_244);
nand U1833 (N_1833,In_274,In_1660);
nor U1834 (N_1834,In_989,In_1050);
or U1835 (N_1835,In_1553,In_110);
nand U1836 (N_1836,In_1093,In_1577);
nor U1837 (N_1837,In_1043,In_1265);
xor U1838 (N_1838,In_1343,In_1335);
nor U1839 (N_1839,In_1017,In_692);
and U1840 (N_1840,In_1391,In_1083);
and U1841 (N_1841,In_220,In_1444);
nand U1842 (N_1842,In_356,In_899);
nand U1843 (N_1843,In_1671,In_1389);
nor U1844 (N_1844,In_429,In_1927);
nand U1845 (N_1845,In_185,In_725);
nand U1846 (N_1846,In_853,In_1225);
or U1847 (N_1847,In_451,In_832);
and U1848 (N_1848,In_914,In_710);
nor U1849 (N_1849,In_1991,In_1438);
xor U1850 (N_1850,In_1354,In_245);
nand U1851 (N_1851,In_353,In_141);
xor U1852 (N_1852,In_697,In_743);
and U1853 (N_1853,In_569,In_1747);
nand U1854 (N_1854,In_1417,In_62);
and U1855 (N_1855,In_1539,In_1545);
xnor U1856 (N_1856,In_1628,In_1467);
nor U1857 (N_1857,In_10,In_342);
and U1858 (N_1858,In_1519,In_1876);
and U1859 (N_1859,In_1227,In_200);
and U1860 (N_1860,In_101,In_617);
xor U1861 (N_1861,In_473,In_1175);
or U1862 (N_1862,In_1737,In_482);
nand U1863 (N_1863,In_1161,In_1342);
xnor U1864 (N_1864,In_409,In_1299);
nor U1865 (N_1865,In_1336,In_979);
nand U1866 (N_1866,In_69,In_1969);
nand U1867 (N_1867,In_101,In_1);
nor U1868 (N_1868,In_1509,In_870);
xnor U1869 (N_1869,In_693,In_1699);
xor U1870 (N_1870,In_1317,In_1621);
nor U1871 (N_1871,In_1733,In_198);
nor U1872 (N_1872,In_1398,In_1409);
xor U1873 (N_1873,In_1820,In_306);
or U1874 (N_1874,In_1253,In_317);
nor U1875 (N_1875,In_173,In_666);
nor U1876 (N_1876,In_663,In_126);
nand U1877 (N_1877,In_172,In_977);
xnor U1878 (N_1878,In_1849,In_720);
or U1879 (N_1879,In_1943,In_681);
and U1880 (N_1880,In_147,In_1216);
nor U1881 (N_1881,In_741,In_1806);
nor U1882 (N_1882,In_1426,In_191);
and U1883 (N_1883,In_503,In_598);
nor U1884 (N_1884,In_825,In_1190);
xnor U1885 (N_1885,In_1921,In_729);
nor U1886 (N_1886,In_107,In_1171);
or U1887 (N_1887,In_1539,In_280);
nand U1888 (N_1888,In_599,In_1339);
nor U1889 (N_1889,In_790,In_1241);
or U1890 (N_1890,In_1703,In_1340);
nand U1891 (N_1891,In_1144,In_282);
nor U1892 (N_1892,In_1691,In_440);
or U1893 (N_1893,In_302,In_1710);
xor U1894 (N_1894,In_555,In_866);
or U1895 (N_1895,In_671,In_1123);
xor U1896 (N_1896,In_633,In_1533);
nand U1897 (N_1897,In_736,In_130);
nor U1898 (N_1898,In_1735,In_1104);
xnor U1899 (N_1899,In_1680,In_1785);
xor U1900 (N_1900,In_1759,In_1450);
nor U1901 (N_1901,In_741,In_1884);
or U1902 (N_1902,In_455,In_489);
and U1903 (N_1903,In_1945,In_1242);
xor U1904 (N_1904,In_246,In_1378);
and U1905 (N_1905,In_541,In_79);
xor U1906 (N_1906,In_1758,In_190);
xor U1907 (N_1907,In_548,In_364);
xor U1908 (N_1908,In_1440,In_1573);
or U1909 (N_1909,In_800,In_1469);
and U1910 (N_1910,In_1804,In_361);
or U1911 (N_1911,In_1805,In_49);
and U1912 (N_1912,In_1460,In_941);
or U1913 (N_1913,In_110,In_1990);
nand U1914 (N_1914,In_1111,In_455);
and U1915 (N_1915,In_302,In_1146);
nand U1916 (N_1916,In_370,In_340);
xor U1917 (N_1917,In_731,In_1616);
nand U1918 (N_1918,In_113,In_287);
nor U1919 (N_1919,In_898,In_1483);
nor U1920 (N_1920,In_969,In_661);
nand U1921 (N_1921,In_1913,In_180);
nor U1922 (N_1922,In_1140,In_1159);
nor U1923 (N_1923,In_236,In_1113);
xor U1924 (N_1924,In_820,In_1079);
nand U1925 (N_1925,In_1974,In_1682);
nand U1926 (N_1926,In_344,In_1032);
nand U1927 (N_1927,In_754,In_1266);
and U1928 (N_1928,In_229,In_1077);
and U1929 (N_1929,In_1560,In_917);
or U1930 (N_1930,In_1101,In_1666);
and U1931 (N_1931,In_1224,In_1445);
nand U1932 (N_1932,In_503,In_1109);
nand U1933 (N_1933,In_36,In_1262);
and U1934 (N_1934,In_1809,In_1671);
xnor U1935 (N_1935,In_1380,In_1829);
nand U1936 (N_1936,In_593,In_1354);
nor U1937 (N_1937,In_156,In_1680);
nor U1938 (N_1938,In_1702,In_876);
xor U1939 (N_1939,In_1930,In_740);
or U1940 (N_1940,In_1029,In_248);
xor U1941 (N_1941,In_1619,In_209);
and U1942 (N_1942,In_819,In_1746);
or U1943 (N_1943,In_1264,In_39);
or U1944 (N_1944,In_837,In_1040);
or U1945 (N_1945,In_103,In_795);
xnor U1946 (N_1946,In_590,In_739);
nand U1947 (N_1947,In_141,In_327);
xor U1948 (N_1948,In_564,In_173);
xor U1949 (N_1949,In_1419,In_45);
nand U1950 (N_1950,In_883,In_1507);
or U1951 (N_1951,In_839,In_732);
nor U1952 (N_1952,In_1594,In_667);
or U1953 (N_1953,In_622,In_1511);
and U1954 (N_1954,In_534,In_925);
or U1955 (N_1955,In_829,In_1745);
xnor U1956 (N_1956,In_1391,In_649);
nor U1957 (N_1957,In_1547,In_1015);
xnor U1958 (N_1958,In_1344,In_641);
nand U1959 (N_1959,In_1741,In_357);
or U1960 (N_1960,In_1424,In_20);
or U1961 (N_1961,In_1743,In_1473);
nand U1962 (N_1962,In_964,In_1297);
nand U1963 (N_1963,In_92,In_320);
or U1964 (N_1964,In_1011,In_511);
and U1965 (N_1965,In_1762,In_589);
nand U1966 (N_1966,In_197,In_1909);
xnor U1967 (N_1967,In_1787,In_562);
or U1968 (N_1968,In_1410,In_1164);
xor U1969 (N_1969,In_531,In_1822);
or U1970 (N_1970,In_1756,In_1445);
nor U1971 (N_1971,In_1378,In_338);
xor U1972 (N_1972,In_1319,In_90);
and U1973 (N_1973,In_598,In_1332);
xor U1974 (N_1974,In_135,In_1923);
or U1975 (N_1975,In_1721,In_1011);
nand U1976 (N_1976,In_1701,In_1199);
xor U1977 (N_1977,In_1199,In_1378);
nor U1978 (N_1978,In_154,In_703);
xnor U1979 (N_1979,In_1556,In_956);
nor U1980 (N_1980,In_1037,In_1536);
or U1981 (N_1981,In_1917,In_840);
xor U1982 (N_1982,In_871,In_1240);
xnor U1983 (N_1983,In_1976,In_179);
or U1984 (N_1984,In_915,In_1338);
nor U1985 (N_1985,In_393,In_202);
nor U1986 (N_1986,In_891,In_133);
and U1987 (N_1987,In_1672,In_405);
nor U1988 (N_1988,In_1505,In_885);
or U1989 (N_1989,In_1849,In_1777);
xor U1990 (N_1990,In_337,In_759);
xnor U1991 (N_1991,In_1913,In_1675);
xor U1992 (N_1992,In_130,In_1274);
xnor U1993 (N_1993,In_329,In_1364);
nor U1994 (N_1994,In_1239,In_642);
and U1995 (N_1995,In_1418,In_1724);
nor U1996 (N_1996,In_1085,In_157);
nor U1997 (N_1997,In_1674,In_1098);
or U1998 (N_1998,In_1426,In_1767);
or U1999 (N_1999,In_837,In_428);
or U2000 (N_2000,In_1284,In_512);
nand U2001 (N_2001,In_1127,In_1082);
or U2002 (N_2002,In_770,In_443);
and U2003 (N_2003,In_1539,In_299);
or U2004 (N_2004,In_386,In_1445);
nand U2005 (N_2005,In_1394,In_1428);
or U2006 (N_2006,In_355,In_249);
and U2007 (N_2007,In_1399,In_1665);
or U2008 (N_2008,In_746,In_1160);
nor U2009 (N_2009,In_110,In_1950);
and U2010 (N_2010,In_885,In_880);
xor U2011 (N_2011,In_1723,In_1928);
xnor U2012 (N_2012,In_1697,In_889);
nor U2013 (N_2013,In_1255,In_185);
and U2014 (N_2014,In_1098,In_662);
and U2015 (N_2015,In_202,In_1738);
nor U2016 (N_2016,In_399,In_912);
xor U2017 (N_2017,In_1422,In_454);
or U2018 (N_2018,In_1069,In_1922);
nor U2019 (N_2019,In_198,In_919);
nor U2020 (N_2020,In_1177,In_1057);
nand U2021 (N_2021,In_1465,In_959);
or U2022 (N_2022,In_1230,In_1618);
xor U2023 (N_2023,In_1101,In_1596);
and U2024 (N_2024,In_1469,In_1416);
nand U2025 (N_2025,In_1827,In_46);
or U2026 (N_2026,In_1261,In_742);
or U2027 (N_2027,In_1306,In_137);
or U2028 (N_2028,In_458,In_793);
xor U2029 (N_2029,In_1236,In_609);
and U2030 (N_2030,In_550,In_1662);
nor U2031 (N_2031,In_1387,In_1468);
and U2032 (N_2032,In_1408,In_592);
xnor U2033 (N_2033,In_1072,In_1656);
and U2034 (N_2034,In_1972,In_1892);
nor U2035 (N_2035,In_12,In_1164);
xor U2036 (N_2036,In_1589,In_1420);
xor U2037 (N_2037,In_1427,In_1181);
and U2038 (N_2038,In_983,In_776);
or U2039 (N_2039,In_890,In_120);
and U2040 (N_2040,In_1620,In_748);
nand U2041 (N_2041,In_1838,In_1652);
and U2042 (N_2042,In_865,In_1884);
nor U2043 (N_2043,In_1245,In_1548);
xnor U2044 (N_2044,In_973,In_1945);
or U2045 (N_2045,In_355,In_514);
nor U2046 (N_2046,In_817,In_341);
or U2047 (N_2047,In_468,In_1131);
or U2048 (N_2048,In_1017,In_10);
xnor U2049 (N_2049,In_1355,In_1687);
or U2050 (N_2050,In_1690,In_1818);
xor U2051 (N_2051,In_1465,In_1552);
or U2052 (N_2052,In_665,In_1361);
or U2053 (N_2053,In_624,In_643);
or U2054 (N_2054,In_656,In_553);
and U2055 (N_2055,In_414,In_1885);
nor U2056 (N_2056,In_1484,In_384);
nand U2057 (N_2057,In_47,In_1727);
xnor U2058 (N_2058,In_768,In_1094);
and U2059 (N_2059,In_884,In_377);
nor U2060 (N_2060,In_1250,In_1783);
and U2061 (N_2061,In_1655,In_204);
or U2062 (N_2062,In_1994,In_1068);
xnor U2063 (N_2063,In_591,In_667);
or U2064 (N_2064,In_749,In_276);
or U2065 (N_2065,In_809,In_1396);
and U2066 (N_2066,In_1081,In_925);
and U2067 (N_2067,In_1213,In_599);
and U2068 (N_2068,In_1363,In_1130);
and U2069 (N_2069,In_1760,In_898);
or U2070 (N_2070,In_269,In_1822);
and U2071 (N_2071,In_1188,In_910);
and U2072 (N_2072,In_960,In_396);
nor U2073 (N_2073,In_596,In_949);
nor U2074 (N_2074,In_1807,In_347);
or U2075 (N_2075,In_482,In_1180);
xor U2076 (N_2076,In_706,In_764);
nor U2077 (N_2077,In_390,In_257);
nor U2078 (N_2078,In_443,In_238);
nor U2079 (N_2079,In_780,In_302);
nand U2080 (N_2080,In_1617,In_1143);
or U2081 (N_2081,In_1421,In_119);
nor U2082 (N_2082,In_80,In_1437);
xor U2083 (N_2083,In_855,In_24);
and U2084 (N_2084,In_143,In_595);
or U2085 (N_2085,In_1441,In_1948);
nor U2086 (N_2086,In_497,In_255);
and U2087 (N_2087,In_1538,In_701);
and U2088 (N_2088,In_989,In_1489);
and U2089 (N_2089,In_1260,In_1392);
nand U2090 (N_2090,In_1508,In_1200);
or U2091 (N_2091,In_24,In_406);
nor U2092 (N_2092,In_1881,In_1556);
nand U2093 (N_2093,In_541,In_671);
xnor U2094 (N_2094,In_1079,In_1784);
xnor U2095 (N_2095,In_1982,In_295);
or U2096 (N_2096,In_469,In_619);
nor U2097 (N_2097,In_416,In_349);
xor U2098 (N_2098,In_1354,In_96);
or U2099 (N_2099,In_1980,In_1348);
xor U2100 (N_2100,In_1274,In_1836);
nand U2101 (N_2101,In_741,In_478);
nand U2102 (N_2102,In_1134,In_1484);
nor U2103 (N_2103,In_1968,In_503);
nand U2104 (N_2104,In_172,In_373);
nor U2105 (N_2105,In_118,In_375);
and U2106 (N_2106,In_683,In_1874);
and U2107 (N_2107,In_688,In_233);
nand U2108 (N_2108,In_1496,In_1873);
and U2109 (N_2109,In_1593,In_1482);
nand U2110 (N_2110,In_201,In_138);
nor U2111 (N_2111,In_1051,In_1973);
or U2112 (N_2112,In_1587,In_744);
nand U2113 (N_2113,In_880,In_151);
or U2114 (N_2114,In_54,In_352);
nor U2115 (N_2115,In_1343,In_1553);
nand U2116 (N_2116,In_1679,In_1084);
or U2117 (N_2117,In_708,In_1730);
xnor U2118 (N_2118,In_240,In_163);
xnor U2119 (N_2119,In_1259,In_1733);
nand U2120 (N_2120,In_1952,In_649);
nor U2121 (N_2121,In_243,In_882);
nand U2122 (N_2122,In_1310,In_274);
and U2123 (N_2123,In_1110,In_1895);
or U2124 (N_2124,In_1027,In_1270);
nor U2125 (N_2125,In_582,In_848);
or U2126 (N_2126,In_645,In_238);
nor U2127 (N_2127,In_1443,In_356);
xor U2128 (N_2128,In_1544,In_1337);
xnor U2129 (N_2129,In_1910,In_1017);
nand U2130 (N_2130,In_374,In_1978);
or U2131 (N_2131,In_403,In_1772);
nand U2132 (N_2132,In_877,In_1727);
and U2133 (N_2133,In_330,In_1120);
nor U2134 (N_2134,In_100,In_53);
nand U2135 (N_2135,In_1134,In_124);
xnor U2136 (N_2136,In_1449,In_1095);
nand U2137 (N_2137,In_354,In_47);
nand U2138 (N_2138,In_1466,In_122);
or U2139 (N_2139,In_125,In_1374);
or U2140 (N_2140,In_967,In_1999);
xor U2141 (N_2141,In_1899,In_967);
or U2142 (N_2142,In_612,In_1352);
nand U2143 (N_2143,In_864,In_1801);
or U2144 (N_2144,In_1895,In_1498);
nor U2145 (N_2145,In_1224,In_197);
nor U2146 (N_2146,In_1997,In_1414);
or U2147 (N_2147,In_1504,In_1645);
and U2148 (N_2148,In_1718,In_1041);
nor U2149 (N_2149,In_383,In_1489);
nand U2150 (N_2150,In_1076,In_329);
nor U2151 (N_2151,In_1377,In_1498);
xnor U2152 (N_2152,In_1490,In_1318);
xor U2153 (N_2153,In_1606,In_971);
nor U2154 (N_2154,In_1194,In_1380);
xor U2155 (N_2155,In_254,In_711);
and U2156 (N_2156,In_1643,In_709);
or U2157 (N_2157,In_1193,In_1460);
nor U2158 (N_2158,In_904,In_1626);
or U2159 (N_2159,In_1415,In_651);
or U2160 (N_2160,In_615,In_830);
or U2161 (N_2161,In_483,In_607);
and U2162 (N_2162,In_1718,In_1496);
or U2163 (N_2163,In_268,In_1409);
xor U2164 (N_2164,In_467,In_654);
and U2165 (N_2165,In_1685,In_1471);
nor U2166 (N_2166,In_155,In_737);
nor U2167 (N_2167,In_1727,In_435);
nor U2168 (N_2168,In_1702,In_1364);
or U2169 (N_2169,In_149,In_56);
nand U2170 (N_2170,In_1938,In_1069);
xnor U2171 (N_2171,In_486,In_1965);
nand U2172 (N_2172,In_1690,In_1799);
xnor U2173 (N_2173,In_1339,In_751);
and U2174 (N_2174,In_1338,In_653);
nand U2175 (N_2175,In_1537,In_1613);
nor U2176 (N_2176,In_962,In_1564);
nor U2177 (N_2177,In_11,In_1992);
nand U2178 (N_2178,In_1184,In_1147);
nand U2179 (N_2179,In_1726,In_59);
nand U2180 (N_2180,In_1252,In_480);
and U2181 (N_2181,In_957,In_1959);
xor U2182 (N_2182,In_322,In_1797);
or U2183 (N_2183,In_508,In_618);
nor U2184 (N_2184,In_1165,In_591);
nand U2185 (N_2185,In_808,In_1066);
or U2186 (N_2186,In_411,In_1561);
nor U2187 (N_2187,In_1929,In_1909);
and U2188 (N_2188,In_1216,In_14);
or U2189 (N_2189,In_1781,In_424);
nand U2190 (N_2190,In_24,In_1503);
nor U2191 (N_2191,In_784,In_465);
or U2192 (N_2192,In_980,In_840);
xnor U2193 (N_2193,In_939,In_732);
or U2194 (N_2194,In_425,In_651);
nor U2195 (N_2195,In_1363,In_254);
or U2196 (N_2196,In_1877,In_899);
xor U2197 (N_2197,In_1145,In_1220);
or U2198 (N_2198,In_819,In_480);
nor U2199 (N_2199,In_454,In_904);
xor U2200 (N_2200,In_1602,In_751);
or U2201 (N_2201,In_1680,In_1555);
or U2202 (N_2202,In_1519,In_123);
xor U2203 (N_2203,In_1088,In_1391);
nor U2204 (N_2204,In_95,In_561);
nand U2205 (N_2205,In_841,In_1139);
nor U2206 (N_2206,In_882,In_1870);
and U2207 (N_2207,In_1194,In_1542);
nand U2208 (N_2208,In_952,In_530);
and U2209 (N_2209,In_1844,In_791);
xor U2210 (N_2210,In_166,In_383);
nor U2211 (N_2211,In_1133,In_1598);
xnor U2212 (N_2212,In_758,In_126);
nand U2213 (N_2213,In_326,In_1782);
nand U2214 (N_2214,In_49,In_359);
and U2215 (N_2215,In_1988,In_367);
nor U2216 (N_2216,In_233,In_1443);
nand U2217 (N_2217,In_429,In_302);
xnor U2218 (N_2218,In_1829,In_665);
or U2219 (N_2219,In_622,In_1888);
or U2220 (N_2220,In_1893,In_109);
or U2221 (N_2221,In_171,In_910);
nand U2222 (N_2222,In_642,In_750);
nand U2223 (N_2223,In_305,In_643);
xnor U2224 (N_2224,In_1380,In_1066);
or U2225 (N_2225,In_382,In_1663);
xor U2226 (N_2226,In_1743,In_243);
or U2227 (N_2227,In_311,In_1489);
and U2228 (N_2228,In_992,In_1918);
nand U2229 (N_2229,In_823,In_1319);
and U2230 (N_2230,In_1843,In_1278);
nand U2231 (N_2231,In_1705,In_1856);
nor U2232 (N_2232,In_1256,In_1253);
or U2233 (N_2233,In_1816,In_653);
xnor U2234 (N_2234,In_1668,In_160);
or U2235 (N_2235,In_1328,In_267);
and U2236 (N_2236,In_850,In_844);
nand U2237 (N_2237,In_1385,In_476);
nand U2238 (N_2238,In_444,In_325);
nand U2239 (N_2239,In_805,In_388);
xnor U2240 (N_2240,In_855,In_1587);
xnor U2241 (N_2241,In_832,In_966);
nand U2242 (N_2242,In_1469,In_490);
or U2243 (N_2243,In_545,In_300);
and U2244 (N_2244,In_1232,In_1047);
or U2245 (N_2245,In_1428,In_1288);
nand U2246 (N_2246,In_405,In_594);
nand U2247 (N_2247,In_1573,In_1346);
and U2248 (N_2248,In_1783,In_1808);
nor U2249 (N_2249,In_1383,In_1371);
nand U2250 (N_2250,In_1929,In_170);
nor U2251 (N_2251,In_433,In_93);
nand U2252 (N_2252,In_1737,In_1328);
nor U2253 (N_2253,In_1401,In_1755);
nor U2254 (N_2254,In_626,In_197);
xor U2255 (N_2255,In_87,In_426);
nor U2256 (N_2256,In_218,In_1690);
nor U2257 (N_2257,In_859,In_464);
and U2258 (N_2258,In_910,In_1859);
nor U2259 (N_2259,In_274,In_986);
xor U2260 (N_2260,In_151,In_288);
and U2261 (N_2261,In_400,In_824);
xnor U2262 (N_2262,In_1581,In_1757);
nor U2263 (N_2263,In_1203,In_1054);
nor U2264 (N_2264,In_1214,In_1320);
xnor U2265 (N_2265,In_928,In_450);
xnor U2266 (N_2266,In_548,In_1931);
xor U2267 (N_2267,In_477,In_1993);
nor U2268 (N_2268,In_224,In_523);
nand U2269 (N_2269,In_1000,In_1399);
nand U2270 (N_2270,In_311,In_774);
nor U2271 (N_2271,In_1437,In_575);
and U2272 (N_2272,In_700,In_1580);
nand U2273 (N_2273,In_1916,In_4);
or U2274 (N_2274,In_1910,In_500);
and U2275 (N_2275,In_1191,In_1130);
or U2276 (N_2276,In_666,In_542);
nand U2277 (N_2277,In_1377,In_765);
nor U2278 (N_2278,In_1520,In_1042);
xnor U2279 (N_2279,In_1234,In_352);
nand U2280 (N_2280,In_820,In_1565);
nand U2281 (N_2281,In_1406,In_631);
nand U2282 (N_2282,In_1568,In_546);
or U2283 (N_2283,In_1843,In_198);
and U2284 (N_2284,In_1174,In_1182);
and U2285 (N_2285,In_1172,In_947);
nor U2286 (N_2286,In_74,In_663);
nor U2287 (N_2287,In_28,In_1675);
nand U2288 (N_2288,In_151,In_1419);
and U2289 (N_2289,In_953,In_760);
xor U2290 (N_2290,In_671,In_1055);
or U2291 (N_2291,In_581,In_1987);
xnor U2292 (N_2292,In_1340,In_1671);
and U2293 (N_2293,In_950,In_1035);
and U2294 (N_2294,In_772,In_1903);
or U2295 (N_2295,In_943,In_709);
xnor U2296 (N_2296,In_1283,In_1821);
xnor U2297 (N_2297,In_1109,In_663);
nand U2298 (N_2298,In_508,In_1368);
nor U2299 (N_2299,In_1845,In_86);
or U2300 (N_2300,In_891,In_982);
and U2301 (N_2301,In_1765,In_1938);
or U2302 (N_2302,In_1817,In_1265);
nand U2303 (N_2303,In_1218,In_410);
nor U2304 (N_2304,In_881,In_406);
xor U2305 (N_2305,In_441,In_29);
and U2306 (N_2306,In_1810,In_984);
or U2307 (N_2307,In_1689,In_1783);
or U2308 (N_2308,In_849,In_863);
xnor U2309 (N_2309,In_265,In_817);
or U2310 (N_2310,In_1245,In_55);
nor U2311 (N_2311,In_991,In_200);
nand U2312 (N_2312,In_486,In_608);
and U2313 (N_2313,In_620,In_136);
nand U2314 (N_2314,In_1719,In_635);
and U2315 (N_2315,In_172,In_1101);
nand U2316 (N_2316,In_1151,In_298);
or U2317 (N_2317,In_274,In_1001);
and U2318 (N_2318,In_177,In_641);
xor U2319 (N_2319,In_805,In_1021);
and U2320 (N_2320,In_23,In_1195);
nor U2321 (N_2321,In_894,In_463);
or U2322 (N_2322,In_30,In_1002);
and U2323 (N_2323,In_1587,In_1460);
nand U2324 (N_2324,In_1149,In_176);
xnor U2325 (N_2325,In_776,In_910);
and U2326 (N_2326,In_646,In_705);
nor U2327 (N_2327,In_888,In_893);
nor U2328 (N_2328,In_617,In_337);
nor U2329 (N_2329,In_267,In_1895);
nand U2330 (N_2330,In_59,In_1147);
nand U2331 (N_2331,In_222,In_115);
nor U2332 (N_2332,In_1580,In_1331);
or U2333 (N_2333,In_139,In_1642);
or U2334 (N_2334,In_1492,In_584);
or U2335 (N_2335,In_542,In_308);
nor U2336 (N_2336,In_1233,In_74);
nand U2337 (N_2337,In_1985,In_413);
or U2338 (N_2338,In_1261,In_1347);
xnor U2339 (N_2339,In_600,In_142);
and U2340 (N_2340,In_787,In_1484);
and U2341 (N_2341,In_752,In_1469);
nor U2342 (N_2342,In_1768,In_1289);
nor U2343 (N_2343,In_1887,In_1593);
nor U2344 (N_2344,In_8,In_926);
and U2345 (N_2345,In_1741,In_1354);
and U2346 (N_2346,In_443,In_1188);
nor U2347 (N_2347,In_717,In_902);
nor U2348 (N_2348,In_1958,In_1235);
or U2349 (N_2349,In_1088,In_1311);
and U2350 (N_2350,In_1742,In_1817);
nand U2351 (N_2351,In_827,In_324);
nor U2352 (N_2352,In_360,In_461);
xnor U2353 (N_2353,In_988,In_828);
and U2354 (N_2354,In_914,In_284);
nand U2355 (N_2355,In_727,In_1608);
and U2356 (N_2356,In_933,In_903);
xnor U2357 (N_2357,In_94,In_1240);
nor U2358 (N_2358,In_387,In_1025);
and U2359 (N_2359,In_13,In_725);
and U2360 (N_2360,In_29,In_1782);
nor U2361 (N_2361,In_523,In_1035);
xor U2362 (N_2362,In_1407,In_1360);
xor U2363 (N_2363,In_1561,In_237);
xnor U2364 (N_2364,In_927,In_795);
nand U2365 (N_2365,In_1116,In_1306);
or U2366 (N_2366,In_1364,In_168);
or U2367 (N_2367,In_671,In_1658);
xor U2368 (N_2368,In_1625,In_1440);
and U2369 (N_2369,In_1125,In_1058);
nand U2370 (N_2370,In_1269,In_1856);
nor U2371 (N_2371,In_1872,In_673);
and U2372 (N_2372,In_1124,In_503);
or U2373 (N_2373,In_140,In_402);
xor U2374 (N_2374,In_360,In_1733);
or U2375 (N_2375,In_1428,In_709);
and U2376 (N_2376,In_774,In_124);
nor U2377 (N_2377,In_1335,In_1702);
xor U2378 (N_2378,In_1352,In_493);
or U2379 (N_2379,In_874,In_1609);
nor U2380 (N_2380,In_235,In_1299);
nand U2381 (N_2381,In_164,In_377);
nor U2382 (N_2382,In_202,In_1886);
and U2383 (N_2383,In_1304,In_1086);
and U2384 (N_2384,In_1271,In_575);
xnor U2385 (N_2385,In_436,In_977);
and U2386 (N_2386,In_719,In_522);
xnor U2387 (N_2387,In_974,In_752);
and U2388 (N_2388,In_1994,In_571);
and U2389 (N_2389,In_594,In_1847);
or U2390 (N_2390,In_1449,In_648);
or U2391 (N_2391,In_384,In_1334);
xor U2392 (N_2392,In_188,In_1133);
nor U2393 (N_2393,In_380,In_207);
nand U2394 (N_2394,In_1665,In_466);
xnor U2395 (N_2395,In_1187,In_570);
nand U2396 (N_2396,In_1637,In_899);
nor U2397 (N_2397,In_1013,In_411);
xnor U2398 (N_2398,In_1788,In_161);
or U2399 (N_2399,In_792,In_1975);
nand U2400 (N_2400,In_1537,In_748);
nand U2401 (N_2401,In_1908,In_1686);
or U2402 (N_2402,In_186,In_589);
nor U2403 (N_2403,In_1524,In_678);
nand U2404 (N_2404,In_231,In_1250);
nor U2405 (N_2405,In_1441,In_1986);
nand U2406 (N_2406,In_1175,In_579);
and U2407 (N_2407,In_1917,In_1775);
or U2408 (N_2408,In_397,In_1025);
nor U2409 (N_2409,In_34,In_1895);
or U2410 (N_2410,In_1146,In_1136);
xor U2411 (N_2411,In_847,In_1204);
or U2412 (N_2412,In_755,In_1812);
xor U2413 (N_2413,In_242,In_662);
or U2414 (N_2414,In_1084,In_1860);
nor U2415 (N_2415,In_359,In_411);
nand U2416 (N_2416,In_531,In_681);
or U2417 (N_2417,In_440,In_161);
nand U2418 (N_2418,In_590,In_430);
nand U2419 (N_2419,In_996,In_1173);
nand U2420 (N_2420,In_478,In_91);
nand U2421 (N_2421,In_1196,In_453);
nand U2422 (N_2422,In_1013,In_301);
nand U2423 (N_2423,In_426,In_946);
nand U2424 (N_2424,In_1847,In_62);
nand U2425 (N_2425,In_1395,In_1787);
or U2426 (N_2426,In_447,In_766);
and U2427 (N_2427,In_17,In_82);
and U2428 (N_2428,In_1880,In_1225);
or U2429 (N_2429,In_309,In_1483);
nand U2430 (N_2430,In_267,In_859);
xor U2431 (N_2431,In_449,In_788);
xor U2432 (N_2432,In_1699,In_187);
or U2433 (N_2433,In_1435,In_1281);
nand U2434 (N_2434,In_1605,In_1606);
nor U2435 (N_2435,In_920,In_1781);
xnor U2436 (N_2436,In_1733,In_100);
nor U2437 (N_2437,In_188,In_585);
or U2438 (N_2438,In_1150,In_1132);
and U2439 (N_2439,In_189,In_1627);
or U2440 (N_2440,In_388,In_1197);
and U2441 (N_2441,In_1491,In_123);
nand U2442 (N_2442,In_1035,In_1674);
nand U2443 (N_2443,In_554,In_849);
and U2444 (N_2444,In_1942,In_87);
or U2445 (N_2445,In_958,In_774);
nand U2446 (N_2446,In_294,In_849);
xnor U2447 (N_2447,In_489,In_400);
and U2448 (N_2448,In_263,In_1648);
nor U2449 (N_2449,In_1682,In_1356);
nor U2450 (N_2450,In_1056,In_571);
nand U2451 (N_2451,In_1049,In_1754);
nand U2452 (N_2452,In_1472,In_1480);
nand U2453 (N_2453,In_1588,In_761);
nand U2454 (N_2454,In_451,In_1334);
xor U2455 (N_2455,In_179,In_1058);
nor U2456 (N_2456,In_1755,In_1954);
xnor U2457 (N_2457,In_422,In_348);
or U2458 (N_2458,In_601,In_520);
or U2459 (N_2459,In_1561,In_1206);
or U2460 (N_2460,In_833,In_704);
and U2461 (N_2461,In_567,In_1696);
or U2462 (N_2462,In_1269,In_1295);
or U2463 (N_2463,In_176,In_49);
xnor U2464 (N_2464,In_971,In_1230);
and U2465 (N_2465,In_1378,In_9);
xnor U2466 (N_2466,In_568,In_987);
nor U2467 (N_2467,In_1612,In_1239);
xnor U2468 (N_2468,In_1802,In_1494);
or U2469 (N_2469,In_1856,In_1022);
nor U2470 (N_2470,In_1337,In_1888);
and U2471 (N_2471,In_383,In_1069);
nor U2472 (N_2472,In_1680,In_782);
nor U2473 (N_2473,In_472,In_657);
and U2474 (N_2474,In_682,In_492);
nand U2475 (N_2475,In_541,In_714);
nand U2476 (N_2476,In_1300,In_1033);
xnor U2477 (N_2477,In_1734,In_1594);
and U2478 (N_2478,In_587,In_945);
nor U2479 (N_2479,In_385,In_803);
nor U2480 (N_2480,In_1425,In_218);
nand U2481 (N_2481,In_1806,In_1313);
and U2482 (N_2482,In_642,In_1033);
or U2483 (N_2483,In_41,In_1288);
and U2484 (N_2484,In_1695,In_925);
or U2485 (N_2485,In_1346,In_399);
nand U2486 (N_2486,In_406,In_1712);
nand U2487 (N_2487,In_1235,In_1084);
nor U2488 (N_2488,In_974,In_1051);
nand U2489 (N_2489,In_358,In_645);
nor U2490 (N_2490,In_1544,In_385);
nor U2491 (N_2491,In_1448,In_286);
xnor U2492 (N_2492,In_1771,In_1360);
nor U2493 (N_2493,In_1480,In_80);
nor U2494 (N_2494,In_1795,In_1191);
nand U2495 (N_2495,In_1138,In_622);
and U2496 (N_2496,In_399,In_1012);
and U2497 (N_2497,In_1468,In_909);
nor U2498 (N_2498,In_368,In_803);
or U2499 (N_2499,In_1579,In_1185);
nor U2500 (N_2500,In_1154,In_412);
nor U2501 (N_2501,In_416,In_291);
and U2502 (N_2502,In_948,In_353);
and U2503 (N_2503,In_1915,In_1031);
nor U2504 (N_2504,In_1217,In_720);
and U2505 (N_2505,In_1360,In_1440);
or U2506 (N_2506,In_898,In_892);
nand U2507 (N_2507,In_847,In_753);
xnor U2508 (N_2508,In_461,In_199);
xnor U2509 (N_2509,In_229,In_1246);
and U2510 (N_2510,In_1910,In_937);
nand U2511 (N_2511,In_1205,In_620);
nor U2512 (N_2512,In_1698,In_1324);
or U2513 (N_2513,In_229,In_1225);
and U2514 (N_2514,In_232,In_1552);
and U2515 (N_2515,In_1031,In_849);
or U2516 (N_2516,In_1736,In_1130);
nand U2517 (N_2517,In_785,In_752);
nor U2518 (N_2518,In_1614,In_990);
nand U2519 (N_2519,In_601,In_497);
nand U2520 (N_2520,In_1675,In_1251);
nand U2521 (N_2521,In_124,In_1718);
or U2522 (N_2522,In_1085,In_72);
and U2523 (N_2523,In_947,In_1256);
nor U2524 (N_2524,In_1770,In_873);
nor U2525 (N_2525,In_1018,In_1814);
nor U2526 (N_2526,In_827,In_1812);
xnor U2527 (N_2527,In_156,In_1193);
xnor U2528 (N_2528,In_491,In_1050);
xnor U2529 (N_2529,In_1491,In_665);
xor U2530 (N_2530,In_556,In_67);
nand U2531 (N_2531,In_405,In_472);
nor U2532 (N_2532,In_1465,In_1155);
nor U2533 (N_2533,In_823,In_1465);
nor U2534 (N_2534,In_250,In_780);
xor U2535 (N_2535,In_1851,In_752);
nor U2536 (N_2536,In_1239,In_1894);
nand U2537 (N_2537,In_722,In_122);
nor U2538 (N_2538,In_987,In_44);
nor U2539 (N_2539,In_495,In_717);
or U2540 (N_2540,In_1534,In_1246);
nor U2541 (N_2541,In_98,In_1069);
nand U2542 (N_2542,In_804,In_1091);
nand U2543 (N_2543,In_25,In_1264);
or U2544 (N_2544,In_663,In_1702);
nand U2545 (N_2545,In_34,In_1575);
xnor U2546 (N_2546,In_473,In_665);
nand U2547 (N_2547,In_585,In_1694);
nand U2548 (N_2548,In_471,In_970);
nor U2549 (N_2549,In_1961,In_7);
and U2550 (N_2550,In_1331,In_1072);
or U2551 (N_2551,In_972,In_1199);
nand U2552 (N_2552,In_1514,In_1067);
and U2553 (N_2553,In_1705,In_439);
nand U2554 (N_2554,In_132,In_574);
xnor U2555 (N_2555,In_1670,In_1328);
or U2556 (N_2556,In_1287,In_1512);
or U2557 (N_2557,In_642,In_781);
nand U2558 (N_2558,In_1798,In_957);
nor U2559 (N_2559,In_563,In_991);
xnor U2560 (N_2560,In_1524,In_493);
nor U2561 (N_2561,In_1108,In_391);
or U2562 (N_2562,In_589,In_643);
and U2563 (N_2563,In_173,In_1040);
or U2564 (N_2564,In_1301,In_589);
xnor U2565 (N_2565,In_497,In_428);
nand U2566 (N_2566,In_185,In_1980);
nand U2567 (N_2567,In_1389,In_983);
xor U2568 (N_2568,In_912,In_663);
nand U2569 (N_2569,In_1621,In_78);
xor U2570 (N_2570,In_1995,In_52);
nor U2571 (N_2571,In_274,In_1736);
nand U2572 (N_2572,In_1367,In_1603);
nor U2573 (N_2573,In_1884,In_1097);
xor U2574 (N_2574,In_1831,In_1486);
or U2575 (N_2575,In_480,In_1470);
and U2576 (N_2576,In_84,In_1739);
or U2577 (N_2577,In_865,In_1783);
nor U2578 (N_2578,In_1623,In_1107);
and U2579 (N_2579,In_331,In_1583);
or U2580 (N_2580,In_168,In_416);
xor U2581 (N_2581,In_171,In_1520);
or U2582 (N_2582,In_576,In_895);
nor U2583 (N_2583,In_203,In_778);
nor U2584 (N_2584,In_1433,In_51);
nor U2585 (N_2585,In_999,In_829);
nand U2586 (N_2586,In_1345,In_428);
or U2587 (N_2587,In_1396,In_54);
nor U2588 (N_2588,In_429,In_229);
nand U2589 (N_2589,In_1899,In_135);
xor U2590 (N_2590,In_550,In_419);
or U2591 (N_2591,In_1786,In_505);
or U2592 (N_2592,In_1786,In_808);
and U2593 (N_2593,In_797,In_72);
nand U2594 (N_2594,In_1501,In_1590);
and U2595 (N_2595,In_1712,In_1509);
and U2596 (N_2596,In_696,In_1901);
or U2597 (N_2597,In_1713,In_424);
xor U2598 (N_2598,In_379,In_687);
nand U2599 (N_2599,In_823,In_1326);
and U2600 (N_2600,In_1403,In_1442);
and U2601 (N_2601,In_1936,In_935);
nor U2602 (N_2602,In_1182,In_1921);
and U2603 (N_2603,In_1860,In_503);
or U2604 (N_2604,In_1671,In_1495);
nand U2605 (N_2605,In_895,In_1952);
nand U2606 (N_2606,In_734,In_234);
nor U2607 (N_2607,In_1507,In_1908);
nand U2608 (N_2608,In_876,In_944);
nand U2609 (N_2609,In_1656,In_1490);
or U2610 (N_2610,In_768,In_1905);
and U2611 (N_2611,In_1622,In_55);
or U2612 (N_2612,In_198,In_721);
and U2613 (N_2613,In_1866,In_1825);
xnor U2614 (N_2614,In_388,In_243);
xor U2615 (N_2615,In_1854,In_334);
nand U2616 (N_2616,In_475,In_1385);
and U2617 (N_2617,In_606,In_115);
and U2618 (N_2618,In_1929,In_1679);
and U2619 (N_2619,In_1791,In_1090);
nor U2620 (N_2620,In_1547,In_621);
or U2621 (N_2621,In_1202,In_782);
or U2622 (N_2622,In_359,In_1382);
and U2623 (N_2623,In_561,In_1939);
xnor U2624 (N_2624,In_1264,In_1581);
and U2625 (N_2625,In_456,In_844);
xor U2626 (N_2626,In_957,In_1108);
nor U2627 (N_2627,In_393,In_1038);
xnor U2628 (N_2628,In_1218,In_1641);
nand U2629 (N_2629,In_424,In_1183);
and U2630 (N_2630,In_680,In_768);
nor U2631 (N_2631,In_1733,In_83);
or U2632 (N_2632,In_946,In_1934);
and U2633 (N_2633,In_878,In_1205);
nand U2634 (N_2634,In_722,In_194);
nand U2635 (N_2635,In_1762,In_159);
nand U2636 (N_2636,In_788,In_1154);
and U2637 (N_2637,In_671,In_1403);
nor U2638 (N_2638,In_938,In_1178);
or U2639 (N_2639,In_1223,In_1519);
nand U2640 (N_2640,In_1291,In_949);
nor U2641 (N_2641,In_738,In_1581);
nor U2642 (N_2642,In_293,In_1356);
xor U2643 (N_2643,In_918,In_1003);
nand U2644 (N_2644,In_647,In_679);
and U2645 (N_2645,In_1812,In_816);
and U2646 (N_2646,In_714,In_580);
or U2647 (N_2647,In_878,In_1427);
nor U2648 (N_2648,In_3,In_1731);
or U2649 (N_2649,In_1700,In_584);
xnor U2650 (N_2650,In_1257,In_1544);
or U2651 (N_2651,In_893,In_471);
and U2652 (N_2652,In_959,In_429);
nor U2653 (N_2653,In_888,In_408);
nor U2654 (N_2654,In_23,In_681);
nor U2655 (N_2655,In_1162,In_269);
or U2656 (N_2656,In_1350,In_1910);
and U2657 (N_2657,In_619,In_1204);
xnor U2658 (N_2658,In_896,In_1518);
or U2659 (N_2659,In_890,In_1671);
nor U2660 (N_2660,In_1378,In_113);
nor U2661 (N_2661,In_1161,In_1312);
xor U2662 (N_2662,In_1077,In_1975);
xor U2663 (N_2663,In_1553,In_1392);
or U2664 (N_2664,In_453,In_1230);
nand U2665 (N_2665,In_610,In_1683);
and U2666 (N_2666,In_721,In_940);
nand U2667 (N_2667,In_1796,In_498);
nor U2668 (N_2668,In_1366,In_1830);
xnor U2669 (N_2669,In_1642,In_88);
or U2670 (N_2670,In_356,In_982);
or U2671 (N_2671,In_675,In_1484);
xnor U2672 (N_2672,In_1957,In_1457);
or U2673 (N_2673,In_1580,In_880);
and U2674 (N_2674,In_644,In_1913);
and U2675 (N_2675,In_1879,In_315);
nor U2676 (N_2676,In_1528,In_952);
nand U2677 (N_2677,In_6,In_1861);
nor U2678 (N_2678,In_1811,In_1416);
nor U2679 (N_2679,In_137,In_135);
and U2680 (N_2680,In_143,In_1152);
and U2681 (N_2681,In_760,In_1816);
nor U2682 (N_2682,In_756,In_1207);
nor U2683 (N_2683,In_1706,In_1582);
nand U2684 (N_2684,In_809,In_1086);
and U2685 (N_2685,In_1075,In_314);
nor U2686 (N_2686,In_1469,In_1872);
xnor U2687 (N_2687,In_912,In_939);
nand U2688 (N_2688,In_674,In_1140);
xnor U2689 (N_2689,In_649,In_216);
or U2690 (N_2690,In_1695,In_1807);
nand U2691 (N_2691,In_1796,In_45);
or U2692 (N_2692,In_1095,In_1723);
and U2693 (N_2693,In_1399,In_1815);
xor U2694 (N_2694,In_1249,In_1346);
or U2695 (N_2695,In_1043,In_879);
nor U2696 (N_2696,In_218,In_1090);
or U2697 (N_2697,In_858,In_1108);
nor U2698 (N_2698,In_1818,In_290);
or U2699 (N_2699,In_1502,In_893);
and U2700 (N_2700,In_1925,In_1907);
xnor U2701 (N_2701,In_188,In_716);
xor U2702 (N_2702,In_1321,In_1836);
nor U2703 (N_2703,In_812,In_1596);
nor U2704 (N_2704,In_1530,In_99);
nand U2705 (N_2705,In_214,In_1112);
nor U2706 (N_2706,In_1742,In_1699);
and U2707 (N_2707,In_1996,In_577);
or U2708 (N_2708,In_1010,In_824);
or U2709 (N_2709,In_664,In_75);
nor U2710 (N_2710,In_1121,In_1901);
or U2711 (N_2711,In_1129,In_1080);
or U2712 (N_2712,In_822,In_1718);
xor U2713 (N_2713,In_24,In_1352);
and U2714 (N_2714,In_1790,In_1307);
nand U2715 (N_2715,In_1142,In_123);
xor U2716 (N_2716,In_1002,In_424);
nand U2717 (N_2717,In_613,In_1563);
and U2718 (N_2718,In_1850,In_1059);
or U2719 (N_2719,In_1887,In_1741);
and U2720 (N_2720,In_82,In_1090);
nor U2721 (N_2721,In_698,In_1064);
or U2722 (N_2722,In_181,In_1670);
nand U2723 (N_2723,In_1569,In_709);
nor U2724 (N_2724,In_673,In_834);
nand U2725 (N_2725,In_1921,In_81);
or U2726 (N_2726,In_1653,In_1661);
xor U2727 (N_2727,In_1880,In_1465);
xnor U2728 (N_2728,In_853,In_1534);
nand U2729 (N_2729,In_140,In_1251);
nand U2730 (N_2730,In_176,In_937);
xnor U2731 (N_2731,In_911,In_1458);
nand U2732 (N_2732,In_1109,In_274);
xor U2733 (N_2733,In_1037,In_1542);
nor U2734 (N_2734,In_1,In_760);
nor U2735 (N_2735,In_1121,In_465);
nand U2736 (N_2736,In_1812,In_586);
and U2737 (N_2737,In_758,In_1361);
nor U2738 (N_2738,In_594,In_1202);
and U2739 (N_2739,In_292,In_1313);
and U2740 (N_2740,In_323,In_417);
or U2741 (N_2741,In_73,In_698);
and U2742 (N_2742,In_196,In_493);
xnor U2743 (N_2743,In_679,In_999);
and U2744 (N_2744,In_935,In_449);
nand U2745 (N_2745,In_1541,In_1843);
and U2746 (N_2746,In_1551,In_1230);
xor U2747 (N_2747,In_245,In_894);
or U2748 (N_2748,In_1530,In_1678);
nor U2749 (N_2749,In_157,In_1632);
nor U2750 (N_2750,In_620,In_1283);
xnor U2751 (N_2751,In_738,In_1279);
and U2752 (N_2752,In_1330,In_1951);
or U2753 (N_2753,In_1308,In_1398);
or U2754 (N_2754,In_1356,In_402);
nor U2755 (N_2755,In_521,In_1526);
xnor U2756 (N_2756,In_1197,In_1646);
xnor U2757 (N_2757,In_1176,In_1079);
nor U2758 (N_2758,In_2,In_1779);
xnor U2759 (N_2759,In_1860,In_1352);
or U2760 (N_2760,In_1519,In_1954);
xnor U2761 (N_2761,In_765,In_1907);
and U2762 (N_2762,In_73,In_1139);
or U2763 (N_2763,In_1361,In_1953);
and U2764 (N_2764,In_1996,In_1243);
nor U2765 (N_2765,In_296,In_1233);
or U2766 (N_2766,In_946,In_669);
and U2767 (N_2767,In_1113,In_341);
or U2768 (N_2768,In_30,In_718);
xor U2769 (N_2769,In_670,In_1077);
or U2770 (N_2770,In_1119,In_705);
and U2771 (N_2771,In_405,In_1537);
and U2772 (N_2772,In_1602,In_1524);
xor U2773 (N_2773,In_1388,In_1600);
xnor U2774 (N_2774,In_1633,In_490);
xor U2775 (N_2775,In_248,In_154);
or U2776 (N_2776,In_642,In_1971);
nor U2777 (N_2777,In_1082,In_1018);
and U2778 (N_2778,In_1775,In_1326);
or U2779 (N_2779,In_566,In_1297);
or U2780 (N_2780,In_676,In_550);
nor U2781 (N_2781,In_502,In_186);
and U2782 (N_2782,In_611,In_1013);
nand U2783 (N_2783,In_1006,In_1044);
and U2784 (N_2784,In_121,In_1372);
and U2785 (N_2785,In_361,In_8);
or U2786 (N_2786,In_781,In_1587);
and U2787 (N_2787,In_485,In_1553);
or U2788 (N_2788,In_619,In_548);
nor U2789 (N_2789,In_917,In_1628);
xnor U2790 (N_2790,In_957,In_1594);
nor U2791 (N_2791,In_866,In_228);
nor U2792 (N_2792,In_818,In_216);
and U2793 (N_2793,In_1373,In_468);
nor U2794 (N_2794,In_662,In_94);
or U2795 (N_2795,In_1486,In_693);
nand U2796 (N_2796,In_995,In_1161);
or U2797 (N_2797,In_1804,In_1178);
xor U2798 (N_2798,In_361,In_417);
nand U2799 (N_2799,In_1969,In_799);
and U2800 (N_2800,In_1973,In_1258);
or U2801 (N_2801,In_1160,In_304);
or U2802 (N_2802,In_407,In_275);
xor U2803 (N_2803,In_1159,In_1871);
and U2804 (N_2804,In_688,In_1905);
xnor U2805 (N_2805,In_1463,In_1726);
or U2806 (N_2806,In_221,In_1278);
or U2807 (N_2807,In_1159,In_1024);
nor U2808 (N_2808,In_1514,In_207);
nand U2809 (N_2809,In_680,In_1094);
xor U2810 (N_2810,In_85,In_1540);
and U2811 (N_2811,In_1817,In_711);
xnor U2812 (N_2812,In_548,In_770);
nand U2813 (N_2813,In_1053,In_54);
nor U2814 (N_2814,In_458,In_134);
nand U2815 (N_2815,In_182,In_50);
nor U2816 (N_2816,In_709,In_1649);
or U2817 (N_2817,In_1201,In_107);
or U2818 (N_2818,In_1910,In_1682);
nand U2819 (N_2819,In_1085,In_1195);
and U2820 (N_2820,In_782,In_1065);
xor U2821 (N_2821,In_1805,In_1100);
nor U2822 (N_2822,In_1109,In_1917);
and U2823 (N_2823,In_1168,In_1035);
nand U2824 (N_2824,In_993,In_1205);
or U2825 (N_2825,In_1042,In_356);
xor U2826 (N_2826,In_952,In_1639);
and U2827 (N_2827,In_1481,In_1997);
or U2828 (N_2828,In_179,In_768);
nand U2829 (N_2829,In_1282,In_1775);
nand U2830 (N_2830,In_1585,In_742);
nor U2831 (N_2831,In_1732,In_1809);
and U2832 (N_2832,In_228,In_1154);
xor U2833 (N_2833,In_1451,In_172);
xnor U2834 (N_2834,In_26,In_1776);
or U2835 (N_2835,In_1018,In_372);
xor U2836 (N_2836,In_1612,In_201);
xnor U2837 (N_2837,In_631,In_1603);
nand U2838 (N_2838,In_1332,In_48);
xnor U2839 (N_2839,In_929,In_357);
or U2840 (N_2840,In_208,In_1768);
nor U2841 (N_2841,In_179,In_1793);
nor U2842 (N_2842,In_229,In_889);
and U2843 (N_2843,In_1680,In_191);
and U2844 (N_2844,In_1475,In_637);
or U2845 (N_2845,In_31,In_1650);
nand U2846 (N_2846,In_1699,In_19);
nor U2847 (N_2847,In_621,In_1914);
or U2848 (N_2848,In_1131,In_1992);
or U2849 (N_2849,In_262,In_778);
or U2850 (N_2850,In_1883,In_354);
nor U2851 (N_2851,In_687,In_950);
and U2852 (N_2852,In_630,In_1065);
nand U2853 (N_2853,In_70,In_644);
or U2854 (N_2854,In_1471,In_351);
nand U2855 (N_2855,In_1758,In_1939);
xnor U2856 (N_2856,In_870,In_971);
or U2857 (N_2857,In_180,In_343);
nor U2858 (N_2858,In_694,In_429);
xnor U2859 (N_2859,In_987,In_1624);
and U2860 (N_2860,In_1752,In_1650);
and U2861 (N_2861,In_1187,In_1261);
nand U2862 (N_2862,In_1712,In_1416);
and U2863 (N_2863,In_1457,In_341);
nand U2864 (N_2864,In_1172,In_1971);
xnor U2865 (N_2865,In_1857,In_1193);
xnor U2866 (N_2866,In_1775,In_1921);
nor U2867 (N_2867,In_1268,In_711);
and U2868 (N_2868,In_993,In_659);
nor U2869 (N_2869,In_1685,In_396);
xor U2870 (N_2870,In_556,In_89);
xnor U2871 (N_2871,In_1190,In_1577);
nor U2872 (N_2872,In_1490,In_884);
nor U2873 (N_2873,In_1702,In_226);
or U2874 (N_2874,In_920,In_520);
nor U2875 (N_2875,In_1121,In_951);
or U2876 (N_2876,In_702,In_984);
nor U2877 (N_2877,In_134,In_487);
xor U2878 (N_2878,In_904,In_1042);
nand U2879 (N_2879,In_1602,In_162);
xor U2880 (N_2880,In_1963,In_439);
and U2881 (N_2881,In_1677,In_1727);
or U2882 (N_2882,In_867,In_411);
or U2883 (N_2883,In_1163,In_261);
nor U2884 (N_2884,In_1937,In_31);
nand U2885 (N_2885,In_435,In_246);
nor U2886 (N_2886,In_1265,In_460);
nor U2887 (N_2887,In_1691,In_877);
xnor U2888 (N_2888,In_1448,In_304);
xnor U2889 (N_2889,In_400,In_884);
nor U2890 (N_2890,In_467,In_522);
and U2891 (N_2891,In_228,In_568);
nand U2892 (N_2892,In_555,In_358);
nand U2893 (N_2893,In_651,In_1240);
nand U2894 (N_2894,In_201,In_1954);
nor U2895 (N_2895,In_81,In_1957);
or U2896 (N_2896,In_583,In_1212);
nor U2897 (N_2897,In_1710,In_1723);
nor U2898 (N_2898,In_44,In_1875);
nor U2899 (N_2899,In_839,In_295);
nor U2900 (N_2900,In_1289,In_734);
and U2901 (N_2901,In_1946,In_1193);
and U2902 (N_2902,In_1787,In_928);
xnor U2903 (N_2903,In_1482,In_599);
or U2904 (N_2904,In_901,In_110);
xnor U2905 (N_2905,In_97,In_279);
or U2906 (N_2906,In_1737,In_878);
nor U2907 (N_2907,In_1564,In_1292);
nor U2908 (N_2908,In_1747,In_1827);
and U2909 (N_2909,In_1843,In_1703);
nand U2910 (N_2910,In_1678,In_1151);
nor U2911 (N_2911,In_761,In_924);
nor U2912 (N_2912,In_1674,In_1102);
nand U2913 (N_2913,In_1032,In_747);
nor U2914 (N_2914,In_1432,In_1282);
and U2915 (N_2915,In_566,In_1426);
nor U2916 (N_2916,In_1738,In_1047);
and U2917 (N_2917,In_741,In_430);
nor U2918 (N_2918,In_1709,In_1458);
xnor U2919 (N_2919,In_1549,In_1672);
nand U2920 (N_2920,In_1995,In_870);
nor U2921 (N_2921,In_1786,In_1433);
or U2922 (N_2922,In_1136,In_610);
xor U2923 (N_2923,In_1452,In_169);
nor U2924 (N_2924,In_1074,In_679);
nand U2925 (N_2925,In_183,In_616);
nand U2926 (N_2926,In_158,In_1303);
and U2927 (N_2927,In_847,In_1618);
xor U2928 (N_2928,In_1631,In_436);
xor U2929 (N_2929,In_707,In_608);
and U2930 (N_2930,In_1264,In_727);
xnor U2931 (N_2931,In_272,In_1403);
nor U2932 (N_2932,In_1544,In_483);
xnor U2933 (N_2933,In_1155,In_1788);
xnor U2934 (N_2934,In_1091,In_1690);
nor U2935 (N_2935,In_40,In_1657);
or U2936 (N_2936,In_860,In_35);
or U2937 (N_2937,In_404,In_287);
nor U2938 (N_2938,In_557,In_997);
nand U2939 (N_2939,In_800,In_1128);
xor U2940 (N_2940,In_721,In_687);
xnor U2941 (N_2941,In_705,In_1896);
and U2942 (N_2942,In_739,In_1755);
xor U2943 (N_2943,In_1644,In_1910);
nor U2944 (N_2944,In_541,In_701);
and U2945 (N_2945,In_1391,In_1750);
or U2946 (N_2946,In_1854,In_554);
nand U2947 (N_2947,In_382,In_505);
nand U2948 (N_2948,In_1166,In_20);
nor U2949 (N_2949,In_1837,In_1061);
or U2950 (N_2950,In_780,In_562);
nand U2951 (N_2951,In_27,In_88);
and U2952 (N_2952,In_523,In_1969);
nand U2953 (N_2953,In_1940,In_1114);
nand U2954 (N_2954,In_1531,In_659);
nor U2955 (N_2955,In_1297,In_656);
or U2956 (N_2956,In_1191,In_1402);
nand U2957 (N_2957,In_152,In_239);
xnor U2958 (N_2958,In_1464,In_900);
xnor U2959 (N_2959,In_1895,In_1641);
and U2960 (N_2960,In_60,In_1630);
nand U2961 (N_2961,In_1615,In_326);
nor U2962 (N_2962,In_1899,In_1689);
xor U2963 (N_2963,In_930,In_292);
nand U2964 (N_2964,In_1946,In_33);
or U2965 (N_2965,In_1244,In_1165);
nor U2966 (N_2966,In_115,In_1924);
nor U2967 (N_2967,In_1918,In_836);
xor U2968 (N_2968,In_808,In_1528);
nand U2969 (N_2969,In_1781,In_115);
or U2970 (N_2970,In_1901,In_1514);
nor U2971 (N_2971,In_1745,In_1626);
or U2972 (N_2972,In_61,In_1941);
nand U2973 (N_2973,In_547,In_1856);
nand U2974 (N_2974,In_772,In_262);
nand U2975 (N_2975,In_1519,In_988);
nand U2976 (N_2976,In_69,In_351);
nand U2977 (N_2977,In_324,In_1970);
xor U2978 (N_2978,In_821,In_904);
and U2979 (N_2979,In_1740,In_40);
nand U2980 (N_2980,In_1270,In_448);
nor U2981 (N_2981,In_1785,In_1820);
and U2982 (N_2982,In_1472,In_815);
and U2983 (N_2983,In_915,In_106);
nand U2984 (N_2984,In_774,In_1879);
xor U2985 (N_2985,In_1293,In_719);
xor U2986 (N_2986,In_754,In_1962);
nor U2987 (N_2987,In_829,In_1087);
and U2988 (N_2988,In_1382,In_1331);
and U2989 (N_2989,In_523,In_1944);
nor U2990 (N_2990,In_1614,In_957);
xor U2991 (N_2991,In_1624,In_1187);
xnor U2992 (N_2992,In_174,In_1224);
or U2993 (N_2993,In_1604,In_284);
nor U2994 (N_2994,In_466,In_813);
or U2995 (N_2995,In_901,In_1442);
xor U2996 (N_2996,In_502,In_539);
nor U2997 (N_2997,In_1277,In_1);
xor U2998 (N_2998,In_1101,In_1463);
and U2999 (N_2999,In_574,In_1278);
and U3000 (N_3000,In_1369,In_409);
or U3001 (N_3001,In_1539,In_833);
xor U3002 (N_3002,In_252,In_529);
nor U3003 (N_3003,In_643,In_1007);
or U3004 (N_3004,In_1794,In_1819);
or U3005 (N_3005,In_24,In_1654);
nor U3006 (N_3006,In_1953,In_1538);
and U3007 (N_3007,In_1157,In_1038);
nand U3008 (N_3008,In_313,In_1349);
nor U3009 (N_3009,In_1740,In_671);
xnor U3010 (N_3010,In_1568,In_769);
nand U3011 (N_3011,In_601,In_616);
xnor U3012 (N_3012,In_1636,In_627);
nand U3013 (N_3013,In_641,In_1741);
or U3014 (N_3014,In_1991,In_1466);
and U3015 (N_3015,In_198,In_697);
or U3016 (N_3016,In_784,In_1229);
or U3017 (N_3017,In_123,In_1801);
nor U3018 (N_3018,In_1578,In_144);
xnor U3019 (N_3019,In_1782,In_1484);
xor U3020 (N_3020,In_1771,In_1576);
xnor U3021 (N_3021,In_1667,In_940);
and U3022 (N_3022,In_1522,In_462);
xnor U3023 (N_3023,In_479,In_1945);
or U3024 (N_3024,In_384,In_1180);
nor U3025 (N_3025,In_1687,In_874);
or U3026 (N_3026,In_1584,In_214);
nor U3027 (N_3027,In_239,In_1014);
and U3028 (N_3028,In_652,In_102);
nand U3029 (N_3029,In_1688,In_1304);
xor U3030 (N_3030,In_1811,In_1733);
nand U3031 (N_3031,In_1797,In_18);
and U3032 (N_3032,In_1487,In_757);
nor U3033 (N_3033,In_1615,In_1726);
nand U3034 (N_3034,In_169,In_532);
and U3035 (N_3035,In_1927,In_613);
nor U3036 (N_3036,In_24,In_204);
and U3037 (N_3037,In_887,In_292);
nor U3038 (N_3038,In_143,In_41);
or U3039 (N_3039,In_1255,In_581);
and U3040 (N_3040,In_753,In_115);
or U3041 (N_3041,In_670,In_1528);
xnor U3042 (N_3042,In_1163,In_1231);
and U3043 (N_3043,In_848,In_1010);
nand U3044 (N_3044,In_1633,In_1258);
and U3045 (N_3045,In_1319,In_1580);
xor U3046 (N_3046,In_1847,In_230);
nor U3047 (N_3047,In_340,In_657);
xor U3048 (N_3048,In_90,In_1196);
xor U3049 (N_3049,In_796,In_442);
nor U3050 (N_3050,In_1237,In_563);
and U3051 (N_3051,In_102,In_1328);
and U3052 (N_3052,In_312,In_196);
nor U3053 (N_3053,In_1962,In_1045);
nor U3054 (N_3054,In_1902,In_1483);
xnor U3055 (N_3055,In_1424,In_652);
nor U3056 (N_3056,In_451,In_1961);
nand U3057 (N_3057,In_51,In_436);
nand U3058 (N_3058,In_467,In_1085);
or U3059 (N_3059,In_1473,In_196);
xnor U3060 (N_3060,In_1865,In_1685);
nand U3061 (N_3061,In_1046,In_1584);
or U3062 (N_3062,In_734,In_961);
nand U3063 (N_3063,In_1233,In_1565);
xnor U3064 (N_3064,In_1392,In_1666);
xor U3065 (N_3065,In_739,In_1677);
and U3066 (N_3066,In_838,In_132);
nand U3067 (N_3067,In_902,In_1434);
nand U3068 (N_3068,In_227,In_342);
xor U3069 (N_3069,In_718,In_1823);
nand U3070 (N_3070,In_1003,In_893);
and U3071 (N_3071,In_1790,In_1942);
and U3072 (N_3072,In_955,In_1656);
xnor U3073 (N_3073,In_149,In_1388);
xnor U3074 (N_3074,In_286,In_652);
and U3075 (N_3075,In_1278,In_123);
nor U3076 (N_3076,In_1651,In_1967);
xnor U3077 (N_3077,In_1401,In_15);
and U3078 (N_3078,In_860,In_1349);
nor U3079 (N_3079,In_973,In_1557);
and U3080 (N_3080,In_1685,In_1436);
nor U3081 (N_3081,In_1075,In_508);
nand U3082 (N_3082,In_1272,In_100);
xor U3083 (N_3083,In_68,In_1661);
or U3084 (N_3084,In_1822,In_691);
and U3085 (N_3085,In_1231,In_1011);
nand U3086 (N_3086,In_408,In_1831);
and U3087 (N_3087,In_1413,In_973);
xnor U3088 (N_3088,In_602,In_1474);
nor U3089 (N_3089,In_730,In_506);
nor U3090 (N_3090,In_79,In_10);
xnor U3091 (N_3091,In_82,In_812);
xor U3092 (N_3092,In_686,In_1867);
xor U3093 (N_3093,In_108,In_1737);
nor U3094 (N_3094,In_1651,In_131);
and U3095 (N_3095,In_1268,In_1332);
nor U3096 (N_3096,In_1127,In_830);
nor U3097 (N_3097,In_566,In_1183);
and U3098 (N_3098,In_546,In_1761);
and U3099 (N_3099,In_558,In_44);
nor U3100 (N_3100,In_365,In_808);
and U3101 (N_3101,In_706,In_456);
xor U3102 (N_3102,In_1953,In_417);
xnor U3103 (N_3103,In_1376,In_276);
xor U3104 (N_3104,In_157,In_599);
xnor U3105 (N_3105,In_1609,In_1724);
xnor U3106 (N_3106,In_553,In_1403);
xor U3107 (N_3107,In_1313,In_143);
and U3108 (N_3108,In_412,In_335);
nand U3109 (N_3109,In_1285,In_1543);
and U3110 (N_3110,In_1774,In_296);
and U3111 (N_3111,In_877,In_1564);
and U3112 (N_3112,In_189,In_1667);
and U3113 (N_3113,In_1857,In_385);
nor U3114 (N_3114,In_781,In_1720);
xnor U3115 (N_3115,In_103,In_1366);
and U3116 (N_3116,In_1898,In_1811);
or U3117 (N_3117,In_413,In_918);
or U3118 (N_3118,In_1656,In_1189);
nand U3119 (N_3119,In_669,In_431);
and U3120 (N_3120,In_51,In_1375);
nor U3121 (N_3121,In_1755,In_2);
xor U3122 (N_3122,In_408,In_832);
nor U3123 (N_3123,In_285,In_1908);
and U3124 (N_3124,In_1770,In_991);
xnor U3125 (N_3125,In_807,In_478);
or U3126 (N_3126,In_1359,In_1063);
and U3127 (N_3127,In_415,In_1813);
and U3128 (N_3128,In_1431,In_1633);
and U3129 (N_3129,In_432,In_1003);
nor U3130 (N_3130,In_1117,In_1401);
and U3131 (N_3131,In_988,In_1944);
and U3132 (N_3132,In_1876,In_1637);
nor U3133 (N_3133,In_381,In_268);
nor U3134 (N_3134,In_1314,In_509);
and U3135 (N_3135,In_1658,In_318);
and U3136 (N_3136,In_60,In_506);
or U3137 (N_3137,In_678,In_646);
or U3138 (N_3138,In_1750,In_483);
xor U3139 (N_3139,In_1372,In_54);
nand U3140 (N_3140,In_402,In_1880);
or U3141 (N_3141,In_1300,In_77);
and U3142 (N_3142,In_783,In_1315);
or U3143 (N_3143,In_440,In_924);
and U3144 (N_3144,In_1573,In_233);
nand U3145 (N_3145,In_1714,In_1676);
and U3146 (N_3146,In_581,In_1018);
or U3147 (N_3147,In_1484,In_877);
xnor U3148 (N_3148,In_1768,In_770);
nor U3149 (N_3149,In_355,In_200);
nand U3150 (N_3150,In_214,In_1489);
xor U3151 (N_3151,In_588,In_1353);
or U3152 (N_3152,In_1934,In_755);
nand U3153 (N_3153,In_1163,In_118);
xnor U3154 (N_3154,In_260,In_763);
nor U3155 (N_3155,In_890,In_1352);
nand U3156 (N_3156,In_509,In_1143);
xor U3157 (N_3157,In_1146,In_523);
xor U3158 (N_3158,In_508,In_1074);
and U3159 (N_3159,In_366,In_1498);
xor U3160 (N_3160,In_1002,In_1055);
and U3161 (N_3161,In_495,In_186);
xor U3162 (N_3162,In_1499,In_1342);
xor U3163 (N_3163,In_1211,In_890);
nor U3164 (N_3164,In_1709,In_513);
and U3165 (N_3165,In_1734,In_1912);
nand U3166 (N_3166,In_779,In_1173);
and U3167 (N_3167,In_1977,In_1631);
nand U3168 (N_3168,In_1637,In_1134);
or U3169 (N_3169,In_183,In_1885);
and U3170 (N_3170,In_1931,In_1359);
and U3171 (N_3171,In_119,In_426);
or U3172 (N_3172,In_1734,In_199);
or U3173 (N_3173,In_1615,In_1410);
or U3174 (N_3174,In_1153,In_1149);
nor U3175 (N_3175,In_847,In_608);
xnor U3176 (N_3176,In_1313,In_647);
nor U3177 (N_3177,In_920,In_1151);
xnor U3178 (N_3178,In_1023,In_1862);
nor U3179 (N_3179,In_1700,In_451);
or U3180 (N_3180,In_928,In_1136);
and U3181 (N_3181,In_1997,In_1188);
xor U3182 (N_3182,In_664,In_290);
and U3183 (N_3183,In_956,In_239);
and U3184 (N_3184,In_64,In_1361);
nor U3185 (N_3185,In_355,In_1434);
nor U3186 (N_3186,In_27,In_1179);
xnor U3187 (N_3187,In_1752,In_1811);
or U3188 (N_3188,In_970,In_1632);
xnor U3189 (N_3189,In_1769,In_1301);
xnor U3190 (N_3190,In_957,In_1397);
nand U3191 (N_3191,In_976,In_1327);
and U3192 (N_3192,In_1855,In_317);
xnor U3193 (N_3193,In_637,In_1400);
nand U3194 (N_3194,In_247,In_112);
nor U3195 (N_3195,In_1468,In_1565);
and U3196 (N_3196,In_1795,In_1404);
or U3197 (N_3197,In_1416,In_1102);
xnor U3198 (N_3198,In_1263,In_1989);
xor U3199 (N_3199,In_152,In_148);
xnor U3200 (N_3200,In_127,In_1482);
nor U3201 (N_3201,In_1346,In_717);
and U3202 (N_3202,In_1939,In_1893);
and U3203 (N_3203,In_255,In_516);
and U3204 (N_3204,In_790,In_1849);
xor U3205 (N_3205,In_1986,In_1333);
and U3206 (N_3206,In_395,In_1144);
nor U3207 (N_3207,In_408,In_1562);
xnor U3208 (N_3208,In_1497,In_1404);
nand U3209 (N_3209,In_1670,In_607);
nor U3210 (N_3210,In_1106,In_196);
and U3211 (N_3211,In_230,In_942);
nor U3212 (N_3212,In_468,In_1350);
xor U3213 (N_3213,In_736,In_1320);
nand U3214 (N_3214,In_337,In_1164);
or U3215 (N_3215,In_1437,In_726);
and U3216 (N_3216,In_1692,In_1653);
xor U3217 (N_3217,In_656,In_513);
or U3218 (N_3218,In_774,In_951);
and U3219 (N_3219,In_1379,In_899);
or U3220 (N_3220,In_1641,In_804);
nor U3221 (N_3221,In_1808,In_1716);
nor U3222 (N_3222,In_1460,In_1800);
and U3223 (N_3223,In_570,In_274);
or U3224 (N_3224,In_1208,In_1954);
nand U3225 (N_3225,In_459,In_391);
nand U3226 (N_3226,In_544,In_405);
nand U3227 (N_3227,In_1685,In_323);
nand U3228 (N_3228,In_1618,In_272);
or U3229 (N_3229,In_1822,In_1452);
and U3230 (N_3230,In_777,In_978);
or U3231 (N_3231,In_1357,In_925);
or U3232 (N_3232,In_703,In_1025);
nor U3233 (N_3233,In_1693,In_247);
and U3234 (N_3234,In_1388,In_1559);
and U3235 (N_3235,In_1961,In_1782);
or U3236 (N_3236,In_1118,In_1668);
nand U3237 (N_3237,In_1595,In_1900);
xor U3238 (N_3238,In_528,In_1410);
nor U3239 (N_3239,In_816,In_958);
xnor U3240 (N_3240,In_1155,In_1148);
nor U3241 (N_3241,In_1308,In_256);
nor U3242 (N_3242,In_1399,In_41);
nor U3243 (N_3243,In_1236,In_1391);
or U3244 (N_3244,In_1743,In_1672);
nor U3245 (N_3245,In_250,In_449);
xnor U3246 (N_3246,In_548,In_525);
nor U3247 (N_3247,In_56,In_1788);
and U3248 (N_3248,In_983,In_1606);
nor U3249 (N_3249,In_861,In_1439);
and U3250 (N_3250,In_1783,In_1178);
xnor U3251 (N_3251,In_392,In_213);
nor U3252 (N_3252,In_1004,In_1386);
and U3253 (N_3253,In_580,In_442);
xor U3254 (N_3254,In_1952,In_738);
or U3255 (N_3255,In_1328,In_898);
and U3256 (N_3256,In_1187,In_1000);
nand U3257 (N_3257,In_1019,In_476);
nor U3258 (N_3258,In_1308,In_1450);
xor U3259 (N_3259,In_113,In_1904);
and U3260 (N_3260,In_1925,In_516);
nand U3261 (N_3261,In_460,In_1578);
nor U3262 (N_3262,In_1600,In_30);
or U3263 (N_3263,In_1774,In_1878);
xnor U3264 (N_3264,In_161,In_289);
nor U3265 (N_3265,In_692,In_121);
nand U3266 (N_3266,In_1020,In_899);
nor U3267 (N_3267,In_595,In_609);
and U3268 (N_3268,In_1219,In_1095);
nand U3269 (N_3269,In_934,In_1053);
and U3270 (N_3270,In_1367,In_1057);
nand U3271 (N_3271,In_439,In_378);
and U3272 (N_3272,In_1587,In_1677);
or U3273 (N_3273,In_1270,In_1508);
nand U3274 (N_3274,In_1432,In_1860);
xnor U3275 (N_3275,In_1533,In_1277);
nor U3276 (N_3276,In_1569,In_1729);
nand U3277 (N_3277,In_597,In_527);
xor U3278 (N_3278,In_1052,In_1704);
xnor U3279 (N_3279,In_984,In_775);
nand U3280 (N_3280,In_1998,In_1204);
xnor U3281 (N_3281,In_1223,In_478);
and U3282 (N_3282,In_872,In_1451);
nor U3283 (N_3283,In_682,In_807);
or U3284 (N_3284,In_970,In_1972);
or U3285 (N_3285,In_497,In_220);
xor U3286 (N_3286,In_978,In_1672);
xnor U3287 (N_3287,In_377,In_1);
nor U3288 (N_3288,In_1985,In_994);
or U3289 (N_3289,In_298,In_1709);
xnor U3290 (N_3290,In_526,In_797);
nor U3291 (N_3291,In_1958,In_638);
and U3292 (N_3292,In_880,In_1708);
xor U3293 (N_3293,In_1463,In_692);
xor U3294 (N_3294,In_749,In_1164);
nor U3295 (N_3295,In_603,In_449);
nor U3296 (N_3296,In_1262,In_1188);
or U3297 (N_3297,In_19,In_1103);
or U3298 (N_3298,In_1604,In_680);
nand U3299 (N_3299,In_1854,In_325);
nor U3300 (N_3300,In_1895,In_440);
nor U3301 (N_3301,In_584,In_1520);
or U3302 (N_3302,In_1903,In_208);
xor U3303 (N_3303,In_527,In_1930);
xnor U3304 (N_3304,In_1994,In_353);
xor U3305 (N_3305,In_648,In_631);
xnor U3306 (N_3306,In_1691,In_1622);
nand U3307 (N_3307,In_695,In_715);
nor U3308 (N_3308,In_1354,In_1343);
or U3309 (N_3309,In_224,In_808);
or U3310 (N_3310,In_611,In_438);
or U3311 (N_3311,In_1728,In_1058);
nand U3312 (N_3312,In_524,In_1315);
nand U3313 (N_3313,In_328,In_972);
or U3314 (N_3314,In_1998,In_340);
or U3315 (N_3315,In_1567,In_925);
or U3316 (N_3316,In_1063,In_628);
nand U3317 (N_3317,In_876,In_1947);
nand U3318 (N_3318,In_1843,In_193);
and U3319 (N_3319,In_271,In_343);
xnor U3320 (N_3320,In_1951,In_26);
nand U3321 (N_3321,In_1988,In_1628);
and U3322 (N_3322,In_991,In_288);
nand U3323 (N_3323,In_1252,In_77);
or U3324 (N_3324,In_469,In_1568);
and U3325 (N_3325,In_1923,In_588);
nor U3326 (N_3326,In_458,In_337);
or U3327 (N_3327,In_254,In_639);
nand U3328 (N_3328,In_179,In_1751);
or U3329 (N_3329,In_673,In_1842);
or U3330 (N_3330,In_1238,In_612);
nor U3331 (N_3331,In_1322,In_976);
nor U3332 (N_3332,In_461,In_1279);
nand U3333 (N_3333,In_1954,In_1059);
nor U3334 (N_3334,In_1497,In_1157);
or U3335 (N_3335,In_1547,In_857);
xor U3336 (N_3336,In_1006,In_1744);
nand U3337 (N_3337,In_625,In_840);
or U3338 (N_3338,In_627,In_998);
nor U3339 (N_3339,In_882,In_802);
nand U3340 (N_3340,In_795,In_1803);
or U3341 (N_3341,In_840,In_990);
nor U3342 (N_3342,In_1357,In_150);
or U3343 (N_3343,In_332,In_1819);
nand U3344 (N_3344,In_1321,In_1246);
nor U3345 (N_3345,In_1604,In_1009);
nor U3346 (N_3346,In_1442,In_800);
and U3347 (N_3347,In_1485,In_174);
nor U3348 (N_3348,In_315,In_478);
or U3349 (N_3349,In_1895,In_1888);
xor U3350 (N_3350,In_1588,In_19);
and U3351 (N_3351,In_80,In_1431);
or U3352 (N_3352,In_403,In_149);
nor U3353 (N_3353,In_835,In_395);
nor U3354 (N_3354,In_1214,In_1979);
nor U3355 (N_3355,In_196,In_1304);
xor U3356 (N_3356,In_1954,In_1345);
nand U3357 (N_3357,In_1273,In_1085);
or U3358 (N_3358,In_1970,In_516);
nor U3359 (N_3359,In_927,In_943);
nor U3360 (N_3360,In_1139,In_1544);
nand U3361 (N_3361,In_653,In_1639);
and U3362 (N_3362,In_1996,In_373);
and U3363 (N_3363,In_1074,In_301);
xnor U3364 (N_3364,In_233,In_1088);
nor U3365 (N_3365,In_458,In_520);
nor U3366 (N_3366,In_1443,In_273);
and U3367 (N_3367,In_811,In_753);
nor U3368 (N_3368,In_1598,In_1755);
or U3369 (N_3369,In_1332,In_1551);
and U3370 (N_3370,In_699,In_1447);
nand U3371 (N_3371,In_1748,In_620);
nand U3372 (N_3372,In_364,In_937);
xor U3373 (N_3373,In_1736,In_1673);
xnor U3374 (N_3374,In_1237,In_1268);
or U3375 (N_3375,In_1599,In_1238);
and U3376 (N_3376,In_84,In_369);
nand U3377 (N_3377,In_1890,In_1153);
nand U3378 (N_3378,In_678,In_1671);
nor U3379 (N_3379,In_1075,In_1499);
and U3380 (N_3380,In_454,In_698);
or U3381 (N_3381,In_858,In_886);
or U3382 (N_3382,In_1196,In_197);
or U3383 (N_3383,In_886,In_181);
xor U3384 (N_3384,In_1778,In_1696);
and U3385 (N_3385,In_847,In_1614);
xor U3386 (N_3386,In_1476,In_342);
xor U3387 (N_3387,In_1299,In_1850);
xor U3388 (N_3388,In_228,In_846);
xnor U3389 (N_3389,In_249,In_1425);
and U3390 (N_3390,In_339,In_1752);
xor U3391 (N_3391,In_1457,In_1609);
or U3392 (N_3392,In_157,In_1476);
xnor U3393 (N_3393,In_1411,In_1986);
or U3394 (N_3394,In_209,In_511);
nor U3395 (N_3395,In_231,In_819);
or U3396 (N_3396,In_746,In_109);
and U3397 (N_3397,In_1395,In_1119);
xnor U3398 (N_3398,In_124,In_840);
or U3399 (N_3399,In_457,In_467);
and U3400 (N_3400,In_633,In_1709);
and U3401 (N_3401,In_147,In_1909);
xor U3402 (N_3402,In_270,In_1999);
or U3403 (N_3403,In_1676,In_1253);
nor U3404 (N_3404,In_1113,In_770);
nor U3405 (N_3405,In_1363,In_281);
nor U3406 (N_3406,In_654,In_845);
nor U3407 (N_3407,In_1528,In_1322);
nand U3408 (N_3408,In_349,In_1829);
nor U3409 (N_3409,In_1022,In_1305);
xor U3410 (N_3410,In_506,In_1739);
nand U3411 (N_3411,In_330,In_1135);
nor U3412 (N_3412,In_1496,In_496);
and U3413 (N_3413,In_1970,In_700);
xor U3414 (N_3414,In_206,In_938);
or U3415 (N_3415,In_1222,In_1394);
or U3416 (N_3416,In_1158,In_814);
and U3417 (N_3417,In_956,In_1647);
or U3418 (N_3418,In_1228,In_1629);
and U3419 (N_3419,In_526,In_670);
and U3420 (N_3420,In_1005,In_567);
xnor U3421 (N_3421,In_575,In_1556);
or U3422 (N_3422,In_1899,In_1264);
xor U3423 (N_3423,In_1883,In_1522);
and U3424 (N_3424,In_429,In_1404);
nor U3425 (N_3425,In_1502,In_1237);
and U3426 (N_3426,In_1655,In_269);
nor U3427 (N_3427,In_89,In_1337);
or U3428 (N_3428,In_702,In_179);
nand U3429 (N_3429,In_57,In_771);
nor U3430 (N_3430,In_1792,In_1857);
or U3431 (N_3431,In_688,In_549);
and U3432 (N_3432,In_187,In_1778);
nor U3433 (N_3433,In_1126,In_1652);
xnor U3434 (N_3434,In_1793,In_1443);
xnor U3435 (N_3435,In_946,In_432);
or U3436 (N_3436,In_1216,In_1377);
and U3437 (N_3437,In_539,In_205);
or U3438 (N_3438,In_1209,In_83);
and U3439 (N_3439,In_1458,In_1128);
xnor U3440 (N_3440,In_752,In_535);
or U3441 (N_3441,In_1616,In_632);
nand U3442 (N_3442,In_267,In_757);
or U3443 (N_3443,In_1677,In_1277);
nand U3444 (N_3444,In_102,In_1793);
nor U3445 (N_3445,In_1963,In_103);
or U3446 (N_3446,In_1769,In_1927);
nor U3447 (N_3447,In_1639,In_1757);
and U3448 (N_3448,In_1716,In_69);
and U3449 (N_3449,In_1974,In_511);
xor U3450 (N_3450,In_1105,In_1812);
xor U3451 (N_3451,In_946,In_1175);
or U3452 (N_3452,In_1460,In_294);
xor U3453 (N_3453,In_1952,In_1671);
nand U3454 (N_3454,In_45,In_1513);
and U3455 (N_3455,In_1259,In_1740);
or U3456 (N_3456,In_794,In_655);
nand U3457 (N_3457,In_1702,In_481);
nand U3458 (N_3458,In_368,In_872);
nand U3459 (N_3459,In_529,In_563);
or U3460 (N_3460,In_878,In_990);
xnor U3461 (N_3461,In_1068,In_800);
xor U3462 (N_3462,In_184,In_1890);
nand U3463 (N_3463,In_1298,In_895);
or U3464 (N_3464,In_1975,In_252);
or U3465 (N_3465,In_1333,In_907);
nand U3466 (N_3466,In_196,In_1600);
or U3467 (N_3467,In_1648,In_599);
and U3468 (N_3468,In_891,In_950);
or U3469 (N_3469,In_689,In_299);
nor U3470 (N_3470,In_1437,In_351);
or U3471 (N_3471,In_1104,In_1768);
and U3472 (N_3472,In_454,In_1784);
nor U3473 (N_3473,In_1373,In_1634);
and U3474 (N_3474,In_1338,In_1490);
or U3475 (N_3475,In_1262,In_1019);
or U3476 (N_3476,In_323,In_1281);
and U3477 (N_3477,In_140,In_635);
nand U3478 (N_3478,In_1583,In_1158);
nor U3479 (N_3479,In_1679,In_1090);
xor U3480 (N_3480,In_1395,In_1517);
and U3481 (N_3481,In_1934,In_1405);
nor U3482 (N_3482,In_1786,In_1216);
nor U3483 (N_3483,In_947,In_1998);
nor U3484 (N_3484,In_661,In_563);
and U3485 (N_3485,In_643,In_1154);
and U3486 (N_3486,In_1403,In_1579);
or U3487 (N_3487,In_546,In_235);
xnor U3488 (N_3488,In_512,In_1208);
and U3489 (N_3489,In_272,In_1659);
nand U3490 (N_3490,In_504,In_437);
nor U3491 (N_3491,In_1822,In_1911);
nand U3492 (N_3492,In_290,In_1446);
and U3493 (N_3493,In_916,In_975);
and U3494 (N_3494,In_767,In_1117);
nor U3495 (N_3495,In_1515,In_664);
and U3496 (N_3496,In_1900,In_1350);
xor U3497 (N_3497,In_1114,In_202);
or U3498 (N_3498,In_1035,In_1915);
xor U3499 (N_3499,In_1920,In_828);
nand U3500 (N_3500,In_1602,In_1168);
nand U3501 (N_3501,In_1495,In_1886);
xnor U3502 (N_3502,In_1447,In_786);
nor U3503 (N_3503,In_386,In_405);
xnor U3504 (N_3504,In_879,In_1391);
nand U3505 (N_3505,In_364,In_1620);
nor U3506 (N_3506,In_1593,In_1709);
and U3507 (N_3507,In_1357,In_1294);
and U3508 (N_3508,In_52,In_1365);
xnor U3509 (N_3509,In_919,In_1932);
nand U3510 (N_3510,In_1835,In_1022);
xnor U3511 (N_3511,In_951,In_1417);
or U3512 (N_3512,In_127,In_1102);
and U3513 (N_3513,In_352,In_818);
xnor U3514 (N_3514,In_1032,In_877);
and U3515 (N_3515,In_1010,In_1344);
and U3516 (N_3516,In_1887,In_403);
nand U3517 (N_3517,In_1942,In_1766);
and U3518 (N_3518,In_1877,In_1756);
xor U3519 (N_3519,In_1080,In_1002);
or U3520 (N_3520,In_1752,In_1467);
xor U3521 (N_3521,In_349,In_453);
nand U3522 (N_3522,In_468,In_616);
nand U3523 (N_3523,In_1877,In_1043);
nor U3524 (N_3524,In_577,In_223);
or U3525 (N_3525,In_1644,In_1580);
nand U3526 (N_3526,In_1670,In_31);
nand U3527 (N_3527,In_1042,In_1337);
nand U3528 (N_3528,In_1591,In_727);
nor U3529 (N_3529,In_1494,In_1034);
xnor U3530 (N_3530,In_1043,In_159);
nor U3531 (N_3531,In_529,In_1107);
nor U3532 (N_3532,In_1350,In_1272);
and U3533 (N_3533,In_382,In_1052);
xor U3534 (N_3534,In_1125,In_339);
nand U3535 (N_3535,In_382,In_1158);
xnor U3536 (N_3536,In_44,In_210);
and U3537 (N_3537,In_727,In_1355);
and U3538 (N_3538,In_564,In_1598);
nand U3539 (N_3539,In_1185,In_619);
xnor U3540 (N_3540,In_1110,In_337);
xor U3541 (N_3541,In_65,In_405);
and U3542 (N_3542,In_714,In_1786);
xnor U3543 (N_3543,In_1715,In_819);
xor U3544 (N_3544,In_1905,In_1319);
xnor U3545 (N_3545,In_1275,In_738);
nor U3546 (N_3546,In_1173,In_75);
or U3547 (N_3547,In_1934,In_344);
nor U3548 (N_3548,In_343,In_183);
xnor U3549 (N_3549,In_332,In_1411);
nor U3550 (N_3550,In_1944,In_571);
and U3551 (N_3551,In_429,In_1764);
nand U3552 (N_3552,In_101,In_1435);
nor U3553 (N_3553,In_373,In_1746);
nor U3554 (N_3554,In_1353,In_1736);
nor U3555 (N_3555,In_1393,In_519);
and U3556 (N_3556,In_1983,In_1713);
or U3557 (N_3557,In_1190,In_1580);
nor U3558 (N_3558,In_549,In_1827);
or U3559 (N_3559,In_1128,In_45);
or U3560 (N_3560,In_407,In_1356);
nand U3561 (N_3561,In_1617,In_1068);
nand U3562 (N_3562,In_1649,In_1391);
xor U3563 (N_3563,In_920,In_1765);
nand U3564 (N_3564,In_1868,In_416);
and U3565 (N_3565,In_928,In_116);
or U3566 (N_3566,In_1852,In_218);
or U3567 (N_3567,In_519,In_1359);
or U3568 (N_3568,In_1835,In_1268);
xor U3569 (N_3569,In_1495,In_1873);
and U3570 (N_3570,In_836,In_773);
or U3571 (N_3571,In_1857,In_1880);
or U3572 (N_3572,In_348,In_1325);
and U3573 (N_3573,In_927,In_632);
nand U3574 (N_3574,In_1315,In_555);
and U3575 (N_3575,In_1137,In_494);
nor U3576 (N_3576,In_1791,In_394);
and U3577 (N_3577,In_1328,In_1733);
nor U3578 (N_3578,In_566,In_1838);
nor U3579 (N_3579,In_70,In_1782);
xnor U3580 (N_3580,In_30,In_626);
and U3581 (N_3581,In_1391,In_1055);
and U3582 (N_3582,In_364,In_1298);
and U3583 (N_3583,In_978,In_656);
nand U3584 (N_3584,In_1074,In_938);
nand U3585 (N_3585,In_993,In_527);
and U3586 (N_3586,In_642,In_864);
and U3587 (N_3587,In_441,In_1448);
and U3588 (N_3588,In_370,In_1744);
or U3589 (N_3589,In_1384,In_1869);
and U3590 (N_3590,In_976,In_1794);
or U3591 (N_3591,In_1644,In_1010);
nor U3592 (N_3592,In_1452,In_895);
and U3593 (N_3593,In_297,In_255);
or U3594 (N_3594,In_849,In_543);
and U3595 (N_3595,In_1951,In_330);
and U3596 (N_3596,In_1020,In_723);
and U3597 (N_3597,In_1055,In_577);
nor U3598 (N_3598,In_63,In_1480);
and U3599 (N_3599,In_1840,In_415);
or U3600 (N_3600,In_204,In_881);
and U3601 (N_3601,In_422,In_78);
or U3602 (N_3602,In_912,In_899);
nand U3603 (N_3603,In_1387,In_1681);
nor U3604 (N_3604,In_27,In_401);
or U3605 (N_3605,In_989,In_947);
or U3606 (N_3606,In_1850,In_1218);
xor U3607 (N_3607,In_1730,In_1491);
and U3608 (N_3608,In_228,In_1733);
and U3609 (N_3609,In_1415,In_1196);
xnor U3610 (N_3610,In_926,In_236);
or U3611 (N_3611,In_962,In_1143);
and U3612 (N_3612,In_1441,In_1854);
and U3613 (N_3613,In_471,In_838);
or U3614 (N_3614,In_1607,In_942);
xnor U3615 (N_3615,In_228,In_185);
and U3616 (N_3616,In_1411,In_1930);
and U3617 (N_3617,In_1155,In_629);
nand U3618 (N_3618,In_1791,In_1587);
nor U3619 (N_3619,In_1569,In_313);
nor U3620 (N_3620,In_709,In_1851);
nand U3621 (N_3621,In_489,In_210);
and U3622 (N_3622,In_900,In_1714);
nand U3623 (N_3623,In_1306,In_67);
nand U3624 (N_3624,In_1024,In_1444);
nand U3625 (N_3625,In_693,In_996);
xor U3626 (N_3626,In_204,In_1770);
xnor U3627 (N_3627,In_649,In_796);
and U3628 (N_3628,In_816,In_1343);
or U3629 (N_3629,In_1183,In_1918);
nand U3630 (N_3630,In_998,In_1113);
or U3631 (N_3631,In_496,In_1965);
xnor U3632 (N_3632,In_663,In_573);
xnor U3633 (N_3633,In_405,In_275);
or U3634 (N_3634,In_467,In_1238);
nor U3635 (N_3635,In_444,In_1970);
and U3636 (N_3636,In_1784,In_1640);
nor U3637 (N_3637,In_464,In_1228);
or U3638 (N_3638,In_206,In_1971);
and U3639 (N_3639,In_529,In_928);
nor U3640 (N_3640,In_1669,In_993);
nor U3641 (N_3641,In_71,In_329);
or U3642 (N_3642,In_138,In_738);
nand U3643 (N_3643,In_1723,In_1599);
xor U3644 (N_3644,In_607,In_1880);
and U3645 (N_3645,In_791,In_1386);
xor U3646 (N_3646,In_312,In_909);
nand U3647 (N_3647,In_868,In_1183);
xnor U3648 (N_3648,In_1056,In_190);
xor U3649 (N_3649,In_492,In_1418);
or U3650 (N_3650,In_1232,In_1306);
xnor U3651 (N_3651,In_695,In_306);
xor U3652 (N_3652,In_917,In_325);
and U3653 (N_3653,In_951,In_1683);
xnor U3654 (N_3654,In_1576,In_973);
nor U3655 (N_3655,In_988,In_1682);
nor U3656 (N_3656,In_216,In_793);
xor U3657 (N_3657,In_962,In_945);
nor U3658 (N_3658,In_599,In_360);
xnor U3659 (N_3659,In_564,In_680);
and U3660 (N_3660,In_68,In_1478);
nor U3661 (N_3661,In_1479,In_1075);
xor U3662 (N_3662,In_1927,In_914);
nand U3663 (N_3663,In_110,In_474);
xnor U3664 (N_3664,In_1852,In_1991);
nor U3665 (N_3665,In_250,In_274);
nor U3666 (N_3666,In_213,In_1407);
nand U3667 (N_3667,In_779,In_1742);
and U3668 (N_3668,In_741,In_894);
nand U3669 (N_3669,In_783,In_1125);
xnor U3670 (N_3670,In_231,In_895);
and U3671 (N_3671,In_28,In_1433);
xor U3672 (N_3672,In_1798,In_923);
xnor U3673 (N_3673,In_1771,In_1714);
or U3674 (N_3674,In_268,In_396);
nand U3675 (N_3675,In_297,In_1054);
and U3676 (N_3676,In_229,In_367);
xnor U3677 (N_3677,In_1257,In_917);
nand U3678 (N_3678,In_794,In_813);
xnor U3679 (N_3679,In_286,In_1997);
xor U3680 (N_3680,In_1746,In_1098);
nor U3681 (N_3681,In_1742,In_1724);
xor U3682 (N_3682,In_1440,In_695);
or U3683 (N_3683,In_1840,In_417);
and U3684 (N_3684,In_1094,In_1476);
and U3685 (N_3685,In_1508,In_249);
xor U3686 (N_3686,In_666,In_1485);
nor U3687 (N_3687,In_1773,In_335);
and U3688 (N_3688,In_1747,In_1305);
xnor U3689 (N_3689,In_1470,In_658);
nor U3690 (N_3690,In_758,In_1338);
xnor U3691 (N_3691,In_1006,In_1652);
nor U3692 (N_3692,In_1911,In_1539);
nor U3693 (N_3693,In_677,In_1977);
nand U3694 (N_3694,In_1947,In_1146);
and U3695 (N_3695,In_195,In_1999);
and U3696 (N_3696,In_1144,In_783);
nand U3697 (N_3697,In_1129,In_1112);
nor U3698 (N_3698,In_1322,In_529);
and U3699 (N_3699,In_1095,In_1113);
nor U3700 (N_3700,In_183,In_887);
or U3701 (N_3701,In_1152,In_1346);
and U3702 (N_3702,In_935,In_216);
nand U3703 (N_3703,In_782,In_1292);
and U3704 (N_3704,In_1382,In_1373);
nand U3705 (N_3705,In_756,In_172);
or U3706 (N_3706,In_546,In_1033);
nand U3707 (N_3707,In_29,In_1111);
xor U3708 (N_3708,In_1860,In_1138);
xor U3709 (N_3709,In_1689,In_1458);
xnor U3710 (N_3710,In_1202,In_1484);
nor U3711 (N_3711,In_262,In_239);
or U3712 (N_3712,In_297,In_21);
xor U3713 (N_3713,In_194,In_1039);
nor U3714 (N_3714,In_938,In_1213);
or U3715 (N_3715,In_370,In_1885);
or U3716 (N_3716,In_705,In_1940);
nor U3717 (N_3717,In_1291,In_1331);
nand U3718 (N_3718,In_1298,In_133);
nor U3719 (N_3719,In_1258,In_494);
or U3720 (N_3720,In_660,In_251);
nand U3721 (N_3721,In_159,In_128);
nor U3722 (N_3722,In_1407,In_1980);
and U3723 (N_3723,In_557,In_1869);
or U3724 (N_3724,In_1553,In_895);
nand U3725 (N_3725,In_145,In_1869);
nor U3726 (N_3726,In_1170,In_947);
nand U3727 (N_3727,In_1288,In_262);
xnor U3728 (N_3728,In_979,In_1944);
nor U3729 (N_3729,In_316,In_1458);
xnor U3730 (N_3730,In_32,In_704);
xnor U3731 (N_3731,In_1266,In_1226);
or U3732 (N_3732,In_161,In_439);
nand U3733 (N_3733,In_544,In_768);
xor U3734 (N_3734,In_1553,In_1635);
nand U3735 (N_3735,In_1674,In_1308);
or U3736 (N_3736,In_29,In_99);
nand U3737 (N_3737,In_1468,In_260);
xnor U3738 (N_3738,In_1051,In_1502);
xor U3739 (N_3739,In_560,In_826);
or U3740 (N_3740,In_1584,In_948);
xnor U3741 (N_3741,In_557,In_656);
nand U3742 (N_3742,In_1779,In_1700);
nor U3743 (N_3743,In_229,In_21);
nand U3744 (N_3744,In_825,In_1634);
or U3745 (N_3745,In_1969,In_914);
nand U3746 (N_3746,In_1285,In_1157);
and U3747 (N_3747,In_1937,In_629);
or U3748 (N_3748,In_235,In_33);
nor U3749 (N_3749,In_991,In_1800);
xnor U3750 (N_3750,In_1882,In_992);
nor U3751 (N_3751,In_1914,In_120);
and U3752 (N_3752,In_533,In_433);
nor U3753 (N_3753,In_269,In_1627);
nand U3754 (N_3754,In_1337,In_1390);
xor U3755 (N_3755,In_643,In_372);
and U3756 (N_3756,In_1200,In_771);
and U3757 (N_3757,In_341,In_1417);
xor U3758 (N_3758,In_1840,In_1833);
nor U3759 (N_3759,In_1861,In_761);
and U3760 (N_3760,In_1975,In_1398);
nand U3761 (N_3761,In_1713,In_1309);
xnor U3762 (N_3762,In_1391,In_715);
nand U3763 (N_3763,In_569,In_400);
and U3764 (N_3764,In_899,In_1743);
or U3765 (N_3765,In_1670,In_1491);
nor U3766 (N_3766,In_134,In_49);
nor U3767 (N_3767,In_64,In_124);
nor U3768 (N_3768,In_859,In_1473);
nor U3769 (N_3769,In_940,In_1436);
and U3770 (N_3770,In_1627,In_1662);
xor U3771 (N_3771,In_459,In_340);
or U3772 (N_3772,In_1,In_975);
or U3773 (N_3773,In_216,In_624);
nor U3774 (N_3774,In_327,In_1309);
and U3775 (N_3775,In_871,In_1725);
nand U3776 (N_3776,In_646,In_1779);
and U3777 (N_3777,In_1889,In_1967);
and U3778 (N_3778,In_1896,In_1215);
and U3779 (N_3779,In_1720,In_829);
nor U3780 (N_3780,In_1356,In_1589);
nand U3781 (N_3781,In_186,In_328);
nor U3782 (N_3782,In_1053,In_1782);
and U3783 (N_3783,In_821,In_1627);
and U3784 (N_3784,In_1855,In_353);
and U3785 (N_3785,In_167,In_930);
and U3786 (N_3786,In_293,In_193);
and U3787 (N_3787,In_21,In_73);
nor U3788 (N_3788,In_34,In_803);
or U3789 (N_3789,In_238,In_825);
or U3790 (N_3790,In_1713,In_109);
nand U3791 (N_3791,In_875,In_620);
nor U3792 (N_3792,In_1128,In_2);
nor U3793 (N_3793,In_1589,In_1932);
nor U3794 (N_3794,In_1844,In_1444);
nor U3795 (N_3795,In_376,In_1549);
and U3796 (N_3796,In_133,In_939);
nand U3797 (N_3797,In_1582,In_1587);
and U3798 (N_3798,In_530,In_19);
xnor U3799 (N_3799,In_1389,In_415);
nor U3800 (N_3800,In_1886,In_1919);
nand U3801 (N_3801,In_932,In_1626);
and U3802 (N_3802,In_1967,In_453);
xor U3803 (N_3803,In_1621,In_484);
and U3804 (N_3804,In_1109,In_1591);
nor U3805 (N_3805,In_1886,In_438);
xnor U3806 (N_3806,In_297,In_739);
xnor U3807 (N_3807,In_73,In_1988);
and U3808 (N_3808,In_1181,In_1790);
xor U3809 (N_3809,In_1338,In_891);
nand U3810 (N_3810,In_185,In_1426);
nand U3811 (N_3811,In_448,In_1767);
and U3812 (N_3812,In_1259,In_130);
nand U3813 (N_3813,In_708,In_1496);
nand U3814 (N_3814,In_9,In_1261);
or U3815 (N_3815,In_226,In_1905);
nor U3816 (N_3816,In_1796,In_67);
xnor U3817 (N_3817,In_1765,In_293);
nor U3818 (N_3818,In_703,In_1762);
and U3819 (N_3819,In_1241,In_652);
nand U3820 (N_3820,In_771,In_1143);
nor U3821 (N_3821,In_386,In_789);
nor U3822 (N_3822,In_75,In_1066);
nor U3823 (N_3823,In_911,In_1232);
nor U3824 (N_3824,In_1521,In_277);
nand U3825 (N_3825,In_835,In_456);
or U3826 (N_3826,In_1239,In_1981);
or U3827 (N_3827,In_1486,In_1452);
nor U3828 (N_3828,In_150,In_1993);
xnor U3829 (N_3829,In_295,In_1134);
and U3830 (N_3830,In_1570,In_291);
nor U3831 (N_3831,In_1437,In_1645);
xor U3832 (N_3832,In_1040,In_374);
nor U3833 (N_3833,In_90,In_945);
xnor U3834 (N_3834,In_449,In_870);
nor U3835 (N_3835,In_1503,In_1686);
nand U3836 (N_3836,In_1827,In_199);
and U3837 (N_3837,In_312,In_1415);
nor U3838 (N_3838,In_1781,In_1144);
and U3839 (N_3839,In_1588,In_1521);
nand U3840 (N_3840,In_1775,In_870);
nand U3841 (N_3841,In_768,In_1312);
or U3842 (N_3842,In_1011,In_931);
or U3843 (N_3843,In_510,In_896);
and U3844 (N_3844,In_488,In_502);
and U3845 (N_3845,In_96,In_1274);
or U3846 (N_3846,In_1134,In_583);
or U3847 (N_3847,In_407,In_1592);
nor U3848 (N_3848,In_1495,In_283);
xor U3849 (N_3849,In_1071,In_1348);
nand U3850 (N_3850,In_1698,In_1111);
nor U3851 (N_3851,In_979,In_350);
nand U3852 (N_3852,In_417,In_704);
nand U3853 (N_3853,In_15,In_1865);
and U3854 (N_3854,In_1325,In_447);
xnor U3855 (N_3855,In_481,In_431);
or U3856 (N_3856,In_1767,In_1494);
xnor U3857 (N_3857,In_636,In_1559);
or U3858 (N_3858,In_393,In_1473);
xnor U3859 (N_3859,In_458,In_1179);
and U3860 (N_3860,In_1028,In_1850);
xor U3861 (N_3861,In_1004,In_1725);
and U3862 (N_3862,In_700,In_1615);
nor U3863 (N_3863,In_1097,In_1892);
nand U3864 (N_3864,In_1045,In_1711);
or U3865 (N_3865,In_1833,In_739);
and U3866 (N_3866,In_639,In_1186);
xor U3867 (N_3867,In_824,In_1880);
xor U3868 (N_3868,In_302,In_482);
xor U3869 (N_3869,In_787,In_918);
xor U3870 (N_3870,In_1139,In_1804);
xnor U3871 (N_3871,In_1343,In_1288);
xnor U3872 (N_3872,In_492,In_1048);
nand U3873 (N_3873,In_653,In_738);
xnor U3874 (N_3874,In_1267,In_569);
and U3875 (N_3875,In_449,In_1784);
xnor U3876 (N_3876,In_561,In_11);
xor U3877 (N_3877,In_874,In_594);
nand U3878 (N_3878,In_703,In_592);
or U3879 (N_3879,In_1828,In_546);
and U3880 (N_3880,In_950,In_1718);
and U3881 (N_3881,In_1173,In_237);
nand U3882 (N_3882,In_1678,In_1083);
or U3883 (N_3883,In_824,In_252);
and U3884 (N_3884,In_628,In_113);
nor U3885 (N_3885,In_1254,In_837);
xnor U3886 (N_3886,In_1621,In_153);
nand U3887 (N_3887,In_1021,In_1344);
and U3888 (N_3888,In_1507,In_188);
nand U3889 (N_3889,In_1908,In_1022);
nand U3890 (N_3890,In_854,In_1127);
xor U3891 (N_3891,In_1895,In_658);
and U3892 (N_3892,In_942,In_955);
and U3893 (N_3893,In_1690,In_1037);
and U3894 (N_3894,In_1126,In_95);
or U3895 (N_3895,In_1533,In_711);
xor U3896 (N_3896,In_230,In_1688);
nor U3897 (N_3897,In_311,In_265);
nor U3898 (N_3898,In_1146,In_1852);
nand U3899 (N_3899,In_638,In_446);
xnor U3900 (N_3900,In_585,In_1157);
and U3901 (N_3901,In_692,In_1057);
xor U3902 (N_3902,In_150,In_1116);
or U3903 (N_3903,In_792,In_415);
or U3904 (N_3904,In_1255,In_392);
or U3905 (N_3905,In_1227,In_1281);
nor U3906 (N_3906,In_189,In_1050);
or U3907 (N_3907,In_1012,In_1229);
or U3908 (N_3908,In_1189,In_738);
and U3909 (N_3909,In_251,In_1874);
nand U3910 (N_3910,In_227,In_1489);
xnor U3911 (N_3911,In_1504,In_1819);
nand U3912 (N_3912,In_1321,In_928);
and U3913 (N_3913,In_699,In_1182);
and U3914 (N_3914,In_753,In_916);
nor U3915 (N_3915,In_122,In_942);
or U3916 (N_3916,In_121,In_34);
nor U3917 (N_3917,In_518,In_1103);
nand U3918 (N_3918,In_1386,In_983);
xor U3919 (N_3919,In_408,In_1118);
nand U3920 (N_3920,In_1959,In_1948);
nand U3921 (N_3921,In_1989,In_814);
nor U3922 (N_3922,In_1910,In_1614);
and U3923 (N_3923,In_1895,In_215);
and U3924 (N_3924,In_1206,In_1897);
nor U3925 (N_3925,In_622,In_607);
xnor U3926 (N_3926,In_1720,In_321);
nor U3927 (N_3927,In_1258,In_269);
and U3928 (N_3928,In_1674,In_1121);
or U3929 (N_3929,In_1787,In_147);
nand U3930 (N_3930,In_535,In_518);
xnor U3931 (N_3931,In_558,In_1892);
nand U3932 (N_3932,In_1979,In_853);
xnor U3933 (N_3933,In_1751,In_1902);
or U3934 (N_3934,In_1845,In_844);
nand U3935 (N_3935,In_1585,In_1572);
or U3936 (N_3936,In_1274,In_1665);
nor U3937 (N_3937,In_991,In_267);
or U3938 (N_3938,In_292,In_653);
xor U3939 (N_3939,In_1001,In_1);
nor U3940 (N_3940,In_185,In_291);
xor U3941 (N_3941,In_805,In_940);
nor U3942 (N_3942,In_849,In_1913);
xnor U3943 (N_3943,In_413,In_634);
xnor U3944 (N_3944,In_956,In_1705);
nand U3945 (N_3945,In_1236,In_1560);
and U3946 (N_3946,In_1605,In_402);
nand U3947 (N_3947,In_692,In_687);
nor U3948 (N_3948,In_1806,In_382);
or U3949 (N_3949,In_1714,In_1915);
xor U3950 (N_3950,In_1182,In_978);
nand U3951 (N_3951,In_1046,In_1371);
or U3952 (N_3952,In_1592,In_1338);
nand U3953 (N_3953,In_1009,In_778);
nand U3954 (N_3954,In_1887,In_1444);
and U3955 (N_3955,In_912,In_754);
xor U3956 (N_3956,In_1483,In_1643);
or U3957 (N_3957,In_829,In_1214);
nor U3958 (N_3958,In_1926,In_1245);
nand U3959 (N_3959,In_260,In_477);
or U3960 (N_3960,In_203,In_320);
nor U3961 (N_3961,In_1312,In_703);
or U3962 (N_3962,In_634,In_510);
or U3963 (N_3963,In_1652,In_452);
or U3964 (N_3964,In_579,In_1288);
nor U3965 (N_3965,In_1502,In_246);
and U3966 (N_3966,In_242,In_1350);
xnor U3967 (N_3967,In_1090,In_1285);
nor U3968 (N_3968,In_255,In_1853);
or U3969 (N_3969,In_1476,In_1475);
or U3970 (N_3970,In_130,In_544);
or U3971 (N_3971,In_1694,In_1728);
and U3972 (N_3972,In_1957,In_1710);
or U3973 (N_3973,In_11,In_1081);
or U3974 (N_3974,In_136,In_472);
nor U3975 (N_3975,In_692,In_1784);
and U3976 (N_3976,In_515,In_609);
and U3977 (N_3977,In_192,In_1471);
xor U3978 (N_3978,In_511,In_1920);
nand U3979 (N_3979,In_369,In_1617);
and U3980 (N_3980,In_1026,In_594);
or U3981 (N_3981,In_1831,In_1841);
xor U3982 (N_3982,In_515,In_1450);
nor U3983 (N_3983,In_1425,In_1477);
nor U3984 (N_3984,In_759,In_1989);
nand U3985 (N_3985,In_1046,In_1044);
xor U3986 (N_3986,In_577,In_572);
nor U3987 (N_3987,In_1131,In_364);
or U3988 (N_3988,In_1013,In_1079);
nor U3989 (N_3989,In_992,In_1349);
and U3990 (N_3990,In_316,In_707);
nand U3991 (N_3991,In_489,In_1263);
nor U3992 (N_3992,In_619,In_1903);
xor U3993 (N_3993,In_167,In_733);
and U3994 (N_3994,In_205,In_1312);
xor U3995 (N_3995,In_1212,In_727);
xor U3996 (N_3996,In_826,In_1346);
nand U3997 (N_3997,In_1272,In_1136);
nor U3998 (N_3998,In_1854,In_1342);
nor U3999 (N_3999,In_967,In_1079);
and U4000 (N_4000,N_1072,N_60);
nor U4001 (N_4001,N_1156,N_2560);
nand U4002 (N_4002,N_2482,N_1470);
nand U4003 (N_4003,N_3583,N_163);
nor U4004 (N_4004,N_1360,N_807);
nor U4005 (N_4005,N_3767,N_240);
and U4006 (N_4006,N_663,N_2373);
nor U4007 (N_4007,N_1339,N_2627);
or U4008 (N_4008,N_702,N_186);
or U4009 (N_4009,N_3410,N_2648);
or U4010 (N_4010,N_3632,N_3238);
and U4011 (N_4011,N_2147,N_608);
or U4012 (N_4012,N_3021,N_2315);
nor U4013 (N_4013,N_1755,N_100);
and U4014 (N_4014,N_1050,N_2811);
or U4015 (N_4015,N_2410,N_3352);
and U4016 (N_4016,N_3622,N_2472);
nor U4017 (N_4017,N_2612,N_952);
xor U4018 (N_4018,N_3903,N_937);
and U4019 (N_4019,N_618,N_2586);
xor U4020 (N_4020,N_3557,N_2501);
nand U4021 (N_4021,N_888,N_2747);
nor U4022 (N_4022,N_2975,N_3842);
nor U4023 (N_4023,N_1611,N_2992);
or U4024 (N_4024,N_954,N_2351);
or U4025 (N_4025,N_1956,N_3653);
and U4026 (N_4026,N_1902,N_1461);
xor U4027 (N_4027,N_569,N_1653);
or U4028 (N_4028,N_3506,N_2773);
and U4029 (N_4029,N_1307,N_1509);
or U4030 (N_4030,N_2121,N_2706);
or U4031 (N_4031,N_2398,N_2141);
nand U4032 (N_4032,N_1354,N_2758);
or U4033 (N_4033,N_1092,N_3912);
or U4034 (N_4034,N_2205,N_2190);
and U4035 (N_4035,N_3642,N_2647);
nor U4036 (N_4036,N_238,N_3971);
xnor U4037 (N_4037,N_1585,N_510);
or U4038 (N_4038,N_3727,N_2071);
nor U4039 (N_4039,N_3533,N_3830);
and U4040 (N_4040,N_3709,N_2316);
xnor U4041 (N_4041,N_3977,N_1166);
and U4042 (N_4042,N_103,N_1679);
nor U4043 (N_4043,N_1448,N_3525);
and U4044 (N_4044,N_2726,N_1034);
or U4045 (N_4045,N_1086,N_3423);
and U4046 (N_4046,N_1052,N_158);
nor U4047 (N_4047,N_675,N_3705);
xor U4048 (N_4048,N_1669,N_3334);
and U4049 (N_4049,N_3820,N_3587);
nand U4050 (N_4050,N_2259,N_3065);
and U4051 (N_4051,N_2452,N_381);
nor U4052 (N_4052,N_1382,N_275);
xor U4053 (N_4053,N_3174,N_3079);
and U4054 (N_4054,N_3791,N_97);
and U4055 (N_4055,N_2120,N_1202);
or U4056 (N_4056,N_1950,N_263);
nor U4057 (N_4057,N_19,N_1140);
xor U4058 (N_4058,N_3414,N_3737);
nand U4059 (N_4059,N_1248,N_1649);
nand U4060 (N_4060,N_3845,N_742);
nor U4061 (N_4061,N_3764,N_11);
and U4062 (N_4062,N_2962,N_1845);
nor U4063 (N_4063,N_3985,N_351);
xnor U4064 (N_4064,N_2495,N_1278);
or U4065 (N_4065,N_1466,N_2709);
nor U4066 (N_4066,N_2300,N_3937);
or U4067 (N_4067,N_3678,N_3413);
nor U4068 (N_4068,N_288,N_2078);
nand U4069 (N_4069,N_2053,N_2035);
and U4070 (N_4070,N_3169,N_3800);
xor U4071 (N_4071,N_5,N_2793);
and U4072 (N_4072,N_10,N_162);
and U4073 (N_4073,N_985,N_2052);
or U4074 (N_4074,N_2260,N_1229);
nand U4075 (N_4075,N_2087,N_1502);
nand U4076 (N_4076,N_208,N_141);
nor U4077 (N_4077,N_328,N_3735);
nand U4078 (N_4078,N_339,N_3429);
xor U4079 (N_4079,N_1594,N_3476);
xor U4080 (N_4080,N_611,N_154);
nor U4081 (N_4081,N_2295,N_3383);
xor U4082 (N_4082,N_2320,N_2307);
nand U4083 (N_4083,N_3955,N_1690);
xnor U4084 (N_4084,N_1384,N_2425);
or U4085 (N_4085,N_3904,N_703);
nand U4086 (N_4086,N_684,N_413);
xor U4087 (N_4087,N_2613,N_1519);
nor U4088 (N_4088,N_3640,N_3324);
or U4089 (N_4089,N_2220,N_649);
nor U4090 (N_4090,N_3217,N_2717);
xor U4091 (N_4091,N_2817,N_532);
nand U4092 (N_4092,N_197,N_1582);
nand U4093 (N_4093,N_3014,N_1393);
or U4094 (N_4094,N_3939,N_2572);
nand U4095 (N_4095,N_358,N_229);
and U4096 (N_4096,N_3726,N_1249);
xor U4097 (N_4097,N_2886,N_1077);
nand U4098 (N_4098,N_2231,N_3952);
and U4099 (N_4099,N_610,N_1122);
nand U4100 (N_4100,N_2303,N_2840);
xor U4101 (N_4101,N_1378,N_1213);
and U4102 (N_4102,N_3976,N_3436);
or U4103 (N_4103,N_1473,N_1480);
xnor U4104 (N_4104,N_193,N_55);
nor U4105 (N_4105,N_1988,N_2085);
or U4106 (N_4106,N_2302,N_1503);
nand U4107 (N_4107,N_3629,N_272);
and U4108 (N_4108,N_3284,N_1369);
xnor U4109 (N_4109,N_1621,N_2249);
nor U4110 (N_4110,N_2856,N_2241);
or U4111 (N_4111,N_1557,N_3356);
and U4112 (N_4112,N_3793,N_1697);
nand U4113 (N_4113,N_2099,N_111);
nand U4114 (N_4114,N_735,N_2702);
or U4115 (N_4115,N_1628,N_803);
nand U4116 (N_4116,N_1962,N_2167);
nor U4117 (N_4117,N_753,N_741);
nor U4118 (N_4118,N_1830,N_2601);
nor U4119 (N_4119,N_3080,N_1525);
nor U4120 (N_4120,N_947,N_1179);
xnor U4121 (N_4121,N_3692,N_1313);
and U4122 (N_4122,N_1280,N_3431);
or U4123 (N_4123,N_565,N_1260);
and U4124 (N_4124,N_3005,N_2211);
nor U4125 (N_4125,N_91,N_2779);
xor U4126 (N_4126,N_3,N_1689);
nand U4127 (N_4127,N_1153,N_646);
and U4128 (N_4128,N_3201,N_1042);
xor U4129 (N_4129,N_2748,N_1693);
xor U4130 (N_4130,N_3092,N_2377);
or U4131 (N_4131,N_2872,N_2730);
nand U4132 (N_4132,N_3670,N_586);
xnor U4133 (N_4133,N_1859,N_3087);
nand U4134 (N_4134,N_2182,N_310);
or U4135 (N_4135,N_1985,N_3913);
nand U4136 (N_4136,N_18,N_1625);
and U4137 (N_4137,N_845,N_1612);
or U4138 (N_4138,N_879,N_463);
xnor U4139 (N_4139,N_2384,N_2072);
xnor U4140 (N_4140,N_830,N_1678);
and U4141 (N_4141,N_2937,N_3321);
nor U4142 (N_4142,N_713,N_3567);
nor U4143 (N_4143,N_1265,N_3287);
nor U4144 (N_4144,N_731,N_2809);
nor U4145 (N_4145,N_698,N_2226);
nand U4146 (N_4146,N_2844,N_1294);
or U4147 (N_4147,N_3975,N_299);
nand U4148 (N_4148,N_3105,N_3991);
xor U4149 (N_4149,N_2764,N_1275);
nor U4150 (N_4150,N_3887,N_2196);
nor U4151 (N_4151,N_266,N_1381);
nand U4152 (N_4152,N_3927,N_1102);
nand U4153 (N_4153,N_605,N_552);
xnor U4154 (N_4154,N_2789,N_3712);
and U4155 (N_4155,N_2026,N_655);
and U4156 (N_4156,N_82,N_3848);
and U4157 (N_4157,N_222,N_1814);
or U4158 (N_4158,N_2331,N_250);
nand U4159 (N_4159,N_3051,N_3535);
nand U4160 (N_4160,N_1416,N_933);
nand U4161 (N_4161,N_2381,N_3390);
xnor U4162 (N_4162,N_2993,N_1090);
nor U4163 (N_4163,N_789,N_1259);
and U4164 (N_4164,N_1289,N_1074);
and U4165 (N_4165,N_3035,N_1844);
xnor U4166 (N_4166,N_699,N_1719);
xor U4167 (N_4167,N_1107,N_87);
and U4168 (N_4168,N_750,N_2914);
nor U4169 (N_4169,N_2973,N_3886);
or U4170 (N_4170,N_2057,N_1626);
or U4171 (N_4171,N_3029,N_2503);
xor U4172 (N_4172,N_3716,N_3624);
xor U4173 (N_4173,N_1131,N_466);
or U4174 (N_4174,N_2642,N_1959);
and U4175 (N_4175,N_3209,N_3697);
and U4176 (N_4176,N_2998,N_3953);
nand U4177 (N_4177,N_828,N_2909);
or U4178 (N_4178,N_2589,N_1565);
or U4179 (N_4179,N_1539,N_3561);
and U4180 (N_4180,N_817,N_3440);
and U4181 (N_4181,N_1918,N_3126);
and U4182 (N_4182,N_28,N_2261);
or U4183 (N_4183,N_923,N_1775);
xor U4184 (N_4184,N_2860,N_3833);
and U4185 (N_4185,N_376,N_3290);
xnor U4186 (N_4186,N_1475,N_264);
or U4187 (N_4187,N_1934,N_3569);
nand U4188 (N_4188,N_3187,N_3817);
nor U4189 (N_4189,N_3838,N_1663);
and U4190 (N_4190,N_1896,N_1367);
or U4191 (N_4191,N_2294,N_1891);
or U4192 (N_4192,N_783,N_2752);
or U4193 (N_4193,N_855,N_829);
and U4194 (N_4194,N_3689,N_3402);
or U4195 (N_4195,N_259,N_1766);
nand U4196 (N_4196,N_2610,N_3344);
xor U4197 (N_4197,N_693,N_812);
or U4198 (N_4198,N_2930,N_387);
xnor U4199 (N_4199,N_3407,N_1426);
xnor U4200 (N_4200,N_770,N_1496);
nand U4201 (N_4201,N_2327,N_848);
xor U4202 (N_4202,N_1610,N_2942);
nand U4203 (N_4203,N_1435,N_1136);
xor U4204 (N_4204,N_3925,N_178);
or U4205 (N_4205,N_48,N_945);
nand U4206 (N_4206,N_1269,N_3828);
nor U4207 (N_4207,N_316,N_3122);
nor U4208 (N_4208,N_631,N_3175);
nand U4209 (N_4209,N_2804,N_3313);
nor U4210 (N_4210,N_896,N_1331);
and U4211 (N_4211,N_1930,N_1262);
or U4212 (N_4212,N_1320,N_1075);
xor U4213 (N_4213,N_2558,N_3456);
xor U4214 (N_4214,N_3672,N_276);
or U4215 (N_4215,N_2280,N_479);
or U4216 (N_4216,N_2563,N_1838);
or U4217 (N_4217,N_1698,N_2518);
xor U4218 (N_4218,N_2927,N_2101);
nand U4219 (N_4219,N_2898,N_718);
and U4220 (N_4220,N_2476,N_279);
nor U4221 (N_4221,N_2511,N_2439);
or U4222 (N_4222,N_1364,N_786);
xor U4223 (N_4223,N_497,N_194);
or U4224 (N_4224,N_3522,N_710);
or U4225 (N_4225,N_3552,N_3969);
or U4226 (N_4226,N_2899,N_3545);
or U4227 (N_4227,N_3192,N_1195);
or U4228 (N_4228,N_995,N_2375);
or U4229 (N_4229,N_2150,N_3097);
and U4230 (N_4230,N_3465,N_3031);
or U4231 (N_4231,N_2913,N_2352);
and U4232 (N_4232,N_2311,N_174);
nor U4233 (N_4233,N_1334,N_1807);
xor U4234 (N_4234,N_508,N_634);
and U4235 (N_4235,N_3154,N_1318);
nor U4236 (N_4236,N_2948,N_1846);
nand U4237 (N_4237,N_2434,N_20);
and U4238 (N_4238,N_143,N_984);
or U4239 (N_4239,N_555,N_1065);
xor U4240 (N_4240,N_3933,N_2370);
nor U4241 (N_4241,N_3544,N_3929);
or U4242 (N_4242,N_3426,N_1476);
or U4243 (N_4243,N_2416,N_3781);
nand U4244 (N_4244,N_3164,N_577);
nand U4245 (N_4245,N_2215,N_1728);
and U4246 (N_4246,N_2578,N_116);
nand U4247 (N_4247,N_2812,N_3990);
xor U4248 (N_4248,N_3481,N_3259);
and U4249 (N_4249,N_325,N_2060);
nor U4250 (N_4250,N_57,N_775);
xnor U4251 (N_4251,N_2639,N_1429);
and U4252 (N_4252,N_3064,N_725);
or U4253 (N_4253,N_2005,N_3314);
or U4254 (N_4254,N_1252,N_223);
nand U4255 (N_4255,N_1404,N_1425);
nand U4256 (N_4256,N_1457,N_1613);
xnor U4257 (N_4257,N_2820,N_1040);
and U4258 (N_4258,N_382,N_2049);
xnor U4259 (N_4259,N_2624,N_2509);
nor U4260 (N_4260,N_2798,N_2710);
and U4261 (N_4261,N_758,N_1178);
and U4262 (N_4262,N_1058,N_2712);
or U4263 (N_4263,N_2704,N_1355);
or U4264 (N_4264,N_2194,N_777);
nand U4265 (N_4265,N_1589,N_3478);
and U4266 (N_4266,N_152,N_424);
or U4267 (N_4267,N_2502,N_3158);
or U4268 (N_4268,N_1304,N_588);
or U4269 (N_4269,N_2739,N_3996);
and U4270 (N_4270,N_2172,N_365);
and U4271 (N_4271,N_2939,N_258);
nand U4272 (N_4272,N_3568,N_1823);
and U4273 (N_4273,N_3112,N_2534);
and U4274 (N_4274,N_2688,N_734);
nand U4275 (N_4275,N_253,N_909);
nor U4276 (N_4276,N_1813,N_681);
and U4277 (N_4277,N_3186,N_2659);
xnor U4278 (N_4278,N_3227,N_1633);
nand U4279 (N_4279,N_391,N_3542);
xor U4280 (N_4280,N_1438,N_3754);
xor U4281 (N_4281,N_2359,N_3684);
and U4282 (N_4282,N_760,N_2990);
or U4283 (N_4283,N_3494,N_2137);
nand U4284 (N_4284,N_1054,N_2514);
and U4285 (N_4285,N_3056,N_2091);
nand U4286 (N_4286,N_654,N_1270);
and U4287 (N_4287,N_261,N_1149);
nor U4288 (N_4288,N_502,N_3289);
nor U4289 (N_4289,N_1939,N_1338);
and U4290 (N_4290,N_1321,N_1251);
or U4291 (N_4291,N_335,N_3068);
xor U4292 (N_4292,N_2247,N_948);
or U4293 (N_4293,N_1029,N_3450);
xnor U4294 (N_4294,N_2403,N_2274);
nand U4295 (N_4295,N_3523,N_3381);
xnor U4296 (N_4296,N_2737,N_360);
and U4297 (N_4297,N_2841,N_334);
xnor U4298 (N_4298,N_274,N_2879);
xnor U4299 (N_4299,N_2979,N_314);
nor U4300 (N_4300,N_1279,N_723);
or U4301 (N_4301,N_2611,N_242);
xnor U4302 (N_4302,N_1507,N_2915);
or U4303 (N_4303,N_1699,N_2614);
and U4304 (N_4304,N_2014,N_341);
or U4305 (N_4305,N_2385,N_721);
nand U4306 (N_4306,N_1007,N_2228);
and U4307 (N_4307,N_2458,N_1783);
xnor U4308 (N_4308,N_1449,N_3309);
or U4309 (N_4309,N_3878,N_1508);
and U4310 (N_4310,N_68,N_875);
and U4311 (N_4311,N_99,N_1949);
and U4312 (N_4312,N_2036,N_3173);
nor U4313 (N_4313,N_2781,N_2650);
and U4314 (N_4314,N_3802,N_3272);
and U4315 (N_4315,N_3947,N_2623);
and U4316 (N_4316,N_2594,N_3536);
nor U4317 (N_4317,N_648,N_2634);
and U4318 (N_4318,N_970,N_1973);
and U4319 (N_4319,N_868,N_2869);
xnor U4320 (N_4320,N_2082,N_1704);
xor U4321 (N_4321,N_1944,N_3411);
and U4322 (N_4322,N_1932,N_776);
nand U4323 (N_4323,N_3916,N_2109);
or U4324 (N_4324,N_873,N_3212);
and U4325 (N_4325,N_1277,N_2009);
nor U4326 (N_4326,N_773,N_1484);
xor U4327 (N_4327,N_2891,N_214);
nor U4328 (N_4328,N_1247,N_2209);
xnor U4329 (N_4329,N_3497,N_3255);
nand U4330 (N_4330,N_3214,N_109);
nand U4331 (N_4331,N_269,N_2148);
xor U4332 (N_4332,N_3090,N_1998);
nand U4333 (N_4333,N_3325,N_3063);
and U4334 (N_4334,N_762,N_3531);
nand U4335 (N_4335,N_3503,N_2124);
nor U4336 (N_4336,N_1544,N_963);
nand U4337 (N_4337,N_1601,N_3801);
and U4338 (N_4338,N_920,N_1722);
nand U4339 (N_4339,N_3905,N_2003);
nor U4340 (N_4340,N_877,N_2007);
and U4341 (N_4341,N_988,N_3576);
and U4342 (N_4342,N_1729,N_460);
or U4343 (N_4343,N_1895,N_2483);
nand U4344 (N_4344,N_231,N_3472);
nand U4345 (N_4345,N_632,N_2636);
xor U4346 (N_4346,N_1041,N_3138);
nand U4347 (N_4347,N_2571,N_2606);
xnor U4348 (N_4348,N_487,N_2751);
nor U4349 (N_4349,N_2644,N_1657);
or U4350 (N_4350,N_1917,N_3194);
and U4351 (N_4351,N_1927,N_3308);
nand U4352 (N_4352,N_1422,N_607);
xor U4353 (N_4353,N_622,N_3637);
or U4354 (N_4354,N_1397,N_3824);
xor U4355 (N_4355,N_3039,N_2631);
or U4356 (N_4356,N_2536,N_2976);
and U4357 (N_4357,N_3085,N_1142);
or U4358 (N_4358,N_3807,N_1769);
nor U4359 (N_4359,N_2881,N_305);
nor U4360 (N_4360,N_1417,N_512);
or U4361 (N_4361,N_54,N_1410);
nor U4362 (N_4362,N_980,N_1855);
nand U4363 (N_4363,N_3070,N_3621);
nor U4364 (N_4364,N_45,N_3302);
nand U4365 (N_4365,N_1744,N_3455);
nor U4366 (N_4366,N_2761,N_1455);
or U4367 (N_4367,N_2023,N_2853);
and U4368 (N_4368,N_159,N_2532);
xor U4369 (N_4369,N_129,N_3796);
nor U4370 (N_4370,N_1586,N_1716);
xor U4371 (N_4371,N_1608,N_2964);
nand U4372 (N_4372,N_1680,N_620);
xnor U4373 (N_4373,N_336,N_3384);
nor U4374 (N_4374,N_972,N_3220);
nand U4375 (N_4375,N_480,N_834);
xor U4376 (N_4376,N_1991,N_2662);
xnor U4377 (N_4377,N_541,N_2897);
or U4378 (N_4378,N_2689,N_2197);
and U4379 (N_4379,N_1365,N_551);
nor U4380 (N_4380,N_267,N_2332);
nor U4381 (N_4381,N_120,N_1066);
or U4382 (N_4382,N_3123,N_3140);
and U4383 (N_4383,N_885,N_1151);
or U4384 (N_4384,N_1208,N_3119);
nor U4385 (N_4385,N_1627,N_801);
or U4386 (N_4386,N_239,N_1309);
nor U4387 (N_4387,N_3020,N_2718);
or U4388 (N_4388,N_3677,N_1462);
xnor U4389 (N_4389,N_1647,N_2441);
xor U4390 (N_4390,N_2920,N_233);
xor U4391 (N_4391,N_412,N_1977);
nor U4392 (N_4392,N_384,N_1616);
nor U4393 (N_4393,N_792,N_2873);
and U4394 (N_4394,N_691,N_2770);
xnor U4395 (N_4395,N_1199,N_2986);
and U4396 (N_4396,N_1812,N_2774);
and U4397 (N_4397,N_3775,N_150);
nand U4398 (N_4398,N_2165,N_943);
or U4399 (N_4399,N_2790,N_567);
or U4400 (N_4400,N_1568,N_3028);
nand U4401 (N_4401,N_3299,N_1184);
nand U4402 (N_4402,N_3498,N_3009);
nor U4403 (N_4403,N_2666,N_346);
or U4404 (N_4404,N_3691,N_3513);
nor U4405 (N_4405,N_1150,N_2004);
xor U4406 (N_4406,N_3364,N_1025);
nor U4407 (N_4407,N_543,N_678);
nor U4408 (N_4408,N_1474,N_1648);
nor U4409 (N_4409,N_547,N_851);
xor U4410 (N_4410,N_3759,N_1407);
and U4411 (N_4411,N_1730,N_3846);
or U4412 (N_4412,N_2158,N_2668);
xor U4413 (N_4413,N_2168,N_3616);
nand U4414 (N_4414,N_1112,N_3271);
and U4415 (N_4415,N_3151,N_1827);
or U4416 (N_4416,N_1560,N_1695);
nor U4417 (N_4417,N_540,N_635);
xor U4418 (N_4418,N_1447,N_2866);
nand U4419 (N_4419,N_2599,N_3841);
or U4420 (N_4420,N_2508,N_2991);
nand U4421 (N_4421,N_3600,N_3508);
and U4422 (N_4422,N_1121,N_3419);
and U4423 (N_4423,N_3331,N_983);
nand U4424 (N_4424,N_1287,N_3100);
nor U4425 (N_4425,N_3141,N_2839);
or U4426 (N_4426,N_1546,N_1774);
nor U4427 (N_4427,N_3137,N_1794);
nor U4428 (N_4428,N_921,N_633);
or U4429 (N_4429,N_3815,N_369);
xor U4430 (N_4430,N_729,N_31);
or U4431 (N_4431,N_1444,N_3311);
nor U4432 (N_4432,N_2025,N_444);
and U4433 (N_4433,N_3091,N_1933);
and U4434 (N_4434,N_3128,N_2728);
and U4435 (N_4435,N_1808,N_534);
nand U4436 (N_4436,N_578,N_3294);
nor U4437 (N_4437,N_2341,N_3917);
xor U4438 (N_4438,N_533,N_3556);
or U4439 (N_4439,N_142,N_371);
and U4440 (N_4440,N_1893,N_374);
nand U4441 (N_4441,N_494,N_1456);
xnor U4442 (N_4442,N_243,N_628);
nor U4443 (N_4443,N_1315,N_473);
nand U4444 (N_4444,N_668,N_3708);
nor U4445 (N_4445,N_308,N_1227);
or U4446 (N_4446,N_3062,N_1796);
or U4447 (N_4447,N_1352,N_166);
nor U4448 (N_4448,N_138,N_3291);
xnor U4449 (N_4449,N_3747,N_1734);
nand U4450 (N_4450,N_630,N_2616);
and U4451 (N_4451,N_132,N_1116);
or U4452 (N_4452,N_484,N_2116);
and U4453 (N_4453,N_1293,N_2479);
nor U4454 (N_4454,N_1976,N_1316);
and U4455 (N_4455,N_673,N_2780);
or U4456 (N_4456,N_2823,N_3923);
nor U4457 (N_4457,N_3093,N_70);
nand U4458 (N_4458,N_3627,N_1314);
or U4459 (N_4459,N_1220,N_2922);
or U4460 (N_4460,N_3773,N_396);
or U4461 (N_4461,N_2095,N_126);
nand U4462 (N_4462,N_1530,N_3260);
nor U4463 (N_4463,N_2454,N_2400);
nor U4464 (N_4464,N_3644,N_3385);
xnor U4465 (N_4465,N_3379,N_2837);
nand U4466 (N_4466,N_3840,N_2608);
xor U4467 (N_4467,N_1618,N_2587);
nand U4468 (N_4468,N_2336,N_993);
xor U4469 (N_4469,N_451,N_3349);
and U4470 (N_4470,N_2402,N_405);
or U4471 (N_4471,N_836,N_1520);
or U4472 (N_4472,N_626,N_1712);
nand U4473 (N_4473,N_1688,N_3441);
xor U4474 (N_4474,N_2225,N_3537);
nor U4475 (N_4475,N_538,N_3286);
xnor U4476 (N_4476,N_2064,N_175);
xnor U4477 (N_4477,N_2696,N_2640);
nor U4478 (N_4478,N_1747,N_661);
nand U4479 (N_4479,N_3191,N_2234);
and U4480 (N_4480,N_1971,N_1573);
nor U4481 (N_4481,N_3563,N_1708);
and U4482 (N_4482,N_2544,N_2633);
or U4483 (N_4483,N_3618,N_1014);
nand U4484 (N_4484,N_3589,N_1261);
and U4485 (N_4485,N_80,N_2040);
nand U4486 (N_4486,N_2554,N_2622);
nand U4487 (N_4487,N_2667,N_1442);
xnor U4488 (N_4488,N_1996,N_2264);
xnor U4489 (N_4489,N_1181,N_869);
nor U4490 (N_4490,N_65,N_2609);
nor U4491 (N_4491,N_2772,N_3844);
nor U4492 (N_4492,N_1987,N_3857);
and U4493 (N_4493,N_592,N_1088);
xnor U4494 (N_4494,N_2230,N_1068);
nand U4495 (N_4495,N_3715,N_2451);
xor U4496 (N_4496,N_640,N_3517);
xor U4497 (N_4497,N_2192,N_2255);
and U4498 (N_4498,N_2801,N_2900);
and U4499 (N_4499,N_2133,N_1776);
nand U4500 (N_4500,N_3662,N_481);
xor U4501 (N_4501,N_260,N_2619);
xor U4502 (N_4502,N_2821,N_1761);
xnor U4503 (N_4503,N_2440,N_1010);
nand U4504 (N_4504,N_1490,N_2232);
nor U4505 (N_4505,N_2177,N_3185);
nor U4506 (N_4506,N_2677,N_1782);
xor U4507 (N_4507,N_3347,N_3771);
and U4508 (N_4508,N_1403,N_3647);
or U4509 (N_4509,N_1076,N_2815);
xnor U4510 (N_4510,N_3425,N_3739);
nor U4511 (N_4511,N_977,N_3106);
and U4512 (N_4512,N_3433,N_1886);
nand U4513 (N_4513,N_3117,N_2288);
nor U4514 (N_4514,N_2119,N_361);
or U4515 (N_4515,N_1528,N_3515);
and U4516 (N_4516,N_3327,N_1370);
and U4517 (N_4517,N_3250,N_3693);
or U4518 (N_4518,N_232,N_1185);
and U4519 (N_4519,N_1471,N_3211);
nor U4520 (N_4520,N_3477,N_3551);
nor U4521 (N_4521,N_2724,N_2545);
and U4522 (N_4522,N_3701,N_201);
and U4523 (N_4523,N_959,N_2328);
nor U4524 (N_4524,N_1336,N_286);
nand U4525 (N_4525,N_3306,N_1070);
xnor U4526 (N_4526,N_2673,N_2256);
nand U4527 (N_4527,N_2059,N_2354);
or U4528 (N_4528,N_2523,N_2000);
nor U4529 (N_4529,N_3908,N_2769);
xor U4530 (N_4530,N_955,N_2074);
or U4531 (N_4531,N_364,N_771);
nand U4532 (N_4532,N_2916,N_1201);
and U4533 (N_4533,N_1562,N_2442);
nor U4534 (N_4534,N_3084,N_3046);
nor U4535 (N_4535,N_1922,N_2965);
nor U4536 (N_4536,N_2768,N_3707);
or U4537 (N_4537,N_2428,N_1436);
or U4538 (N_4538,N_2491,N_2902);
nor U4539 (N_4539,N_2314,N_2334);
xnor U4540 (N_4540,N_2157,N_1593);
or U4541 (N_4541,N_1175,N_989);
nor U4542 (N_4542,N_3574,N_3361);
and U4543 (N_4543,N_3110,N_826);
xnor U4544 (N_4544,N_456,N_3510);
and U4545 (N_4545,N_2367,N_813);
or U4546 (N_4546,N_690,N_3876);
or U4547 (N_4547,N_1888,N_1351);
nand U4548 (N_4548,N_3918,N_301);
or U4549 (N_4549,N_997,N_3251);
xor U4550 (N_4550,N_3412,N_2546);
and U4551 (N_4551,N_2982,N_2016);
or U4552 (N_4552,N_32,N_1296);
nand U4553 (N_4553,N_1214,N_3353);
nor U4554 (N_4554,N_3959,N_3505);
xnor U4555 (N_4555,N_3017,N_3532);
xnor U4556 (N_4556,N_1898,N_1291);
nor U4557 (N_4557,N_3659,N_3835);
nor U4558 (N_4558,N_3585,N_724);
xor U4559 (N_4559,N_2675,N_3466);
nand U4560 (N_4560,N_2421,N_515);
xnor U4561 (N_4561,N_3495,N_3631);
nor U4562 (N_4562,N_659,N_2203);
xnor U4563 (N_4563,N_1592,N_3276);
or U4564 (N_4564,N_3258,N_1432);
nor U4565 (N_4565,N_3825,N_3898);
and U4566 (N_4566,N_3706,N_3668);
xor U4567 (N_4567,N_2178,N_759);
xor U4568 (N_4568,N_825,N_778);
nor U4569 (N_4569,N_3579,N_603);
xnor U4570 (N_4570,N_787,N_1083);
xnor U4571 (N_4571,N_3954,N_3555);
nor U4572 (N_4572,N_859,N_2061);
xor U4573 (N_4573,N_1062,N_1521);
nor U4574 (N_4574,N_1118,N_1754);
nor U4575 (N_4575,N_3245,N_2921);
xnor U4576 (N_4576,N_2374,N_1824);
or U4577 (N_4577,N_2955,N_2830);
nand U4578 (N_4578,N_1746,N_1743);
xor U4579 (N_4579,N_2173,N_1767);
xor U4580 (N_4580,N_3232,N_1505);
nor U4581 (N_4581,N_3964,N_1243);
nor U4582 (N_4582,N_3373,N_1709);
nor U4583 (N_4583,N_1552,N_674);
or U4584 (N_4584,N_612,N_1867);
or U4585 (N_4585,N_53,N_905);
nor U4586 (N_4586,N_1975,N_447);
or U4587 (N_4587,N_224,N_3671);
and U4588 (N_4588,N_1146,N_3605);
xor U4589 (N_4589,N_2233,N_3602);
and U4590 (N_4590,N_315,N_165);
nand U4591 (N_4591,N_319,N_2713);
nand U4592 (N_4592,N_1974,N_815);
or U4593 (N_4593,N_3152,N_2073);
nor U4594 (N_4594,N_906,N_1598);
and U4595 (N_4595,N_2753,N_1488);
and U4596 (N_4596,N_1760,N_3511);
xnor U4597 (N_4597,N_3502,N_282);
and U4598 (N_4598,N_1402,N_3518);
nor U4599 (N_4599,N_1551,N_3619);
nand U4600 (N_4600,N_3703,N_3116);
or U4601 (N_4601,N_2360,N_2176);
or U4602 (N_4602,N_2826,N_1452);
and U4603 (N_4603,N_2489,N_3399);
nor U4604 (N_4604,N_1952,N_3060);
and U4605 (N_4605,N_205,N_671);
and U4606 (N_4606,N_1132,N_3277);
nand U4607 (N_4607,N_2788,N_1602);
nand U4608 (N_4608,N_455,N_1089);
nor U4609 (N_4609,N_2574,N_3680);
xnor U4610 (N_4610,N_774,N_135);
xor U4611 (N_4611,N_85,N_3667);
and U4612 (N_4612,N_1597,N_2814);
or U4613 (N_4613,N_1000,N_3957);
nor U4614 (N_4614,N_2940,N_3998);
xnor U4615 (N_4615,N_2834,N_953);
or U4616 (N_4616,N_3463,N_1591);
and U4617 (N_4617,N_931,N_3658);
xnor U4618 (N_4618,N_2784,N_2522);
nand U4619 (N_4619,N_1285,N_1720);
xnor U4620 (N_4620,N_248,N_1931);
nand U4621 (N_4621,N_3491,N_1174);
and U4622 (N_4622,N_69,N_968);
xor U4623 (N_4623,N_13,N_1940);
xnor U4624 (N_4624,N_951,N_372);
nor U4625 (N_4625,N_1753,N_658);
xor U4626 (N_4626,N_3673,N_2304);
nand U4627 (N_4627,N_2654,N_3422);
nor U4628 (N_4628,N_2024,N_206);
xnor U4629 (N_4629,N_1312,N_3088);
nand U4630 (N_4630,N_472,N_3714);
nand U4631 (N_4631,N_573,N_523);
or U4632 (N_4632,N_1854,N_2281);
xnor U4633 (N_4633,N_1696,N_2286);
or U4634 (N_4634,N_255,N_1815);
and U4635 (N_4635,N_3749,N_3880);
and U4636 (N_4636,N_2340,N_228);
nor U4637 (N_4637,N_3696,N_2047);
nand U4638 (N_4638,N_1599,N_3124);
and U4639 (N_4639,N_1873,N_2858);
nor U4640 (N_4640,N_3592,N_856);
xnor U4641 (N_4641,N_331,N_2419);
or U4642 (N_4642,N_3333,N_3166);
nor U4643 (N_4643,N_1777,N_914);
xnor U4644 (N_4644,N_3252,N_385);
and U4645 (N_4645,N_2754,N_296);
xnor U4646 (N_4646,N_2765,N_3235);
and U4647 (N_4647,N_797,N_471);
xor U4648 (N_4648,N_3649,N_410);
nor U4649 (N_4649,N_3883,N_732);
nand U4650 (N_4650,N_642,N_3394);
and U4651 (N_4651,N_3165,N_2020);
or U4652 (N_4652,N_1206,N_1885);
nor U4653 (N_4653,N_280,N_2658);
xor U4654 (N_4654,N_295,N_2567);
nor U4655 (N_4655,N_3650,N_1263);
nand U4656 (N_4656,N_3906,N_670);
xor U4657 (N_4657,N_1009,N_207);
and U4658 (N_4658,N_772,N_3058);
nand U4659 (N_4659,N_3590,N_1994);
xor U4660 (N_4660,N_991,N_378);
and U4661 (N_4661,N_2252,N_584);
nand U4662 (N_4662,N_35,N_2457);
xor U4663 (N_4663,N_16,N_1479);
nor U4664 (N_4664,N_1392,N_1955);
nor U4665 (N_4665,N_1938,N_134);
or U4666 (N_4666,N_998,N_894);
xnor U4667 (N_4667,N_3439,N_749);
or U4668 (N_4668,N_3504,N_3266);
and U4669 (N_4669,N_1330,N_3045);
xnor U4670 (N_4670,N_3922,N_922);
nor U4671 (N_4671,N_1325,N_1832);
or U4672 (N_4672,N_3179,N_2051);
nor U4673 (N_4673,N_1234,N_1138);
nand U4674 (N_4674,N_1135,N_3030);
nor U4675 (N_4675,N_736,N_2722);
nand U4676 (N_4676,N_2951,N_3388);
nor U4677 (N_4677,N_3866,N_940);
nand U4678 (N_4678,N_589,N_3882);
nor U4679 (N_4679,N_3340,N_2732);
or U4680 (N_4680,N_1604,N_306);
and U4681 (N_4681,N_907,N_1023);
or U4682 (N_4682,N_1759,N_1139);
or U4683 (N_4683,N_1806,N_950);
nand U4684 (N_4684,N_225,N_1851);
xor U4685 (N_4685,N_59,N_3961);
nand U4686 (N_4686,N_604,N_1344);
nor U4687 (N_4687,N_76,N_2130);
and U4688 (N_4688,N_3948,N_1590);
xnor U4689 (N_4689,N_2980,N_1387);
xor U4690 (N_4690,N_1123,N_3121);
nor U4691 (N_4691,N_3473,N_3139);
xnor U4692 (N_4692,N_2660,N_513);
xor U4693 (N_4693,N_3591,N_1250);
or U4694 (N_4694,N_469,N_3687);
or U4695 (N_4695,N_2632,N_1550);
nor U4696 (N_4696,N_1506,N_283);
xnor U4697 (N_4697,N_2656,N_3669);
or U4698 (N_4698,N_3042,N_3521);
xnor U4699 (N_4699,N_215,N_1577);
and U4700 (N_4700,N_1238,N_3626);
xor U4701 (N_4701,N_2468,N_2235);
nand U4702 (N_4702,N_1347,N_298);
and U4703 (N_4703,N_1230,N_1523);
and U4704 (N_4704,N_2427,N_3889);
nor U4705 (N_4705,N_2144,N_2607);
or U4706 (N_4706,N_625,N_2595);
xnor U4707 (N_4707,N_957,N_404);
nor U4708 (N_4708,N_1576,N_58);
xor U4709 (N_4709,N_161,N_3558);
or U4710 (N_4710,N_140,N_409);
and U4711 (N_4711,N_1152,N_1226);
nand U4712 (N_4712,N_1069,N_445);
or U4713 (N_4713,N_2720,N_1271);
and U4714 (N_4714,N_839,N_2653);
nor U4715 (N_4715,N_1644,N_352);
xnor U4716 (N_4716,N_2012,N_1856);
nand U4717 (N_4717,N_2156,N_1908);
or U4718 (N_4718,N_2615,N_338);
nor U4719 (N_4719,N_2933,N_2393);
or U4720 (N_4720,N_2655,N_454);
xor U4721 (N_4721,N_3443,N_3012);
nor U4722 (N_4722,N_2800,N_474);
nand U4723 (N_4723,N_916,N_1822);
and U4724 (N_4724,N_872,N_781);
xor U4725 (N_4725,N_2911,N_880);
nand U4726 (N_4726,N_3725,N_3720);
nor U4727 (N_4727,N_2776,N_2716);
or U4728 (N_4728,N_1276,N_291);
nor U4729 (N_4729,N_3114,N_1624);
or U4730 (N_4730,N_3218,N_1835);
or U4731 (N_4731,N_2832,N_3928);
or U4732 (N_4732,N_342,N_1943);
and U4733 (N_4733,N_226,N_244);
or U4734 (N_4734,N_322,N_1948);
nand U4735 (N_4735,N_990,N_2347);
xor U4736 (N_4736,N_170,N_1019);
xnor U4737 (N_4737,N_1379,N_2464);
or U4738 (N_4738,N_1481,N_1966);
nor U4739 (N_4739,N_3978,N_2516);
or U4740 (N_4740,N_1820,N_1163);
xor U4741 (N_4741,N_3417,N_3983);
nor U4742 (N_4742,N_3623,N_3358);
or U4743 (N_4743,N_247,N_1833);
or U4744 (N_4744,N_3500,N_490);
xnor U4745 (N_4745,N_1482,N_2828);
or U4746 (N_4746,N_1522,N_96);
xor U4747 (N_4747,N_1636,N_1798);
and U4748 (N_4748,N_2778,N_1458);
nor U4749 (N_4749,N_52,N_3868);
nand U4750 (N_4750,N_1567,N_1772);
nor U4751 (N_4751,N_2847,N_3044);
xnor U4752 (N_4752,N_521,N_1332);
or U4753 (N_4753,N_2691,N_430);
and U4754 (N_4754,N_2944,N_660);
and U4755 (N_4755,N_3520,N_2649);
xnor U4756 (N_4756,N_1553,N_3885);
or U4757 (N_4757,N_1324,N_2013);
nor U4758 (N_4758,N_3528,N_1642);
or U4759 (N_4759,N_2743,N_400);
and U4760 (N_4760,N_1128,N_3595);
or U4761 (N_4761,N_946,N_2698);
xor U4762 (N_4762,N_2070,N_1095);
xnor U4763 (N_4763,N_1190,N_2941);
nor U4764 (N_4764,N_2863,N_3172);
and U4765 (N_4765,N_2905,N_3613);
nor U4766 (N_4766,N_401,N_917);
and U4767 (N_4767,N_3965,N_3095);
nor U4768 (N_4768,N_1431,N_2960);
nand U4769 (N_4769,N_1028,N_1006);
nand U4770 (N_4770,N_2076,N_3695);
xor U4771 (N_4771,N_2257,N_173);
xor U4772 (N_4772,N_3318,N_1752);
nand U4773 (N_4773,N_1751,N_1561);
xor U4774 (N_4774,N_437,N_714);
and U4775 (N_4775,N_256,N_353);
nand U4776 (N_4776,N_1450,N_2248);
nor U4777 (N_4777,N_426,N_2305);
nor U4778 (N_4778,N_1899,N_1273);
or U4779 (N_4779,N_3267,N_1638);
nor U4780 (N_4780,N_1736,N_75);
nand U4781 (N_4781,N_956,N_2582);
xor U4782 (N_4782,N_373,N_3480);
and U4783 (N_4783,N_2422,N_2436);
nor U4784 (N_4784,N_3052,N_613);
or U4785 (N_4785,N_2426,N_1839);
or U4786 (N_4786,N_1540,N_3972);
or U4787 (N_4787,N_1868,N_2846);
and U4788 (N_4788,N_822,N_3549);
or U4789 (N_4789,N_3120,N_478);
nand U4790 (N_4790,N_1740,N_1104);
or U4791 (N_4791,N_3683,N_1606);
nor U4792 (N_4792,N_1701,N_3874);
and U4793 (N_4793,N_3810,N_3899);
nand U4794 (N_4794,N_2456,N_1641);
nor U4795 (N_4795,N_903,N_3050);
nor U4796 (N_4796,N_1511,N_419);
xor U4797 (N_4797,N_2700,N_3832);
or U4798 (N_4798,N_3171,N_3546);
nor U4799 (N_4799,N_2810,N_3823);
nor U4800 (N_4800,N_1645,N_2394);
nand U4801 (N_4801,N_2345,N_23);
xor U4802 (N_4802,N_2139,N_2603);
or U4803 (N_4803,N_865,N_9);
xor U4804 (N_4804,N_2657,N_2127);
nand U4805 (N_4805,N_3307,N_3776);
or U4806 (N_4806,N_3809,N_185);
and U4807 (N_4807,N_1394,N_3843);
or U4808 (N_4808,N_1013,N_2851);
or U4809 (N_4809,N_304,N_2399);
xnor U4810 (N_4810,N_1614,N_3392);
nand U4811 (N_4811,N_2350,N_619);
nor U4812 (N_4812,N_727,N_870);
nor U4813 (N_4813,N_2027,N_2746);
and U4814 (N_4814,N_245,N_3198);
nand U4815 (N_4815,N_3096,N_705);
nand U4816 (N_4816,N_2184,N_2272);
and U4817 (N_4817,N_1997,N_3966);
or U4818 (N_4818,N_1780,N_290);
and U4819 (N_4819,N_976,N_695);
nor U4820 (N_4820,N_3748,N_3445);
or U4821 (N_4821,N_2131,N_1862);
nor U4822 (N_4822,N_1526,N_3733);
xnor U4823 (N_4823,N_1717,N_583);
nor U4824 (N_4824,N_102,N_591);
nor U4825 (N_4825,N_1803,N_1840);
and U4826 (N_4826,N_90,N_199);
xnor U4827 (N_4827,N_2323,N_2423);
or U4828 (N_4828,N_1346,N_3200);
or U4829 (N_4829,N_137,N_39);
xnor U4830 (N_4830,N_2547,N_704);
nor U4831 (N_4831,N_3493,N_2861);
nor U4832 (N_4832,N_2415,N_3283);
nand U4833 (N_4833,N_1119,N_1257);
nor U4834 (N_4834,N_2039,N_2474);
nor U4835 (N_4835,N_1295,N_1853);
and U4836 (N_4836,N_3620,N_3345);
or U4837 (N_4837,N_2564,N_3420);
nand U4838 (N_4838,N_3719,N_468);
nand U4839 (N_4839,N_2443,N_1874);
xnor U4840 (N_4840,N_2310,N_516);
or U4841 (N_4841,N_665,N_1099);
nand U4842 (N_4842,N_536,N_2693);
nor U4843 (N_4843,N_2510,N_2605);
nor U4844 (N_4844,N_1084,N_849);
nand U4845 (N_4845,N_974,N_2349);
xor U4846 (N_4846,N_130,N_0);
nand U4847 (N_4847,N_144,N_2486);
xnor U4848 (N_4848,N_2229,N_2238);
or U4849 (N_4849,N_3249,N_2200);
and U4850 (N_4850,N_2299,N_3547);
and U4851 (N_4851,N_2371,N_730);
nor U4852 (N_4852,N_1818,N_380);
nand U4853 (N_4853,N_2412,N_2690);
and U4854 (N_4854,N_3073,N_2217);
nand U4855 (N_4855,N_1305,N_1549);
xor U4856 (N_4856,N_3132,N_1329);
or U4857 (N_4857,N_3125,N_1587);
or U4858 (N_4858,N_2189,N_558);
xor U4859 (N_4859,N_436,N_3337);
nor U4860 (N_4860,N_2202,N_3034);
nand U4861 (N_4861,N_1489,N_1267);
and U4862 (N_4862,N_1858,N_3543);
xor U4863 (N_4863,N_1881,N_1756);
xnor U4864 (N_4864,N_2684,N_3113);
nor U4865 (N_4865,N_271,N_2104);
and U4866 (N_4866,N_21,N_1529);
nor U4867 (N_4867,N_2505,N_278);
nor U4868 (N_4868,N_3753,N_2355);
or U4869 (N_4869,N_3393,N_987);
xnor U4870 (N_4870,N_106,N_1548);
and U4871 (N_4871,N_3409,N_3367);
and U4872 (N_4872,N_3951,N_2882);
nor U4873 (N_4873,N_2597,N_183);
xnor U4874 (N_4874,N_1018,N_2110);
and U4875 (N_4875,N_3241,N_1377);
and U4876 (N_4876,N_1935,N_81);
xnor U4877 (N_4877,N_2848,N_3025);
xnor U4878 (N_4878,N_3675,N_576);
nand U4879 (N_4879,N_3881,N_3049);
xnor U4880 (N_4880,N_1900,N_1857);
nor U4881 (N_4881,N_3943,N_1723);
nand U4882 (N_4882,N_2265,N_2223);
and U4883 (N_4883,N_1433,N_2430);
and U4884 (N_4884,N_3156,N_2625);
xor U4885 (N_4885,N_3679,N_3451);
nor U4886 (N_4886,N_2807,N_1274);
xnor U4887 (N_4887,N_1210,N_1323);
nor U4888 (N_4888,N_785,N_1129);
and U4889 (N_4889,N_2585,N_3133);
and U4890 (N_4890,N_3934,N_3902);
or U4891 (N_4891,N_636,N_3341);
xnor U4892 (N_4892,N_3682,N_3580);
nor U4893 (N_4893,N_3295,N_3148);
nand U4894 (N_4894,N_2835,N_2420);
and U4895 (N_4895,N_1120,N_2208);
and U4896 (N_4896,N_606,N_2473);
nand U4897 (N_4897,N_1096,N_3798);
or U4898 (N_4898,N_1919,N_688);
or U4899 (N_4899,N_1510,N_3037);
nor U4900 (N_4900,N_1579,N_1225);
xnor U4901 (N_4901,N_1045,N_181);
nand U4902 (N_4902,N_3573,N_2292);
xnor U4903 (N_4903,N_2296,N_2333);
nand U4904 (N_4904,N_590,N_3674);
nand U4905 (N_4905,N_2335,N_1143);
xnor U4906 (N_4906,N_669,N_1983);
nand U4907 (N_4907,N_1515,N_2525);
nand U4908 (N_4908,N_2596,N_1564);
xnor U4909 (N_4909,N_2031,N_1008);
xnor U4910 (N_4910,N_1493,N_395);
nand U4911 (N_4911,N_2741,N_887);
xnor U4912 (N_4912,N_3509,N_2890);
and U4913 (N_4913,N_2604,N_2028);
or U4914 (N_4914,N_3630,N_210);
nand U4915 (N_4915,N_50,N_2910);
or U4916 (N_4916,N_644,N_2135);
xnor U4917 (N_4917,N_2321,N_66);
nor U4918 (N_4918,N_3242,N_898);
nand U4919 (N_4919,N_1563,N_2829);
xor U4920 (N_4920,N_594,N_556);
nor U4921 (N_4921,N_2723,N_3779);
xnor U4922 (N_4922,N_2850,N_1860);
or U4923 (N_4923,N_967,N_2170);
or U4924 (N_4924,N_2322,N_1787);
nand U4925 (N_4925,N_446,N_1517);
nand U4926 (N_4926,N_2263,N_2708);
nor U4927 (N_4927,N_2187,N_209);
or U4928 (N_4928,N_2816,N_3081);
nor U4929 (N_4929,N_2729,N_212);
or U4930 (N_4930,N_249,N_3278);
or U4931 (N_4931,N_932,N_526);
nor U4932 (N_4932,N_3661,N_1993);
and U4933 (N_4933,N_3921,N_2358);
and U4934 (N_4934,N_3772,N_2107);
xor U4935 (N_4935,N_3813,N_1232);
and U4936 (N_4936,N_2297,N_2978);
or U4937 (N_4937,N_1258,N_3288);
or U4938 (N_4938,N_3010,N_938);
xnor U4939 (N_4939,N_64,N_2204);
and U4940 (N_4940,N_2467,N_3656);
xnor U4941 (N_4941,N_349,N_2048);
nand U4942 (N_4942,N_1578,N_561);
or U4943 (N_4943,N_2090,N_3736);
nand U4944 (N_4944,N_2151,N_2543);
nand U4945 (N_4945,N_2282,N_1714);
nand U4946 (N_4946,N_1834,N_3257);
nand U4947 (N_4947,N_3372,N_236);
or U4948 (N_4948,N_1080,N_2727);
nand U4949 (N_4949,N_443,N_1038);
nor U4950 (N_4950,N_2542,N_1097);
nand U4951 (N_4951,N_3572,N_1368);
and U4952 (N_4952,N_3988,N_3766);
xor U4953 (N_4953,N_1419,N_1821);
and U4954 (N_4954,N_2929,N_978);
xnor U4955 (N_4955,N_2892,N_2160);
and U4956 (N_4956,N_657,N_285);
nor U4957 (N_4957,N_3945,N_824);
and U4958 (N_4958,N_2733,N_1303);
or U4959 (N_4959,N_986,N_841);
nand U4960 (N_4960,N_461,N_1093);
and U4961 (N_4961,N_3819,N_2959);
or U4962 (N_4962,N_1194,N_2731);
nor U4963 (N_4963,N_2069,N_3024);
or U4964 (N_4964,N_2529,N_1581);
nor U4965 (N_4965,N_2775,N_2527);
nand U4966 (N_4966,N_939,N_397);
nand U4967 (N_4967,N_3755,N_1731);
or U4968 (N_4968,N_2470,N_1925);
and U4969 (N_4969,N_1487,N_2669);
or U4970 (N_4970,N_763,N_2870);
or U4971 (N_4971,N_2984,N_1785);
or U4972 (N_4972,N_3941,N_3131);
or U4973 (N_4973,N_3486,N_1837);
xor U4974 (N_4974,N_2626,N_624);
and U4975 (N_4975,N_1547,N_1327);
and U4976 (N_4976,N_1191,N_1073);
nand U4977 (N_4977,N_3236,N_2538);
xor U4978 (N_4978,N_2932,N_3946);
or U4979 (N_4979,N_3963,N_2348);
nor U4980 (N_4980,N_2871,N_1147);
xnor U4981 (N_4981,N_1335,N_2058);
xor U4982 (N_4982,N_155,N_3007);
or U4983 (N_4983,N_503,N_440);
or U4984 (N_4984,N_3646,N_3195);
and U4985 (N_4985,N_1861,N_3507);
and U4986 (N_4986,N_1726,N_3237);
and U4987 (N_4987,N_3449,N_3471);
nor U4988 (N_4988,N_1634,N_2550);
nor U4989 (N_4989,N_164,N_3860);
nor U4990 (N_4990,N_2843,N_1750);
and U4991 (N_4991,N_3228,N_3207);
nand U4992 (N_4992,N_2268,N_3304);
nand U4993 (N_4993,N_843,N_464);
nand U4994 (N_4994,N_2045,N_1739);
nand U4995 (N_4995,N_107,N_3538);
and U4996 (N_4996,N_2903,N_3666);
nor U4997 (N_4997,N_2140,N_2961);
nand U4998 (N_4998,N_3911,N_1188);
nand U4999 (N_4999,N_3723,N_2346);
or U5000 (N_5000,N_1406,N_3761);
xnor U5001 (N_5001,N_1114,N_3664);
or U5002 (N_5002,N_715,N_3803);
and U5003 (N_5003,N_3297,N_420);
xnor U5004 (N_5004,N_190,N_1216);
xor U5005 (N_5005,N_549,N_1666);
nand U5006 (N_5006,N_3821,N_2273);
xnor U5007 (N_5007,N_3109,N_434);
or U5008 (N_5008,N_597,N_832);
nand U5009 (N_5009,N_768,N_3261);
or U5010 (N_5010,N_1326,N_2408);
nand U5011 (N_5011,N_1792,N_982);
nand U5012 (N_5012,N_709,N_1137);
and U5013 (N_5013,N_151,N_3718);
nand U5014 (N_5014,N_581,N_890);
xor U5015 (N_5015,N_3322,N_429);
nand U5016 (N_5016,N_2096,N_3438);
xor U5017 (N_5017,N_3280,N_1144);
nand U5018 (N_5018,N_2018,N_1607);
nor U5019 (N_5019,N_2466,N_2862);
and U5020 (N_5020,N_3888,N_2191);
and U5021 (N_5021,N_2520,N_2113);
nor U5022 (N_5022,N_2431,N_294);
xnor U5023 (N_5023,N_554,N_2163);
nor U5024 (N_5024,N_2138,N_2617);
xor U5025 (N_5025,N_449,N_518);
or U5026 (N_5026,N_2487,N_1682);
nor U5027 (N_5027,N_1990,N_1459);
xnor U5028 (N_5028,N_337,N_2098);
nor U5029 (N_5029,N_417,N_1036);
nand U5030 (N_5030,N_2771,N_2246);
nand U5031 (N_5031,N_2132,N_3746);
xor U5032 (N_5032,N_2488,N_2490);
or U5033 (N_5033,N_399,N_3987);
and U5034 (N_5034,N_3982,N_1411);
nor U5035 (N_5035,N_1498,N_1619);
xnor U5036 (N_5036,N_1639,N_268);
xor U5037 (N_5037,N_572,N_3434);
nor U5038 (N_5038,N_1061,N_3146);
nand U5039 (N_5039,N_808,N_3596);
xor U5040 (N_5040,N_3416,N_2777);
and U5041 (N_5041,N_1501,N_3816);
nand U5042 (N_5042,N_38,N_3270);
and U5043 (N_5043,N_1883,N_2206);
nor U5044 (N_5044,N_3593,N_2183);
xor U5045 (N_5045,N_2437,N_3273);
or U5046 (N_5046,N_1534,N_2171);
xor U5047 (N_5047,N_3282,N_1674);
or U5048 (N_5048,N_2118,N_3594);
xnor U5049 (N_5049,N_2212,N_2888);
or U5050 (N_5050,N_864,N_3994);
xor U5051 (N_5051,N_3740,N_816);
or U5052 (N_5052,N_3300,N_3002);
xor U5053 (N_5053,N_2063,N_398);
xnor U5054 (N_5054,N_2561,N_531);
or U5055 (N_5055,N_146,N_761);
and U5056 (N_5056,N_2290,N_2808);
and U5057 (N_5057,N_2549,N_1972);
and U5058 (N_5058,N_2376,N_1961);
xnor U5059 (N_5059,N_277,N_408);
and U5060 (N_5060,N_835,N_582);
xnor U5061 (N_5061,N_652,N_1391);
and U5062 (N_5062,N_685,N_2989);
or U5063 (N_5063,N_1913,N_2880);
and U5064 (N_5064,N_3335,N_2240);
or U5065 (N_5065,N_3490,N_627);
nor U5066 (N_5066,N_3265,N_960);
nand U5067 (N_5067,N_936,N_1172);
xor U5068 (N_5068,N_1707,N_2361);
nor U5069 (N_5069,N_1085,N_629);
nand U5070 (N_5070,N_728,N_1103);
xor U5071 (N_5071,N_530,N_176);
and U5072 (N_5072,N_2043,N_2919);
nor U5073 (N_5073,N_1060,N_320);
xor U5074 (N_5074,N_423,N_913);
and U5075 (N_5075,N_3981,N_580);
xor U5076 (N_5076,N_3222,N_559);
and U5077 (N_5077,N_1288,N_545);
xnor U5078 (N_5078,N_1852,N_3458);
xnor U5079 (N_5079,N_2438,N_3206);
nand U5080 (N_5080,N_2065,N_1681);
nand U5081 (N_5081,N_1451,N_1483);
xnor U5082 (N_5082,N_3645,N_3163);
and U5083 (N_5083,N_1504,N_964);
nand U5084 (N_5084,N_1371,N_1236);
xor U5085 (N_5085,N_1514,N_2838);
or U5086 (N_5086,N_2312,N_477);
nor U5087 (N_5087,N_2313,N_1667);
nand U5088 (N_5088,N_1725,N_1843);
xor U5089 (N_5089,N_2565,N_3094);
xnor U5090 (N_5090,N_1801,N_3873);
xnor U5091 (N_5091,N_3183,N_2357);
or U5092 (N_5092,N_2389,N_254);
nand U5093 (N_5093,N_3488,N_2153);
and U5094 (N_5094,N_3858,N_3459);
or U5095 (N_5095,N_958,N_3326);
xor U5096 (N_5096,N_15,N_3129);
nand U5097 (N_5097,N_2931,N_3870);
and U5098 (N_5098,N_2418,N_3636);
and U5099 (N_5099,N_1424,N_1283);
nor U5100 (N_5100,N_3865,N_3281);
xor U5101 (N_5101,N_2799,N_3118);
xor U5102 (N_5102,N_1907,N_3986);
xnor U5103 (N_5103,N_2901,N_574);
xor U5104 (N_5104,N_1390,N_1741);
xnor U5105 (N_5105,N_2629,N_17);
nand U5106 (N_5106,N_1890,N_1871);
or U5107 (N_5107,N_3435,N_1713);
xnor U5108 (N_5108,N_3919,N_47);
nand U5109 (N_5109,N_2526,N_88);
xor U5110 (N_5110,N_1969,N_2949);
nand U5111 (N_5111,N_2738,N_1603);
nor U5112 (N_5112,N_1958,N_3785);
nand U5113 (N_5113,N_3197,N_949);
xor U5114 (N_5114,N_191,N_1005);
nor U5115 (N_5115,N_1477,N_3699);
and U5116 (N_5116,N_1640,N_3849);
xor U5117 (N_5117,N_3262,N_1909);
nand U5118 (N_5118,N_1901,N_457);
nand U5119 (N_5119,N_1850,N_2513);
nor U5120 (N_5120,N_2122,N_3348);
nand U5121 (N_5121,N_769,N_2792);
xnor U5122 (N_5122,N_3914,N_84);
or U5123 (N_5123,N_889,N_2553);
and U5124 (N_5124,N_415,N_3512);
nand U5125 (N_5125,N_651,N_1453);
and U5126 (N_5126,N_63,N_3728);
or U5127 (N_5127,N_3421,N_1535);
and U5128 (N_5128,N_2267,N_168);
and U5129 (N_5129,N_1497,N_465);
xor U5130 (N_5130,N_2188,N_2971);
nand U5131 (N_5131,N_2719,N_831);
and U5132 (N_5132,N_3055,N_2435);
nor U5133 (N_5133,N_3611,N_1763);
nor U5134 (N_5134,N_3711,N_3758);
or U5135 (N_5135,N_867,N_2638);
xor U5136 (N_5136,N_1427,N_3405);
nand U5137 (N_5137,N_1395,N_641);
nor U5138 (N_5138,N_3665,N_3053);
nand U5139 (N_5139,N_2287,N_3962);
and U5140 (N_5140,N_1133,N_1322);
nand U5141 (N_5141,N_2062,N_1711);
xor U5142 (N_5142,N_3315,N_2056);
nand U5143 (N_5143,N_1349,N_318);
and U5144 (N_5144,N_265,N_2692);
or U5145 (N_5145,N_3279,N_1875);
xor U5146 (N_5146,N_2066,N_3320);
nand U5147 (N_5147,N_664,N_220);
nor U5148 (N_5148,N_1485,N_3408);
xnor U5149 (N_5149,N_3713,N_14);
nor U5150 (N_5150,N_3208,N_1702);
xor U5151 (N_5151,N_2956,N_1584);
and U5152 (N_5152,N_708,N_3980);
or U5153 (N_5153,N_406,N_2106);
or U5154 (N_5154,N_3292,N_3751);
nand U5155 (N_5155,N_2824,N_3818);
and U5156 (N_5156,N_2997,N_427);
nand U5157 (N_5157,N_3368,N_507);
nand U5158 (N_5158,N_748,N_1572);
and U5159 (N_5159,N_897,N_216);
or U5160 (N_5160,N_3893,N_2444);
nor U5161 (N_5161,N_779,N_324);
xnor U5162 (N_5162,N_1180,N_579);
nor U5163 (N_5163,N_3360,N_1467);
xor U5164 (N_5164,N_2030,N_2382);
nand U5165 (N_5165,N_2972,N_1665);
nor U5166 (N_5166,N_1884,N_1957);
and U5167 (N_5167,N_219,N_1253);
nand U5168 (N_5168,N_2480,N_3298);
and U5169 (N_5169,N_2683,N_2876);
nor U5170 (N_5170,N_421,N_3784);
nor U5171 (N_5171,N_3376,N_3470);
and U5172 (N_5172,N_3127,N_1037);
xnor U5173 (N_5173,N_2559,N_823);
or U5174 (N_5174,N_1317,N_403);
nand U5175 (N_5175,N_751,N_1380);
xor U5176 (N_5176,N_2950,N_131);
and U5177 (N_5177,N_616,N_411);
nor U5178 (N_5178,N_1308,N_2337);
or U5179 (N_5179,N_1004,N_2041);
nor U5180 (N_5180,N_1664,N_2338);
nor U5181 (N_5181,N_3167,N_83);
or U5182 (N_5182,N_1710,N_1600);
and U5183 (N_5183,N_3915,N_2339);
nor U5184 (N_5184,N_407,N_1003);
and U5185 (N_5185,N_3794,N_2540);
or U5186 (N_5186,N_3487,N_287);
nand U5187 (N_5187,N_467,N_3762);
or U5188 (N_5188,N_1024,N_3374);
nand U5189 (N_5189,N_2996,N_1903);
nor U5190 (N_5190,N_2001,N_928);
and U5191 (N_5191,N_2796,N_2181);
and U5192 (N_5192,N_2580,N_1866);
or U5193 (N_5193,N_1655,N_3231);
or U5194 (N_5194,N_1984,N_72);
nand U5195 (N_5195,N_2579,N_2411);
or U5196 (N_5196,N_2363,N_3685);
nor U5197 (N_5197,N_2562,N_2159);
or U5198 (N_5198,N_3189,N_1797);
and U5199 (N_5199,N_2938,N_499);
or U5200 (N_5200,N_2037,N_453);
and U5201 (N_5201,N_1361,N_204);
and U5202 (N_5202,N_2519,N_3454);
and U5203 (N_5203,N_1623,N_3196);
or U5204 (N_5204,N_347,N_388);
and U5205 (N_5205,N_2236,N_1389);
nand U5206 (N_5206,N_2895,N_2068);
nand U5207 (N_5207,N_566,N_3026);
nor U5208 (N_5208,N_2029,N_2934);
xor U5209 (N_5209,N_386,N_966);
or U5210 (N_5210,N_1828,N_1804);
and U5211 (N_5211,N_3950,N_297);
nand U5212 (N_5212,N_2102,N_863);
nand U5213 (N_5213,N_2067,N_74);
xor U5214 (N_5214,N_2714,N_1651);
and U5215 (N_5215,N_2266,N_2954);
xnor U5216 (N_5216,N_1995,N_12);
nand U5217 (N_5217,N_3688,N_1192);
or U5218 (N_5218,N_2952,N_1923);
and U5219 (N_5219,N_2372,N_3910);
xnor U5220 (N_5220,N_3564,N_3831);
nand U5221 (N_5221,N_2,N_1079);
or U5222 (N_5222,N_1173,N_746);
or U5223 (N_5223,N_2088,N_1203);
nor U5224 (N_5224,N_3015,N_356);
and U5225 (N_5225,N_2551,N_392);
and U5226 (N_5226,N_598,N_1176);
or U5227 (N_5227,N_2957,N_1609);
nand U5228 (N_5228,N_127,N_999);
xnor U5229 (N_5229,N_2661,N_791);
nor U5230 (N_5230,N_3432,N_2977);
nor U5231 (N_5231,N_707,N_1703);
nand U5232 (N_5232,N_692,N_3332);
xnor U5233 (N_5233,N_934,N_2484);
nor U5234 (N_5234,N_2498,N_2143);
xor U5235 (N_5235,N_840,N_1383);
or U5236 (N_5236,N_2893,N_3805);
nor U5237 (N_5237,N_1171,N_2618);
nand U5238 (N_5238,N_2859,N_2742);
nand U5239 (N_5239,N_1802,N_902);
and U5240 (N_5240,N_289,N_30);
and U5241 (N_5241,N_3710,N_3215);
nor U5242 (N_5242,N_2134,N_3464);
nor U5243 (N_5243,N_3365,N_3635);
nand U5244 (N_5244,N_3305,N_1947);
nand U5245 (N_5245,N_1637,N_2042);
or U5246 (N_5246,N_3071,N_3475);
and U5247 (N_5247,N_1558,N_1359);
and U5248 (N_5248,N_2904,N_3721);
nor U5249 (N_5249,N_3075,N_2289);
xor U5250 (N_5250,N_3526,N_3757);
nand U5251 (N_5251,N_3048,N_177);
and U5252 (N_5252,N_1894,N_3160);
or U5253 (N_5253,N_67,N_1187);
nor U5254 (N_5254,N_3248,N_1662);
nand U5255 (N_5255,N_1048,N_1015);
xnor U5256 (N_5256,N_1622,N_172);
xor U5257 (N_5257,N_1878,N_321);
nor U5258 (N_5258,N_853,N_2864);
nor U5259 (N_5259,N_377,N_3199);
or U5260 (N_5260,N_1113,N_51);
and U5261 (N_5261,N_1672,N_1002);
nor U5262 (N_5262,N_1343,N_3442);
nand U5263 (N_5263,N_2469,N_3006);
and U5264 (N_5264,N_1569,N_2600);
and U5265 (N_5265,N_910,N_1212);
nor U5266 (N_5266,N_722,N_2149);
xor U5267 (N_5267,N_3244,N_2787);
and U5268 (N_5268,N_1495,N_438);
nor U5269 (N_5269,N_192,N_1668);
or U5270 (N_5270,N_861,N_3704);
and U5271 (N_5271,N_3851,N_3836);
and U5272 (N_5272,N_389,N_3742);
xnor U5273 (N_5273,N_2278,N_1762);
nor U5274 (N_5274,N_486,N_1167);
or U5275 (N_5275,N_383,N_1571);
nand U5276 (N_5276,N_696,N_3240);
nor U5277 (N_5277,N_3895,N_33);
or U5278 (N_5278,N_1677,N_1675);
nor U5279 (N_5279,N_1745,N_930);
or U5280 (N_5280,N_3744,N_878);
and U5281 (N_5281,N_148,N_169);
xnor U5282 (N_5282,N_585,N_1968);
and U5283 (N_5283,N_1366,N_3655);
or U5284 (N_5284,N_1,N_3243);
xnor U5285 (N_5285,N_2515,N_2054);
and U5286 (N_5286,N_809,N_3275);
and U5287 (N_5287,N_2878,N_3743);
xor U5288 (N_5288,N_3492,N_211);
and U5289 (N_5289,N_1964,N_3098);
nand U5290 (N_5290,N_2857,N_706);
and U5291 (N_5291,N_1233,N_3362);
nand U5292 (N_5292,N_3799,N_246);
nor U5293 (N_5293,N_1541,N_414);
nor U5294 (N_5294,N_1660,N_3054);
nor U5295 (N_5295,N_1570,N_599);
nor U5296 (N_5296,N_2330,N_3524);
xnor U5297 (N_5297,N_2325,N_3853);
and U5298 (N_5298,N_1319,N_637);
and U5299 (N_5299,N_767,N_2046);
or U5300 (N_5300,N_509,N_1825);
nor U5301 (N_5301,N_355,N_1465);
or U5302 (N_5302,N_1237,N_2089);
or U5303 (N_5303,N_1398,N_2097);
nand U5304 (N_5304,N_2852,N_719);
nand U5305 (N_5305,N_683,N_804);
and U5306 (N_5306,N_3949,N_2557);
and U5307 (N_5307,N_2276,N_1652);
and U5308 (N_5308,N_2874,N_3023);
or U5309 (N_5309,N_1771,N_27);
xnor U5310 (N_5310,N_3534,N_428);
nand U5311 (N_5311,N_1911,N_3724);
or U5312 (N_5312,N_3357,N_2987);
or U5313 (N_5313,N_764,N_3188);
nor U5314 (N_5314,N_1980,N_2449);
nor U5315 (N_5315,N_147,N_3074);
and U5316 (N_5316,N_2237,N_3484);
and U5317 (N_5317,N_716,N_3760);
or U5318 (N_5318,N_3792,N_1299);
or U5319 (N_5319,N_2086,N_7);
nor U5320 (N_5320,N_1297,N_3852);
nand U5321 (N_5321,N_2271,N_2478);
xor U5322 (N_5322,N_3604,N_623);
nor U5323 (N_5323,N_3936,N_149);
nand U5324 (N_5324,N_3553,N_2258);
nor U5325 (N_5325,N_1375,N_1399);
nand U5326 (N_5326,N_3274,N_1235);
or U5327 (N_5327,N_935,N_2983);
and U5328 (N_5328,N_2401,N_2963);
nor U5329 (N_5329,N_1412,N_3686);
and U5330 (N_5330,N_3999,N_1357);
xnor U5331 (N_5331,N_2242,N_3256);
and U5332 (N_5332,N_2887,N_1415);
nor U5333 (N_5333,N_3403,N_866);
nor U5334 (N_5334,N_1348,N_3690);
or U5335 (N_5335,N_498,N_1282);
xor U5336 (N_5336,N_1869,N_1421);
or U5337 (N_5337,N_2050,N_3346);
nor U5338 (N_5338,N_814,N_2010);
or U5339 (N_5339,N_3370,N_3924);
or U5340 (N_5340,N_1057,N_2044);
and U5341 (N_5341,N_3389,N_439);
nor U5342 (N_5342,N_3752,N_1039);
nor U5343 (N_5343,N_1218,N_1460);
nor U5344 (N_5344,N_3301,N_3447);
nor U5345 (N_5345,N_1486,N_1272);
nand U5346 (N_5346,N_2763,N_1244);
or U5347 (N_5347,N_1228,N_2908);
and U5348 (N_5348,N_3369,N_3224);
nor U5349 (N_5349,N_94,N_180);
xor U5350 (N_5350,N_493,N_2369);
nor U5351 (N_5351,N_3001,N_237);
xor U5352 (N_5352,N_3234,N_3777);
xor U5353 (N_5353,N_818,N_697);
nor U5354 (N_5354,N_726,N_2496);
nor U5355 (N_5355,N_3316,N_3061);
nand U5356 (N_5356,N_1385,N_3397);
nand U5357 (N_5357,N_806,N_3229);
xor U5358 (N_5358,N_1454,N_3391);
xor U5359 (N_5359,N_2269,N_522);
nor U5360 (N_5360,N_251,N_3253);
nand U5361 (N_5361,N_2117,N_1531);
or U5362 (N_5362,N_3729,N_1816);
nand U5363 (N_5363,N_2105,N_1765);
or U5364 (N_5364,N_1559,N_3681);
nand U5365 (N_5365,N_3581,N_794);
or U5366 (N_5366,N_838,N_3654);
xnor U5367 (N_5367,N_800,N_2154);
nand U5368 (N_5368,N_145,N_3453);
and U5369 (N_5369,N_108,N_973);
nor U5370 (N_5370,N_93,N_2083);
nor U5371 (N_5371,N_1437,N_542);
nand U5372 (N_5372,N_2943,N_1162);
and U5373 (N_5373,N_2705,N_1463);
or U5374 (N_5374,N_1953,N_125);
and U5375 (N_5375,N_3168,N_3788);
nor U5376 (N_5376,N_2465,N_3578);
nor U5377 (N_5377,N_4,N_2926);
xor U5378 (N_5378,N_3527,N_262);
nor U5379 (N_5379,N_900,N_3750);
xor U5380 (N_5380,N_3418,N_2279);
nor U5381 (N_5381,N_929,N_2537);
or U5382 (N_5382,N_363,N_448);
nand U5383 (N_5383,N_996,N_1445);
and U5384 (N_5384,N_2199,N_78);
or U5385 (N_5385,N_852,N_2250);
nor U5386 (N_5386,N_492,N_195);
nor U5387 (N_5387,N_3702,N_2497);
nand U5388 (N_5388,N_2448,N_1124);
nor U5389 (N_5389,N_2755,N_2591);
nor U5390 (N_5390,N_3115,N_2988);
xor U5391 (N_5391,N_2008,N_1341);
nand U5392 (N_5392,N_3970,N_3328);
or U5393 (N_5393,N_2463,N_3479);
or U5394 (N_5394,N_3586,N_311);
xnor U5395 (N_5395,N_2680,N_2925);
nor U5396 (N_5396,N_2136,N_876);
or U5397 (N_5397,N_511,N_1478);
xor U5398 (N_5398,N_1937,N_819);
nor U5399 (N_5399,N_3516,N_1595);
or U5400 (N_5400,N_3452,N_3780);
and U5401 (N_5401,N_3462,N_1186);
nor U5402 (N_5402,N_3424,N_1847);
or U5403 (N_5403,N_3609,N_1941);
or U5404 (N_5404,N_1356,N_979);
nand U5405 (N_5405,N_3387,N_6);
nand U5406 (N_5406,N_3177,N_3329);
and U5407 (N_5407,N_2865,N_883);
nand U5408 (N_5408,N_2663,N_3648);
xnor U5409 (N_5409,N_1981,N_2767);
or U5410 (N_5410,N_2011,N_1268);
nor U5411 (N_5411,N_1685,N_3153);
xor U5412 (N_5412,N_527,N_3018);
nor U5413 (N_5413,N_2664,N_871);
or U5414 (N_5414,N_2174,N_46);
or U5415 (N_5415,N_3571,N_621);
or U5416 (N_5416,N_3827,N_1044);
nand U5417 (N_5417,N_3808,N_1468);
or U5418 (N_5418,N_926,N_1512);
xnor U5419 (N_5419,N_1145,N_367);
or U5420 (N_5420,N_156,N_1518);
or U5421 (N_5421,N_3930,N_3223);
nor U5422 (N_5422,N_1718,N_1914);
xnor U5423 (N_5423,N_3269,N_3013);
and U5424 (N_5424,N_3401,N_1081);
nor U5425 (N_5425,N_1245,N_975);
and U5426 (N_5426,N_2678,N_3770);
xor U5427 (N_5427,N_2021,N_3371);
nand U5428 (N_5428,N_307,N_105);
and U5429 (N_5429,N_901,N_2576);
or U5430 (N_5430,N_1298,N_345);
xnor U5431 (N_5431,N_3778,N_911);
nor U5432 (N_5432,N_962,N_483);
xnor U5433 (N_5433,N_2445,N_2679);
and U5434 (N_5434,N_2507,N_3339);
xor U5435 (N_5435,N_3427,N_3812);
and U5436 (N_5436,N_2917,N_1778);
or U5437 (N_5437,N_2080,N_2499);
nor U5438 (N_5438,N_1342,N_3501);
nor U5439 (N_5439,N_1632,N_1063);
or U5440 (N_5440,N_3147,N_2894);
nand U5441 (N_5441,N_1605,N_2362);
or U5442 (N_5442,N_647,N_1001);
nor U5443 (N_5443,N_519,N_2573);
and U5444 (N_5444,N_1781,N_1805);
or U5445 (N_5445,N_3603,N_458);
xor U5446 (N_5446,N_1643,N_915);
or U5447 (N_5447,N_1491,N_2699);
or U5448 (N_5448,N_62,N_2356);
nor U5449 (N_5449,N_2344,N_1727);
and U5450 (N_5450,N_1516,N_3539);
or U5451 (N_5451,N_3958,N_2575);
or U5452 (N_5452,N_1705,N_3396);
nor U5453 (N_5453,N_3734,N_1989);
and U5454 (N_5454,N_3355,N_2652);
nor U5455 (N_5455,N_489,N_1363);
nand U5456 (N_5456,N_2306,N_2707);
or U5457 (N_5457,N_2492,N_1217);
nand U5458 (N_5458,N_3900,N_788);
xor U5459 (N_5459,N_687,N_1524);
or U5460 (N_5460,N_2676,N_3213);
and U5461 (N_5461,N_3565,N_912);
nand U5462 (N_5462,N_701,N_680);
nor U5463 (N_5463,N_366,N_653);
and U5464 (N_5464,N_1231,N_3869);
or U5465 (N_5465,N_850,N_1472);
and U5466 (N_5466,N_3359,N_1301);
and U5467 (N_5467,N_1016,N_2485);
nor U5468 (N_5468,N_2946,N_1784);
nand U5469 (N_5469,N_609,N_3901);
or U5470 (N_5470,N_3786,N_798);
xnor U5471 (N_5471,N_1239,N_2782);
xor U5472 (N_5472,N_981,N_2687);
nor U5473 (N_5473,N_3446,N_3363);
xnor U5474 (N_5474,N_666,N_2849);
nand U5475 (N_5475,N_1094,N_3057);
or U5476 (N_5476,N_2409,N_3829);
nor U5477 (N_5477,N_2155,N_2584);
nor U5478 (N_5478,N_329,N_3041);
xnor U5479 (N_5479,N_2672,N_393);
and U5480 (N_5480,N_1819,N_2129);
nand U5481 (N_5481,N_1177,N_2912);
nor U5482 (N_5482,N_117,N_1376);
or U5483 (N_5483,N_2379,N_2855);
and U5484 (N_5484,N_3203,N_941);
or U5485 (N_5485,N_3319,N_1786);
nor U5486 (N_5486,N_1809,N_1536);
and U5487 (N_5487,N_1700,N_1936);
nand U5488 (N_5488,N_3474,N_3130);
or U5489 (N_5489,N_2783,N_1737);
xor U5490 (N_5490,N_3086,N_2111);
and U5491 (N_5491,N_1768,N_1631);
or U5492 (N_5492,N_1951,N_124);
and U5493 (N_5493,N_3350,N_765);
xnor U5494 (N_5494,N_1205,N_617);
or U5495 (N_5495,N_553,N_1100);
and U5496 (N_5496,N_1223,N_2974);
or U5497 (N_5497,N_2006,N_784);
or U5498 (N_5498,N_3867,N_3892);
and U5499 (N_5499,N_2245,N_128);
or U5500 (N_5500,N_755,N_343);
xor U5501 (N_5501,N_1887,N_2711);
nor U5502 (N_5502,N_924,N_766);
nor U5503 (N_5503,N_118,N_733);
nand U5504 (N_5504,N_1877,N_3157);
nor U5505 (N_5505,N_1916,N_2022);
xnor U5506 (N_5506,N_2740,N_2588);
or U5507 (N_5507,N_1965,N_2461);
nand U5508 (N_5508,N_795,N_2854);
nor U5509 (N_5509,N_491,N_745);
and U5510 (N_5510,N_1800,N_884);
and U5511 (N_5511,N_2651,N_3584);
nor U5512 (N_5512,N_3343,N_1033);
nor U5513 (N_5513,N_3303,N_3107);
nand U5514 (N_5514,N_1915,N_811);
nor U5515 (N_5515,N_2760,N_198);
or U5516 (N_5516,N_1733,N_3082);
xnor U5517 (N_5517,N_1182,N_3448);
and U5518 (N_5518,N_112,N_3182);
nor U5519 (N_5519,N_3625,N_3717);
and U5520 (N_5520,N_2504,N_2500);
xor U5521 (N_5521,N_3855,N_418);
or U5522 (N_5522,N_2524,N_3066);
or U5523 (N_5523,N_601,N_2270);
nand U5524 (N_5524,N_1125,N_3864);
or U5525 (N_5525,N_26,N_1630);
xnor U5526 (N_5526,N_218,N_3103);
and U5527 (N_5527,N_1266,N_1056);
or U5528 (N_5528,N_3657,N_1992);
nand U5529 (N_5529,N_2100,N_3783);
or U5530 (N_5530,N_711,N_2298);
nor U5531 (N_5531,N_3854,N_3377);
nand U5532 (N_5532,N_1169,N_3676);
nor U5533 (N_5533,N_3460,N_252);
and U5534 (N_5534,N_3588,N_1198);
and U5535 (N_5535,N_2391,N_2593);
or U5536 (N_5536,N_3730,N_2162);
or U5537 (N_5537,N_1059,N_919);
nand U5538 (N_5538,N_184,N_2079);
nor U5539 (N_5539,N_3822,N_1742);
xor U5540 (N_5540,N_3926,N_2958);
nand U5541 (N_5541,N_2386,N_2896);
xor U5542 (N_5542,N_1091,N_1328);
or U5543 (N_5543,N_2293,N_2981);
nand U5544 (N_5544,N_1910,N_2213);
nand U5545 (N_5545,N_571,N_1204);
or U5546 (N_5546,N_98,N_79);
or U5547 (N_5547,N_3400,N_123);
nor U5548 (N_5548,N_744,N_189);
nand U5549 (N_5549,N_3226,N_2628);
and U5550 (N_5550,N_2831,N_882);
and U5551 (N_5551,N_1870,N_115);
or U5552 (N_5552,N_3960,N_42);
xnor U5553 (N_5553,N_638,N_2433);
xnor U5554 (N_5554,N_333,N_3894);
nand U5555 (N_5555,N_1545,N_36);
nor U5556 (N_5556,N_1799,N_187);
xor U5557 (N_5557,N_927,N_537);
and U5558 (N_5558,N_431,N_1021);
or U5559 (N_5559,N_3877,N_2166);
nand U5560 (N_5560,N_1646,N_2103);
and U5561 (N_5561,N_1101,N_1694);
or U5562 (N_5562,N_3310,N_1043);
xnor U5563 (N_5563,N_2033,N_2216);
and U5564 (N_5564,N_1388,N_3268);
or U5565 (N_5565,N_1358,N_3638);
xnor U5566 (N_5566,N_686,N_3731);
xnor U5567 (N_5567,N_1692,N_1340);
nand U5568 (N_5568,N_593,N_844);
xor U5569 (N_5569,N_3634,N_1942);
or U5570 (N_5570,N_672,N_1904);
or U5571 (N_5571,N_1982,N_2539);
nor U5572 (N_5572,N_8,N_3790);
nor U5573 (N_5573,N_217,N_136);
nand U5574 (N_5574,N_3935,N_2019);
or U5575 (N_5575,N_1588,N_1789);
xor U5576 (N_5576,N_203,N_2759);
nand U5577 (N_5577,N_854,N_3967);
xor U5578 (N_5578,N_485,N_2077);
and U5579 (N_5579,N_171,N_348);
nor U5580 (N_5580,N_1513,N_857);
nor U5581 (N_5581,N_1154,N_2309);
or U5582 (N_5582,N_3428,N_2198);
or U5583 (N_5583,N_3022,N_1017);
nand U5584 (N_5584,N_2734,N_2665);
xor U5585 (N_5585,N_3142,N_1160);
or U5586 (N_5586,N_2745,N_2969);
nor U5587 (N_5587,N_1110,N_3597);
nand U5588 (N_5588,N_2462,N_2414);
or U5589 (N_5589,N_309,N_3102);
and U5590 (N_5590,N_1671,N_2342);
or U5591 (N_5591,N_548,N_546);
or U5592 (N_5592,N_2413,N_435);
nand U5593 (N_5593,N_676,N_24);
nand U5594 (N_5594,N_2889,N_2806);
or U5595 (N_5595,N_1064,N_1055);
nor U5596 (N_5596,N_3992,N_782);
and U5597 (N_5597,N_3660,N_3003);
and U5598 (N_5598,N_3811,N_514);
xnor U5599 (N_5599,N_2535,N_3847);
and U5600 (N_5600,N_2646,N_2239);
nor U5601 (N_5601,N_862,N_874);
and U5602 (N_5602,N_359,N_1543);
and U5603 (N_5603,N_1246,N_104);
nand U5604 (N_5604,N_1554,N_3839);
or U5605 (N_5605,N_3317,N_1928);
xnor U5606 (N_5606,N_293,N_1408);
nand U5607 (N_5607,N_3530,N_1848);
or U5608 (N_5608,N_501,N_528);
nor U5609 (N_5609,N_1400,N_1673);
nor U5610 (N_5610,N_3607,N_562);
or U5611 (N_5611,N_2907,N_1157);
and U5612 (N_5612,N_3482,N_1764);
or U5613 (N_5613,N_273,N_3264);
xnor U5614 (N_5614,N_29,N_1292);
nand U5615 (N_5615,N_41,N_3932);
or U5616 (N_5616,N_2343,N_1757);
nand U5617 (N_5617,N_2947,N_2995);
nor U5618 (N_5618,N_3202,N_2126);
or U5619 (N_5619,N_1963,N_1396);
nand U5620 (N_5620,N_92,N_881);
nor U5621 (N_5621,N_95,N_500);
nor U5622 (N_5622,N_3834,N_682);
or U5623 (N_5623,N_3529,N_3768);
nand U5624 (N_5624,N_1434,N_756);
nand U5625 (N_5625,N_2936,N_2868);
or U5626 (N_5626,N_1115,N_2766);
nand U5627 (N_5627,N_3378,N_3144);
nor U5628 (N_5628,N_3612,N_2407);
or U5629 (N_5629,N_3974,N_1032);
and U5630 (N_5630,N_568,N_1574);
or U5631 (N_5631,N_2084,N_432);
nor U5632 (N_5632,N_1423,N_2884);
and U5633 (N_5633,N_2570,N_2552);
nand U5634 (N_5634,N_2002,N_3738);
or U5635 (N_5635,N_662,N_1256);
and U5636 (N_5636,N_496,N_2924);
or U5637 (N_5637,N_1889,N_1011);
or U5638 (N_5638,N_2548,N_1926);
or U5639 (N_5639,N_2918,N_375);
nor U5640 (N_5640,N_3263,N_3859);
or U5641 (N_5641,N_1409,N_3469);
xor U5642 (N_5642,N_2319,N_656);
and U5643 (N_5643,N_2146,N_2108);
nand U5644 (N_5644,N_1161,N_1687);
or U5645 (N_5645,N_747,N_895);
nand U5646 (N_5646,N_1051,N_3559);
nor U5647 (N_5647,N_1047,N_2637);
and U5648 (N_5648,N_1770,N_3863);
and U5649 (N_5649,N_1492,N_643);
nor U5650 (N_5650,N_677,N_689);
xnor U5651 (N_5651,N_1721,N_3230);
and U5652 (N_5652,N_1464,N_3221);
xnor U5653 (N_5653,N_1067,N_1430);
and U5654 (N_5654,N_3850,N_2115);
nor U5655 (N_5655,N_3047,N_1158);
and U5656 (N_5656,N_2645,N_1620);
and U5657 (N_5657,N_1500,N_1880);
nand U5658 (N_5658,N_971,N_441);
xnor U5659 (N_5659,N_2055,N_2756);
xnor U5660 (N_5660,N_1566,N_2475);
nor U5661 (N_5661,N_602,N_2885);
nand U5662 (N_5662,N_73,N_904);
or U5663 (N_5663,N_450,N_2092);
or U5664 (N_5664,N_182,N_2392);
nand U5665 (N_5665,N_1078,N_3000);
and U5666 (N_5666,N_2566,N_394);
and U5667 (N_5667,N_1732,N_2365);
and U5668 (N_5668,N_1978,N_1960);
or U5669 (N_5669,N_2317,N_3599);
and U5670 (N_5670,N_504,N_860);
xor U5671 (N_5671,N_313,N_3920);
and U5672 (N_5672,N_2744,N_2813);
nand U5673 (N_5673,N_213,N_2635);
xnor U5674 (N_5674,N_1046,N_1945);
xnor U5675 (N_5675,N_1022,N_3879);
xor U5676 (N_5676,N_2877,N_3382);
nand U5677 (N_5677,N_908,N_2517);
nand U5678 (N_5678,N_3444,N_3342);
nor U5679 (N_5679,N_3149,N_3582);
nor U5680 (N_5680,N_2406,N_524);
and U5681 (N_5681,N_2725,N_2785);
nand U5682 (N_5682,N_1735,N_810);
and U5683 (N_5683,N_2404,N_3246);
and U5684 (N_5684,N_1035,N_2512);
and U5685 (N_5685,N_720,N_3027);
or U5686 (N_5686,N_1221,N_133);
xor U5687 (N_5687,N_2695,N_2218);
nand U5688 (N_5688,N_1795,N_77);
or U5689 (N_5689,N_1790,N_2283);
xor U5690 (N_5690,N_3826,N_1026);
and U5691 (N_5691,N_2175,N_3404);
or U5692 (N_5692,N_3089,N_3216);
xor U5693 (N_5693,N_3763,N_3104);
nand U5694 (N_5694,N_539,N_886);
xnor U5695 (N_5695,N_2251,N_2396);
xor U5696 (N_5696,N_535,N_2583);
nand U5697 (N_5697,N_292,N_1306);
and U5698 (N_5698,N_520,N_3296);
xor U5699 (N_5699,N_827,N_442);
and U5700 (N_5700,N_37,N_1538);
xor U5701 (N_5701,N_3797,N_3101);
nand U5702 (N_5702,N_2038,N_459);
nor U5703 (N_5703,N_3038,N_3004);
or U5704 (N_5704,N_3722,N_2833);
and U5705 (N_5705,N_1499,N_3993);
or U5706 (N_5706,N_2193,N_2494);
or U5707 (N_5707,N_821,N_1290);
and U5708 (N_5708,N_3083,N_3540);
and U5709 (N_5709,N_2528,N_416);
and U5710 (N_5710,N_2697,N_3550);
xnor U5711 (N_5711,N_2592,N_2999);
or U5712 (N_5712,N_3745,N_114);
nor U5713 (N_5713,N_1615,N_969);
and U5714 (N_5714,N_3437,N_1345);
or U5715 (N_5715,N_3554,N_3483);
xnor U5716 (N_5716,N_754,N_600);
xor U5717 (N_5717,N_1920,N_1580);
xor U5718 (N_5718,N_1012,N_2447);
nand U5719 (N_5719,N_3059,N_805);
nor U5720 (N_5720,N_1373,N_3225);
nor U5721 (N_5721,N_2968,N_2284);
xor U5722 (N_5722,N_563,N_2577);
or U5723 (N_5723,N_1286,N_1658);
xor U5724 (N_5724,N_379,N_1527);
xnor U5725 (N_5725,N_3756,N_2875);
nand U5726 (N_5726,N_3909,N_1240);
nor U5727 (N_5727,N_740,N_3485);
nor U5728 (N_5728,N_3134,N_893);
or U5729 (N_5729,N_3997,N_505);
or U5730 (N_5730,N_1706,N_2994);
nand U5731 (N_5731,N_737,N_3940);
or U5732 (N_5732,N_1650,N_1864);
and U5733 (N_5733,N_113,N_1405);
or U5734 (N_5734,N_3184,N_1532);
and U5735 (N_5735,N_2794,N_344);
nor U5736 (N_5736,N_1469,N_3938);
nor U5737 (N_5737,N_1193,N_3011);
xor U5738 (N_5738,N_1443,N_2555);
nand U5739 (N_5739,N_595,N_1281);
or U5740 (N_5740,N_550,N_2405);
and U5741 (N_5741,N_101,N_3067);
nand U5742 (N_5742,N_3285,N_2842);
nand U5743 (N_5743,N_3562,N_1826);
nand U5744 (N_5744,N_575,N_1105);
nor U5745 (N_5745,N_2114,N_3336);
nand U5746 (N_5746,N_2590,N_557);
nand U5747 (N_5747,N_2432,N_679);
nand U5748 (N_5748,N_2459,N_3239);
and U5749 (N_5749,N_1302,N_1082);
and U5750 (N_5750,N_303,N_350);
nor U5751 (N_5751,N_1418,N_1071);
or U5752 (N_5752,N_596,N_1255);
xor U5753 (N_5753,N_1108,N_1661);
xnor U5754 (N_5754,N_2291,N_3615);
nand U5755 (N_5755,N_1811,N_1954);
nor U5756 (N_5756,N_1863,N_1779);
nor U5757 (N_5757,N_639,N_3694);
or U5758 (N_5758,N_1207,N_3135);
nand U5759 (N_5759,N_3468,N_2308);
and U5760 (N_5760,N_2602,N_3643);
and U5761 (N_5761,N_488,N_3312);
xnor U5762 (N_5762,N_2195,N_2797);
or U5763 (N_5763,N_757,N_2819);
and U5764 (N_5764,N_717,N_2923);
nand U5765 (N_5765,N_2201,N_2366);
xnor U5766 (N_5766,N_3795,N_1196);
or U5767 (N_5767,N_2541,N_2224);
or U5768 (N_5768,N_3323,N_2152);
xnor U5769 (N_5769,N_2533,N_25);
nand U5770 (N_5770,N_3178,N_3601);
xnor U5771 (N_5771,N_2329,N_3732);
nor U5772 (N_5772,N_1841,N_167);
nand U5773 (N_5773,N_994,N_1773);
and U5774 (N_5774,N_56,N_1111);
or U5775 (N_5775,N_1109,N_858);
nand U5776 (N_5776,N_2219,N_2395);
or U5777 (N_5777,N_1020,N_1130);
and U5778 (N_5778,N_1141,N_1310);
nor U5779 (N_5779,N_2142,N_3019);
nand U5780 (N_5780,N_3036,N_1892);
and U5781 (N_5781,N_3610,N_3204);
or U5782 (N_5782,N_462,N_3598);
nand U5783 (N_5783,N_1882,N_1686);
xor U5784 (N_5784,N_2836,N_3496);
xnor U5785 (N_5785,N_2081,N_891);
or U5786 (N_5786,N_2210,N_1242);
nor U5787 (N_5787,N_3942,N_2318);
and U5788 (N_5788,N_2453,N_2380);
nor U5789 (N_5789,N_2277,N_3663);
or U5790 (N_5790,N_2032,N_3457);
nor U5791 (N_5791,N_3956,N_89);
nand U5792 (N_5792,N_799,N_2169);
nand U5793 (N_5793,N_2324,N_2424);
and U5794 (N_5794,N_1946,N_1912);
nor U5795 (N_5795,N_1817,N_780);
nand U5796 (N_5796,N_1556,N_3351);
or U5797 (N_5797,N_837,N_560);
and U5798 (N_5798,N_694,N_1337);
nor U5799 (N_5799,N_362,N_1106);
xnor U5800 (N_5800,N_1159,N_3406);
or U5801 (N_5801,N_2802,N_3176);
and U5802 (N_5802,N_1670,N_2827);
and U5803 (N_5803,N_1831,N_402);
nor U5804 (N_5804,N_2701,N_3338);
nor U5805 (N_5805,N_1197,N_2953);
nand U5806 (N_5806,N_2161,N_2388);
and U5807 (N_5807,N_1254,N_2670);
xnor U5808 (N_5808,N_3769,N_2285);
xor U5809 (N_5809,N_157,N_2446);
nand U5810 (N_5810,N_2568,N_1533);
or U5811 (N_5811,N_1222,N_1087);
xor U5812 (N_5812,N_2227,N_3293);
and U5813 (N_5813,N_357,N_270);
and U5814 (N_5814,N_2075,N_1865);
nand U5815 (N_5815,N_614,N_3170);
nand U5816 (N_5816,N_2556,N_3155);
xor U5817 (N_5817,N_1905,N_3566);
and U5818 (N_5818,N_570,N_2721);
and U5819 (N_5819,N_2825,N_61);
xor U5820 (N_5820,N_1872,N_3884);
or U5821 (N_5821,N_1117,N_2935);
and U5822 (N_5822,N_3247,N_2686);
xnor U5823 (N_5823,N_3233,N_300);
nand U5824 (N_5824,N_1494,N_340);
xor U5825 (N_5825,N_1876,N_918);
nor U5826 (N_5826,N_820,N_257);
nor U5827 (N_5827,N_3032,N_71);
or U5828 (N_5828,N_738,N_1353);
or U5829 (N_5829,N_1842,N_3380);
nand U5830 (N_5830,N_2390,N_2985);
nor U5831 (N_5831,N_234,N_3143);
or U5832 (N_5832,N_1350,N_752);
or U5833 (N_5833,N_712,N_284);
or U5834 (N_5834,N_188,N_2254);
nand U5835 (N_5835,N_2179,N_2417);
nor U5836 (N_5836,N_452,N_3161);
or U5837 (N_5837,N_1209,N_2387);
nand U5838 (N_5838,N_790,N_1738);
nand U5839 (N_5839,N_2125,N_3741);
and U5840 (N_5840,N_1170,N_899);
nand U5841 (N_5841,N_1446,N_3639);
nor U5842 (N_5842,N_2243,N_3541);
nand U5843 (N_5843,N_2630,N_3984);
and U5844 (N_5844,N_2906,N_1575);
or U5845 (N_5845,N_3254,N_1683);
and U5846 (N_5846,N_2450,N_2506);
nand U5847 (N_5847,N_230,N_3989);
nand U5848 (N_5848,N_3430,N_3782);
and U5849 (N_5849,N_110,N_1189);
xor U5850 (N_5850,N_2805,N_1027);
nor U5851 (N_5851,N_3099,N_1986);
nor U5852 (N_5852,N_3386,N_1684);
nor U5853 (N_5853,N_2867,N_1979);
xnor U5854 (N_5854,N_332,N_3614);
nand U5855 (N_5855,N_2803,N_2015);
and U5856 (N_5856,N_3136,N_422);
xor U5857 (N_5857,N_3606,N_2383);
or U5858 (N_5858,N_3608,N_1715);
xor U5859 (N_5859,N_3008,N_3575);
and U5860 (N_5860,N_3897,N_3219);
and U5861 (N_5861,N_2145,N_3069);
nor U5862 (N_5862,N_3570,N_3514);
and U5863 (N_5863,N_22,N_1829);
nor U5864 (N_5864,N_847,N_3641);
nand U5865 (N_5865,N_221,N_2735);
or U5866 (N_5866,N_2703,N_476);
nand U5867 (N_5867,N_667,N_2671);
or U5868 (N_5868,N_2353,N_1031);
nand U5869 (N_5869,N_3330,N_1542);
or U5870 (N_5870,N_1793,N_2262);
or U5871 (N_5871,N_1333,N_3415);
nand U5872 (N_5872,N_2694,N_3180);
nor U5873 (N_5873,N_2791,N_119);
nor U5874 (N_5874,N_529,N_2970);
nand U5875 (N_5875,N_3890,N_965);
and U5876 (N_5876,N_739,N_1836);
xnor U5877 (N_5877,N_3787,N_833);
xnor U5878 (N_5878,N_1165,N_2253);
xor U5879 (N_5879,N_3150,N_743);
nand U5880 (N_5880,N_645,N_1183);
and U5881 (N_5881,N_1967,N_3931);
nand U5882 (N_5882,N_1211,N_2786);
and U5883 (N_5883,N_2493,N_2750);
and U5884 (N_5884,N_3652,N_3043);
nand U5885 (N_5885,N_1724,N_1401);
or U5886 (N_5886,N_2845,N_3193);
nor U5887 (N_5887,N_2736,N_793);
nand U5888 (N_5888,N_3145,N_3210);
or U5889 (N_5889,N_2094,N_1168);
or U5890 (N_5890,N_3108,N_121);
and U5891 (N_5891,N_330,N_3461);
nor U5892 (N_5892,N_179,N_153);
and U5893 (N_5893,N_2569,N_2017);
xnor U5894 (N_5894,N_2945,N_1555);
or U5895 (N_5895,N_122,N_1264);
xnor U5896 (N_5896,N_86,N_3700);
xor U5897 (N_5897,N_1629,N_1030);
or U5898 (N_5898,N_3489,N_2641);
nor U5899 (N_5899,N_2164,N_1126);
nand U5900 (N_5900,N_1134,N_1999);
and U5901 (N_5901,N_160,N_3375);
or U5902 (N_5902,N_40,N_43);
nor U5903 (N_5903,N_1215,N_3698);
nand U5904 (N_5904,N_1155,N_2364);
nand U5905 (N_5905,N_544,N_327);
or U5906 (N_5906,N_1428,N_942);
nand U5907 (N_5907,N_3076,N_1791);
xor U5908 (N_5908,N_3395,N_3862);
nor U5909 (N_5909,N_2244,N_2326);
xnor U5910 (N_5910,N_1897,N_1148);
xor U5911 (N_5911,N_587,N_1810);
or U5912 (N_5912,N_2180,N_1386);
or U5913 (N_5913,N_1596,N_2368);
nand U5914 (N_5914,N_475,N_2397);
or U5915 (N_5915,N_2521,N_49);
nand U5916 (N_5916,N_1758,N_3856);
nor U5917 (N_5917,N_139,N_2034);
or U5918 (N_5918,N_3871,N_1049);
xor U5919 (N_5919,N_196,N_200);
and U5920 (N_5920,N_1929,N_3907);
xnor U5921 (N_5921,N_2186,N_1300);
nor U5922 (N_5922,N_2757,N_1439);
xnor U5923 (N_5923,N_525,N_202);
and U5924 (N_5924,N_3995,N_3467);
xor U5925 (N_5925,N_1362,N_3651);
nand U5926 (N_5926,N_2214,N_961);
nand U5927 (N_5927,N_3111,N_2822);
xor U5928 (N_5928,N_1200,N_3789);
nand U5929 (N_5929,N_390,N_517);
and U5930 (N_5930,N_2795,N_3765);
xor U5931 (N_5931,N_3077,N_3804);
or U5932 (N_5932,N_235,N_944);
and U5933 (N_5933,N_1654,N_796);
or U5934 (N_5934,N_1311,N_1413);
and U5935 (N_5935,N_992,N_1241);
or U5936 (N_5936,N_1921,N_368);
xor U5937 (N_5937,N_2620,N_3891);
and U5938 (N_5938,N_1659,N_1098);
or U5939 (N_5939,N_1924,N_2682);
nor U5940 (N_5940,N_3861,N_3633);
or U5941 (N_5941,N_2715,N_1849);
xor U5942 (N_5942,N_1372,N_3875);
xnor U5943 (N_5943,N_3837,N_317);
nor U5944 (N_5944,N_3872,N_506);
or U5945 (N_5945,N_3896,N_470);
or U5946 (N_5946,N_3499,N_2429);
and U5947 (N_5947,N_482,N_925);
xnor U5948 (N_5948,N_44,N_2455);
or U5949 (N_5949,N_3072,N_564);
nand U5950 (N_5950,N_3398,N_370);
or U5951 (N_5951,N_2685,N_2128);
and U5952 (N_5952,N_1224,N_2531);
and U5953 (N_5953,N_1656,N_2818);
or U5954 (N_5954,N_2185,N_3774);
nor U5955 (N_5955,N_1748,N_3806);
or U5956 (N_5956,N_2967,N_802);
and U5957 (N_5957,N_354,N_495);
or U5958 (N_5958,N_2530,N_1583);
xnor U5959 (N_5959,N_3162,N_3577);
nand U5960 (N_5960,N_2207,N_3181);
nor U5961 (N_5961,N_1441,N_2112);
and U5962 (N_5962,N_2928,N_241);
xor U5963 (N_5963,N_433,N_2681);
xor U5964 (N_5964,N_3040,N_2093);
or U5965 (N_5965,N_2966,N_2674);
and U5966 (N_5966,N_227,N_1879);
and U5967 (N_5967,N_3205,N_650);
and U5968 (N_5968,N_326,N_846);
or U5969 (N_5969,N_2471,N_2581);
nor U5970 (N_5970,N_2460,N_3814);
nand U5971 (N_5971,N_2598,N_3519);
nand U5972 (N_5972,N_1420,N_1788);
and U5973 (N_5973,N_892,N_1749);
xnor U5974 (N_5974,N_842,N_2222);
and U5975 (N_5975,N_3078,N_2221);
nor U5976 (N_5976,N_3628,N_1970);
xor U5977 (N_5977,N_323,N_1906);
nand U5978 (N_5978,N_2378,N_1676);
nand U5979 (N_5979,N_2123,N_3617);
nor U5980 (N_5980,N_1284,N_1127);
xor U5981 (N_5981,N_3979,N_700);
nor U5982 (N_5982,N_302,N_3159);
nand U5983 (N_5983,N_312,N_2481);
nor U5984 (N_5984,N_3366,N_615);
nor U5985 (N_5985,N_1053,N_3190);
nand U5986 (N_5986,N_1635,N_1374);
xor U5987 (N_5987,N_3968,N_3354);
nor U5988 (N_5988,N_1537,N_2275);
or U5989 (N_5989,N_1617,N_281);
xnor U5990 (N_5990,N_1164,N_3560);
or U5991 (N_5991,N_2477,N_425);
or U5992 (N_5992,N_3944,N_3016);
xnor U5993 (N_5993,N_2621,N_2762);
nand U5994 (N_5994,N_1691,N_3033);
and U5995 (N_5995,N_2883,N_34);
and U5996 (N_5996,N_2749,N_2301);
xor U5997 (N_5997,N_1440,N_3973);
nor U5998 (N_5998,N_1414,N_3548);
and U5999 (N_5999,N_1219,N_2643);
or U6000 (N_6000,N_563,N_1401);
and U6001 (N_6001,N_2211,N_2262);
nor U6002 (N_6002,N_3040,N_1715);
or U6003 (N_6003,N_3194,N_3407);
and U6004 (N_6004,N_2465,N_3973);
nor U6005 (N_6005,N_3764,N_315);
xor U6006 (N_6006,N_192,N_664);
xnor U6007 (N_6007,N_763,N_2864);
nand U6008 (N_6008,N_1489,N_2298);
and U6009 (N_6009,N_3682,N_1695);
xor U6010 (N_6010,N_3475,N_1814);
nor U6011 (N_6011,N_2777,N_504);
and U6012 (N_6012,N_2547,N_3642);
xor U6013 (N_6013,N_3682,N_2592);
xnor U6014 (N_6014,N_294,N_3371);
nand U6015 (N_6015,N_902,N_1826);
nor U6016 (N_6016,N_3107,N_3332);
nand U6017 (N_6017,N_1351,N_579);
and U6018 (N_6018,N_2943,N_1715);
xnor U6019 (N_6019,N_3180,N_2408);
nand U6020 (N_6020,N_553,N_3671);
nand U6021 (N_6021,N_2046,N_1308);
nor U6022 (N_6022,N_3055,N_343);
and U6023 (N_6023,N_819,N_3956);
xor U6024 (N_6024,N_3350,N_188);
nand U6025 (N_6025,N_1190,N_1011);
and U6026 (N_6026,N_2395,N_1511);
nor U6027 (N_6027,N_1669,N_3270);
nand U6028 (N_6028,N_3785,N_3078);
nor U6029 (N_6029,N_1701,N_2364);
nand U6030 (N_6030,N_1888,N_741);
xor U6031 (N_6031,N_2826,N_2383);
xnor U6032 (N_6032,N_852,N_3270);
xor U6033 (N_6033,N_716,N_3800);
and U6034 (N_6034,N_3314,N_1191);
nand U6035 (N_6035,N_1344,N_2897);
nand U6036 (N_6036,N_728,N_32);
nor U6037 (N_6037,N_3658,N_757);
nand U6038 (N_6038,N_687,N_3837);
or U6039 (N_6039,N_3707,N_3189);
or U6040 (N_6040,N_268,N_2423);
nand U6041 (N_6041,N_2525,N_2013);
and U6042 (N_6042,N_1188,N_2640);
or U6043 (N_6043,N_1009,N_187);
nand U6044 (N_6044,N_2196,N_1698);
and U6045 (N_6045,N_2509,N_2409);
and U6046 (N_6046,N_3419,N_2356);
xnor U6047 (N_6047,N_1980,N_2337);
xnor U6048 (N_6048,N_645,N_2672);
or U6049 (N_6049,N_1807,N_163);
nor U6050 (N_6050,N_3031,N_3065);
and U6051 (N_6051,N_2350,N_1942);
nand U6052 (N_6052,N_3738,N_2422);
and U6053 (N_6053,N_1636,N_2238);
nor U6054 (N_6054,N_2969,N_1955);
and U6055 (N_6055,N_936,N_3831);
nand U6056 (N_6056,N_1059,N_3180);
or U6057 (N_6057,N_3576,N_394);
and U6058 (N_6058,N_2263,N_1865);
and U6059 (N_6059,N_2923,N_1405);
nand U6060 (N_6060,N_3470,N_85);
or U6061 (N_6061,N_2905,N_3541);
or U6062 (N_6062,N_3505,N_1341);
nand U6063 (N_6063,N_3085,N_3649);
nor U6064 (N_6064,N_2223,N_2061);
nor U6065 (N_6065,N_1563,N_1715);
nor U6066 (N_6066,N_2805,N_1295);
xor U6067 (N_6067,N_2537,N_3545);
nor U6068 (N_6068,N_3744,N_3436);
xnor U6069 (N_6069,N_245,N_1250);
and U6070 (N_6070,N_3832,N_3764);
and U6071 (N_6071,N_2532,N_3046);
or U6072 (N_6072,N_3995,N_2502);
or U6073 (N_6073,N_1491,N_3126);
xnor U6074 (N_6074,N_813,N_54);
nand U6075 (N_6075,N_1923,N_3952);
nor U6076 (N_6076,N_3739,N_3342);
xor U6077 (N_6077,N_1878,N_2691);
and U6078 (N_6078,N_1875,N_858);
xor U6079 (N_6079,N_399,N_1556);
xnor U6080 (N_6080,N_2146,N_3869);
or U6081 (N_6081,N_2450,N_32);
and U6082 (N_6082,N_3723,N_2417);
nand U6083 (N_6083,N_485,N_1752);
xnor U6084 (N_6084,N_3501,N_1892);
or U6085 (N_6085,N_2456,N_3216);
xor U6086 (N_6086,N_631,N_1390);
nor U6087 (N_6087,N_1110,N_1900);
or U6088 (N_6088,N_939,N_2775);
and U6089 (N_6089,N_1736,N_3773);
and U6090 (N_6090,N_3224,N_767);
and U6091 (N_6091,N_2612,N_2108);
nand U6092 (N_6092,N_2021,N_97);
nand U6093 (N_6093,N_1770,N_3599);
nor U6094 (N_6094,N_1621,N_1572);
xnor U6095 (N_6095,N_2914,N_457);
and U6096 (N_6096,N_2042,N_1601);
nor U6097 (N_6097,N_3401,N_232);
and U6098 (N_6098,N_32,N_719);
xor U6099 (N_6099,N_1452,N_3768);
and U6100 (N_6100,N_2419,N_1493);
nand U6101 (N_6101,N_2000,N_994);
or U6102 (N_6102,N_1194,N_1164);
or U6103 (N_6103,N_441,N_3998);
nand U6104 (N_6104,N_1111,N_1303);
xnor U6105 (N_6105,N_107,N_1682);
nor U6106 (N_6106,N_2015,N_2592);
nand U6107 (N_6107,N_3027,N_1508);
and U6108 (N_6108,N_513,N_224);
or U6109 (N_6109,N_1760,N_208);
nand U6110 (N_6110,N_2097,N_179);
nor U6111 (N_6111,N_2033,N_727);
nand U6112 (N_6112,N_3545,N_3380);
and U6113 (N_6113,N_1277,N_2578);
or U6114 (N_6114,N_590,N_2235);
xor U6115 (N_6115,N_3847,N_547);
and U6116 (N_6116,N_3964,N_3686);
nor U6117 (N_6117,N_2623,N_873);
and U6118 (N_6118,N_2810,N_3601);
xnor U6119 (N_6119,N_199,N_2733);
nor U6120 (N_6120,N_1462,N_3655);
nor U6121 (N_6121,N_1191,N_892);
nand U6122 (N_6122,N_2653,N_486);
nor U6123 (N_6123,N_2618,N_1305);
xnor U6124 (N_6124,N_3827,N_2553);
xor U6125 (N_6125,N_413,N_3199);
or U6126 (N_6126,N_212,N_3972);
or U6127 (N_6127,N_1120,N_1193);
and U6128 (N_6128,N_2616,N_901);
and U6129 (N_6129,N_3146,N_840);
or U6130 (N_6130,N_2474,N_1422);
nor U6131 (N_6131,N_3823,N_2358);
or U6132 (N_6132,N_3420,N_3170);
and U6133 (N_6133,N_133,N_3554);
nand U6134 (N_6134,N_292,N_3630);
xnor U6135 (N_6135,N_1466,N_446);
or U6136 (N_6136,N_3321,N_2216);
and U6137 (N_6137,N_1481,N_2847);
or U6138 (N_6138,N_3222,N_1495);
xor U6139 (N_6139,N_813,N_740);
nand U6140 (N_6140,N_3,N_3577);
xnor U6141 (N_6141,N_498,N_3628);
nor U6142 (N_6142,N_2469,N_1879);
xnor U6143 (N_6143,N_129,N_3349);
nand U6144 (N_6144,N_2638,N_48);
nand U6145 (N_6145,N_3992,N_2554);
xnor U6146 (N_6146,N_2764,N_1054);
nand U6147 (N_6147,N_316,N_86);
and U6148 (N_6148,N_2034,N_3010);
and U6149 (N_6149,N_3672,N_659);
xor U6150 (N_6150,N_3823,N_250);
or U6151 (N_6151,N_3646,N_3576);
nand U6152 (N_6152,N_975,N_149);
xor U6153 (N_6153,N_2383,N_3988);
nor U6154 (N_6154,N_1585,N_1651);
and U6155 (N_6155,N_926,N_519);
nand U6156 (N_6156,N_3621,N_1012);
and U6157 (N_6157,N_2646,N_2434);
xnor U6158 (N_6158,N_3148,N_1983);
or U6159 (N_6159,N_3207,N_701);
xor U6160 (N_6160,N_1121,N_2451);
and U6161 (N_6161,N_3379,N_3633);
xnor U6162 (N_6162,N_125,N_1432);
xnor U6163 (N_6163,N_1263,N_3588);
nand U6164 (N_6164,N_221,N_3018);
nand U6165 (N_6165,N_863,N_1313);
xor U6166 (N_6166,N_1376,N_2460);
nor U6167 (N_6167,N_768,N_3071);
xnor U6168 (N_6168,N_2278,N_1352);
nand U6169 (N_6169,N_2984,N_3771);
and U6170 (N_6170,N_2142,N_3028);
nand U6171 (N_6171,N_2258,N_2912);
and U6172 (N_6172,N_2882,N_2165);
nor U6173 (N_6173,N_422,N_2254);
or U6174 (N_6174,N_723,N_658);
and U6175 (N_6175,N_3690,N_2961);
nand U6176 (N_6176,N_2089,N_568);
or U6177 (N_6177,N_789,N_3075);
xor U6178 (N_6178,N_1666,N_805);
nand U6179 (N_6179,N_2666,N_2170);
or U6180 (N_6180,N_392,N_1023);
and U6181 (N_6181,N_40,N_1260);
xnor U6182 (N_6182,N_303,N_3295);
nor U6183 (N_6183,N_3514,N_1556);
nor U6184 (N_6184,N_161,N_1734);
or U6185 (N_6185,N_1989,N_1991);
xor U6186 (N_6186,N_525,N_579);
nor U6187 (N_6187,N_305,N_3064);
and U6188 (N_6188,N_2003,N_529);
nand U6189 (N_6189,N_2507,N_2711);
or U6190 (N_6190,N_1632,N_63);
nand U6191 (N_6191,N_3467,N_1069);
or U6192 (N_6192,N_664,N_727);
nand U6193 (N_6193,N_1122,N_3509);
nand U6194 (N_6194,N_2975,N_3497);
or U6195 (N_6195,N_1117,N_419);
xor U6196 (N_6196,N_3361,N_2798);
xnor U6197 (N_6197,N_1292,N_1259);
or U6198 (N_6198,N_77,N_486);
and U6199 (N_6199,N_3150,N_3950);
and U6200 (N_6200,N_3736,N_3206);
and U6201 (N_6201,N_1912,N_183);
and U6202 (N_6202,N_708,N_1980);
nand U6203 (N_6203,N_1582,N_879);
xnor U6204 (N_6204,N_1160,N_3635);
or U6205 (N_6205,N_3845,N_3786);
and U6206 (N_6206,N_2034,N_1598);
and U6207 (N_6207,N_143,N_1235);
and U6208 (N_6208,N_646,N_415);
and U6209 (N_6209,N_3319,N_3630);
or U6210 (N_6210,N_841,N_3502);
or U6211 (N_6211,N_641,N_80);
or U6212 (N_6212,N_850,N_1075);
nand U6213 (N_6213,N_1789,N_12);
or U6214 (N_6214,N_1375,N_1240);
or U6215 (N_6215,N_2007,N_3819);
and U6216 (N_6216,N_3050,N_1166);
nand U6217 (N_6217,N_1165,N_662);
or U6218 (N_6218,N_2302,N_3134);
or U6219 (N_6219,N_1983,N_2228);
nor U6220 (N_6220,N_2102,N_3670);
xor U6221 (N_6221,N_1684,N_3820);
nor U6222 (N_6222,N_1208,N_2344);
and U6223 (N_6223,N_3578,N_3255);
or U6224 (N_6224,N_2448,N_3428);
xor U6225 (N_6225,N_3112,N_980);
nor U6226 (N_6226,N_497,N_2449);
xnor U6227 (N_6227,N_1050,N_3441);
nor U6228 (N_6228,N_1401,N_3091);
and U6229 (N_6229,N_1312,N_3740);
or U6230 (N_6230,N_43,N_2585);
or U6231 (N_6231,N_3251,N_2530);
nor U6232 (N_6232,N_3285,N_691);
xnor U6233 (N_6233,N_381,N_2807);
nand U6234 (N_6234,N_1736,N_1635);
and U6235 (N_6235,N_262,N_732);
and U6236 (N_6236,N_3276,N_1218);
and U6237 (N_6237,N_3881,N_227);
nor U6238 (N_6238,N_1366,N_2085);
or U6239 (N_6239,N_2167,N_219);
xnor U6240 (N_6240,N_1977,N_2785);
or U6241 (N_6241,N_1720,N_902);
or U6242 (N_6242,N_264,N_378);
nand U6243 (N_6243,N_1093,N_1825);
xor U6244 (N_6244,N_225,N_3838);
xor U6245 (N_6245,N_632,N_3614);
nand U6246 (N_6246,N_2887,N_2286);
or U6247 (N_6247,N_1088,N_2695);
nand U6248 (N_6248,N_1357,N_3734);
and U6249 (N_6249,N_2300,N_2968);
or U6250 (N_6250,N_2340,N_1823);
or U6251 (N_6251,N_3149,N_3637);
or U6252 (N_6252,N_2185,N_252);
nand U6253 (N_6253,N_353,N_3399);
or U6254 (N_6254,N_1749,N_1045);
xor U6255 (N_6255,N_2273,N_186);
or U6256 (N_6256,N_1657,N_1635);
nor U6257 (N_6257,N_1729,N_1316);
xnor U6258 (N_6258,N_1969,N_965);
or U6259 (N_6259,N_3812,N_1519);
xnor U6260 (N_6260,N_1272,N_1213);
or U6261 (N_6261,N_3533,N_2781);
and U6262 (N_6262,N_3026,N_72);
and U6263 (N_6263,N_3900,N_1397);
and U6264 (N_6264,N_3192,N_1017);
or U6265 (N_6265,N_1232,N_2187);
and U6266 (N_6266,N_1012,N_2972);
xor U6267 (N_6267,N_2806,N_173);
nor U6268 (N_6268,N_238,N_2834);
nor U6269 (N_6269,N_2123,N_1674);
or U6270 (N_6270,N_222,N_2274);
or U6271 (N_6271,N_3052,N_2170);
and U6272 (N_6272,N_2582,N_1982);
xor U6273 (N_6273,N_3107,N_2086);
xor U6274 (N_6274,N_134,N_3118);
and U6275 (N_6275,N_352,N_3784);
or U6276 (N_6276,N_2966,N_1271);
and U6277 (N_6277,N_2116,N_3227);
or U6278 (N_6278,N_294,N_3860);
xnor U6279 (N_6279,N_2549,N_34);
or U6280 (N_6280,N_1159,N_1496);
or U6281 (N_6281,N_3140,N_449);
nand U6282 (N_6282,N_1818,N_1637);
and U6283 (N_6283,N_912,N_2378);
and U6284 (N_6284,N_3165,N_821);
and U6285 (N_6285,N_1669,N_216);
nor U6286 (N_6286,N_1554,N_1726);
xor U6287 (N_6287,N_2583,N_3683);
or U6288 (N_6288,N_2723,N_1048);
nor U6289 (N_6289,N_1018,N_1633);
xnor U6290 (N_6290,N_2267,N_1857);
xor U6291 (N_6291,N_940,N_1623);
and U6292 (N_6292,N_3363,N_2708);
or U6293 (N_6293,N_2901,N_3924);
and U6294 (N_6294,N_1395,N_1307);
nor U6295 (N_6295,N_1079,N_2711);
or U6296 (N_6296,N_622,N_1812);
xor U6297 (N_6297,N_2411,N_1024);
nand U6298 (N_6298,N_1506,N_3468);
or U6299 (N_6299,N_2487,N_1846);
nor U6300 (N_6300,N_2175,N_14);
xnor U6301 (N_6301,N_2767,N_1146);
or U6302 (N_6302,N_2080,N_2708);
nand U6303 (N_6303,N_183,N_2004);
xor U6304 (N_6304,N_2126,N_121);
or U6305 (N_6305,N_2203,N_2384);
or U6306 (N_6306,N_609,N_2145);
xor U6307 (N_6307,N_2015,N_69);
and U6308 (N_6308,N_2995,N_3436);
nor U6309 (N_6309,N_3203,N_3071);
xor U6310 (N_6310,N_3097,N_3011);
nand U6311 (N_6311,N_2987,N_1708);
nand U6312 (N_6312,N_2234,N_1397);
and U6313 (N_6313,N_2210,N_1416);
xnor U6314 (N_6314,N_1400,N_3864);
and U6315 (N_6315,N_2432,N_2787);
and U6316 (N_6316,N_1059,N_1196);
xnor U6317 (N_6317,N_3154,N_1134);
xor U6318 (N_6318,N_2169,N_3152);
nor U6319 (N_6319,N_1872,N_1443);
xnor U6320 (N_6320,N_1114,N_784);
and U6321 (N_6321,N_409,N_254);
nand U6322 (N_6322,N_2093,N_1611);
nor U6323 (N_6323,N_2715,N_2639);
or U6324 (N_6324,N_2950,N_318);
xor U6325 (N_6325,N_469,N_2888);
nand U6326 (N_6326,N_1301,N_3843);
or U6327 (N_6327,N_840,N_2374);
xnor U6328 (N_6328,N_1755,N_524);
or U6329 (N_6329,N_1297,N_363);
xor U6330 (N_6330,N_3793,N_119);
nand U6331 (N_6331,N_2648,N_3967);
and U6332 (N_6332,N_1364,N_1495);
nor U6333 (N_6333,N_3994,N_3675);
or U6334 (N_6334,N_2971,N_1320);
xor U6335 (N_6335,N_2774,N_3035);
nand U6336 (N_6336,N_1078,N_3357);
or U6337 (N_6337,N_2058,N_504);
or U6338 (N_6338,N_1439,N_2886);
and U6339 (N_6339,N_1241,N_961);
and U6340 (N_6340,N_1808,N_2825);
and U6341 (N_6341,N_1889,N_3591);
xor U6342 (N_6342,N_3869,N_1296);
xor U6343 (N_6343,N_3680,N_2587);
and U6344 (N_6344,N_54,N_3249);
nor U6345 (N_6345,N_406,N_1975);
and U6346 (N_6346,N_160,N_905);
and U6347 (N_6347,N_1731,N_2349);
xnor U6348 (N_6348,N_286,N_3179);
nor U6349 (N_6349,N_557,N_3113);
xnor U6350 (N_6350,N_1294,N_681);
or U6351 (N_6351,N_111,N_3775);
xor U6352 (N_6352,N_1106,N_3479);
and U6353 (N_6353,N_2217,N_1340);
xnor U6354 (N_6354,N_2457,N_1155);
or U6355 (N_6355,N_3900,N_3458);
and U6356 (N_6356,N_2357,N_2739);
xor U6357 (N_6357,N_1875,N_2335);
nor U6358 (N_6358,N_3554,N_3775);
nand U6359 (N_6359,N_1408,N_2639);
or U6360 (N_6360,N_1394,N_1843);
and U6361 (N_6361,N_1077,N_2661);
and U6362 (N_6362,N_2770,N_2362);
or U6363 (N_6363,N_441,N_3565);
or U6364 (N_6364,N_1234,N_2504);
or U6365 (N_6365,N_3691,N_1865);
and U6366 (N_6366,N_2012,N_143);
or U6367 (N_6367,N_2998,N_25);
nand U6368 (N_6368,N_745,N_1015);
nor U6369 (N_6369,N_374,N_316);
or U6370 (N_6370,N_270,N_753);
or U6371 (N_6371,N_2516,N_481);
or U6372 (N_6372,N_2972,N_3344);
or U6373 (N_6373,N_1272,N_2747);
nand U6374 (N_6374,N_1813,N_827);
and U6375 (N_6375,N_1727,N_1679);
xor U6376 (N_6376,N_2402,N_1832);
and U6377 (N_6377,N_2760,N_1490);
xnor U6378 (N_6378,N_3242,N_3882);
or U6379 (N_6379,N_710,N_119);
and U6380 (N_6380,N_3451,N_2246);
nand U6381 (N_6381,N_3739,N_350);
nand U6382 (N_6382,N_829,N_2290);
nor U6383 (N_6383,N_3987,N_1524);
nand U6384 (N_6384,N_3604,N_1520);
or U6385 (N_6385,N_12,N_2741);
or U6386 (N_6386,N_3466,N_1690);
or U6387 (N_6387,N_1610,N_385);
xor U6388 (N_6388,N_2060,N_2517);
nor U6389 (N_6389,N_103,N_3544);
and U6390 (N_6390,N_1124,N_1375);
and U6391 (N_6391,N_315,N_2833);
or U6392 (N_6392,N_1924,N_3411);
nand U6393 (N_6393,N_992,N_1767);
nor U6394 (N_6394,N_325,N_170);
or U6395 (N_6395,N_2118,N_261);
xor U6396 (N_6396,N_2946,N_298);
nand U6397 (N_6397,N_771,N_2887);
xnor U6398 (N_6398,N_3341,N_1884);
or U6399 (N_6399,N_517,N_3970);
xnor U6400 (N_6400,N_3303,N_530);
or U6401 (N_6401,N_1316,N_1708);
xnor U6402 (N_6402,N_2472,N_275);
or U6403 (N_6403,N_3491,N_3129);
nor U6404 (N_6404,N_788,N_2859);
and U6405 (N_6405,N_1440,N_249);
nand U6406 (N_6406,N_182,N_3581);
or U6407 (N_6407,N_1044,N_1417);
and U6408 (N_6408,N_2049,N_1766);
and U6409 (N_6409,N_257,N_3003);
xnor U6410 (N_6410,N_622,N_2044);
nand U6411 (N_6411,N_1154,N_2742);
and U6412 (N_6412,N_3458,N_2554);
nand U6413 (N_6413,N_379,N_1923);
xnor U6414 (N_6414,N_1388,N_2218);
or U6415 (N_6415,N_591,N_3730);
nand U6416 (N_6416,N_1173,N_2678);
xnor U6417 (N_6417,N_2648,N_868);
nand U6418 (N_6418,N_66,N_38);
nor U6419 (N_6419,N_3054,N_614);
xnor U6420 (N_6420,N_93,N_2026);
and U6421 (N_6421,N_38,N_3169);
nand U6422 (N_6422,N_518,N_2061);
or U6423 (N_6423,N_3325,N_945);
nand U6424 (N_6424,N_1123,N_1266);
nand U6425 (N_6425,N_2530,N_1325);
nand U6426 (N_6426,N_3330,N_1693);
nor U6427 (N_6427,N_2843,N_1489);
and U6428 (N_6428,N_2415,N_104);
nand U6429 (N_6429,N_3133,N_2347);
and U6430 (N_6430,N_3591,N_1026);
and U6431 (N_6431,N_2925,N_2764);
and U6432 (N_6432,N_1719,N_243);
nor U6433 (N_6433,N_2424,N_1863);
nand U6434 (N_6434,N_1383,N_120);
or U6435 (N_6435,N_3979,N_3481);
nand U6436 (N_6436,N_881,N_375);
nor U6437 (N_6437,N_201,N_1186);
xnor U6438 (N_6438,N_2442,N_3246);
xnor U6439 (N_6439,N_3862,N_2477);
nor U6440 (N_6440,N_2357,N_1696);
nor U6441 (N_6441,N_808,N_2145);
nor U6442 (N_6442,N_3385,N_3822);
or U6443 (N_6443,N_506,N_2225);
and U6444 (N_6444,N_1256,N_3929);
nor U6445 (N_6445,N_225,N_3022);
and U6446 (N_6446,N_2174,N_920);
xor U6447 (N_6447,N_2776,N_559);
nand U6448 (N_6448,N_3075,N_890);
and U6449 (N_6449,N_2097,N_1126);
nor U6450 (N_6450,N_2894,N_1726);
nand U6451 (N_6451,N_3856,N_213);
or U6452 (N_6452,N_3195,N_1012);
nor U6453 (N_6453,N_369,N_1005);
nor U6454 (N_6454,N_1806,N_2351);
nor U6455 (N_6455,N_65,N_3885);
and U6456 (N_6456,N_1877,N_2252);
nand U6457 (N_6457,N_1082,N_3590);
nand U6458 (N_6458,N_2430,N_3409);
and U6459 (N_6459,N_1180,N_2956);
nor U6460 (N_6460,N_1996,N_2150);
nor U6461 (N_6461,N_1965,N_450);
nand U6462 (N_6462,N_3044,N_1450);
nor U6463 (N_6463,N_2071,N_363);
or U6464 (N_6464,N_3245,N_1136);
and U6465 (N_6465,N_3106,N_621);
or U6466 (N_6466,N_1646,N_502);
and U6467 (N_6467,N_1928,N_2638);
xnor U6468 (N_6468,N_3580,N_1298);
xnor U6469 (N_6469,N_3208,N_3729);
nand U6470 (N_6470,N_955,N_2374);
nor U6471 (N_6471,N_1681,N_2510);
and U6472 (N_6472,N_257,N_2593);
and U6473 (N_6473,N_3443,N_205);
or U6474 (N_6474,N_3817,N_3387);
xnor U6475 (N_6475,N_2635,N_1563);
or U6476 (N_6476,N_1450,N_322);
xor U6477 (N_6477,N_2711,N_1777);
and U6478 (N_6478,N_634,N_457);
nor U6479 (N_6479,N_711,N_2073);
xnor U6480 (N_6480,N_1355,N_3886);
or U6481 (N_6481,N_1574,N_2905);
nand U6482 (N_6482,N_1710,N_1912);
nor U6483 (N_6483,N_1695,N_1195);
xnor U6484 (N_6484,N_2839,N_3946);
or U6485 (N_6485,N_958,N_1676);
nor U6486 (N_6486,N_743,N_607);
nand U6487 (N_6487,N_3246,N_159);
xnor U6488 (N_6488,N_1130,N_647);
or U6489 (N_6489,N_2921,N_3530);
nand U6490 (N_6490,N_1548,N_3827);
nor U6491 (N_6491,N_1303,N_3316);
or U6492 (N_6492,N_901,N_3729);
nand U6493 (N_6493,N_1523,N_1512);
and U6494 (N_6494,N_929,N_2284);
or U6495 (N_6495,N_1003,N_5);
nor U6496 (N_6496,N_2117,N_2454);
or U6497 (N_6497,N_730,N_233);
nand U6498 (N_6498,N_2181,N_2180);
nor U6499 (N_6499,N_265,N_1601);
nor U6500 (N_6500,N_1507,N_3659);
nor U6501 (N_6501,N_2000,N_880);
and U6502 (N_6502,N_2478,N_3844);
nor U6503 (N_6503,N_1936,N_3937);
or U6504 (N_6504,N_3948,N_2677);
and U6505 (N_6505,N_3348,N_2940);
nand U6506 (N_6506,N_1690,N_2780);
xor U6507 (N_6507,N_315,N_3309);
and U6508 (N_6508,N_80,N_2460);
and U6509 (N_6509,N_2240,N_1336);
nand U6510 (N_6510,N_2020,N_1708);
nand U6511 (N_6511,N_2103,N_2780);
or U6512 (N_6512,N_326,N_675);
and U6513 (N_6513,N_2604,N_2137);
nor U6514 (N_6514,N_2154,N_608);
nor U6515 (N_6515,N_3242,N_2906);
and U6516 (N_6516,N_803,N_1632);
xnor U6517 (N_6517,N_880,N_416);
nor U6518 (N_6518,N_597,N_1156);
nor U6519 (N_6519,N_2888,N_353);
or U6520 (N_6520,N_3215,N_3660);
or U6521 (N_6521,N_1333,N_887);
nor U6522 (N_6522,N_181,N_760);
and U6523 (N_6523,N_1387,N_317);
or U6524 (N_6524,N_1041,N_2747);
nor U6525 (N_6525,N_1234,N_2944);
or U6526 (N_6526,N_3063,N_2740);
and U6527 (N_6527,N_3037,N_1422);
nand U6528 (N_6528,N_3488,N_3009);
nand U6529 (N_6529,N_3773,N_3946);
xnor U6530 (N_6530,N_484,N_568);
nand U6531 (N_6531,N_1358,N_2698);
and U6532 (N_6532,N_3901,N_254);
or U6533 (N_6533,N_1136,N_2339);
or U6534 (N_6534,N_2144,N_3797);
and U6535 (N_6535,N_1258,N_1631);
xor U6536 (N_6536,N_333,N_2487);
or U6537 (N_6537,N_2986,N_760);
or U6538 (N_6538,N_3810,N_2007);
and U6539 (N_6539,N_1128,N_2986);
nand U6540 (N_6540,N_1894,N_373);
xnor U6541 (N_6541,N_3186,N_740);
xor U6542 (N_6542,N_1892,N_3333);
or U6543 (N_6543,N_1236,N_196);
or U6544 (N_6544,N_2722,N_1194);
nand U6545 (N_6545,N_3794,N_427);
nor U6546 (N_6546,N_2522,N_2215);
nand U6547 (N_6547,N_2453,N_2185);
and U6548 (N_6548,N_2503,N_472);
and U6549 (N_6549,N_1393,N_1912);
xnor U6550 (N_6550,N_3180,N_3138);
nand U6551 (N_6551,N_3755,N_2708);
and U6552 (N_6552,N_2465,N_2226);
or U6553 (N_6553,N_2488,N_1472);
xnor U6554 (N_6554,N_2552,N_2556);
and U6555 (N_6555,N_1896,N_3518);
or U6556 (N_6556,N_2972,N_1124);
nand U6557 (N_6557,N_1019,N_2473);
or U6558 (N_6558,N_2220,N_2158);
nand U6559 (N_6559,N_2922,N_1054);
nor U6560 (N_6560,N_1882,N_541);
xnor U6561 (N_6561,N_1315,N_1114);
and U6562 (N_6562,N_110,N_3849);
and U6563 (N_6563,N_32,N_1439);
or U6564 (N_6564,N_2732,N_3560);
and U6565 (N_6565,N_2253,N_3070);
nor U6566 (N_6566,N_1266,N_1277);
nor U6567 (N_6567,N_1670,N_2771);
and U6568 (N_6568,N_3454,N_1012);
xnor U6569 (N_6569,N_2364,N_1291);
nor U6570 (N_6570,N_1857,N_3613);
nand U6571 (N_6571,N_7,N_1169);
or U6572 (N_6572,N_3297,N_1093);
nand U6573 (N_6573,N_864,N_1029);
nor U6574 (N_6574,N_1517,N_787);
xnor U6575 (N_6575,N_1880,N_2067);
or U6576 (N_6576,N_2436,N_1544);
and U6577 (N_6577,N_1590,N_3834);
or U6578 (N_6578,N_2899,N_872);
nand U6579 (N_6579,N_2466,N_376);
nor U6580 (N_6580,N_2558,N_3690);
nand U6581 (N_6581,N_684,N_2525);
and U6582 (N_6582,N_2190,N_464);
and U6583 (N_6583,N_3740,N_1573);
or U6584 (N_6584,N_3269,N_3153);
nor U6585 (N_6585,N_3502,N_3448);
or U6586 (N_6586,N_2875,N_3409);
and U6587 (N_6587,N_2478,N_2512);
nand U6588 (N_6588,N_1694,N_2616);
xor U6589 (N_6589,N_3302,N_2323);
nor U6590 (N_6590,N_2947,N_169);
and U6591 (N_6591,N_1029,N_2917);
xor U6592 (N_6592,N_624,N_3809);
or U6593 (N_6593,N_3369,N_2923);
xor U6594 (N_6594,N_1982,N_466);
nand U6595 (N_6595,N_358,N_1954);
and U6596 (N_6596,N_3223,N_3641);
xor U6597 (N_6597,N_2009,N_3559);
xor U6598 (N_6598,N_1383,N_1850);
nor U6599 (N_6599,N_3254,N_3973);
nand U6600 (N_6600,N_495,N_709);
and U6601 (N_6601,N_1690,N_533);
and U6602 (N_6602,N_1904,N_1622);
nor U6603 (N_6603,N_866,N_2850);
nor U6604 (N_6604,N_537,N_111);
nand U6605 (N_6605,N_2601,N_2334);
nand U6606 (N_6606,N_381,N_122);
xnor U6607 (N_6607,N_2698,N_1722);
nand U6608 (N_6608,N_3295,N_899);
and U6609 (N_6609,N_2343,N_137);
xor U6610 (N_6610,N_2893,N_540);
nor U6611 (N_6611,N_245,N_2210);
nand U6612 (N_6612,N_870,N_357);
or U6613 (N_6613,N_1658,N_1937);
or U6614 (N_6614,N_530,N_252);
nor U6615 (N_6615,N_1878,N_1838);
nor U6616 (N_6616,N_1517,N_3701);
nand U6617 (N_6617,N_2307,N_3124);
xor U6618 (N_6618,N_1592,N_3959);
and U6619 (N_6619,N_1500,N_3488);
xnor U6620 (N_6620,N_1607,N_3394);
nor U6621 (N_6621,N_2922,N_3623);
or U6622 (N_6622,N_1421,N_974);
and U6623 (N_6623,N_3438,N_686);
xor U6624 (N_6624,N_467,N_1917);
nand U6625 (N_6625,N_2825,N_481);
xor U6626 (N_6626,N_1853,N_1077);
xnor U6627 (N_6627,N_111,N_387);
and U6628 (N_6628,N_3858,N_3379);
nand U6629 (N_6629,N_1015,N_2261);
nand U6630 (N_6630,N_3210,N_682);
nor U6631 (N_6631,N_3829,N_3457);
xor U6632 (N_6632,N_1117,N_1231);
or U6633 (N_6633,N_1828,N_3433);
xnor U6634 (N_6634,N_1393,N_612);
or U6635 (N_6635,N_3154,N_3414);
or U6636 (N_6636,N_1519,N_2184);
nand U6637 (N_6637,N_955,N_56);
and U6638 (N_6638,N_1238,N_3445);
nor U6639 (N_6639,N_1605,N_3700);
xor U6640 (N_6640,N_2149,N_2549);
xnor U6641 (N_6641,N_977,N_1760);
xnor U6642 (N_6642,N_780,N_2609);
xor U6643 (N_6643,N_2339,N_3498);
or U6644 (N_6644,N_541,N_3323);
and U6645 (N_6645,N_3419,N_1855);
nor U6646 (N_6646,N_946,N_1472);
or U6647 (N_6647,N_3670,N_828);
nor U6648 (N_6648,N_3563,N_3057);
or U6649 (N_6649,N_2805,N_2573);
nor U6650 (N_6650,N_2548,N_1879);
xnor U6651 (N_6651,N_1977,N_2100);
nand U6652 (N_6652,N_3361,N_3387);
or U6653 (N_6653,N_1886,N_2383);
nand U6654 (N_6654,N_726,N_701);
nor U6655 (N_6655,N_3271,N_3782);
xor U6656 (N_6656,N_2308,N_338);
xnor U6657 (N_6657,N_3605,N_3493);
nand U6658 (N_6658,N_2402,N_1060);
and U6659 (N_6659,N_754,N_2778);
nor U6660 (N_6660,N_3604,N_1202);
and U6661 (N_6661,N_3001,N_1563);
xor U6662 (N_6662,N_3133,N_826);
nor U6663 (N_6663,N_1766,N_2693);
or U6664 (N_6664,N_3352,N_1841);
nor U6665 (N_6665,N_1744,N_2673);
nand U6666 (N_6666,N_3890,N_550);
nor U6667 (N_6667,N_3832,N_1531);
or U6668 (N_6668,N_29,N_121);
xnor U6669 (N_6669,N_2545,N_1085);
nand U6670 (N_6670,N_2899,N_521);
and U6671 (N_6671,N_3227,N_2231);
and U6672 (N_6672,N_2196,N_1811);
nand U6673 (N_6673,N_2880,N_3825);
xor U6674 (N_6674,N_1706,N_2002);
or U6675 (N_6675,N_3391,N_1396);
nor U6676 (N_6676,N_2886,N_3482);
nor U6677 (N_6677,N_2075,N_1970);
nand U6678 (N_6678,N_2354,N_960);
and U6679 (N_6679,N_1545,N_2364);
nand U6680 (N_6680,N_1344,N_3337);
or U6681 (N_6681,N_2,N_102);
nand U6682 (N_6682,N_2540,N_2574);
or U6683 (N_6683,N_3277,N_2779);
nor U6684 (N_6684,N_2788,N_399);
nand U6685 (N_6685,N_2951,N_1761);
nor U6686 (N_6686,N_3371,N_2155);
xor U6687 (N_6687,N_1222,N_2114);
xnor U6688 (N_6688,N_3521,N_2158);
or U6689 (N_6689,N_1425,N_3469);
and U6690 (N_6690,N_1570,N_1883);
nand U6691 (N_6691,N_2659,N_83);
xnor U6692 (N_6692,N_252,N_1866);
nand U6693 (N_6693,N_3801,N_2856);
nor U6694 (N_6694,N_1159,N_2915);
and U6695 (N_6695,N_278,N_507);
or U6696 (N_6696,N_3990,N_213);
nand U6697 (N_6697,N_721,N_2138);
nor U6698 (N_6698,N_1811,N_616);
nor U6699 (N_6699,N_2972,N_2211);
xor U6700 (N_6700,N_2948,N_1994);
nand U6701 (N_6701,N_2744,N_2111);
nand U6702 (N_6702,N_1005,N_3856);
xnor U6703 (N_6703,N_1119,N_3944);
xor U6704 (N_6704,N_3037,N_3691);
nor U6705 (N_6705,N_3455,N_1933);
or U6706 (N_6706,N_3534,N_3798);
nor U6707 (N_6707,N_3147,N_2260);
and U6708 (N_6708,N_714,N_72);
xor U6709 (N_6709,N_618,N_3347);
nor U6710 (N_6710,N_2478,N_1941);
nor U6711 (N_6711,N_1732,N_2664);
or U6712 (N_6712,N_3489,N_1662);
nor U6713 (N_6713,N_2546,N_2561);
xor U6714 (N_6714,N_3953,N_3389);
and U6715 (N_6715,N_3930,N_3608);
and U6716 (N_6716,N_107,N_2530);
or U6717 (N_6717,N_2568,N_3747);
or U6718 (N_6718,N_778,N_39);
and U6719 (N_6719,N_2140,N_2097);
nand U6720 (N_6720,N_969,N_1353);
nand U6721 (N_6721,N_1373,N_209);
or U6722 (N_6722,N_1272,N_3308);
xor U6723 (N_6723,N_1795,N_1508);
and U6724 (N_6724,N_1942,N_667);
or U6725 (N_6725,N_790,N_1297);
and U6726 (N_6726,N_1726,N_1464);
and U6727 (N_6727,N_3479,N_1133);
nand U6728 (N_6728,N_2990,N_3164);
or U6729 (N_6729,N_3404,N_2010);
or U6730 (N_6730,N_2404,N_3710);
and U6731 (N_6731,N_1716,N_1905);
nand U6732 (N_6732,N_2888,N_3197);
or U6733 (N_6733,N_3687,N_1365);
nor U6734 (N_6734,N_1445,N_418);
nand U6735 (N_6735,N_3665,N_3919);
or U6736 (N_6736,N_979,N_1741);
nand U6737 (N_6737,N_823,N_2123);
and U6738 (N_6738,N_1432,N_2173);
or U6739 (N_6739,N_1710,N_3640);
xnor U6740 (N_6740,N_1485,N_1673);
or U6741 (N_6741,N_2235,N_1931);
nor U6742 (N_6742,N_3015,N_3037);
and U6743 (N_6743,N_139,N_1383);
nand U6744 (N_6744,N_3228,N_2703);
xnor U6745 (N_6745,N_1911,N_1655);
and U6746 (N_6746,N_785,N_3572);
or U6747 (N_6747,N_3426,N_2109);
nand U6748 (N_6748,N_3860,N_3263);
xnor U6749 (N_6749,N_1698,N_1099);
nand U6750 (N_6750,N_455,N_1055);
nand U6751 (N_6751,N_3576,N_236);
nand U6752 (N_6752,N_3121,N_201);
or U6753 (N_6753,N_1600,N_2462);
nand U6754 (N_6754,N_267,N_958);
or U6755 (N_6755,N_493,N_914);
or U6756 (N_6756,N_3133,N_906);
and U6757 (N_6757,N_3757,N_3253);
nor U6758 (N_6758,N_469,N_992);
xnor U6759 (N_6759,N_895,N_1165);
or U6760 (N_6760,N_3353,N_2122);
or U6761 (N_6761,N_1892,N_3807);
or U6762 (N_6762,N_1394,N_3998);
xnor U6763 (N_6763,N_1589,N_3835);
nor U6764 (N_6764,N_2907,N_3406);
or U6765 (N_6765,N_2951,N_2724);
nand U6766 (N_6766,N_1205,N_373);
nor U6767 (N_6767,N_2653,N_3205);
nor U6768 (N_6768,N_3663,N_2969);
xor U6769 (N_6769,N_1128,N_1551);
nor U6770 (N_6770,N_1813,N_1940);
and U6771 (N_6771,N_802,N_2048);
and U6772 (N_6772,N_791,N_2800);
nand U6773 (N_6773,N_131,N_1182);
and U6774 (N_6774,N_1765,N_1630);
and U6775 (N_6775,N_2637,N_3478);
nor U6776 (N_6776,N_598,N_1025);
nand U6777 (N_6777,N_2799,N_3515);
and U6778 (N_6778,N_2216,N_3967);
nand U6779 (N_6779,N_1381,N_1855);
and U6780 (N_6780,N_2294,N_2448);
nand U6781 (N_6781,N_1573,N_1427);
xor U6782 (N_6782,N_1145,N_3346);
nand U6783 (N_6783,N_3969,N_3210);
nor U6784 (N_6784,N_1569,N_3856);
nor U6785 (N_6785,N_1610,N_11);
and U6786 (N_6786,N_1761,N_1478);
xnor U6787 (N_6787,N_2390,N_3714);
nor U6788 (N_6788,N_2533,N_1261);
nand U6789 (N_6789,N_2653,N_1038);
nand U6790 (N_6790,N_2863,N_3187);
nand U6791 (N_6791,N_3657,N_2668);
and U6792 (N_6792,N_2678,N_1055);
and U6793 (N_6793,N_3615,N_158);
and U6794 (N_6794,N_824,N_3410);
or U6795 (N_6795,N_3712,N_1710);
nand U6796 (N_6796,N_3132,N_133);
nand U6797 (N_6797,N_572,N_964);
xor U6798 (N_6798,N_3126,N_3114);
and U6799 (N_6799,N_1686,N_3816);
nand U6800 (N_6800,N_1553,N_1317);
nor U6801 (N_6801,N_1107,N_3545);
or U6802 (N_6802,N_1397,N_1388);
nand U6803 (N_6803,N_2604,N_11);
nand U6804 (N_6804,N_2315,N_1319);
nand U6805 (N_6805,N_954,N_2749);
nand U6806 (N_6806,N_2725,N_2044);
or U6807 (N_6807,N_442,N_2779);
xnor U6808 (N_6808,N_1049,N_264);
xnor U6809 (N_6809,N_2231,N_3957);
nor U6810 (N_6810,N_1627,N_3598);
nor U6811 (N_6811,N_646,N_1072);
nor U6812 (N_6812,N_1080,N_3075);
xnor U6813 (N_6813,N_708,N_2311);
nand U6814 (N_6814,N_535,N_2412);
xnor U6815 (N_6815,N_662,N_3913);
or U6816 (N_6816,N_2171,N_2029);
and U6817 (N_6817,N_1995,N_711);
nor U6818 (N_6818,N_3618,N_3015);
nor U6819 (N_6819,N_945,N_1105);
nor U6820 (N_6820,N_1532,N_159);
and U6821 (N_6821,N_291,N_825);
xnor U6822 (N_6822,N_2980,N_3207);
xnor U6823 (N_6823,N_650,N_2093);
and U6824 (N_6824,N_1129,N_578);
xnor U6825 (N_6825,N_2225,N_2245);
and U6826 (N_6826,N_3897,N_1795);
xnor U6827 (N_6827,N_3380,N_1911);
nand U6828 (N_6828,N_1098,N_1374);
nand U6829 (N_6829,N_2428,N_422);
or U6830 (N_6830,N_3083,N_3626);
and U6831 (N_6831,N_2284,N_71);
nor U6832 (N_6832,N_2494,N_3667);
nand U6833 (N_6833,N_1809,N_136);
or U6834 (N_6834,N_2926,N_1843);
and U6835 (N_6835,N_982,N_3341);
nand U6836 (N_6836,N_3318,N_2065);
or U6837 (N_6837,N_1190,N_2615);
and U6838 (N_6838,N_2645,N_1047);
nand U6839 (N_6839,N_874,N_3204);
nand U6840 (N_6840,N_183,N_1418);
or U6841 (N_6841,N_1010,N_2643);
or U6842 (N_6842,N_502,N_1953);
nand U6843 (N_6843,N_270,N_2357);
nand U6844 (N_6844,N_3423,N_2783);
nor U6845 (N_6845,N_2305,N_785);
xnor U6846 (N_6846,N_49,N_1494);
nand U6847 (N_6847,N_2319,N_2494);
or U6848 (N_6848,N_294,N_933);
or U6849 (N_6849,N_1771,N_2201);
or U6850 (N_6850,N_1865,N_1019);
nor U6851 (N_6851,N_3822,N_3958);
nand U6852 (N_6852,N_3104,N_3962);
or U6853 (N_6853,N_948,N_728);
xor U6854 (N_6854,N_3820,N_731);
nand U6855 (N_6855,N_1618,N_3985);
nor U6856 (N_6856,N_2537,N_672);
and U6857 (N_6857,N_1957,N_3663);
and U6858 (N_6858,N_345,N_2498);
or U6859 (N_6859,N_1411,N_2700);
nand U6860 (N_6860,N_651,N_1827);
and U6861 (N_6861,N_1993,N_2795);
and U6862 (N_6862,N_3872,N_1762);
and U6863 (N_6863,N_2738,N_1951);
nor U6864 (N_6864,N_968,N_876);
and U6865 (N_6865,N_3925,N_3295);
nor U6866 (N_6866,N_1397,N_3435);
xor U6867 (N_6867,N_2686,N_7);
xnor U6868 (N_6868,N_3068,N_3045);
xor U6869 (N_6869,N_3362,N_1229);
nand U6870 (N_6870,N_3044,N_2841);
xor U6871 (N_6871,N_3436,N_587);
nand U6872 (N_6872,N_3477,N_1553);
and U6873 (N_6873,N_1322,N_3867);
nand U6874 (N_6874,N_1921,N_2283);
nor U6875 (N_6875,N_2402,N_297);
nor U6876 (N_6876,N_2628,N_120);
nor U6877 (N_6877,N_1326,N_1460);
xor U6878 (N_6878,N_735,N_2665);
and U6879 (N_6879,N_1946,N_1162);
xor U6880 (N_6880,N_1974,N_2773);
or U6881 (N_6881,N_1530,N_2494);
or U6882 (N_6882,N_665,N_3604);
nand U6883 (N_6883,N_3530,N_939);
and U6884 (N_6884,N_316,N_1132);
xor U6885 (N_6885,N_1270,N_3116);
and U6886 (N_6886,N_94,N_2504);
nand U6887 (N_6887,N_192,N_937);
xor U6888 (N_6888,N_3837,N_1320);
nand U6889 (N_6889,N_870,N_2507);
nor U6890 (N_6890,N_2453,N_3161);
and U6891 (N_6891,N_1018,N_827);
and U6892 (N_6892,N_3115,N_2091);
xnor U6893 (N_6893,N_3578,N_1672);
xnor U6894 (N_6894,N_979,N_1173);
and U6895 (N_6895,N_650,N_1698);
xnor U6896 (N_6896,N_686,N_197);
xnor U6897 (N_6897,N_2925,N_3862);
nand U6898 (N_6898,N_1638,N_1615);
and U6899 (N_6899,N_1921,N_1585);
nor U6900 (N_6900,N_537,N_1510);
or U6901 (N_6901,N_154,N_815);
xor U6902 (N_6902,N_298,N_872);
or U6903 (N_6903,N_3277,N_1906);
and U6904 (N_6904,N_1998,N_2163);
nand U6905 (N_6905,N_3576,N_3345);
nand U6906 (N_6906,N_880,N_2952);
and U6907 (N_6907,N_3519,N_68);
or U6908 (N_6908,N_1367,N_3932);
nand U6909 (N_6909,N_994,N_145);
and U6910 (N_6910,N_1373,N_1692);
nand U6911 (N_6911,N_3214,N_210);
nor U6912 (N_6912,N_1929,N_1720);
or U6913 (N_6913,N_1418,N_322);
xnor U6914 (N_6914,N_1144,N_2844);
or U6915 (N_6915,N_688,N_2488);
nor U6916 (N_6916,N_282,N_2551);
nand U6917 (N_6917,N_1863,N_3904);
or U6918 (N_6918,N_2763,N_2436);
and U6919 (N_6919,N_1390,N_306);
and U6920 (N_6920,N_1963,N_497);
and U6921 (N_6921,N_614,N_149);
nand U6922 (N_6922,N_3864,N_550);
nand U6923 (N_6923,N_910,N_3893);
nor U6924 (N_6924,N_526,N_3920);
and U6925 (N_6925,N_605,N_1374);
and U6926 (N_6926,N_1043,N_3424);
or U6927 (N_6927,N_327,N_3074);
nor U6928 (N_6928,N_3595,N_2823);
or U6929 (N_6929,N_3097,N_2648);
and U6930 (N_6930,N_238,N_3228);
nand U6931 (N_6931,N_534,N_2374);
xor U6932 (N_6932,N_1448,N_2165);
and U6933 (N_6933,N_3332,N_3110);
nor U6934 (N_6934,N_3568,N_2041);
or U6935 (N_6935,N_622,N_1281);
or U6936 (N_6936,N_3645,N_1485);
nor U6937 (N_6937,N_122,N_1006);
nand U6938 (N_6938,N_3313,N_2963);
or U6939 (N_6939,N_2982,N_1414);
nand U6940 (N_6940,N_104,N_3374);
or U6941 (N_6941,N_2252,N_1737);
xor U6942 (N_6942,N_1508,N_1928);
and U6943 (N_6943,N_2286,N_3895);
nand U6944 (N_6944,N_365,N_1384);
xnor U6945 (N_6945,N_903,N_2181);
and U6946 (N_6946,N_761,N_1757);
nand U6947 (N_6947,N_3080,N_2357);
nor U6948 (N_6948,N_3843,N_1832);
nor U6949 (N_6949,N_2284,N_3378);
nand U6950 (N_6950,N_2257,N_2354);
xor U6951 (N_6951,N_1131,N_629);
nor U6952 (N_6952,N_2126,N_3500);
or U6953 (N_6953,N_2001,N_1059);
nand U6954 (N_6954,N_3005,N_669);
and U6955 (N_6955,N_3019,N_1357);
xor U6956 (N_6956,N_487,N_1271);
xnor U6957 (N_6957,N_230,N_3918);
or U6958 (N_6958,N_481,N_3398);
and U6959 (N_6959,N_3384,N_3082);
xor U6960 (N_6960,N_2571,N_275);
nand U6961 (N_6961,N_935,N_2231);
nand U6962 (N_6962,N_3335,N_3830);
or U6963 (N_6963,N_3339,N_2214);
nand U6964 (N_6964,N_3266,N_3064);
and U6965 (N_6965,N_826,N_211);
xnor U6966 (N_6966,N_848,N_2503);
nor U6967 (N_6967,N_1392,N_332);
or U6968 (N_6968,N_1490,N_1171);
or U6969 (N_6969,N_2863,N_2252);
nand U6970 (N_6970,N_3393,N_2342);
xnor U6971 (N_6971,N_1234,N_2362);
and U6972 (N_6972,N_2258,N_3940);
or U6973 (N_6973,N_2432,N_389);
or U6974 (N_6974,N_1487,N_2266);
nor U6975 (N_6975,N_3585,N_2969);
nand U6976 (N_6976,N_2168,N_2555);
and U6977 (N_6977,N_834,N_3697);
nand U6978 (N_6978,N_1016,N_3892);
nand U6979 (N_6979,N_1785,N_2525);
or U6980 (N_6980,N_2205,N_2024);
nor U6981 (N_6981,N_1840,N_118);
and U6982 (N_6982,N_2541,N_1019);
and U6983 (N_6983,N_677,N_73);
xor U6984 (N_6984,N_83,N_2759);
xnor U6985 (N_6985,N_2589,N_1548);
nor U6986 (N_6986,N_1275,N_35);
and U6987 (N_6987,N_766,N_3700);
nor U6988 (N_6988,N_1520,N_3040);
nor U6989 (N_6989,N_3609,N_1101);
or U6990 (N_6990,N_1615,N_2769);
nor U6991 (N_6991,N_3869,N_2091);
nor U6992 (N_6992,N_187,N_3357);
nand U6993 (N_6993,N_3942,N_2093);
nor U6994 (N_6994,N_731,N_2948);
xor U6995 (N_6995,N_3351,N_3023);
nand U6996 (N_6996,N_553,N_3008);
xor U6997 (N_6997,N_3685,N_2850);
xnor U6998 (N_6998,N_172,N_995);
nand U6999 (N_6999,N_2979,N_3422);
nor U7000 (N_7000,N_3789,N_2191);
xnor U7001 (N_7001,N_1403,N_3735);
nand U7002 (N_7002,N_201,N_2686);
xnor U7003 (N_7003,N_2230,N_2431);
or U7004 (N_7004,N_3314,N_2085);
xnor U7005 (N_7005,N_2356,N_667);
xor U7006 (N_7006,N_2158,N_3696);
xnor U7007 (N_7007,N_2535,N_3565);
or U7008 (N_7008,N_700,N_3626);
and U7009 (N_7009,N_3464,N_2540);
nand U7010 (N_7010,N_3495,N_1103);
nor U7011 (N_7011,N_390,N_3036);
or U7012 (N_7012,N_3842,N_2355);
nor U7013 (N_7013,N_2569,N_2308);
or U7014 (N_7014,N_2198,N_2943);
or U7015 (N_7015,N_3619,N_2803);
nand U7016 (N_7016,N_2364,N_533);
and U7017 (N_7017,N_1557,N_3989);
or U7018 (N_7018,N_516,N_1041);
or U7019 (N_7019,N_3569,N_3966);
xor U7020 (N_7020,N_800,N_30);
nand U7021 (N_7021,N_2006,N_2117);
and U7022 (N_7022,N_359,N_1876);
nor U7023 (N_7023,N_2867,N_481);
xnor U7024 (N_7024,N_976,N_1440);
nand U7025 (N_7025,N_182,N_2366);
and U7026 (N_7026,N_231,N_2289);
or U7027 (N_7027,N_1616,N_2442);
or U7028 (N_7028,N_3783,N_1111);
and U7029 (N_7029,N_3561,N_1180);
and U7030 (N_7030,N_2075,N_1877);
and U7031 (N_7031,N_644,N_1976);
or U7032 (N_7032,N_753,N_3605);
xor U7033 (N_7033,N_3896,N_81);
xor U7034 (N_7034,N_1685,N_822);
xnor U7035 (N_7035,N_832,N_3723);
or U7036 (N_7036,N_2264,N_3928);
nor U7037 (N_7037,N_987,N_430);
xor U7038 (N_7038,N_2167,N_276);
xor U7039 (N_7039,N_3682,N_204);
nand U7040 (N_7040,N_934,N_920);
nand U7041 (N_7041,N_2484,N_3307);
and U7042 (N_7042,N_2485,N_990);
nand U7043 (N_7043,N_1999,N_1061);
nor U7044 (N_7044,N_2644,N_3066);
nand U7045 (N_7045,N_2106,N_601);
or U7046 (N_7046,N_1450,N_3446);
nand U7047 (N_7047,N_710,N_472);
or U7048 (N_7048,N_3687,N_1867);
nand U7049 (N_7049,N_2686,N_1307);
xnor U7050 (N_7050,N_2037,N_2681);
xnor U7051 (N_7051,N_800,N_3807);
nand U7052 (N_7052,N_787,N_3128);
nor U7053 (N_7053,N_3963,N_1937);
nor U7054 (N_7054,N_327,N_3769);
and U7055 (N_7055,N_3146,N_576);
nand U7056 (N_7056,N_525,N_3726);
nor U7057 (N_7057,N_33,N_1767);
nand U7058 (N_7058,N_3699,N_1375);
nor U7059 (N_7059,N_885,N_844);
or U7060 (N_7060,N_1781,N_2290);
and U7061 (N_7061,N_929,N_1917);
nand U7062 (N_7062,N_1574,N_2148);
or U7063 (N_7063,N_873,N_3373);
nand U7064 (N_7064,N_3164,N_2646);
nor U7065 (N_7065,N_820,N_2905);
nor U7066 (N_7066,N_2377,N_2926);
and U7067 (N_7067,N_3367,N_588);
xor U7068 (N_7068,N_2048,N_2347);
nor U7069 (N_7069,N_3374,N_3590);
nand U7070 (N_7070,N_3785,N_3496);
and U7071 (N_7071,N_2475,N_1880);
nor U7072 (N_7072,N_2351,N_1572);
nor U7073 (N_7073,N_2232,N_862);
xnor U7074 (N_7074,N_3563,N_1352);
or U7075 (N_7075,N_718,N_3609);
or U7076 (N_7076,N_1925,N_2937);
nand U7077 (N_7077,N_1513,N_730);
and U7078 (N_7078,N_3917,N_2731);
nor U7079 (N_7079,N_3695,N_667);
and U7080 (N_7080,N_2835,N_2389);
or U7081 (N_7081,N_331,N_2202);
nand U7082 (N_7082,N_42,N_1097);
and U7083 (N_7083,N_2472,N_3927);
nor U7084 (N_7084,N_2189,N_3831);
and U7085 (N_7085,N_917,N_1229);
nand U7086 (N_7086,N_3753,N_959);
or U7087 (N_7087,N_3408,N_1473);
xnor U7088 (N_7088,N_3069,N_1597);
nand U7089 (N_7089,N_3610,N_488);
xnor U7090 (N_7090,N_1071,N_2702);
nand U7091 (N_7091,N_2492,N_145);
or U7092 (N_7092,N_1181,N_2146);
nand U7093 (N_7093,N_1613,N_1709);
nand U7094 (N_7094,N_2677,N_1811);
nor U7095 (N_7095,N_492,N_926);
and U7096 (N_7096,N_2567,N_3311);
or U7097 (N_7097,N_3018,N_1427);
or U7098 (N_7098,N_3944,N_2415);
nor U7099 (N_7099,N_2911,N_3519);
nor U7100 (N_7100,N_3510,N_3156);
nand U7101 (N_7101,N_32,N_3325);
and U7102 (N_7102,N_1631,N_1915);
and U7103 (N_7103,N_351,N_308);
or U7104 (N_7104,N_1793,N_1943);
nor U7105 (N_7105,N_89,N_374);
and U7106 (N_7106,N_88,N_506);
or U7107 (N_7107,N_1132,N_430);
xor U7108 (N_7108,N_3220,N_1806);
xnor U7109 (N_7109,N_3878,N_1113);
xnor U7110 (N_7110,N_1050,N_646);
nand U7111 (N_7111,N_3417,N_3652);
or U7112 (N_7112,N_3344,N_77);
nand U7113 (N_7113,N_344,N_2765);
nor U7114 (N_7114,N_3928,N_877);
or U7115 (N_7115,N_254,N_638);
xor U7116 (N_7116,N_1842,N_2324);
nand U7117 (N_7117,N_1368,N_3887);
xnor U7118 (N_7118,N_805,N_617);
and U7119 (N_7119,N_3438,N_2951);
xor U7120 (N_7120,N_112,N_3478);
xnor U7121 (N_7121,N_23,N_1003);
and U7122 (N_7122,N_643,N_621);
and U7123 (N_7123,N_2385,N_720);
nor U7124 (N_7124,N_3522,N_2394);
nand U7125 (N_7125,N_2994,N_3024);
and U7126 (N_7126,N_3264,N_2405);
or U7127 (N_7127,N_3729,N_979);
or U7128 (N_7128,N_991,N_2265);
nor U7129 (N_7129,N_2646,N_1080);
or U7130 (N_7130,N_3878,N_1046);
and U7131 (N_7131,N_2634,N_1355);
or U7132 (N_7132,N_2649,N_3659);
nor U7133 (N_7133,N_3979,N_2835);
and U7134 (N_7134,N_475,N_1197);
nand U7135 (N_7135,N_3376,N_3448);
and U7136 (N_7136,N_3223,N_510);
xnor U7137 (N_7137,N_873,N_2532);
or U7138 (N_7138,N_1075,N_382);
xnor U7139 (N_7139,N_1903,N_2326);
or U7140 (N_7140,N_865,N_1294);
and U7141 (N_7141,N_1336,N_3821);
nand U7142 (N_7142,N_2036,N_3772);
nand U7143 (N_7143,N_1483,N_3056);
nor U7144 (N_7144,N_2177,N_1599);
and U7145 (N_7145,N_2271,N_530);
xor U7146 (N_7146,N_2884,N_3846);
xnor U7147 (N_7147,N_3570,N_460);
and U7148 (N_7148,N_321,N_999);
or U7149 (N_7149,N_901,N_1930);
xnor U7150 (N_7150,N_2760,N_3391);
and U7151 (N_7151,N_576,N_2593);
xor U7152 (N_7152,N_1484,N_2674);
or U7153 (N_7153,N_3201,N_2930);
and U7154 (N_7154,N_1714,N_1548);
nand U7155 (N_7155,N_2664,N_3407);
nor U7156 (N_7156,N_2892,N_2745);
nand U7157 (N_7157,N_2758,N_3492);
and U7158 (N_7158,N_3628,N_3661);
or U7159 (N_7159,N_3629,N_74);
or U7160 (N_7160,N_1710,N_662);
or U7161 (N_7161,N_1322,N_838);
nand U7162 (N_7162,N_33,N_3986);
nor U7163 (N_7163,N_3759,N_3884);
xor U7164 (N_7164,N_3924,N_2448);
and U7165 (N_7165,N_1892,N_898);
xnor U7166 (N_7166,N_3466,N_1907);
xnor U7167 (N_7167,N_79,N_2649);
nand U7168 (N_7168,N_3983,N_3465);
xor U7169 (N_7169,N_3270,N_508);
nand U7170 (N_7170,N_1280,N_543);
and U7171 (N_7171,N_1934,N_616);
or U7172 (N_7172,N_3929,N_1795);
nand U7173 (N_7173,N_1790,N_3872);
and U7174 (N_7174,N_2452,N_1118);
nor U7175 (N_7175,N_3903,N_1457);
and U7176 (N_7176,N_2949,N_1379);
and U7177 (N_7177,N_2252,N_2782);
xor U7178 (N_7178,N_3190,N_594);
nand U7179 (N_7179,N_1649,N_2970);
xnor U7180 (N_7180,N_3646,N_1043);
and U7181 (N_7181,N_243,N_2032);
xor U7182 (N_7182,N_3557,N_1498);
or U7183 (N_7183,N_3348,N_2554);
or U7184 (N_7184,N_3532,N_529);
nor U7185 (N_7185,N_1769,N_58);
or U7186 (N_7186,N_3230,N_1205);
or U7187 (N_7187,N_2845,N_3937);
and U7188 (N_7188,N_2649,N_389);
or U7189 (N_7189,N_1076,N_3702);
and U7190 (N_7190,N_199,N_3693);
xor U7191 (N_7191,N_3046,N_1654);
or U7192 (N_7192,N_502,N_3181);
and U7193 (N_7193,N_2111,N_3410);
nor U7194 (N_7194,N_3592,N_977);
nor U7195 (N_7195,N_658,N_1812);
and U7196 (N_7196,N_341,N_886);
nand U7197 (N_7197,N_1004,N_2707);
nor U7198 (N_7198,N_768,N_156);
xnor U7199 (N_7199,N_3491,N_371);
nor U7200 (N_7200,N_2437,N_151);
xor U7201 (N_7201,N_2317,N_1277);
or U7202 (N_7202,N_630,N_631);
or U7203 (N_7203,N_2468,N_2904);
nand U7204 (N_7204,N_3053,N_3577);
nand U7205 (N_7205,N_1089,N_3845);
xor U7206 (N_7206,N_1323,N_1428);
and U7207 (N_7207,N_213,N_1684);
nand U7208 (N_7208,N_3755,N_341);
xnor U7209 (N_7209,N_881,N_1446);
and U7210 (N_7210,N_3434,N_791);
xnor U7211 (N_7211,N_2908,N_2376);
and U7212 (N_7212,N_3694,N_2424);
xnor U7213 (N_7213,N_3311,N_1783);
or U7214 (N_7214,N_2247,N_1641);
nor U7215 (N_7215,N_392,N_3561);
or U7216 (N_7216,N_2103,N_1144);
nand U7217 (N_7217,N_2625,N_2887);
xor U7218 (N_7218,N_773,N_103);
or U7219 (N_7219,N_3988,N_974);
and U7220 (N_7220,N_2248,N_3075);
and U7221 (N_7221,N_1165,N_3911);
and U7222 (N_7222,N_2241,N_316);
nor U7223 (N_7223,N_869,N_2428);
xnor U7224 (N_7224,N_595,N_1115);
xor U7225 (N_7225,N_1098,N_2464);
nand U7226 (N_7226,N_1813,N_97);
and U7227 (N_7227,N_225,N_966);
or U7228 (N_7228,N_1763,N_2413);
and U7229 (N_7229,N_1774,N_1783);
nand U7230 (N_7230,N_1258,N_2234);
nand U7231 (N_7231,N_754,N_1499);
nor U7232 (N_7232,N_3576,N_2634);
nand U7233 (N_7233,N_1818,N_135);
nor U7234 (N_7234,N_2251,N_1488);
xor U7235 (N_7235,N_950,N_1086);
nand U7236 (N_7236,N_1654,N_1582);
xnor U7237 (N_7237,N_3661,N_3866);
xnor U7238 (N_7238,N_840,N_108);
xor U7239 (N_7239,N_3400,N_1265);
nand U7240 (N_7240,N_3488,N_3730);
xor U7241 (N_7241,N_501,N_295);
nand U7242 (N_7242,N_3879,N_455);
and U7243 (N_7243,N_994,N_640);
nor U7244 (N_7244,N_1946,N_3352);
or U7245 (N_7245,N_1230,N_2040);
xor U7246 (N_7246,N_3238,N_3158);
xor U7247 (N_7247,N_377,N_692);
xor U7248 (N_7248,N_3622,N_3997);
xnor U7249 (N_7249,N_1238,N_849);
xor U7250 (N_7250,N_2398,N_2120);
or U7251 (N_7251,N_87,N_1518);
and U7252 (N_7252,N_75,N_2519);
nand U7253 (N_7253,N_23,N_139);
or U7254 (N_7254,N_960,N_832);
nor U7255 (N_7255,N_2967,N_786);
nor U7256 (N_7256,N_2132,N_1511);
and U7257 (N_7257,N_2116,N_3843);
and U7258 (N_7258,N_53,N_1588);
nand U7259 (N_7259,N_1425,N_550);
and U7260 (N_7260,N_2152,N_1321);
nor U7261 (N_7261,N_161,N_37);
nand U7262 (N_7262,N_3130,N_3957);
and U7263 (N_7263,N_3745,N_376);
xnor U7264 (N_7264,N_2523,N_3791);
nand U7265 (N_7265,N_626,N_2593);
nand U7266 (N_7266,N_1766,N_2076);
and U7267 (N_7267,N_2683,N_3634);
nand U7268 (N_7268,N_918,N_1983);
xnor U7269 (N_7269,N_3882,N_2239);
xnor U7270 (N_7270,N_1486,N_1527);
xor U7271 (N_7271,N_479,N_618);
or U7272 (N_7272,N_240,N_189);
xnor U7273 (N_7273,N_3445,N_2655);
and U7274 (N_7274,N_1607,N_2361);
or U7275 (N_7275,N_328,N_762);
nand U7276 (N_7276,N_608,N_3355);
nand U7277 (N_7277,N_3047,N_1929);
xor U7278 (N_7278,N_2217,N_645);
and U7279 (N_7279,N_1029,N_2520);
xnor U7280 (N_7280,N_574,N_1956);
xnor U7281 (N_7281,N_1970,N_323);
nand U7282 (N_7282,N_1342,N_773);
nor U7283 (N_7283,N_1681,N_1659);
nor U7284 (N_7284,N_1044,N_881);
nand U7285 (N_7285,N_2810,N_3964);
xor U7286 (N_7286,N_2107,N_1620);
nand U7287 (N_7287,N_805,N_3101);
and U7288 (N_7288,N_3181,N_1910);
or U7289 (N_7289,N_1190,N_3304);
nor U7290 (N_7290,N_3084,N_2316);
nand U7291 (N_7291,N_2711,N_2102);
nor U7292 (N_7292,N_1917,N_2536);
or U7293 (N_7293,N_1558,N_1973);
nand U7294 (N_7294,N_20,N_803);
nor U7295 (N_7295,N_2802,N_2229);
xor U7296 (N_7296,N_2089,N_2718);
and U7297 (N_7297,N_1937,N_3618);
nand U7298 (N_7298,N_192,N_1411);
xor U7299 (N_7299,N_3400,N_3349);
nand U7300 (N_7300,N_1955,N_1799);
xor U7301 (N_7301,N_1944,N_326);
and U7302 (N_7302,N_2159,N_2558);
or U7303 (N_7303,N_1627,N_3709);
nor U7304 (N_7304,N_1946,N_929);
and U7305 (N_7305,N_2961,N_1751);
and U7306 (N_7306,N_2035,N_2671);
xor U7307 (N_7307,N_152,N_1273);
and U7308 (N_7308,N_1181,N_3407);
and U7309 (N_7309,N_252,N_3656);
and U7310 (N_7310,N_2718,N_3542);
xor U7311 (N_7311,N_912,N_824);
nor U7312 (N_7312,N_3956,N_3336);
xor U7313 (N_7313,N_473,N_3428);
and U7314 (N_7314,N_1304,N_1952);
nor U7315 (N_7315,N_831,N_2857);
nor U7316 (N_7316,N_3222,N_2113);
nor U7317 (N_7317,N_3555,N_2628);
nand U7318 (N_7318,N_1309,N_2065);
nand U7319 (N_7319,N_3291,N_90);
xor U7320 (N_7320,N_1219,N_3511);
nand U7321 (N_7321,N_1960,N_1815);
nor U7322 (N_7322,N_3462,N_3344);
nor U7323 (N_7323,N_1321,N_2499);
and U7324 (N_7324,N_775,N_2963);
or U7325 (N_7325,N_3638,N_3645);
and U7326 (N_7326,N_468,N_1410);
and U7327 (N_7327,N_2251,N_548);
xor U7328 (N_7328,N_2969,N_1222);
nor U7329 (N_7329,N_290,N_463);
and U7330 (N_7330,N_3436,N_2989);
or U7331 (N_7331,N_1926,N_802);
or U7332 (N_7332,N_551,N_231);
nand U7333 (N_7333,N_785,N_3943);
or U7334 (N_7334,N_2204,N_2244);
nor U7335 (N_7335,N_1792,N_3829);
or U7336 (N_7336,N_105,N_1962);
and U7337 (N_7337,N_3217,N_3992);
and U7338 (N_7338,N_2727,N_1008);
nand U7339 (N_7339,N_3260,N_1910);
nand U7340 (N_7340,N_2179,N_614);
nor U7341 (N_7341,N_3423,N_1508);
or U7342 (N_7342,N_2486,N_3887);
and U7343 (N_7343,N_3743,N_415);
nand U7344 (N_7344,N_316,N_3675);
or U7345 (N_7345,N_1319,N_3861);
nand U7346 (N_7346,N_3524,N_1873);
or U7347 (N_7347,N_2517,N_2044);
nand U7348 (N_7348,N_1698,N_77);
nand U7349 (N_7349,N_2608,N_152);
nand U7350 (N_7350,N_392,N_2369);
xnor U7351 (N_7351,N_2900,N_3302);
or U7352 (N_7352,N_518,N_1168);
nor U7353 (N_7353,N_3243,N_3436);
xor U7354 (N_7354,N_1269,N_648);
and U7355 (N_7355,N_3603,N_3306);
or U7356 (N_7356,N_3852,N_1448);
nand U7357 (N_7357,N_3784,N_1846);
nor U7358 (N_7358,N_317,N_3950);
or U7359 (N_7359,N_1773,N_469);
xor U7360 (N_7360,N_586,N_2384);
xor U7361 (N_7361,N_2722,N_2860);
nand U7362 (N_7362,N_46,N_448);
or U7363 (N_7363,N_1925,N_271);
and U7364 (N_7364,N_713,N_2308);
and U7365 (N_7365,N_65,N_3063);
and U7366 (N_7366,N_1116,N_527);
nor U7367 (N_7367,N_2054,N_2280);
nor U7368 (N_7368,N_1244,N_2036);
xor U7369 (N_7369,N_883,N_2258);
and U7370 (N_7370,N_1994,N_1840);
or U7371 (N_7371,N_529,N_276);
or U7372 (N_7372,N_1543,N_1221);
xor U7373 (N_7373,N_2847,N_2882);
or U7374 (N_7374,N_1802,N_979);
and U7375 (N_7375,N_714,N_3854);
or U7376 (N_7376,N_890,N_1774);
xor U7377 (N_7377,N_2994,N_2022);
nor U7378 (N_7378,N_638,N_3336);
and U7379 (N_7379,N_3183,N_2704);
or U7380 (N_7380,N_3827,N_3092);
nor U7381 (N_7381,N_96,N_234);
xor U7382 (N_7382,N_1635,N_3631);
and U7383 (N_7383,N_888,N_876);
nor U7384 (N_7384,N_1846,N_103);
xor U7385 (N_7385,N_1775,N_897);
and U7386 (N_7386,N_1663,N_781);
nand U7387 (N_7387,N_1777,N_554);
xnor U7388 (N_7388,N_2127,N_3666);
nor U7389 (N_7389,N_1229,N_2776);
or U7390 (N_7390,N_3267,N_1881);
nor U7391 (N_7391,N_156,N_2004);
and U7392 (N_7392,N_1945,N_3726);
nor U7393 (N_7393,N_329,N_2605);
nand U7394 (N_7394,N_3024,N_1732);
or U7395 (N_7395,N_673,N_3155);
and U7396 (N_7396,N_2429,N_1644);
nand U7397 (N_7397,N_2745,N_51);
and U7398 (N_7398,N_864,N_3593);
nor U7399 (N_7399,N_1456,N_2149);
xnor U7400 (N_7400,N_3120,N_195);
nand U7401 (N_7401,N_2852,N_1466);
nand U7402 (N_7402,N_447,N_704);
nand U7403 (N_7403,N_1842,N_1426);
nor U7404 (N_7404,N_2806,N_3334);
and U7405 (N_7405,N_302,N_924);
xor U7406 (N_7406,N_851,N_3189);
or U7407 (N_7407,N_3821,N_2038);
or U7408 (N_7408,N_1549,N_1240);
nor U7409 (N_7409,N_3957,N_2857);
and U7410 (N_7410,N_1023,N_3789);
or U7411 (N_7411,N_23,N_747);
nor U7412 (N_7412,N_1903,N_611);
xnor U7413 (N_7413,N_2394,N_1319);
or U7414 (N_7414,N_2528,N_2433);
or U7415 (N_7415,N_2458,N_3573);
nand U7416 (N_7416,N_3299,N_1928);
nand U7417 (N_7417,N_1530,N_181);
or U7418 (N_7418,N_3466,N_1366);
nand U7419 (N_7419,N_1329,N_3054);
or U7420 (N_7420,N_2147,N_2231);
nor U7421 (N_7421,N_3686,N_2899);
nor U7422 (N_7422,N_1703,N_2687);
and U7423 (N_7423,N_114,N_3093);
nand U7424 (N_7424,N_1093,N_2003);
nand U7425 (N_7425,N_2791,N_2269);
nand U7426 (N_7426,N_3723,N_2685);
xnor U7427 (N_7427,N_2328,N_520);
or U7428 (N_7428,N_3066,N_1751);
nand U7429 (N_7429,N_3579,N_2960);
nand U7430 (N_7430,N_916,N_1944);
nand U7431 (N_7431,N_221,N_2871);
nand U7432 (N_7432,N_3480,N_1528);
xnor U7433 (N_7433,N_3086,N_2255);
xnor U7434 (N_7434,N_1323,N_1876);
nor U7435 (N_7435,N_3244,N_3959);
nand U7436 (N_7436,N_1968,N_2597);
nor U7437 (N_7437,N_2756,N_1771);
xor U7438 (N_7438,N_3830,N_2975);
and U7439 (N_7439,N_813,N_3415);
xor U7440 (N_7440,N_3775,N_3490);
and U7441 (N_7441,N_2805,N_1055);
nand U7442 (N_7442,N_1748,N_3378);
nor U7443 (N_7443,N_3680,N_3014);
nand U7444 (N_7444,N_1209,N_2980);
xor U7445 (N_7445,N_820,N_1247);
and U7446 (N_7446,N_3790,N_3356);
xor U7447 (N_7447,N_3711,N_1570);
or U7448 (N_7448,N_328,N_2023);
nand U7449 (N_7449,N_3803,N_147);
nand U7450 (N_7450,N_2876,N_41);
xnor U7451 (N_7451,N_3288,N_2822);
or U7452 (N_7452,N_2323,N_2295);
and U7453 (N_7453,N_946,N_1908);
nand U7454 (N_7454,N_1942,N_7);
xnor U7455 (N_7455,N_644,N_1021);
or U7456 (N_7456,N_737,N_2310);
xor U7457 (N_7457,N_3092,N_2682);
and U7458 (N_7458,N_2604,N_1809);
nand U7459 (N_7459,N_54,N_455);
xnor U7460 (N_7460,N_1951,N_2662);
nand U7461 (N_7461,N_2173,N_3352);
nand U7462 (N_7462,N_2777,N_106);
nor U7463 (N_7463,N_33,N_1237);
xnor U7464 (N_7464,N_2437,N_1827);
nor U7465 (N_7465,N_1909,N_1928);
xnor U7466 (N_7466,N_380,N_434);
xor U7467 (N_7467,N_3079,N_469);
and U7468 (N_7468,N_3442,N_3217);
nor U7469 (N_7469,N_2143,N_677);
nor U7470 (N_7470,N_3851,N_1613);
nor U7471 (N_7471,N_3253,N_238);
nand U7472 (N_7472,N_3646,N_2625);
nand U7473 (N_7473,N_3781,N_3930);
xor U7474 (N_7474,N_971,N_3377);
nor U7475 (N_7475,N_1504,N_3442);
nand U7476 (N_7476,N_2051,N_1114);
and U7477 (N_7477,N_3045,N_3473);
nand U7478 (N_7478,N_2225,N_2775);
or U7479 (N_7479,N_528,N_434);
or U7480 (N_7480,N_2125,N_2334);
nand U7481 (N_7481,N_1531,N_713);
and U7482 (N_7482,N_2450,N_2291);
nand U7483 (N_7483,N_2233,N_2202);
nor U7484 (N_7484,N_1821,N_3829);
nor U7485 (N_7485,N_3484,N_3127);
nand U7486 (N_7486,N_362,N_2433);
nand U7487 (N_7487,N_2866,N_780);
xor U7488 (N_7488,N_3474,N_2960);
nand U7489 (N_7489,N_1408,N_1453);
or U7490 (N_7490,N_3946,N_2830);
nor U7491 (N_7491,N_1817,N_1161);
nor U7492 (N_7492,N_1033,N_1551);
nor U7493 (N_7493,N_3676,N_464);
nand U7494 (N_7494,N_1399,N_357);
xor U7495 (N_7495,N_1408,N_2897);
and U7496 (N_7496,N_1807,N_3573);
nor U7497 (N_7497,N_320,N_1949);
xor U7498 (N_7498,N_728,N_472);
and U7499 (N_7499,N_1967,N_1928);
and U7500 (N_7500,N_672,N_1773);
nor U7501 (N_7501,N_2930,N_1072);
and U7502 (N_7502,N_2230,N_1294);
xnor U7503 (N_7503,N_1319,N_1795);
xor U7504 (N_7504,N_3583,N_821);
nand U7505 (N_7505,N_361,N_854);
nor U7506 (N_7506,N_208,N_3212);
and U7507 (N_7507,N_2546,N_618);
or U7508 (N_7508,N_870,N_3650);
or U7509 (N_7509,N_1534,N_3001);
nor U7510 (N_7510,N_445,N_3188);
xor U7511 (N_7511,N_1582,N_1563);
nor U7512 (N_7512,N_2846,N_3648);
or U7513 (N_7513,N_960,N_55);
nor U7514 (N_7514,N_21,N_117);
and U7515 (N_7515,N_1414,N_2471);
xor U7516 (N_7516,N_2558,N_2964);
nor U7517 (N_7517,N_707,N_3286);
and U7518 (N_7518,N_272,N_1309);
and U7519 (N_7519,N_252,N_321);
nand U7520 (N_7520,N_2707,N_1992);
and U7521 (N_7521,N_3219,N_849);
xor U7522 (N_7522,N_295,N_2985);
or U7523 (N_7523,N_540,N_682);
or U7524 (N_7524,N_1632,N_2522);
nand U7525 (N_7525,N_1608,N_3102);
nand U7526 (N_7526,N_3659,N_2707);
nand U7527 (N_7527,N_2093,N_656);
and U7528 (N_7528,N_1505,N_3827);
nand U7529 (N_7529,N_844,N_294);
or U7530 (N_7530,N_2451,N_1361);
and U7531 (N_7531,N_2910,N_2399);
xor U7532 (N_7532,N_3440,N_778);
or U7533 (N_7533,N_1562,N_3461);
xor U7534 (N_7534,N_655,N_3835);
and U7535 (N_7535,N_3770,N_163);
and U7536 (N_7536,N_3184,N_2282);
nor U7537 (N_7537,N_804,N_3681);
nor U7538 (N_7538,N_1940,N_419);
and U7539 (N_7539,N_3551,N_3936);
xor U7540 (N_7540,N_637,N_501);
or U7541 (N_7541,N_304,N_2086);
nand U7542 (N_7542,N_920,N_3351);
and U7543 (N_7543,N_71,N_1369);
or U7544 (N_7544,N_3042,N_781);
or U7545 (N_7545,N_1531,N_807);
and U7546 (N_7546,N_139,N_861);
nand U7547 (N_7547,N_2011,N_3295);
or U7548 (N_7548,N_3498,N_2532);
nand U7549 (N_7549,N_1185,N_1262);
or U7550 (N_7550,N_2165,N_584);
or U7551 (N_7551,N_1342,N_2218);
or U7552 (N_7552,N_3285,N_479);
nor U7553 (N_7553,N_1086,N_3297);
or U7554 (N_7554,N_3667,N_3310);
or U7555 (N_7555,N_1370,N_1634);
nand U7556 (N_7556,N_3657,N_3904);
nand U7557 (N_7557,N_1070,N_3761);
nand U7558 (N_7558,N_1654,N_2267);
nand U7559 (N_7559,N_3030,N_2821);
and U7560 (N_7560,N_3870,N_2309);
xnor U7561 (N_7561,N_3971,N_1836);
and U7562 (N_7562,N_2080,N_3556);
xnor U7563 (N_7563,N_2809,N_31);
nor U7564 (N_7564,N_3970,N_150);
or U7565 (N_7565,N_1936,N_2540);
nor U7566 (N_7566,N_1751,N_1701);
nand U7567 (N_7567,N_3728,N_878);
or U7568 (N_7568,N_2395,N_1554);
xnor U7569 (N_7569,N_1247,N_644);
or U7570 (N_7570,N_3385,N_2047);
xnor U7571 (N_7571,N_526,N_3027);
xor U7572 (N_7572,N_3416,N_1137);
nand U7573 (N_7573,N_2048,N_1362);
and U7574 (N_7574,N_1896,N_34);
or U7575 (N_7575,N_1465,N_3462);
or U7576 (N_7576,N_3512,N_3551);
and U7577 (N_7577,N_3280,N_3401);
and U7578 (N_7578,N_1909,N_383);
xnor U7579 (N_7579,N_1626,N_1591);
nand U7580 (N_7580,N_2816,N_3481);
nand U7581 (N_7581,N_1400,N_3000);
xor U7582 (N_7582,N_2413,N_3515);
and U7583 (N_7583,N_2170,N_236);
nand U7584 (N_7584,N_1781,N_3723);
or U7585 (N_7585,N_2952,N_3595);
xnor U7586 (N_7586,N_3367,N_3981);
and U7587 (N_7587,N_1776,N_597);
nand U7588 (N_7588,N_3135,N_2107);
or U7589 (N_7589,N_1888,N_2134);
or U7590 (N_7590,N_2395,N_3838);
and U7591 (N_7591,N_1182,N_2134);
xnor U7592 (N_7592,N_2633,N_837);
xnor U7593 (N_7593,N_1504,N_2306);
or U7594 (N_7594,N_100,N_1219);
or U7595 (N_7595,N_3997,N_1861);
nand U7596 (N_7596,N_1944,N_1425);
and U7597 (N_7597,N_1312,N_996);
nor U7598 (N_7598,N_2557,N_938);
and U7599 (N_7599,N_4,N_1267);
nand U7600 (N_7600,N_3262,N_2572);
xor U7601 (N_7601,N_958,N_971);
xnor U7602 (N_7602,N_2846,N_3651);
nor U7603 (N_7603,N_2783,N_648);
xor U7604 (N_7604,N_1765,N_2601);
xor U7605 (N_7605,N_2518,N_117);
nor U7606 (N_7606,N_883,N_3848);
nor U7607 (N_7607,N_915,N_1991);
xor U7608 (N_7608,N_3591,N_2204);
nand U7609 (N_7609,N_3279,N_1786);
and U7610 (N_7610,N_2975,N_830);
or U7611 (N_7611,N_1169,N_3653);
and U7612 (N_7612,N_3925,N_338);
nor U7613 (N_7613,N_3872,N_994);
or U7614 (N_7614,N_3227,N_93);
nor U7615 (N_7615,N_1349,N_2457);
nor U7616 (N_7616,N_3870,N_3389);
nor U7617 (N_7617,N_3544,N_1286);
or U7618 (N_7618,N_2847,N_2502);
and U7619 (N_7619,N_2576,N_911);
nand U7620 (N_7620,N_1937,N_170);
nor U7621 (N_7621,N_1414,N_670);
nand U7622 (N_7622,N_2387,N_295);
nand U7623 (N_7623,N_947,N_1343);
xor U7624 (N_7624,N_3031,N_3115);
xnor U7625 (N_7625,N_387,N_1156);
xor U7626 (N_7626,N_2433,N_3562);
nor U7627 (N_7627,N_2486,N_619);
xor U7628 (N_7628,N_3560,N_1611);
and U7629 (N_7629,N_2222,N_684);
and U7630 (N_7630,N_2983,N_3788);
nor U7631 (N_7631,N_3624,N_1444);
and U7632 (N_7632,N_2999,N_1414);
nor U7633 (N_7633,N_1532,N_1046);
and U7634 (N_7634,N_1562,N_2209);
nand U7635 (N_7635,N_2603,N_2380);
nand U7636 (N_7636,N_298,N_3312);
nand U7637 (N_7637,N_739,N_3645);
or U7638 (N_7638,N_2090,N_1524);
nor U7639 (N_7639,N_1889,N_9);
and U7640 (N_7640,N_948,N_737);
and U7641 (N_7641,N_2895,N_1541);
xnor U7642 (N_7642,N_2594,N_3320);
xnor U7643 (N_7643,N_2155,N_1260);
or U7644 (N_7644,N_821,N_633);
or U7645 (N_7645,N_716,N_1459);
or U7646 (N_7646,N_2308,N_761);
nor U7647 (N_7647,N_1989,N_2846);
and U7648 (N_7648,N_1111,N_184);
xor U7649 (N_7649,N_2408,N_1565);
and U7650 (N_7650,N_2533,N_2375);
nor U7651 (N_7651,N_2351,N_1238);
nor U7652 (N_7652,N_3727,N_3440);
nand U7653 (N_7653,N_3988,N_1934);
or U7654 (N_7654,N_3779,N_3764);
nand U7655 (N_7655,N_2898,N_3853);
xor U7656 (N_7656,N_907,N_1798);
xnor U7657 (N_7657,N_1001,N_3708);
and U7658 (N_7658,N_1766,N_2129);
xnor U7659 (N_7659,N_1151,N_715);
or U7660 (N_7660,N_599,N_1350);
xnor U7661 (N_7661,N_3351,N_1285);
xnor U7662 (N_7662,N_2849,N_1315);
nand U7663 (N_7663,N_1769,N_3812);
or U7664 (N_7664,N_3715,N_308);
nor U7665 (N_7665,N_3049,N_861);
or U7666 (N_7666,N_1234,N_569);
nand U7667 (N_7667,N_3220,N_1899);
and U7668 (N_7668,N_2310,N_2434);
or U7669 (N_7669,N_162,N_2263);
and U7670 (N_7670,N_3163,N_2731);
nand U7671 (N_7671,N_1609,N_600);
or U7672 (N_7672,N_2212,N_3749);
and U7673 (N_7673,N_1678,N_1725);
or U7674 (N_7674,N_335,N_3026);
nand U7675 (N_7675,N_63,N_1664);
or U7676 (N_7676,N_1673,N_3152);
nand U7677 (N_7677,N_0,N_2470);
xnor U7678 (N_7678,N_1128,N_703);
or U7679 (N_7679,N_2889,N_383);
nand U7680 (N_7680,N_3811,N_1565);
or U7681 (N_7681,N_1944,N_657);
and U7682 (N_7682,N_963,N_2248);
nand U7683 (N_7683,N_2188,N_173);
or U7684 (N_7684,N_1690,N_2222);
and U7685 (N_7685,N_3654,N_2909);
nor U7686 (N_7686,N_3578,N_2772);
xnor U7687 (N_7687,N_3201,N_3205);
nor U7688 (N_7688,N_2194,N_1676);
nand U7689 (N_7689,N_3212,N_3345);
nand U7690 (N_7690,N_939,N_265);
xnor U7691 (N_7691,N_1151,N_482);
xor U7692 (N_7692,N_2179,N_3322);
nor U7693 (N_7693,N_488,N_97);
xnor U7694 (N_7694,N_1918,N_3263);
and U7695 (N_7695,N_1652,N_3864);
nor U7696 (N_7696,N_2436,N_2630);
nor U7697 (N_7697,N_1428,N_125);
and U7698 (N_7698,N_3076,N_528);
nand U7699 (N_7699,N_2247,N_1648);
nor U7700 (N_7700,N_3641,N_2554);
and U7701 (N_7701,N_1716,N_3017);
xnor U7702 (N_7702,N_1274,N_3957);
xnor U7703 (N_7703,N_2371,N_3751);
nor U7704 (N_7704,N_3779,N_3511);
nand U7705 (N_7705,N_2192,N_1312);
nor U7706 (N_7706,N_3150,N_2998);
and U7707 (N_7707,N_753,N_3440);
nor U7708 (N_7708,N_621,N_845);
nor U7709 (N_7709,N_3317,N_658);
and U7710 (N_7710,N_1956,N_445);
nand U7711 (N_7711,N_2120,N_220);
xor U7712 (N_7712,N_2051,N_2686);
nand U7713 (N_7713,N_3796,N_389);
or U7714 (N_7714,N_1439,N_2108);
nand U7715 (N_7715,N_2463,N_3141);
xor U7716 (N_7716,N_2194,N_3750);
nor U7717 (N_7717,N_3216,N_3142);
and U7718 (N_7718,N_101,N_2128);
nand U7719 (N_7719,N_3193,N_2480);
nand U7720 (N_7720,N_3662,N_1007);
or U7721 (N_7721,N_1118,N_2268);
nand U7722 (N_7722,N_1579,N_1253);
nand U7723 (N_7723,N_3703,N_1150);
xnor U7724 (N_7724,N_3001,N_2514);
and U7725 (N_7725,N_29,N_355);
and U7726 (N_7726,N_2612,N_621);
xor U7727 (N_7727,N_2462,N_3462);
nor U7728 (N_7728,N_619,N_2140);
and U7729 (N_7729,N_3561,N_2676);
nor U7730 (N_7730,N_3082,N_2945);
xor U7731 (N_7731,N_210,N_3472);
nand U7732 (N_7732,N_2434,N_2112);
nand U7733 (N_7733,N_98,N_2971);
nor U7734 (N_7734,N_283,N_2585);
and U7735 (N_7735,N_2364,N_2014);
nand U7736 (N_7736,N_2336,N_1762);
xnor U7737 (N_7737,N_601,N_2178);
nand U7738 (N_7738,N_670,N_449);
xnor U7739 (N_7739,N_1651,N_3436);
xor U7740 (N_7740,N_2518,N_899);
nor U7741 (N_7741,N_1342,N_3492);
nand U7742 (N_7742,N_3162,N_2889);
xor U7743 (N_7743,N_2986,N_796);
nand U7744 (N_7744,N_1095,N_3335);
or U7745 (N_7745,N_2145,N_423);
nand U7746 (N_7746,N_2167,N_225);
nor U7747 (N_7747,N_3128,N_3238);
nand U7748 (N_7748,N_1147,N_1028);
or U7749 (N_7749,N_1148,N_2098);
nor U7750 (N_7750,N_1872,N_2799);
xor U7751 (N_7751,N_531,N_2562);
xor U7752 (N_7752,N_32,N_832);
nor U7753 (N_7753,N_441,N_3667);
xnor U7754 (N_7754,N_3172,N_1859);
xnor U7755 (N_7755,N_2456,N_2256);
or U7756 (N_7756,N_2749,N_1774);
nand U7757 (N_7757,N_359,N_727);
xnor U7758 (N_7758,N_2569,N_3065);
nand U7759 (N_7759,N_3549,N_2234);
nand U7760 (N_7760,N_2559,N_3940);
nor U7761 (N_7761,N_3363,N_1329);
nor U7762 (N_7762,N_526,N_1294);
nand U7763 (N_7763,N_2151,N_1220);
xor U7764 (N_7764,N_3071,N_309);
nand U7765 (N_7765,N_2684,N_3863);
nor U7766 (N_7766,N_304,N_708);
nand U7767 (N_7767,N_2627,N_3233);
xor U7768 (N_7768,N_2299,N_3323);
or U7769 (N_7769,N_3006,N_326);
or U7770 (N_7770,N_2826,N_688);
xor U7771 (N_7771,N_2421,N_1382);
nand U7772 (N_7772,N_1965,N_3471);
nor U7773 (N_7773,N_891,N_3378);
or U7774 (N_7774,N_2399,N_3648);
nand U7775 (N_7775,N_788,N_3336);
xnor U7776 (N_7776,N_3667,N_600);
nor U7777 (N_7777,N_3661,N_2846);
and U7778 (N_7778,N_3655,N_1750);
xnor U7779 (N_7779,N_1438,N_2966);
or U7780 (N_7780,N_3542,N_1480);
and U7781 (N_7781,N_3365,N_1075);
or U7782 (N_7782,N_615,N_490);
xor U7783 (N_7783,N_2977,N_3753);
or U7784 (N_7784,N_1300,N_847);
or U7785 (N_7785,N_3304,N_593);
nand U7786 (N_7786,N_1693,N_1819);
and U7787 (N_7787,N_949,N_2719);
and U7788 (N_7788,N_2190,N_1704);
and U7789 (N_7789,N_799,N_1934);
or U7790 (N_7790,N_2142,N_998);
or U7791 (N_7791,N_2131,N_1881);
and U7792 (N_7792,N_3670,N_543);
nor U7793 (N_7793,N_346,N_1546);
nand U7794 (N_7794,N_2666,N_2386);
nor U7795 (N_7795,N_673,N_720);
and U7796 (N_7796,N_2802,N_1826);
nand U7797 (N_7797,N_503,N_1803);
xor U7798 (N_7798,N_104,N_2704);
nand U7799 (N_7799,N_2180,N_696);
or U7800 (N_7800,N_3489,N_3451);
and U7801 (N_7801,N_1709,N_2827);
xnor U7802 (N_7802,N_2091,N_3951);
nand U7803 (N_7803,N_1083,N_2001);
nand U7804 (N_7804,N_3925,N_3408);
and U7805 (N_7805,N_1310,N_2515);
nand U7806 (N_7806,N_2006,N_3467);
or U7807 (N_7807,N_210,N_59);
or U7808 (N_7808,N_630,N_2794);
xor U7809 (N_7809,N_326,N_1857);
nor U7810 (N_7810,N_3271,N_573);
and U7811 (N_7811,N_543,N_2664);
xnor U7812 (N_7812,N_2178,N_2406);
and U7813 (N_7813,N_654,N_2313);
and U7814 (N_7814,N_3815,N_2689);
nor U7815 (N_7815,N_29,N_2193);
nor U7816 (N_7816,N_3082,N_1779);
xor U7817 (N_7817,N_382,N_764);
or U7818 (N_7818,N_324,N_1737);
nor U7819 (N_7819,N_3099,N_3370);
nor U7820 (N_7820,N_1313,N_1502);
xor U7821 (N_7821,N_343,N_762);
or U7822 (N_7822,N_445,N_1143);
nor U7823 (N_7823,N_3239,N_3794);
nor U7824 (N_7824,N_1954,N_1564);
xor U7825 (N_7825,N_2695,N_3050);
nor U7826 (N_7826,N_833,N_2223);
xnor U7827 (N_7827,N_3404,N_195);
or U7828 (N_7828,N_1055,N_264);
xnor U7829 (N_7829,N_1689,N_3847);
xnor U7830 (N_7830,N_2758,N_2121);
xor U7831 (N_7831,N_1680,N_1987);
or U7832 (N_7832,N_1315,N_2803);
and U7833 (N_7833,N_3870,N_3098);
nand U7834 (N_7834,N_3243,N_2442);
nand U7835 (N_7835,N_1744,N_3909);
nand U7836 (N_7836,N_3608,N_3504);
and U7837 (N_7837,N_3420,N_570);
xnor U7838 (N_7838,N_1850,N_1529);
xor U7839 (N_7839,N_3078,N_1597);
xor U7840 (N_7840,N_336,N_2231);
or U7841 (N_7841,N_1409,N_1277);
and U7842 (N_7842,N_2576,N_1493);
or U7843 (N_7843,N_688,N_3832);
nor U7844 (N_7844,N_3859,N_2582);
nand U7845 (N_7845,N_1651,N_3049);
and U7846 (N_7846,N_3578,N_3047);
nand U7847 (N_7847,N_2414,N_3771);
or U7848 (N_7848,N_2864,N_3213);
nor U7849 (N_7849,N_466,N_2182);
and U7850 (N_7850,N_1438,N_2353);
xnor U7851 (N_7851,N_3615,N_3700);
or U7852 (N_7852,N_2948,N_3185);
or U7853 (N_7853,N_2833,N_1271);
xnor U7854 (N_7854,N_3850,N_753);
or U7855 (N_7855,N_3467,N_2550);
nor U7856 (N_7856,N_1147,N_587);
nor U7857 (N_7857,N_2466,N_392);
nand U7858 (N_7858,N_436,N_2979);
and U7859 (N_7859,N_3611,N_146);
and U7860 (N_7860,N_1013,N_1119);
and U7861 (N_7861,N_3408,N_2704);
nor U7862 (N_7862,N_2728,N_2224);
or U7863 (N_7863,N_2614,N_1751);
xor U7864 (N_7864,N_2245,N_892);
nand U7865 (N_7865,N_1569,N_919);
or U7866 (N_7866,N_1037,N_1618);
xor U7867 (N_7867,N_276,N_1475);
nor U7868 (N_7868,N_885,N_2849);
nor U7869 (N_7869,N_599,N_162);
xnor U7870 (N_7870,N_2883,N_2017);
xnor U7871 (N_7871,N_342,N_3071);
nand U7872 (N_7872,N_934,N_2101);
and U7873 (N_7873,N_663,N_3014);
and U7874 (N_7874,N_859,N_1703);
nand U7875 (N_7875,N_3168,N_1650);
or U7876 (N_7876,N_2548,N_1246);
nand U7877 (N_7877,N_273,N_3667);
or U7878 (N_7878,N_1237,N_1420);
and U7879 (N_7879,N_296,N_3230);
nand U7880 (N_7880,N_1609,N_2017);
nand U7881 (N_7881,N_1607,N_3174);
nand U7882 (N_7882,N_1550,N_3696);
or U7883 (N_7883,N_1324,N_776);
nor U7884 (N_7884,N_44,N_1863);
or U7885 (N_7885,N_1080,N_1631);
xnor U7886 (N_7886,N_193,N_3740);
nor U7887 (N_7887,N_3449,N_325);
or U7888 (N_7888,N_234,N_3858);
nor U7889 (N_7889,N_2559,N_1505);
nand U7890 (N_7890,N_648,N_734);
xnor U7891 (N_7891,N_3698,N_3066);
nor U7892 (N_7892,N_1399,N_111);
nor U7893 (N_7893,N_3123,N_1632);
nor U7894 (N_7894,N_34,N_3963);
nand U7895 (N_7895,N_178,N_2486);
nand U7896 (N_7896,N_3968,N_1843);
and U7897 (N_7897,N_2323,N_2670);
xnor U7898 (N_7898,N_2631,N_163);
nand U7899 (N_7899,N_3804,N_372);
or U7900 (N_7900,N_3990,N_1588);
and U7901 (N_7901,N_3753,N_1177);
xor U7902 (N_7902,N_1141,N_2527);
or U7903 (N_7903,N_2768,N_1461);
and U7904 (N_7904,N_728,N_2777);
xnor U7905 (N_7905,N_1974,N_3645);
and U7906 (N_7906,N_2726,N_2697);
or U7907 (N_7907,N_3584,N_2885);
nand U7908 (N_7908,N_1158,N_3086);
and U7909 (N_7909,N_313,N_75);
nor U7910 (N_7910,N_1109,N_1517);
or U7911 (N_7911,N_3500,N_1226);
and U7912 (N_7912,N_1211,N_752);
xnor U7913 (N_7913,N_3370,N_1756);
or U7914 (N_7914,N_2782,N_2923);
and U7915 (N_7915,N_1854,N_3478);
and U7916 (N_7916,N_842,N_3247);
nor U7917 (N_7917,N_1017,N_3125);
and U7918 (N_7918,N_1731,N_2324);
or U7919 (N_7919,N_1147,N_3431);
nor U7920 (N_7920,N_874,N_516);
nor U7921 (N_7921,N_2684,N_272);
nand U7922 (N_7922,N_3064,N_2022);
nor U7923 (N_7923,N_1365,N_3614);
nand U7924 (N_7924,N_3738,N_2859);
xnor U7925 (N_7925,N_380,N_527);
and U7926 (N_7926,N_1240,N_3575);
nand U7927 (N_7927,N_2383,N_1708);
nand U7928 (N_7928,N_784,N_1148);
and U7929 (N_7929,N_1262,N_192);
nor U7930 (N_7930,N_1259,N_2356);
xor U7931 (N_7931,N_3646,N_3503);
nand U7932 (N_7932,N_1018,N_857);
nand U7933 (N_7933,N_3964,N_145);
nor U7934 (N_7934,N_1398,N_2029);
or U7935 (N_7935,N_3254,N_2221);
nor U7936 (N_7936,N_2230,N_623);
xor U7937 (N_7937,N_1927,N_1545);
nor U7938 (N_7938,N_2713,N_3320);
nor U7939 (N_7939,N_2885,N_1180);
and U7940 (N_7940,N_1663,N_3002);
nor U7941 (N_7941,N_2443,N_2397);
nor U7942 (N_7942,N_79,N_1331);
nand U7943 (N_7943,N_917,N_2253);
or U7944 (N_7944,N_628,N_3300);
and U7945 (N_7945,N_2327,N_3025);
or U7946 (N_7946,N_2939,N_1066);
nor U7947 (N_7947,N_3447,N_2297);
nand U7948 (N_7948,N_3747,N_3406);
nand U7949 (N_7949,N_3811,N_1423);
or U7950 (N_7950,N_2394,N_2995);
or U7951 (N_7951,N_1284,N_3153);
xnor U7952 (N_7952,N_2654,N_3889);
xor U7953 (N_7953,N_325,N_137);
nor U7954 (N_7954,N_1927,N_2162);
xnor U7955 (N_7955,N_503,N_2602);
xnor U7956 (N_7956,N_2298,N_255);
nand U7957 (N_7957,N_3781,N_3646);
nor U7958 (N_7958,N_3764,N_2524);
nand U7959 (N_7959,N_1745,N_1661);
nand U7960 (N_7960,N_2355,N_1701);
xor U7961 (N_7961,N_3292,N_2386);
or U7962 (N_7962,N_620,N_1764);
or U7963 (N_7963,N_467,N_637);
or U7964 (N_7964,N_1507,N_2862);
nand U7965 (N_7965,N_1644,N_2164);
nor U7966 (N_7966,N_2877,N_1167);
xor U7967 (N_7967,N_762,N_3422);
nand U7968 (N_7968,N_2763,N_794);
and U7969 (N_7969,N_3828,N_2531);
nor U7970 (N_7970,N_1240,N_1260);
or U7971 (N_7971,N_1959,N_757);
and U7972 (N_7972,N_202,N_2210);
or U7973 (N_7973,N_2390,N_840);
or U7974 (N_7974,N_2078,N_427);
and U7975 (N_7975,N_2199,N_3987);
xnor U7976 (N_7976,N_750,N_2634);
nand U7977 (N_7977,N_497,N_2434);
and U7978 (N_7978,N_3924,N_195);
xnor U7979 (N_7979,N_2426,N_2175);
or U7980 (N_7980,N_164,N_616);
nand U7981 (N_7981,N_1495,N_711);
xor U7982 (N_7982,N_473,N_2965);
nand U7983 (N_7983,N_1966,N_1792);
nand U7984 (N_7984,N_2744,N_2976);
nand U7985 (N_7985,N_1512,N_1131);
nor U7986 (N_7986,N_1333,N_638);
nand U7987 (N_7987,N_1010,N_2304);
or U7988 (N_7988,N_1498,N_1557);
and U7989 (N_7989,N_1825,N_3963);
xnor U7990 (N_7990,N_1385,N_41);
or U7991 (N_7991,N_1576,N_704);
or U7992 (N_7992,N_1424,N_3181);
xor U7993 (N_7993,N_2406,N_3871);
xnor U7994 (N_7994,N_1507,N_1615);
and U7995 (N_7995,N_1195,N_2515);
xnor U7996 (N_7996,N_393,N_2248);
xor U7997 (N_7997,N_2513,N_1143);
nand U7998 (N_7998,N_3412,N_2675);
nor U7999 (N_7999,N_3522,N_1854);
nor U8000 (N_8000,N_6392,N_5285);
nand U8001 (N_8001,N_7742,N_7145);
and U8002 (N_8002,N_7795,N_7882);
nor U8003 (N_8003,N_7226,N_4744);
nor U8004 (N_8004,N_4466,N_5232);
or U8005 (N_8005,N_5694,N_6217);
nand U8006 (N_8006,N_6707,N_7392);
nand U8007 (N_8007,N_6274,N_6744);
xor U8008 (N_8008,N_6869,N_5888);
nor U8009 (N_8009,N_7983,N_7540);
or U8010 (N_8010,N_4695,N_7784);
xor U8011 (N_8011,N_7681,N_6405);
or U8012 (N_8012,N_7129,N_6410);
or U8013 (N_8013,N_5481,N_6350);
and U8014 (N_8014,N_5721,N_7611);
and U8015 (N_8015,N_4420,N_5150);
and U8016 (N_8016,N_6070,N_4947);
or U8017 (N_8017,N_5622,N_7080);
and U8018 (N_8018,N_4862,N_4883);
nor U8019 (N_8019,N_4277,N_4388);
and U8020 (N_8020,N_6716,N_5914);
xor U8021 (N_8021,N_5327,N_5455);
nand U8022 (N_8022,N_6829,N_5410);
nor U8023 (N_8023,N_6301,N_5325);
nor U8024 (N_8024,N_5819,N_7230);
nor U8025 (N_8025,N_5445,N_7068);
nor U8026 (N_8026,N_5913,N_5041);
and U8027 (N_8027,N_4007,N_4326);
xor U8028 (N_8028,N_5203,N_7724);
nor U8029 (N_8029,N_4507,N_4151);
and U8030 (N_8030,N_4405,N_7058);
xnor U8031 (N_8031,N_4456,N_6721);
and U8032 (N_8032,N_4557,N_6694);
nand U8033 (N_8033,N_4153,N_7934);
xnor U8034 (N_8034,N_4047,N_7994);
xnor U8035 (N_8035,N_6195,N_4867);
xor U8036 (N_8036,N_5512,N_6962);
xor U8037 (N_8037,N_6881,N_5769);
nand U8038 (N_8038,N_5322,N_6371);
nand U8039 (N_8039,N_6859,N_5526);
xor U8040 (N_8040,N_5818,N_4214);
nor U8041 (N_8041,N_7308,N_6280);
nor U8042 (N_8042,N_6895,N_6130);
and U8043 (N_8043,N_4685,N_5353);
xor U8044 (N_8044,N_7870,N_7001);
and U8045 (N_8045,N_7224,N_5693);
nor U8046 (N_8046,N_6315,N_4457);
xnor U8047 (N_8047,N_4417,N_7964);
xor U8048 (N_8048,N_5376,N_7662);
and U8049 (N_8049,N_5043,N_7028);
nand U8050 (N_8050,N_5534,N_5932);
xnor U8051 (N_8051,N_4999,N_6335);
nand U8052 (N_8052,N_6632,N_5130);
or U8053 (N_8053,N_6206,N_6409);
nand U8054 (N_8054,N_4910,N_7205);
and U8055 (N_8055,N_5848,N_4163);
nand U8056 (N_8056,N_5523,N_5112);
nor U8057 (N_8057,N_5921,N_4485);
and U8058 (N_8058,N_4442,N_7651);
xnor U8059 (N_8059,N_7461,N_6474);
xor U8060 (N_8060,N_7860,N_5415);
and U8061 (N_8061,N_4017,N_4849);
or U8062 (N_8062,N_4034,N_7701);
and U8063 (N_8063,N_5123,N_6913);
nor U8064 (N_8064,N_7568,N_5647);
or U8065 (N_8065,N_5042,N_7546);
and U8066 (N_8066,N_7844,N_6053);
nand U8067 (N_8067,N_6578,N_4187);
or U8068 (N_8068,N_5256,N_4546);
and U8069 (N_8069,N_4336,N_4671);
and U8070 (N_8070,N_4359,N_6509);
xor U8071 (N_8071,N_7897,N_7060);
nand U8072 (N_8072,N_5614,N_7351);
nor U8073 (N_8073,N_4223,N_6990);
xnor U8074 (N_8074,N_5072,N_5566);
nand U8075 (N_8075,N_5413,N_7930);
and U8076 (N_8076,N_6564,N_7604);
nand U8077 (N_8077,N_6450,N_6118);
nor U8078 (N_8078,N_6902,N_7457);
xor U8079 (N_8079,N_6162,N_5795);
or U8080 (N_8080,N_4379,N_4589);
nand U8081 (N_8081,N_7074,N_6739);
nor U8082 (N_8082,N_6670,N_4085);
nand U8083 (N_8083,N_4620,N_6952);
and U8084 (N_8084,N_4448,N_6624);
nor U8085 (N_8085,N_5463,N_7723);
xnor U8086 (N_8086,N_6240,N_6360);
nor U8087 (N_8087,N_6364,N_6877);
nand U8088 (N_8088,N_6215,N_6435);
nor U8089 (N_8089,N_5714,N_5129);
nor U8090 (N_8090,N_6305,N_7082);
or U8091 (N_8091,N_6170,N_6229);
xnor U8092 (N_8092,N_4776,N_5493);
and U8093 (N_8093,N_4675,N_5626);
nand U8094 (N_8094,N_5907,N_4263);
xnor U8095 (N_8095,N_6297,N_5996);
xor U8096 (N_8096,N_7372,N_6674);
xnor U8097 (N_8097,N_5246,N_5135);
and U8098 (N_8098,N_4161,N_6770);
nand U8099 (N_8099,N_5751,N_7585);
nor U8100 (N_8100,N_7209,N_6927);
nand U8101 (N_8101,N_7227,N_7523);
or U8102 (N_8102,N_5800,N_5599);
and U8103 (N_8103,N_4008,N_7279);
nor U8104 (N_8104,N_6664,N_5343);
nand U8105 (N_8105,N_7613,N_7026);
nand U8106 (N_8106,N_4341,N_4015);
nand U8107 (N_8107,N_6768,N_5158);
and U8108 (N_8108,N_5840,N_7039);
nand U8109 (N_8109,N_6306,N_4385);
xor U8110 (N_8110,N_4451,N_7966);
nor U8111 (N_8111,N_5804,N_7879);
nor U8112 (N_8112,N_7922,N_5420);
nand U8113 (N_8113,N_5136,N_7244);
nor U8114 (N_8114,N_7626,N_5990);
nor U8115 (N_8115,N_4073,N_4221);
and U8116 (N_8116,N_5930,N_6749);
nor U8117 (N_8117,N_4583,N_5483);
nor U8118 (N_8118,N_7381,N_6494);
or U8119 (N_8119,N_4256,N_5142);
xor U8120 (N_8120,N_4259,N_4291);
nor U8121 (N_8121,N_7789,N_6958);
nand U8122 (N_8122,N_5598,N_7458);
nand U8123 (N_8123,N_6846,N_4663);
nor U8124 (N_8124,N_7252,N_4817);
xnor U8125 (N_8125,N_6987,N_5014);
or U8126 (N_8126,N_4310,N_4745);
and U8127 (N_8127,N_5211,N_6889);
or U8128 (N_8128,N_7545,N_7929);
and U8129 (N_8129,N_6122,N_7002);
or U8130 (N_8130,N_7534,N_6196);
and U8131 (N_8131,N_7495,N_6650);
and U8132 (N_8132,N_4975,N_4390);
nor U8133 (N_8133,N_7576,N_5497);
and U8134 (N_8134,N_4136,N_6393);
nand U8135 (N_8135,N_4183,N_5374);
xnor U8136 (N_8136,N_7676,N_4660);
nand U8137 (N_8137,N_5633,N_6642);
nand U8138 (N_8138,N_6172,N_6055);
xor U8139 (N_8139,N_5583,N_5385);
nand U8140 (N_8140,N_7283,N_7671);
xor U8141 (N_8141,N_4827,N_5286);
or U8142 (N_8142,N_4866,N_6385);
nor U8143 (N_8143,N_7935,N_7642);
or U8144 (N_8144,N_5931,N_6948);
and U8145 (N_8145,N_5557,N_6953);
or U8146 (N_8146,N_6328,N_4595);
nor U8147 (N_8147,N_4552,N_7905);
or U8148 (N_8148,N_5834,N_5433);
xor U8149 (N_8149,N_7980,N_7618);
nand U8150 (N_8150,N_7407,N_4545);
and U8151 (N_8151,N_4189,N_5838);
or U8152 (N_8152,N_7510,N_4232);
nand U8153 (N_8153,N_6841,N_5744);
nor U8154 (N_8154,N_5520,N_7262);
or U8155 (N_8155,N_6856,N_6411);
xor U8156 (N_8156,N_6531,N_5912);
or U8157 (N_8157,N_5017,N_5046);
and U8158 (N_8158,N_5507,N_5160);
and U8159 (N_8159,N_4544,N_5216);
nand U8160 (N_8160,N_6997,N_4782);
nor U8161 (N_8161,N_6361,N_4218);
or U8162 (N_8162,N_6465,N_4712);
nor U8163 (N_8163,N_4932,N_4972);
nand U8164 (N_8164,N_7218,N_7007);
nor U8165 (N_8165,N_6271,N_5967);
or U8166 (N_8166,N_5812,N_4599);
or U8167 (N_8167,N_5715,N_6822);
nand U8168 (N_8168,N_7959,N_6980);
nor U8169 (N_8169,N_6054,N_6915);
xor U8170 (N_8170,N_6547,N_5839);
nor U8171 (N_8171,N_6384,N_4625);
or U8172 (N_8172,N_4453,N_6710);
nor U8173 (N_8173,N_7997,N_4224);
or U8174 (N_8174,N_6086,N_6837);
xor U8175 (N_8175,N_6662,N_7717);
or U8176 (N_8176,N_4643,N_4918);
nor U8177 (N_8177,N_7264,N_6097);
nand U8178 (N_8178,N_7232,N_5977);
or U8179 (N_8179,N_4115,N_5886);
nand U8180 (N_8180,N_6002,N_7360);
nor U8181 (N_8181,N_5828,N_5151);
xnor U8182 (N_8182,N_5952,N_7962);
or U8183 (N_8183,N_6608,N_6050);
and U8184 (N_8184,N_4195,N_5971);
nor U8185 (N_8185,N_5550,N_6138);
or U8186 (N_8186,N_5779,N_4391);
or U8187 (N_8187,N_4303,N_6545);
nor U8188 (N_8188,N_5960,N_7072);
xor U8189 (N_8189,N_6427,N_6181);
nor U8190 (N_8190,N_6897,N_6141);
and U8191 (N_8191,N_4260,N_7975);
nand U8192 (N_8192,N_4345,N_5891);
nor U8193 (N_8193,N_5350,N_5860);
nor U8194 (N_8194,N_6520,N_5456);
nor U8195 (N_8195,N_6223,N_7559);
nor U8196 (N_8196,N_5597,N_7536);
nand U8197 (N_8197,N_6894,N_7739);
or U8198 (N_8198,N_4812,N_6471);
nor U8199 (N_8199,N_5241,N_6777);
nor U8200 (N_8200,N_4815,N_6066);
or U8201 (N_8201,N_7819,N_7786);
nor U8202 (N_8202,N_4759,N_4309);
and U8203 (N_8203,N_6134,N_4750);
xor U8204 (N_8204,N_5214,N_6688);
nand U8205 (N_8205,N_7791,N_6470);
and U8206 (N_8206,N_6498,N_4031);
nand U8207 (N_8207,N_7910,N_7292);
and U8208 (N_8208,N_7869,N_6575);
or U8209 (N_8209,N_5149,N_4880);
and U8210 (N_8210,N_4297,N_4113);
or U8211 (N_8211,N_4254,N_7606);
nand U8212 (N_8212,N_7765,N_4963);
xor U8213 (N_8213,N_6145,N_5166);
nand U8214 (N_8214,N_4528,N_6728);
xnor U8215 (N_8215,N_6012,N_5352);
nor U8216 (N_8216,N_4874,N_7034);
and U8217 (N_8217,N_7160,N_7364);
nand U8218 (N_8218,N_7688,N_4348);
nand U8219 (N_8219,N_6541,N_4202);
nand U8220 (N_8220,N_6783,N_7537);
xor U8221 (N_8221,N_6221,N_4030);
or U8222 (N_8222,N_4710,N_6318);
nor U8223 (N_8223,N_6584,N_6210);
and U8224 (N_8224,N_7733,N_5293);
nor U8225 (N_8225,N_4861,N_6189);
or U8226 (N_8226,N_4598,N_7104);
and U8227 (N_8227,N_4495,N_6942);
nor U8228 (N_8228,N_5815,N_5096);
or U8229 (N_8229,N_4988,N_4316);
xor U8230 (N_8230,N_5242,N_7615);
xor U8231 (N_8231,N_5106,N_6528);
nand U8232 (N_8232,N_4046,N_4241);
nor U8233 (N_8233,N_5051,N_4220);
or U8234 (N_8234,N_5513,N_7646);
and U8235 (N_8235,N_5746,N_6748);
or U8236 (N_8236,N_5808,N_7259);
nor U8237 (N_8237,N_5857,N_5404);
xor U8238 (N_8238,N_6540,N_6590);
or U8239 (N_8239,N_6092,N_4013);
nor U8240 (N_8240,N_7636,N_6971);
xor U8241 (N_8241,N_5398,N_5425);
or U8242 (N_8242,N_6302,N_4839);
nor U8243 (N_8243,N_6794,N_4038);
nor U8244 (N_8244,N_4936,N_4833);
nor U8245 (N_8245,N_5044,N_4367);
or U8246 (N_8246,N_7533,N_6478);
xor U8247 (N_8247,N_5450,N_7976);
nand U8248 (N_8248,N_4967,N_5058);
or U8249 (N_8249,N_7459,N_5169);
xor U8250 (N_8250,N_4987,N_6787);
and U8251 (N_8251,N_7555,N_5331);
xnor U8252 (N_8252,N_5755,N_5025);
nor U8253 (N_8253,N_7201,N_5358);
nand U8254 (N_8254,N_6563,N_5603);
nand U8255 (N_8255,N_7347,N_5368);
or U8256 (N_8256,N_4826,N_6154);
xnor U8257 (N_8257,N_6451,N_4009);
nor U8258 (N_8258,N_5225,N_6931);
xnor U8259 (N_8259,N_4253,N_7309);
and U8260 (N_8260,N_6703,N_5898);
or U8261 (N_8261,N_7297,N_5627);
or U8262 (N_8262,N_6253,N_4686);
or U8263 (N_8263,N_7320,N_5743);
and U8264 (N_8264,N_7311,N_5654);
nand U8265 (N_8265,N_6544,N_4677);
or U8266 (N_8266,N_7776,N_7951);
nand U8267 (N_8267,N_4271,N_6191);
and U8268 (N_8268,N_4144,N_7720);
nor U8269 (N_8269,N_7690,N_7054);
nor U8270 (N_8270,N_4330,N_4642);
and U8271 (N_8271,N_6916,N_7845);
or U8272 (N_8272,N_6960,N_6135);
and U8273 (N_8273,N_6178,N_4067);
xor U8274 (N_8274,N_6352,N_5069);
and U8275 (N_8275,N_5612,N_4604);
or U8276 (N_8276,N_6665,N_5710);
nand U8277 (N_8277,N_5408,N_5605);
or U8278 (N_8278,N_4701,N_4210);
nor U8279 (N_8279,N_5437,N_6585);
and U8280 (N_8280,N_7734,N_5669);
or U8281 (N_8281,N_4480,N_4505);
xnor U8282 (N_8282,N_4851,N_7186);
nor U8283 (N_8283,N_4740,N_7582);
or U8284 (N_8284,N_7766,N_7917);
nor U8285 (N_8285,N_6651,N_5370);
and U8286 (N_8286,N_6260,N_6398);
xor U8287 (N_8287,N_4538,N_6408);
nand U8288 (N_8288,N_4753,N_4061);
nand U8289 (N_8289,N_7422,N_6853);
nand U8290 (N_8290,N_5298,N_6279);
nor U8291 (N_8291,N_7649,N_7140);
nand U8292 (N_8292,N_4597,N_7208);
nor U8293 (N_8293,N_7063,N_5167);
xnor U8294 (N_8294,N_6255,N_7041);
or U8295 (N_8295,N_7363,N_4895);
or U8296 (N_8296,N_5318,N_4237);
nand U8297 (N_8297,N_7743,N_6803);
nand U8298 (N_8298,N_7065,N_5538);
and U8299 (N_8299,N_4727,N_7949);
and U8300 (N_8300,N_7328,N_6944);
nor U8301 (N_8301,N_6394,N_5110);
xor U8302 (N_8302,N_4818,N_7403);
nand U8303 (N_8303,N_6173,N_4471);
nor U8304 (N_8304,N_4952,N_4509);
xnor U8305 (N_8305,N_7889,N_5998);
nand U8306 (N_8306,N_7829,N_7989);
and U8307 (N_8307,N_6734,N_7076);
or U8308 (N_8308,N_7163,N_6995);
nand U8309 (N_8309,N_7094,N_5790);
or U8310 (N_8310,N_7515,N_4418);
nor U8311 (N_8311,N_6970,N_6036);
nand U8312 (N_8312,N_6359,N_6505);
and U8313 (N_8313,N_6761,N_7056);
nor U8314 (N_8314,N_5011,N_5901);
nand U8315 (N_8315,N_5897,N_5319);
xor U8316 (N_8316,N_4708,N_7553);
or U8317 (N_8317,N_5419,N_7658);
nor U8318 (N_8318,N_5143,N_7118);
nor U8319 (N_8319,N_5787,N_7497);
nand U8320 (N_8320,N_6824,N_6929);
or U8321 (N_8321,N_6375,N_4059);
and U8322 (N_8322,N_7037,N_6506);
nor U8323 (N_8323,N_4487,N_4315);
nand U8324 (N_8324,N_7116,N_5723);
or U8325 (N_8325,N_5561,N_6515);
nand U8326 (N_8326,N_6430,N_6542);
and U8327 (N_8327,N_4321,N_7888);
nand U8328 (N_8328,N_4234,N_4056);
nand U8329 (N_8329,N_5268,N_5986);
nand U8330 (N_8330,N_7302,N_7047);
and U8331 (N_8331,N_4130,N_5024);
or U8332 (N_8332,N_5832,N_6233);
and U8333 (N_8333,N_6552,N_7965);
nor U8334 (N_8334,N_7411,N_6179);
xor U8335 (N_8335,N_4943,N_7077);
nand U8336 (N_8336,N_6556,N_7918);
nor U8337 (N_8337,N_4173,N_6250);
or U8338 (N_8338,N_7324,N_7286);
or U8339 (N_8339,N_7854,N_6197);
nand U8340 (N_8340,N_4617,N_6421);
nor U8341 (N_8341,N_4105,N_7023);
and U8342 (N_8342,N_6898,N_7024);
nand U8343 (N_8343,N_7603,N_7915);
and U8344 (N_8344,N_6914,N_5308);
nand U8345 (N_8345,N_5274,N_5400);
nand U8346 (N_8346,N_7414,N_6938);
or U8347 (N_8347,N_5027,N_4728);
nand U8348 (N_8348,N_4063,N_6730);
xnor U8349 (N_8349,N_4333,N_6756);
xor U8350 (N_8350,N_5066,N_7435);
nand U8351 (N_8351,N_5393,N_5399);
and U8352 (N_8352,N_5426,N_6699);
nand U8353 (N_8353,N_4039,N_6521);
xor U8354 (N_8354,N_7017,N_5661);
xor U8355 (N_8355,N_5681,N_5152);
nor U8356 (N_8356,N_7728,N_6562);
and U8357 (N_8357,N_4486,N_6164);
xnor U8358 (N_8358,N_6968,N_6599);
xnor U8359 (N_8359,N_4872,N_5965);
or U8360 (N_8360,N_6947,N_4689);
or U8361 (N_8361,N_6268,N_6878);
nor U8362 (N_8362,N_6833,N_4317);
or U8363 (N_8363,N_5510,N_6047);
or U8364 (N_8364,N_7702,N_7144);
and U8365 (N_8365,N_5099,N_7345);
nor U8366 (N_8366,N_7756,N_5012);
or U8367 (N_8367,N_4116,N_7652);
nor U8368 (N_8368,N_7294,N_4351);
xor U8369 (N_8369,N_4885,N_6236);
nor U8370 (N_8370,N_4768,N_4879);
and U8371 (N_8371,N_6549,N_6330);
and U8372 (N_8372,N_5397,N_4416);
or U8373 (N_8373,N_6461,N_6501);
xnor U8374 (N_8374,N_7210,N_6941);
and U8375 (N_8375,N_6114,N_4494);
or U8376 (N_8376,N_5192,N_6368);
or U8377 (N_8377,N_6156,N_5488);
or U8378 (N_8378,N_7855,N_6489);
nor U8379 (N_8379,N_6637,N_5013);
or U8380 (N_8380,N_6087,N_4730);
nor U8381 (N_8381,N_6950,N_7638);
nor U8382 (N_8382,N_6443,N_4117);
and U8383 (N_8383,N_7272,N_5973);
nand U8384 (N_8384,N_5444,N_6370);
xnor U8385 (N_8385,N_6083,N_5585);
or U8386 (N_8386,N_6993,N_5029);
or U8387 (N_8387,N_5810,N_7185);
or U8388 (N_8388,N_6152,N_4631);
and U8389 (N_8389,N_4296,N_4697);
or U8390 (N_8390,N_7837,N_5309);
nand U8391 (N_8391,N_6862,N_4215);
nor U8392 (N_8392,N_4962,N_5462);
nor U8393 (N_8393,N_5854,N_5927);
and U8394 (N_8394,N_6992,N_7267);
nand U8395 (N_8395,N_5191,N_5757);
or U8396 (N_8396,N_7327,N_7647);
and U8397 (N_8397,N_7761,N_6157);
and U8398 (N_8398,N_5473,N_6316);
or U8399 (N_8399,N_5826,N_4429);
or U8400 (N_8400,N_6022,N_5972);
or U8401 (N_8401,N_7274,N_5544);
xor U8402 (N_8402,N_4762,N_4363);
xnor U8403 (N_8403,N_5539,N_4981);
and U8404 (N_8404,N_5364,N_4755);
or U8405 (N_8405,N_5489,N_4089);
xnor U8406 (N_8406,N_6533,N_4227);
xnor U8407 (N_8407,N_4562,N_7931);
or U8408 (N_8408,N_7052,N_7531);
nand U8409 (N_8409,N_5611,N_6779);
xor U8410 (N_8410,N_4908,N_7212);
xor U8411 (N_8411,N_5163,N_7035);
nor U8412 (N_8412,N_6733,N_6843);
nor U8413 (N_8413,N_6858,N_6726);
or U8414 (N_8414,N_5357,N_5803);
xnor U8415 (N_8415,N_7549,N_7612);
nor U8416 (N_8416,N_7339,N_6702);
and U8417 (N_8417,N_6340,N_7059);
and U8418 (N_8418,N_7444,N_4257);
xnor U8419 (N_8419,N_4667,N_4725);
nor U8420 (N_8420,N_7207,N_6872);
or U8421 (N_8421,N_7132,N_7925);
nand U8422 (N_8422,N_6034,N_6887);
and U8423 (N_8423,N_7044,N_6742);
nor U8424 (N_8424,N_7386,N_5508);
nand U8425 (N_8425,N_4714,N_7872);
or U8426 (N_8426,N_4892,N_5920);
nand U8427 (N_8427,N_7772,N_7767);
and U8428 (N_8428,N_7600,N_7721);
nor U8429 (N_8429,N_5414,N_6848);
nor U8430 (N_8430,N_4389,N_6077);
xor U8431 (N_8431,N_4177,N_4349);
nand U8432 (N_8432,N_7919,N_4829);
and U8433 (N_8433,N_5401,N_5616);
and U8434 (N_8434,N_5438,N_5396);
nand U8435 (N_8435,N_4150,N_4452);
nand U8436 (N_8436,N_6620,N_6116);
and U8437 (N_8437,N_7004,N_6587);
and U8438 (N_8438,N_6560,N_4353);
and U8439 (N_8439,N_4270,N_6198);
nor U8440 (N_8440,N_6979,N_6937);
or U8441 (N_8441,N_4447,N_7792);
nand U8442 (N_8442,N_4662,N_4930);
or U8443 (N_8443,N_5524,N_5650);
xnor U8444 (N_8444,N_4843,N_4699);
xnor U8445 (N_8445,N_5644,N_4498);
xnor U8446 (N_8446,N_5591,N_4275);
nand U8447 (N_8447,N_5454,N_7171);
nand U8448 (N_8448,N_4915,N_6220);
and U8449 (N_8449,N_5732,N_6883);
xor U8450 (N_8450,N_6446,N_5138);
or U8451 (N_8451,N_4760,N_4541);
or U8452 (N_8452,N_6448,N_7348);
nor U8453 (N_8453,N_6566,N_4683);
nor U8454 (N_8454,N_5219,N_5159);
and U8455 (N_8455,N_7383,N_5125);
nor U8456 (N_8456,N_5625,N_4409);
and U8457 (N_8457,N_4053,N_5252);
nor U8458 (N_8458,N_7202,N_4992);
or U8459 (N_8459,N_5864,N_6462);
nand U8460 (N_8460,N_5894,N_6457);
and U8461 (N_8461,N_6071,N_4157);
nor U8462 (N_8462,N_5359,N_5317);
xnor U8463 (N_8463,N_4884,N_5228);
or U8464 (N_8464,N_6765,N_5060);
or U8465 (N_8465,N_7331,N_6123);
or U8466 (N_8466,N_6378,N_6985);
nor U8467 (N_8467,N_6806,N_5296);
xor U8468 (N_8468,N_6672,N_5080);
and U8469 (N_8469,N_5976,N_7928);
nor U8470 (N_8470,N_6759,N_7590);
xnor U8471 (N_8471,N_7395,N_5435);
xnor U8472 (N_8472,N_6709,N_4294);
nor U8473 (N_8473,N_7012,N_7165);
or U8474 (N_8474,N_7187,N_7969);
xnor U8475 (N_8475,N_5141,N_7599);
xnor U8476 (N_8476,N_6731,N_4968);
nor U8477 (N_8477,N_4567,N_6956);
xor U8478 (N_8478,N_6906,N_7445);
nand U8479 (N_8479,N_5602,N_4900);
nand U8480 (N_8480,N_4190,N_5194);
nor U8481 (N_8481,N_5861,N_6800);
nor U8482 (N_8482,N_5082,N_6463);
nand U8483 (N_8483,N_7946,N_4463);
or U8484 (N_8484,N_4547,N_7305);
nor U8485 (N_8485,N_5428,N_5153);
or U8486 (N_8486,N_5243,N_7030);
or U8487 (N_8487,N_4649,N_7390);
and U8488 (N_8488,N_4431,N_7388);
xnor U8489 (N_8489,N_7261,N_5295);
or U8490 (N_8490,N_5227,N_5073);
and U8491 (N_8491,N_5934,N_4517);
or U8492 (N_8492,N_7130,N_5432);
nor U8493 (N_8493,N_6028,N_7763);
nand U8494 (N_8494,N_4690,N_5290);
xnor U8495 (N_8495,N_6079,N_7238);
nor U8496 (N_8496,N_6063,N_7508);
and U8497 (N_8497,N_5939,N_7117);
nand U8498 (N_8498,N_7033,N_4375);
or U8499 (N_8499,N_5372,N_4112);
nor U8500 (N_8500,N_7374,N_6322);
or U8501 (N_8501,N_6013,N_7581);
or U8502 (N_8502,N_7911,N_7744);
and U8503 (N_8503,N_6850,N_6251);
nand U8504 (N_8504,N_4392,N_4844);
nor U8505 (N_8505,N_5495,N_4939);
nor U8506 (N_8506,N_4558,N_7441);
nor U8507 (N_8507,N_4596,N_4219);
xor U8508 (N_8508,N_6679,N_4796);
nand U8509 (N_8509,N_7750,N_6372);
xor U8510 (N_8510,N_7852,N_6265);
xnor U8511 (N_8511,N_5980,N_5664);
xnor U8512 (N_8512,N_4106,N_6143);
nand U8513 (N_8513,N_7438,N_6230);
nor U8514 (N_8514,N_5412,N_7423);
and U8515 (N_8515,N_5068,N_5119);
and U8516 (N_8516,N_7621,N_4140);
nand U8517 (N_8517,N_4726,N_5686);
and U8518 (N_8518,N_4858,N_6561);
xor U8519 (N_8519,N_7886,N_5629);
or U8520 (N_8520,N_6523,N_6346);
or U8521 (N_8521,N_7830,N_7016);
or U8522 (N_8522,N_6060,N_7511);
nor U8523 (N_8523,N_5558,N_7282);
xor U8524 (N_8524,N_6604,N_4472);
nand U8525 (N_8525,N_4041,N_7704);
and U8526 (N_8526,N_4518,N_4731);
xnor U8527 (N_8527,N_4170,N_6376);
xor U8528 (N_8528,N_6413,N_4191);
xnor U8529 (N_8529,N_5684,N_6631);
or U8530 (N_8530,N_5735,N_5504);
or U8531 (N_8531,N_7166,N_6782);
nand U8532 (N_8532,N_7195,N_4422);
nor U8533 (N_8533,N_4548,N_7115);
xor U8534 (N_8534,N_5292,N_7110);
and U8535 (N_8535,N_6606,N_7516);
nand U8536 (N_8536,N_7982,N_4470);
xor U8537 (N_8537,N_6321,N_6124);
xor U8538 (N_8538,N_4327,N_6508);
nand U8539 (N_8539,N_7101,N_4523);
xor U8540 (N_8540,N_6081,N_6751);
and U8541 (N_8541,N_5574,N_6444);
nand U8542 (N_8542,N_4593,N_7719);
nor U8543 (N_8543,N_4192,N_4290);
xor U8544 (N_8544,N_4790,N_5948);
or U8545 (N_8545,N_6586,N_4159);
or U8546 (N_8546,N_7156,N_5822);
nand U8547 (N_8547,N_7474,N_4743);
xor U8548 (N_8548,N_4983,N_5718);
nand U8549 (N_8549,N_7256,N_4164);
nor U8550 (N_8550,N_6011,N_4870);
nand U8551 (N_8551,N_4933,N_5004);
nor U8552 (N_8552,N_7973,N_4678);
nand U8553 (N_8553,N_7812,N_4914);
nand U8554 (N_8554,N_4581,N_6420);
xnor U8555 (N_8555,N_5395,N_5403);
nand U8556 (N_8556,N_7410,N_5618);
and U8557 (N_8557,N_7316,N_4147);
nand U8558 (N_8558,N_7578,N_6426);
and U8559 (N_8559,N_6177,N_4670);
nor U8560 (N_8560,N_4054,N_6167);
nand U8561 (N_8561,N_5257,N_7278);
nor U8562 (N_8562,N_6468,N_5651);
xor U8563 (N_8563,N_4657,N_7203);
nand U8564 (N_8564,N_5390,N_4739);
and U8565 (N_8565,N_4941,N_4926);
and U8566 (N_8566,N_6555,N_7257);
or U8567 (N_8567,N_4284,N_5230);
or U8568 (N_8568,N_6294,N_6094);
xnor U8569 (N_8569,N_4763,N_7112);
nand U8570 (N_8570,N_4644,N_5262);
or U8571 (N_8571,N_5245,N_4093);
or U8572 (N_8572,N_5758,N_4821);
and U8573 (N_8573,N_6262,N_4916);
nand U8574 (N_8574,N_6597,N_7005);
xnor U8575 (N_8575,N_7818,N_5753);
or U8576 (N_8576,N_5868,N_6784);
nor U8577 (N_8577,N_6010,N_7820);
and U8578 (N_8578,N_5300,N_4446);
xor U8579 (N_8579,N_4415,N_4881);
nand U8580 (N_8580,N_4226,N_6187);
and U8581 (N_8581,N_4907,N_5607);
nand U8582 (N_8582,N_4773,N_7231);
and U8583 (N_8583,N_6401,N_6016);
nand U8584 (N_8584,N_5287,N_4104);
nand U8585 (N_8585,N_6259,N_7142);
nor U8586 (N_8586,N_7943,N_4656);
nor U8587 (N_8587,N_6299,N_4860);
xnor U8588 (N_8588,N_7544,N_7293);
nand U8589 (N_8589,N_4088,N_4361);
nand U8590 (N_8590,N_5460,N_5975);
xor U8591 (N_8591,N_5666,N_7680);
xor U8592 (N_8592,N_4986,N_4311);
nand U8593 (N_8593,N_7214,N_4023);
nor U8594 (N_8594,N_4467,N_7769);
nand U8595 (N_8595,N_7485,N_7689);
and U8596 (N_8596,N_6105,N_7679);
and U8597 (N_8597,N_4329,N_4396);
and U8598 (N_8598,N_7628,N_4792);
nor U8599 (N_8599,N_4090,N_7788);
or U8600 (N_8600,N_7416,N_7757);
and U8601 (N_8601,N_6754,N_6292);
nor U8602 (N_8602,N_5794,N_4929);
nor U8603 (N_8603,N_6589,N_7427);
or U8604 (N_8604,N_4654,N_4394);
nand U8605 (N_8605,N_5623,N_4539);
nand U8606 (N_8606,N_7159,N_4959);
nor U8607 (N_8607,N_5008,N_7365);
and U8608 (N_8608,N_7296,N_6400);
and U8609 (N_8609,N_6963,N_7950);
nor U8610 (N_8610,N_5175,N_4334);
nor U8611 (N_8611,N_5009,N_6311);
or U8612 (N_8612,N_4898,N_5813);
or U8613 (N_8613,N_5678,N_7310);
xor U8614 (N_8614,N_4636,N_4079);
and U8615 (N_8615,N_5471,N_5122);
nand U8616 (N_8616,N_7169,N_5883);
nand U8617 (N_8617,N_6295,N_6065);
or U8618 (N_8618,N_7220,N_7770);
or U8619 (N_8619,N_7807,N_7102);
and U8620 (N_8620,N_5271,N_7298);
xnor U8621 (N_8621,N_6565,N_4927);
and U8622 (N_8622,N_7967,N_6868);
or U8623 (N_8623,N_4107,N_5134);
or U8624 (N_8624,N_5620,N_5464);
nand U8625 (N_8625,N_6329,N_7932);
nand U8626 (N_8626,N_7710,N_7478);
nor U8627 (N_8627,N_4246,N_6453);
nor U8628 (N_8628,N_6341,N_7079);
or U8629 (N_8629,N_7329,N_6404);
xnor U8630 (N_8630,N_4158,N_4798);
or U8631 (N_8631,N_5494,N_7686);
or U8632 (N_8632,N_5181,N_4629);
nor U8633 (N_8633,N_6252,N_4419);
or U8634 (N_8634,N_5760,N_5797);
nor U8635 (N_8635,N_5849,N_4850);
nor U8636 (N_8636,N_5502,N_7822);
nor U8637 (N_8637,N_6827,N_5880);
or U8638 (N_8638,N_7269,N_5811);
nor U8639 (N_8639,N_6419,N_4033);
nand U8640 (N_8640,N_4923,N_7677);
and U8641 (N_8641,N_7509,N_5021);
and U8642 (N_8642,N_4767,N_5668);
and U8643 (N_8643,N_6660,N_5448);
and U8644 (N_8644,N_4269,N_6282);
nor U8645 (N_8645,N_5193,N_7085);
nand U8646 (N_8646,N_5239,N_6414);
and U8647 (N_8647,N_5467,N_5470);
and U8648 (N_8648,N_6551,N_6729);
and U8649 (N_8649,N_4510,N_5083);
and U8650 (N_8650,N_5270,N_6237);
or U8651 (N_8651,N_4771,N_5431);
xnor U8652 (N_8652,N_5312,N_4478);
nand U8653 (N_8653,N_7313,N_7753);
xnor U8654 (N_8654,N_7906,N_4945);
or U8655 (N_8655,N_4188,N_4909);
and U8656 (N_8656,N_7810,N_5517);
nand U8657 (N_8657,N_6991,N_4004);
nand U8658 (N_8658,N_4868,N_5115);
nand U8659 (N_8659,N_5005,N_5018);
nand U8660 (N_8660,N_6256,N_5204);
or U8661 (N_8661,N_5983,N_5212);
or U8662 (N_8662,N_4171,N_6056);
or U8663 (N_8663,N_7098,N_7589);
or U8664 (N_8664,N_5984,N_5146);
nand U8665 (N_8665,N_4942,N_5541);
and U8666 (N_8666,N_4977,N_6625);
nor U8667 (N_8667,N_7440,N_5601);
or U8668 (N_8668,N_4835,N_7685);
or U8669 (N_8669,N_6725,N_4891);
nor U8670 (N_8670,N_6591,N_7245);
nand U8671 (N_8671,N_5105,N_5356);
nand U8672 (N_8672,N_4302,N_4577);
or U8673 (N_8673,N_7119,N_5542);
or U8674 (N_8674,N_6440,N_5802);
or U8675 (N_8675,N_4092,N_5205);
or U8676 (N_8676,N_4582,N_6727);
nand U8677 (N_8677,N_5545,N_6799);
and U8678 (N_8678,N_5348,N_4200);
xnor U8679 (N_8679,N_4435,N_4274);
nand U8680 (N_8680,N_6546,N_4772);
and U8681 (N_8681,N_5982,N_7718);
or U8682 (N_8682,N_5850,N_7491);
nand U8683 (N_8683,N_4247,N_4810);
nand U8684 (N_8684,N_5363,N_6524);
xor U8685 (N_8685,N_4550,N_4848);
and U8686 (N_8686,N_5916,N_6192);
or U8687 (N_8687,N_6692,N_5764);
nor U8688 (N_8688,N_7371,N_6873);
xor U8689 (N_8689,N_4646,N_6242);
or U8690 (N_8690,N_6107,N_4414);
nand U8691 (N_8691,N_6245,N_7237);
and U8692 (N_8692,N_7808,N_6317);
nor U8693 (N_8693,N_4903,N_7806);
and U8694 (N_8694,N_4990,N_6844);
and U8695 (N_8695,N_4255,N_6075);
nor U8696 (N_8696,N_6228,N_4281);
or U8697 (N_8697,N_5747,N_7216);
or U8698 (N_8698,N_7081,N_4166);
xor U8699 (N_8699,N_6793,N_7359);
or U8700 (N_8700,N_6304,N_7805);
xnor U8701 (N_8701,N_4035,N_5168);
or U8702 (N_8702,N_4012,N_7471);
xnor U8703 (N_8703,N_6772,N_7399);
nand U8704 (N_8704,N_4273,N_4238);
xor U8705 (N_8705,N_4250,N_5563);
or U8706 (N_8706,N_5055,N_7018);
and U8707 (N_8707,N_7481,N_4949);
xor U8708 (N_8708,N_6701,N_7151);
xor U8709 (N_8709,N_4563,N_4515);
nand U8710 (N_8710,N_7527,N_7154);
and U8711 (N_8711,N_7687,N_6876);
nor U8712 (N_8712,N_6062,N_7464);
nand U8713 (N_8713,N_7550,N_5624);
nor U8714 (N_8714,N_7779,N_7051);
nand U8715 (N_8715,N_6592,N_5900);
and U8716 (N_8716,N_7401,N_6396);
or U8717 (N_8717,N_4609,N_6852);
nand U8718 (N_8718,N_7513,N_6343);
and U8719 (N_8719,N_6169,N_6325);
xnor U8720 (N_8720,N_7177,N_6798);
xnor U8721 (N_8721,N_5266,N_5736);
and U8722 (N_8722,N_4029,N_5575);
and U8723 (N_8723,N_4010,N_7446);
and U8724 (N_8724,N_6175,N_4174);
xnor U8725 (N_8725,N_4114,N_4803);
or U8726 (N_8726,N_6403,N_6569);
or U8727 (N_8727,N_4213,N_7042);
xnor U8728 (N_8728,N_7378,N_5969);
nor U8729 (N_8729,N_4454,N_6110);
xnor U8730 (N_8730,N_5780,N_4655);
nor U8731 (N_8731,N_5991,N_4354);
nand U8732 (N_8732,N_7814,N_4921);
and U8733 (N_8733,N_7693,N_6042);
xnor U8734 (N_8734,N_4608,N_7565);
and U8735 (N_8735,N_5899,N_5867);
nand U8736 (N_8736,N_7632,N_5717);
nand U8737 (N_8737,N_7057,N_6769);
xnor U8738 (N_8738,N_6273,N_6479);
and U8739 (N_8739,N_7853,N_7175);
or U8740 (N_8740,N_7299,N_6773);
and U8741 (N_8741,N_4110,N_5917);
nor U8742 (N_8742,N_6511,N_5535);
or U8743 (N_8743,N_4672,N_6326);
xnor U8744 (N_8744,N_6723,N_7774);
or U8745 (N_8745,N_7700,N_6548);
nand U8746 (N_8746,N_5062,N_5720);
or U8747 (N_8747,N_4591,N_5781);
and U8748 (N_8748,N_4371,N_5938);
and U8749 (N_8749,N_6493,N_6239);
and U8750 (N_8750,N_4288,N_7190);
nand U8751 (N_8751,N_4324,N_6363);
nor U8752 (N_8752,N_5699,N_6814);
nand U8753 (N_8753,N_6627,N_7344);
xor U8754 (N_8754,N_6024,N_4475);
or U8755 (N_8755,N_5337,N_7794);
or U8756 (N_8756,N_4997,N_7981);
xnor U8757 (N_8757,N_6437,N_5476);
nor U8758 (N_8758,N_6354,N_7655);
nand U8759 (N_8759,N_6819,N_4493);
or U8760 (N_8760,N_4160,N_4713);
nand U8761 (N_8761,N_5562,N_4133);
nor U8762 (N_8762,N_7804,N_7315);
xor U8763 (N_8763,N_7366,N_7176);
nand U8764 (N_8764,N_6476,N_4906);
xor U8765 (N_8765,N_7143,N_6365);
or U8766 (N_8766,N_4308,N_5911);
and U8767 (N_8767,N_4834,N_7715);
nand U8768 (N_8768,N_4101,N_7157);
nor U8769 (N_8769,N_6955,N_7188);
nor U8770 (N_8770,N_6685,N_6510);
or U8771 (N_8771,N_6621,N_6965);
and U8772 (N_8772,N_5798,N_7877);
nand U8773 (N_8773,N_5533,N_7048);
xor U8774 (N_8774,N_4492,N_6460);
nor U8775 (N_8775,N_7862,N_5328);
nor U8776 (N_8776,N_6901,N_7100);
nor U8777 (N_8777,N_7561,N_6909);
and U8778 (N_8778,N_6048,N_7797);
nor U8779 (N_8779,N_4764,N_6922);
nand U8780 (N_8780,N_6683,N_7488);
nand U8781 (N_8781,N_4228,N_5330);
or U8782 (N_8782,N_6717,N_4384);
xor U8783 (N_8783,N_5284,N_5427);
xnor U8784 (N_8784,N_7924,N_6085);
or U8785 (N_8785,N_7583,N_6456);
nor U8786 (N_8786,N_5908,N_6349);
and U8787 (N_8787,N_6386,N_7903);
nand U8788 (N_8788,N_4781,N_5360);
nand U8789 (N_8789,N_4869,N_5974);
nand U8790 (N_8790,N_4863,N_4520);
nor U8791 (N_8791,N_6888,N_6091);
nand U8792 (N_8792,N_5407,N_4468);
or U8793 (N_8793,N_4299,N_5084);
or U8794 (N_8794,N_7179,N_6165);
or U8795 (N_8795,N_6522,N_4532);
or U8796 (N_8796,N_5422,N_4634);
or U8797 (N_8797,N_6964,N_4169);
and U8798 (N_8798,N_6429,N_7174);
and U8799 (N_8799,N_5941,N_7415);
nand U8800 (N_8800,N_6281,N_5411);
and U8801 (N_8801,N_5551,N_6289);
nor U8802 (N_8802,N_5708,N_4614);
xnor U8803 (N_8803,N_7249,N_4749);
xor U8804 (N_8804,N_5173,N_6415);
and U8805 (N_8805,N_4855,N_6319);
and U8806 (N_8806,N_4024,N_7300);
xor U8807 (N_8807,N_5511,N_5178);
xnor U8808 (N_8808,N_7321,N_5197);
xor U8809 (N_8809,N_4616,N_7832);
and U8810 (N_8810,N_7480,N_7518);
and U8811 (N_8811,N_7172,N_4312);
or U8812 (N_8812,N_5316,N_4131);
xor U8813 (N_8813,N_4580,N_7741);
nor U8814 (N_8814,N_4074,N_4286);
and U8815 (N_8815,N_4124,N_4142);
or U8816 (N_8816,N_4248,N_7920);
nand U8817 (N_8817,N_4207,N_4268);
xor U8818 (N_8818,N_6994,N_5436);
or U8819 (N_8819,N_4488,N_7921);
xor U8820 (N_8820,N_7287,N_7684);
or U8821 (N_8821,N_5600,N_4961);
or U8822 (N_8822,N_5392,N_4216);
and U8823 (N_8823,N_4331,N_4167);
xor U8824 (N_8824,N_5750,N_4201);
xor U8825 (N_8825,N_5277,N_5208);
or U8826 (N_8826,N_5334,N_4194);
or U8827 (N_8827,N_5637,N_7735);
xnor U8828 (N_8828,N_4335,N_7221);
or U8829 (N_8829,N_5248,N_5712);
and U8830 (N_8830,N_7437,N_6331);
nand U8831 (N_8831,N_7375,N_4553);
xor U8832 (N_8832,N_4536,N_6379);
nand U8833 (N_8833,N_7998,N_6051);
xnor U8834 (N_8834,N_5690,N_6747);
or U8835 (N_8835,N_5077,N_5947);
nor U8836 (N_8836,N_5993,N_5553);
xor U8837 (N_8837,N_5418,N_7066);
nand U8838 (N_8838,N_5145,N_4619);
or U8839 (N_8839,N_6514,N_4397);
and U8840 (N_8840,N_4836,N_4045);
xor U8841 (N_8841,N_4406,N_5902);
xnor U8842 (N_8842,N_7890,N_5451);
nand U8843 (N_8843,N_5092,N_6700);
nand U8844 (N_8844,N_7198,N_4272);
and U8845 (N_8845,N_6387,N_4469);
nand U8846 (N_8846,N_4381,N_5179);
xnor U8847 (N_8847,N_6810,N_5032);
nor U8848 (N_8848,N_6972,N_7859);
or U8849 (N_8849,N_6188,N_5843);
and U8850 (N_8850,N_5301,N_6283);
nand U8851 (N_8851,N_4083,N_6389);
nor U8852 (N_8852,N_7643,N_5997);
xor U8853 (N_8853,N_5676,N_6383);
xnor U8854 (N_8854,N_7592,N_5490);
nand U8855 (N_8855,N_6472,N_6581);
nor U8856 (N_8856,N_4449,N_7014);
nand U8857 (N_8857,N_6272,N_4724);
xor U8858 (N_8858,N_7986,N_7420);
xnor U8859 (N_8859,N_6432,N_6825);
nand U8860 (N_8860,N_7650,N_5341);
nand U8861 (N_8861,N_5177,N_4332);
xor U8862 (N_8862,N_5478,N_7974);
or U8863 (N_8863,N_6224,N_4888);
or U8864 (N_8864,N_5310,N_4057);
and U8865 (N_8865,N_4779,N_4148);
xnor U8866 (N_8866,N_6832,N_4587);
nor U8867 (N_8867,N_4086,N_4902);
xor U8868 (N_8868,N_4896,N_7640);
xnor U8869 (N_8869,N_7255,N_7598);
nor U8870 (N_8870,N_4700,N_6438);
or U8871 (N_8871,N_5999,N_7706);
and U8872 (N_8872,N_5354,N_7340);
nand U8873 (N_8873,N_5954,N_7878);
xor U8874 (N_8874,N_5617,N_4503);
nor U8875 (N_8875,N_7290,N_7284);
xnor U8876 (N_8876,N_6978,N_6797);
or U8877 (N_8877,N_4793,N_4969);
and U8878 (N_8878,N_7670,N_4820);
xnor U8879 (N_8879,N_7722,N_5332);
and U8880 (N_8880,N_6977,N_6628);
or U8881 (N_8881,N_6666,N_6805);
and U8882 (N_8882,N_7985,N_4521);
nand U8883 (N_8883,N_6069,N_6764);
xnor U8884 (N_8884,N_7954,N_6018);
or U8885 (N_8885,N_7405,N_7124);
xnor U8886 (N_8886,N_7428,N_7839);
and U8887 (N_8887,N_7197,N_4919);
or U8888 (N_8888,N_5133,N_6932);
nand U8889 (N_8889,N_4298,N_5567);
and U8890 (N_8890,N_4890,N_6133);
nand U8891 (N_8891,N_6477,N_6826);
xor U8892 (N_8892,N_7825,N_4682);
or U8893 (N_8893,N_6269,N_6243);
nand U8894 (N_8894,N_4205,N_4687);
and U8895 (N_8895,N_5923,N_5531);
nor U8896 (N_8896,N_5793,N_6458);
nand U8897 (N_8897,N_5559,N_7367);
nor U8898 (N_8898,N_7003,N_7505);
or U8899 (N_8899,N_4240,N_4769);
and U8900 (N_8900,N_6146,N_7709);
nand U8901 (N_8901,N_6218,N_6121);
or U8902 (N_8902,N_5734,N_5656);
nor U8903 (N_8903,N_4134,N_4465);
nand U8904 (N_8904,N_7128,N_4535);
xor U8905 (N_8905,N_4096,N_5371);
nand U8906 (N_8906,N_6641,N_5943);
and U8907 (N_8907,N_6988,N_5703);
or U8908 (N_8908,N_5254,N_6064);
nor U8909 (N_8909,N_5453,N_7755);
nor U8910 (N_8910,N_4421,N_5756);
nor U8911 (N_8911,N_7876,N_7955);
xor U8912 (N_8912,N_4600,N_5737);
or U8913 (N_8913,N_7588,N_5696);
and U8914 (N_8914,N_4575,N_7285);
xor U8915 (N_8915,N_5582,N_5259);
nor U8916 (N_8916,N_4152,N_5198);
nor U8917 (N_8917,N_5253,N_6439);
and U8918 (N_8918,N_5937,N_7473);
or U8919 (N_8919,N_7940,N_4301);
and U8920 (N_8920,N_7450,N_5796);
and U8921 (N_8921,N_4742,N_5196);
nand U8922 (N_8922,N_5064,N_5820);
or U8923 (N_8923,N_5951,N_7126);
and U8924 (N_8924,N_6142,N_7490);
nand U8925 (N_8925,N_5306,N_6495);
nand U8926 (N_8926,N_6983,N_7477);
and U8927 (N_8927,N_7803,N_7824);
xnor U8928 (N_8928,N_7431,N_5632);
and U8929 (N_8929,N_5180,N_5851);
xor U8930 (N_8930,N_7580,N_7926);
xor U8931 (N_8931,N_4516,N_6842);
or U8932 (N_8932,N_4444,N_5516);
or U8933 (N_8933,N_4132,N_7377);
nand U8934 (N_8934,N_6618,N_5157);
nor U8935 (N_8935,N_6766,N_4711);
nand U8936 (N_8936,N_4477,N_4196);
nand U8937 (N_8937,N_6358,N_7970);
xor U8938 (N_8938,N_6532,N_6668);
xor U8939 (N_8939,N_4976,N_4954);
nand U8940 (N_8940,N_6324,N_7349);
and U8941 (N_8941,N_6258,N_5190);
xor U8942 (N_8942,N_7984,N_6078);
nand U8943 (N_8943,N_5869,N_7306);
nand U8944 (N_8944,N_6981,N_7801);
or U8945 (N_8945,N_6235,N_4055);
nand U8946 (N_8946,N_6101,N_6989);
and U8947 (N_8947,N_5554,N_5767);
and U8948 (N_8948,N_6998,N_5429);
nand U8949 (N_8949,N_4957,N_6954);
xnor U8950 (N_8950,N_4612,N_6518);
and U8951 (N_8951,N_6095,N_7433);
and U8952 (N_8952,N_6369,N_4650);
nor U8953 (N_8953,N_6996,N_4368);
or U8954 (N_8954,N_5889,N_7011);
nor U8955 (N_8955,N_4222,N_7809);
and U8956 (N_8956,N_5234,N_7933);
or U8957 (N_8957,N_6636,N_7522);
nor U8958 (N_8958,N_7530,N_7402);
xnor U8959 (N_8959,N_6828,N_6003);
nand U8960 (N_8960,N_5440,N_4679);
and U8961 (N_8961,N_7635,N_4078);
nor U8962 (N_8962,N_6802,N_5754);
or U8963 (N_8963,N_7673,N_6939);
nand U8964 (N_8964,N_4570,N_5648);
and U8965 (N_8965,N_7633,N_6093);
nand U8966 (N_8966,N_4956,N_7745);
or U8967 (N_8967,N_5434,N_6648);
and U8968 (N_8968,N_4809,N_6626);
xnor U8969 (N_8969,N_4393,N_7846);
xnor U8970 (N_8970,N_6940,N_7904);
nand U8971 (N_8971,N_7738,N_4482);
nor U8972 (N_8972,N_7370,N_6649);
nor U8973 (N_8973,N_4378,N_5345);
or U8974 (N_8974,N_6945,N_7192);
and U8975 (N_8975,N_7193,N_6109);
and U8976 (N_8976,N_5050,N_5630);
nor U8977 (N_8977,N_4383,N_7032);
xor U8978 (N_8978,N_4995,N_4193);
nand U8979 (N_8979,N_7182,N_6234);
nand U8980 (N_8980,N_4993,N_6911);
and U8981 (N_8981,N_4676,N_4125);
or U8982 (N_8982,N_5215,N_5870);
nand U8983 (N_8983,N_5565,N_5186);
nand U8984 (N_8984,N_6491,N_7025);
nand U8985 (N_8985,N_6248,N_5817);
xor U8986 (N_8986,N_7936,N_5963);
xor U8987 (N_8987,N_7499,N_7663);
and U8988 (N_8988,N_6613,N_5038);
nor U8989 (N_8989,N_5391,N_4081);
or U8990 (N_8990,N_7268,N_5267);
or U8991 (N_8991,N_4282,N_7152);
xor U8992 (N_8992,N_4489,N_5139);
or U8993 (N_8993,N_4931,N_4703);
nor U8994 (N_8994,N_7713,N_7289);
nand U8995 (N_8995,N_5447,N_5701);
nor U8996 (N_8996,N_5700,N_5581);
nand U8997 (N_8997,N_6231,N_5987);
nor U8998 (N_8998,N_4588,N_4578);
and U8999 (N_8999,N_4323,N_7134);
xnor U9000 (N_9000,N_6257,N_7419);
nor U9001 (N_9001,N_5702,N_7699);
nand U9002 (N_9002,N_6640,N_4832);
and U9003 (N_9003,N_7184,N_5805);
or U9004 (N_9004,N_5091,N_7645);
nor U9005 (N_9005,N_5355,N_7614);
nand U9006 (N_9006,N_6890,N_7708);
and U9007 (N_9007,N_7887,N_4464);
or U9008 (N_9008,N_7627,N_5770);
xor U9009 (N_9009,N_6951,N_4443);
nand U9010 (N_9010,N_6323,N_6082);
nand U9011 (N_9011,N_4242,N_5441);
and U9012 (N_9012,N_6880,N_5915);
and U9013 (N_9013,N_6886,N_7732);
xor U9014 (N_9014,N_5210,N_6866);
or U9015 (N_9015,N_5402,N_7010);
xnor U9016 (N_9016,N_5584,N_4162);
or U9017 (N_9017,N_4300,N_6017);
or U9018 (N_9018,N_6643,N_6149);
nor U9019 (N_9019,N_5381,N_6454);
or U9020 (N_9020,N_4928,N_6760);
xnor U9021 (N_9021,N_7622,N_5200);
nor U9022 (N_9022,N_5837,N_4411);
nand U9023 (N_9023,N_6418,N_7049);
and U9024 (N_9024,N_4018,N_4235);
nor U9025 (N_9025,N_7923,N_6357);
xor U9026 (N_9026,N_7153,N_7916);
nand U9027 (N_9027,N_6790,N_5789);
nand U9028 (N_9028,N_6999,N_5022);
and U9029 (N_9029,N_4555,N_6336);
or U9030 (N_9030,N_4408,N_7532);
xor U9031 (N_9031,N_6583,N_6267);
nand U9032 (N_9032,N_7835,N_5188);
and U9033 (N_9033,N_7661,N_7653);
or U9034 (N_9034,N_4049,N_5093);
nor U9035 (N_9035,N_6959,N_5342);
xor U9036 (N_9036,N_7250,N_6355);
and U9037 (N_9037,N_5047,N_6622);
or U9038 (N_9038,N_7135,N_6108);
nand U9039 (N_9039,N_7291,N_6314);
nor U9040 (N_9040,N_7263,N_5658);
or U9041 (N_9041,N_6128,N_7173);
nor U9042 (N_9042,N_7475,N_6276);
and U9043 (N_9043,N_6923,N_4831);
or U9044 (N_9044,N_7384,N_7842);
nor U9045 (N_9045,N_6708,N_4016);
nor U9046 (N_9046,N_6287,N_7939);
nor U9047 (N_9047,N_5728,N_4149);
or U9048 (N_9048,N_6647,N_6486);
and U9049 (N_9049,N_6127,N_5207);
or U9050 (N_9050,N_7893,N_5010);
or U9051 (N_9051,N_6261,N_6745);
nor U9052 (N_9052,N_7430,N_4590);
and U9053 (N_9053,N_4382,N_4266);
and U9054 (N_9054,N_6184,N_5347);
nor U9055 (N_9055,N_5944,N_6345);
nand U9056 (N_9056,N_4304,N_7666);
and U9057 (N_9057,N_5087,N_7368);
nor U9058 (N_9058,N_7875,N_5683);
or U9059 (N_9059,N_4661,N_7956);
xor U9060 (N_9060,N_7639,N_4971);
or U9061 (N_9061,N_5692,N_4723);
xnor U9062 (N_9062,N_6907,N_6771);
and U9063 (N_9063,N_4267,N_5763);
and U9064 (N_9064,N_5003,N_6513);
xor U9065 (N_9065,N_7892,N_5525);
xnor U9066 (N_9066,N_4857,N_7682);
nor U9067 (N_9067,N_6681,N_6691);
xnor U9068 (N_9068,N_6117,N_6073);
or U9069 (N_9069,N_4665,N_5446);
nand U9070 (N_9070,N_5465,N_5827);
or U9071 (N_9071,N_7730,N_5652);
xnor U9072 (N_9072,N_5094,N_7092);
nand U9073 (N_9073,N_7729,N_7215);
and U9074 (N_9074,N_4122,N_7624);
or U9075 (N_9075,N_4119,N_5529);
xor U9076 (N_9076,N_4154,N_5487);
and U9077 (N_9077,N_7777,N_6639);
nand U9078 (N_9078,N_7019,N_6216);
nor U9079 (N_9079,N_4973,N_4399);
and U9080 (N_9080,N_4533,N_5387);
nand U9081 (N_9081,N_4964,N_7566);
nor U9082 (N_9082,N_7095,N_6007);
nand U9083 (N_9083,N_6174,N_7577);
xor U9084 (N_9084,N_4974,N_4816);
nor U9085 (N_9085,N_4525,N_4736);
or U9086 (N_9086,N_4307,N_6059);
nor U9087 (N_9087,N_4434,N_4455);
and U9088 (N_9088,N_4051,N_6527);
nor U9089 (N_9089,N_7217,N_5189);
nor U9090 (N_9090,N_5821,N_6347);
nand U9091 (N_9091,N_4506,N_5577);
and U9092 (N_9092,N_4607,N_7075);
nand U9093 (N_9093,N_6338,N_5484);
xor U9094 (N_9094,N_7524,N_5634);
and U9095 (N_9095,N_5236,N_4178);
xor U9096 (N_9096,N_6961,N_6129);
nand U9097 (N_9097,N_7996,N_7659);
or U9098 (N_9098,N_5081,N_7139);
nand U9099 (N_9099,N_7409,N_7097);
and U9100 (N_9100,N_4702,N_5323);
nand U9101 (N_9101,N_7979,N_7591);
nor U9102 (N_9102,N_7146,N_5375);
or U9103 (N_9103,N_6638,N_4320);
or U9104 (N_9104,N_6027,N_7385);
xor U9105 (N_9105,N_5056,N_5882);
nand U9106 (N_9106,N_6381,N_5543);
and U9107 (N_9107,N_4630,N_5505);
or U9108 (N_9108,N_7178,N_6576);
or U9109 (N_9109,N_6543,N_6102);
xor U9110 (N_9110,N_4001,N_6910);
or U9111 (N_9111,N_5892,N_6222);
or U9112 (N_9112,N_7191,N_4439);
nor U9113 (N_9113,N_6380,N_6388);
nand U9114 (N_9114,N_4476,N_5054);
or U9115 (N_9115,N_5217,N_6516);
nand U9116 (N_9116,N_7610,N_4225);
nand U9117 (N_9117,N_7335,N_4103);
and U9118 (N_9118,N_4729,N_6882);
or U9119 (N_9119,N_5477,N_7705);
nand U9120 (N_9120,N_7050,N_4576);
nor U9121 (N_9121,N_6057,N_4912);
and U9122 (N_9122,N_4027,N_6037);
or U9123 (N_9123,N_6132,N_6899);
xor U9124 (N_9124,N_7046,N_7771);
xor U9125 (N_9125,N_4775,N_7616);
or U9126 (N_9126,N_5078,N_5045);
nor U9127 (N_9127,N_5250,N_4328);
nor U9128 (N_9128,N_7333,N_4852);
and U9129 (N_9129,N_7447,N_6482);
xnor U9130 (N_9130,N_5877,N_4624);
or U9131 (N_9131,N_6023,N_6776);
or U9132 (N_9132,N_6155,N_4847);
nor U9133 (N_9133,N_4717,N_5663);
or U9134 (N_9134,N_4684,N_4751);
nand U9135 (N_9135,N_4108,N_6840);
nand U9136 (N_9136,N_6752,N_4412);
nand U9137 (N_9137,N_5713,N_6973);
nor U9138 (N_9138,N_6487,N_6616);
nand U9139 (N_9139,N_4741,N_7233);
or U9140 (N_9140,N_6865,N_7972);
xor U9141 (N_9141,N_7605,N_5856);
xnor U9142 (N_9142,N_7235,N_7895);
nor U9143 (N_9143,N_7539,N_7418);
or U9144 (N_9144,N_6818,N_5120);
xor U9145 (N_9145,N_6550,N_4566);
nor U9146 (N_9146,N_7971,N_4846);
nor U9147 (N_9147,N_5871,N_6025);
xor U9148 (N_9148,N_5107,N_6792);
nand U9149 (N_9149,N_5195,N_6005);
and U9150 (N_9150,N_6000,N_7740);
or U9151 (N_9151,N_5170,N_4433);
and U9152 (N_9152,N_7894,N_6148);
or U9153 (N_9153,N_5809,N_4709);
xor U9154 (N_9154,N_4387,N_4043);
nor U9155 (N_9155,N_7361,N_4622);
nor U9156 (N_9156,N_5885,N_6918);
or U9157 (N_9157,N_7090,N_5571);
nor U9158 (N_9158,N_5384,N_5844);
nand U9159 (N_9159,N_4797,N_4006);
nand U9160 (N_9160,N_4984,N_5536);
or U9161 (N_9161,N_6663,N_6052);
or U9162 (N_9162,N_4076,N_7084);
nor U9163 (N_9163,N_6424,N_5479);
xnor U9164 (N_9164,N_7466,N_7498);
nand U9165 (N_9165,N_7489,N_5036);
xnor U9166 (N_9166,N_4126,N_4673);
or U9167 (N_9167,N_4623,N_5492);
nand U9168 (N_9168,N_7891,N_7609);
nor U9169 (N_9169,N_5778,N_6488);
nand U9170 (N_9170,N_6904,N_4365);
or U9171 (N_9171,N_5636,N_5667);
nand U9172 (N_9172,N_5031,N_5366);
and U9173 (N_9173,N_4402,N_5224);
nand U9174 (N_9174,N_6753,N_4789);
nor U9175 (N_9175,N_6032,N_5791);
nor U9176 (N_9176,N_5579,N_7260);
nand U9177 (N_9177,N_5724,N_5935);
nand U9178 (N_9178,N_6351,N_6512);
xor U9179 (N_9179,N_4097,N_5324);
nor U9180 (N_9180,N_5807,N_5307);
or U9181 (N_9181,N_7796,N_4481);
and U9182 (N_9182,N_4830,N_7696);
nor U9183 (N_9183,N_6757,N_7073);
and U9184 (N_9184,N_5570,N_7456);
or U9185 (N_9185,N_7641,N_5156);
nor U9186 (N_9186,N_4980,N_6969);
xor U9187 (N_9187,N_5580,N_4568);
and U9188 (N_9188,N_4720,N_6755);
nand U9189 (N_9189,N_5095,N_4819);
xor U9190 (N_9190,N_5321,N_6500);
and U9191 (N_9191,N_6594,N_5028);
nor U9192 (N_9192,N_5202,N_5280);
nor U9193 (N_9193,N_7567,N_5606);
nor U9194 (N_9194,N_7325,N_4123);
or U9195 (N_9195,N_5727,N_5237);
or U9196 (N_9196,N_4638,N_4982);
or U9197 (N_9197,N_7460,N_4887);
and U9198 (N_9198,N_5336,N_4734);
or U9199 (N_9199,N_7529,N_7322);
or U9200 (N_9200,N_7746,N_6601);
nor U9201 (N_9201,N_7948,N_6845);
nand U9202 (N_9202,N_5707,N_6207);
and U9203 (N_9203,N_7343,N_7694);
nand U9204 (N_9204,N_7021,N_4549);
and U9205 (N_9205,N_5406,N_7463);
nand U9206 (N_9206,N_5970,N_4199);
or U9207 (N_9207,N_7251,N_4652);
xnor U9208 (N_9208,N_7199,N_4864);
nor U9209 (N_9209,N_4249,N_6193);
xnor U9210 (N_9210,N_5098,N_5592);
xnor U9211 (N_9211,N_7695,N_7086);
nor U9212 (N_9212,N_4950,N_7747);
nand U9213 (N_9213,N_6870,N_5311);
or U9214 (N_9214,N_7341,N_7467);
or U9215 (N_9215,N_7907,N_6452);
nor U9216 (N_9216,N_5642,N_4899);
or U9217 (N_9217,N_6353,N_5569);
xor U9218 (N_9218,N_4560,N_7843);
or U9219 (N_9219,N_7127,N_4424);
nand U9220 (N_9220,N_4003,N_5176);
and U9221 (N_9221,N_4287,N_6499);
and U9222 (N_9222,N_7630,N_4694);
nand U9223 (N_9223,N_5086,N_7945);
nand U9224 (N_9224,N_5862,N_7167);
or U9225 (N_9225,N_7020,N_5835);
nand U9226 (N_9226,N_6209,N_6150);
and U9227 (N_9227,N_4019,N_7204);
xnor U9228 (N_9228,N_4551,N_4501);
nand U9229 (N_9229,N_7913,N_7571);
or U9230 (N_9230,N_4129,N_4377);
or U9231 (N_9231,N_7977,N_4497);
or U9232 (N_9232,N_6851,N_4966);
or U9233 (N_9233,N_7525,N_5768);
nor U9234 (N_9234,N_7137,N_5394);
and U9235 (N_9235,N_7136,N_6441);
and U9236 (N_9236,N_7247,N_5788);
and U9237 (N_9237,N_6125,N_7398);
and U9238 (N_9238,N_6653,N_5785);
or U9239 (N_9239,N_5964,N_6241);
nor U9240 (N_9240,N_4920,N_6791);
or U9241 (N_9241,N_6362,N_6153);
nor U9242 (N_9242,N_6630,N_5303);
nor U9243 (N_9243,N_6115,N_4176);
nor U9244 (N_9244,N_6020,N_4423);
nand U9245 (N_9245,N_6786,N_5924);
or U9246 (N_9246,N_5382,N_4380);
and U9247 (N_9247,N_6008,N_5294);
nor U9248 (N_9248,N_7008,N_5549);
nand U9249 (N_9249,N_4693,N_6553);
nand U9250 (N_9250,N_7572,N_6473);
nand U9251 (N_9251,N_4212,N_7353);
nand U9252 (N_9252,N_4783,N_5784);
xnor U9253 (N_9253,N_4064,N_5000);
nand U9254 (N_9254,N_4765,N_4526);
and U9255 (N_9255,N_6160,N_6789);
nor U9256 (N_9256,N_7813,N_7999);
nor U9257 (N_9257,N_6334,N_5830);
xnor U9258 (N_9258,N_5847,N_5509);
nand U9259 (N_9259,N_6483,N_5187);
nand U9260 (N_9260,N_5506,N_5646);
and U9261 (N_9261,N_5587,N_4060);
nand U9262 (N_9262,N_7617,N_4403);
nor U9263 (N_9263,N_5836,N_5226);
or U9264 (N_9264,N_5749,N_7318);
or U9265 (N_9265,N_6120,N_4474);
nor U9266 (N_9266,N_6984,N_6168);
and U9267 (N_9267,N_4068,N_7362);
xor U9268 (N_9268,N_4182,N_7736);
nand U9269 (N_9269,N_5088,N_5161);
or U9270 (N_9270,N_7851,N_5771);
xnor U9271 (N_9271,N_6676,N_7472);
nand U9272 (N_9272,N_6417,N_4985);
xor U9273 (N_9273,N_7558,N_4082);
nand U9274 (N_9274,N_4346,N_7748);
and U9275 (N_9275,N_5966,N_5034);
nor U9276 (N_9276,N_5568,N_7000);
or U9277 (N_9277,N_5065,N_7295);
nand U9278 (N_9278,N_4722,N_4554);
and U9279 (N_9279,N_6030,N_7502);
xnor U9280 (N_9280,N_4000,N_7439);
or U9281 (N_9281,N_7234,N_4951);
and U9282 (N_9282,N_7648,N_4052);
nor U9283 (N_9283,N_6136,N_4648);
or U9284 (N_9284,N_5659,N_4996);
or U9285 (N_9285,N_5383,N_7799);
and U9286 (N_9286,N_6246,N_5076);
or U9287 (N_9287,N_7669,N_4627);
and U9288 (N_9288,N_5388,N_6867);
nand U9289 (N_9289,N_7355,N_7519);
nor U9290 (N_9290,N_4318,N_5209);
nor U9291 (N_9291,N_7601,N_7927);
or U9292 (N_9292,N_4540,N_6015);
nand U9293 (N_9293,N_4785,N_6629);
and U9294 (N_9294,N_7697,N_7664);
nand U9295 (N_9295,N_6208,N_6738);
or U9296 (N_9296,N_6140,N_4666);
xnor U9297 (N_9297,N_4786,N_7968);
or U9298 (N_9298,N_4979,N_4613);
nor U9299 (N_9299,N_5033,N_4934);
nand U9300 (N_9300,N_5858,N_7326);
xor U9301 (N_9301,N_7899,N_6019);
nand U9302 (N_9302,N_5006,N_5773);
and U9303 (N_9303,N_6908,N_5380);
nor U9304 (N_9304,N_7775,N_4306);
or U9305 (N_9305,N_6572,N_7486);
nor U9306 (N_9306,N_4239,N_4758);
xnor U9307 (N_9307,N_6490,N_7782);
nor U9308 (N_9308,N_7357,N_6526);
and U9309 (N_9309,N_6244,N_4404);
nand U9310 (N_9310,N_6434,N_7564);
and U9311 (N_9311,N_4935,N_4343);
and U9312 (N_9312,N_7397,N_6718);
or U9313 (N_9313,N_5329,N_6693);
or U9314 (N_9314,N_7236,N_7436);
or U9315 (N_9315,N_5206,N_5829);
or U9316 (N_9316,N_6615,N_6678);
nor U9317 (N_9317,N_6303,N_7821);
and U9318 (N_9318,N_5945,N_5677);
or U9319 (N_9319,N_4645,N_5879);
xnor U9320 (N_9320,N_7069,N_4777);
nand U9321 (N_9321,N_7714,N_5926);
xnor U9322 (N_9322,N_5468,N_5873);
nand U9323 (N_9323,N_4233,N_7455);
and U9324 (N_9324,N_7040,N_7541);
nand U9325 (N_9325,N_5111,N_7223);
and U9326 (N_9326,N_6646,N_4137);
nor U9327 (N_9327,N_5452,N_6557);
nand U9328 (N_9328,N_7754,N_5833);
nor U9329 (N_9329,N_7995,N_7500);
and U9330 (N_9330,N_5344,N_4340);
nor U9331 (N_9331,N_6342,N_7181);
or U9332 (N_9332,N_6296,N_5199);
and U9333 (N_9333,N_4036,N_6896);
nand U9334 (N_9334,N_6574,N_6740);
or U9335 (N_9335,N_4531,N_6308);
or U9336 (N_9336,N_7547,N_6671);
xor U9337 (N_9337,N_4344,N_7494);
nor U9338 (N_9338,N_5593,N_7276);
nor U9339 (N_9339,N_5799,N_6934);
or U9340 (N_9340,N_6855,N_4635);
nor U9341 (N_9341,N_6686,N_5255);
xnor U9342 (N_9342,N_6126,N_7631);
and U9343 (N_9343,N_6226,N_7105);
nand U9344 (N_9344,N_6785,N_4611);
nor U9345 (N_9345,N_6481,N_4369);
and U9346 (N_9346,N_4209,N_7275);
xor U9347 (N_9347,N_4135,N_5482);
nand U9348 (N_9348,N_5458,N_4953);
and U9349 (N_9349,N_7625,N_7387);
nor U9350 (N_9350,N_4707,N_5846);
xor U9351 (N_9351,N_4084,N_6808);
and U9352 (N_9352,N_4904,N_5532);
xnor U9353 (N_9353,N_5910,N_4026);
nand U9354 (N_9354,N_4674,N_5548);
nor U9355 (N_9355,N_4524,N_6571);
or U9356 (N_9356,N_7802,N_6719);
nor U9357 (N_9357,N_7443,N_7602);
nand U9358 (N_9358,N_7731,N_4198);
xnor U9359 (N_9359,N_5564,N_7113);
or U9360 (N_9360,N_5953,N_5697);
and U9361 (N_9361,N_7958,N_4606);
or U9362 (N_9362,N_6348,N_7332);
nor U9363 (N_9363,N_7225,N_4203);
nand U9364 (N_9364,N_7944,N_7379);
and U9365 (N_9365,N_6137,N_5884);
or U9366 (N_9366,N_5026,N_4565);
xnor U9367 (N_9367,N_6277,N_5745);
and U9368 (N_9368,N_7479,N_5782);
and U9369 (N_9369,N_6924,N_4156);
nor U9370 (N_9370,N_6712,N_5288);
nor U9371 (N_9371,N_4069,N_5079);
and U9372 (N_9372,N_6377,N_6203);
xnor U9373 (N_9373,N_7908,N_6684);
xor U9374 (N_9374,N_6285,N_5859);
xnor U9375 (N_9375,N_4946,N_5023);
nand U9376 (N_9376,N_4180,N_5631);
or U9377 (N_9377,N_6374,N_4400);
or U9378 (N_9378,N_6186,N_6067);
xor U9379 (N_9379,N_5279,N_4823);
and U9380 (N_9380,N_4438,N_7667);
nor U9381 (N_9381,N_4913,N_4795);
or U9382 (N_9382,N_7991,N_4099);
xnor U9383 (N_9383,N_7031,N_7258);
xnor U9384 (N_9384,N_6309,N_4095);
and U9385 (N_9385,N_5377,N_7668);
and U9386 (N_9386,N_4559,N_5461);
and U9387 (N_9387,N_5716,N_6464);
xnor U9388 (N_9388,N_6517,N_6854);
nor U9389 (N_9389,N_5174,N_5588);
xor U9390 (N_9390,N_6967,N_5439);
nand U9391 (N_9391,N_6339,N_5748);
nor U9392 (N_9392,N_7836,N_7953);
nand U9393 (N_9393,N_4040,N_4811);
or U9394 (N_9394,N_4882,N_7514);
and U9395 (N_9395,N_5103,N_5852);
and U9396 (N_9396,N_6058,N_6530);
or U9397 (N_9397,N_4911,N_7787);
xor U9398 (N_9398,N_5604,N_6284);
nor U9399 (N_9399,N_5016,N_6390);
nand U9400 (N_9400,N_5500,N_7902);
or U9401 (N_9401,N_7417,N_6529);
and U9402 (N_9402,N_6497,N_4691);
xor U9403 (N_9403,N_5137,N_7147);
and U9404 (N_9404,N_6158,N_5691);
nand U9405 (N_9405,N_7196,N_7759);
nand U9406 (N_9406,N_6788,N_5333);
and U9407 (N_9407,N_5733,N_5373);
nor U9408 (N_9408,N_6874,N_5313);
or U9409 (N_9409,N_7912,N_7266);
and U9410 (N_9410,N_7336,N_7078);
xor U9411 (N_9411,N_4922,N_4211);
nand U9412 (N_9412,N_7952,N_6654);
and U9413 (N_9413,N_4236,N_4357);
nor U9414 (N_9414,N_7963,N_7593);
nor U9415 (N_9415,N_5346,N_7712);
nand U9416 (N_9416,N_7857,N_7608);
and U9417 (N_9417,N_7053,N_6804);
nor U9418 (N_9418,N_5315,N_5515);
and U9419 (N_9419,N_5722,N_5546);
or U9420 (N_9420,N_4845,N_4989);
nand U9421 (N_9421,N_6382,N_5075);
xor U9422 (N_9422,N_5007,N_6089);
or U9423 (N_9423,N_6778,N_4264);
xnor U9424 (N_9424,N_6603,N_4519);
xor U9425 (N_9425,N_7408,N_6857);
or U9426 (N_9426,N_6762,N_5297);
nor U9427 (N_9427,N_7484,N_7270);
nor U9428 (N_9428,N_5689,N_6428);
xor U9429 (N_9429,N_4261,N_5148);
nor U9430 (N_9430,N_5147,N_5994);
nand U9431 (N_9431,N_4651,N_7623);
nor U9432 (N_9432,N_5814,N_4511);
nor U9433 (N_9433,N_6041,N_5235);
nand U9434 (N_9434,N_6219,N_7620);
xor U9435 (N_9435,N_6467,N_5244);
nand U9436 (N_9436,N_6775,N_6080);
xnor U9437 (N_9437,N_7584,N_5362);
or U9438 (N_9438,N_4262,N_5405);
or U9439 (N_9439,N_4806,N_7482);
or U9440 (N_9440,N_5302,N_5865);
or U9441 (N_9441,N_6706,N_6836);
xor U9442 (N_9442,N_6068,N_6113);
nand U9443 (N_9443,N_6633,N_7158);
nand U9444 (N_9444,N_7562,N_6705);
xor U9445 (N_9445,N_4181,N_4185);
xor U9446 (N_9446,N_7828,N_6879);
nand U9447 (N_9447,N_6644,N_6682);
xor U9448 (N_9448,N_4602,N_6183);
nor U9449 (N_9449,N_7125,N_4428);
nor U9450 (N_9450,N_7785,N_4356);
nor U9451 (N_9451,N_5126,N_6559);
or U9452 (N_9452,N_7992,N_5155);
xor U9453 (N_9453,N_4372,N_5040);
and U9454 (N_9454,N_6657,N_4473);
or U9455 (N_9455,N_4109,N_4011);
nor U9456 (N_9456,N_7678,N_5645);
nand U9457 (N_9457,N_4573,N_7762);
xnor U9458 (N_9458,N_4020,N_6180);
or U9459 (N_9459,N_6416,N_4374);
and U9460 (N_9460,N_6021,N_4659);
nor U9461 (N_9461,N_7790,N_6227);
nand U9462 (N_9462,N_5102,N_4322);
and U9463 (N_9463,N_5472,N_4572);
or U9464 (N_9464,N_4314,N_6275);
xnor U9465 (N_9465,N_4094,N_7654);
nand U9466 (N_9466,N_7656,N_7168);
nand U9467 (N_9467,N_7737,N_5089);
nand U9468 (N_9468,N_4022,N_7535);
nor U9469 (N_9469,N_5121,N_7062);
xor U9470 (N_9470,N_4716,N_7691);
xor U9471 (N_9471,N_7027,N_7096);
nor U9472 (N_9472,N_6503,N_5019);
xnor U9473 (N_9473,N_7961,N_7868);
and U9474 (N_9474,N_4738,N_4653);
or U9475 (N_9475,N_6610,N_4842);
xor U9476 (N_9476,N_6356,N_6864);
nor U9477 (N_9477,N_7242,N_4111);
nor U9478 (N_9478,N_6835,N_6905);
xor U9479 (N_9479,N_4732,N_6986);
and U9480 (N_9480,N_4462,N_7317);
nor U9481 (N_9481,N_6893,N_4229);
nor U9482 (N_9482,N_5114,N_7947);
nand U9483 (N_9483,N_6634,N_6445);
nand U9484 (N_9484,N_7394,N_5572);
nand U9485 (N_9485,N_6737,N_6714);
and U9486 (N_9486,N_5906,N_4155);
nand U9487 (N_9487,N_5905,N_6538);
nand U9488 (N_9488,N_4938,N_7406);
xor U9489 (N_9489,N_6724,N_5131);
nor U9490 (N_9490,N_4994,N_6667);
nand U9491 (N_9491,N_5556,N_5001);
nand U9492 (N_9492,N_5672,N_5108);
nor U9493 (N_9493,N_7476,N_6298);
or U9494 (N_9494,N_7239,N_4143);
and U9495 (N_9495,N_5052,N_6202);
xor U9496 (N_9496,N_4146,N_7885);
xor U9497 (N_9497,N_5709,N_5918);
xor U9498 (N_9498,N_4637,N_7183);
nor U9499 (N_9499,N_6290,N_7901);
nand U9500 (N_9500,N_7453,N_7573);
xnor U9501 (N_9501,N_6656,N_6820);
nand U9502 (N_9502,N_4841,N_6831);
xnor U9503 (N_9503,N_5314,N_6796);
and U9504 (N_9504,N_4172,N_4756);
or U9505 (N_9505,N_4698,N_6286);
nand U9506 (N_9506,N_6695,N_5704);
nand U9507 (N_9507,N_6088,N_6811);
nor U9508 (N_9508,N_5037,N_5144);
or U9509 (N_9509,N_7551,N_5662);
nand U9510 (N_9510,N_6190,N_4688);
nor U9511 (N_9511,N_6205,N_6928);
or U9512 (N_9512,N_5127,N_5922);
nand U9513 (N_9513,N_4940,N_5675);
xnor U9514 (N_9514,N_5231,N_6009);
nor U9515 (N_9515,N_7009,N_6900);
or U9516 (N_9516,N_4490,N_6185);
or U9517 (N_9517,N_4897,N_5118);
nor U9518 (N_9518,N_7241,N_6119);
nand U9519 (N_9519,N_5379,N_6936);
and U9520 (N_9520,N_4633,N_4430);
nand U9521 (N_9521,N_7213,N_6159);
xnor U9522 (N_9522,N_6598,N_7883);
and U9523 (N_9523,N_4278,N_4770);
or U9524 (N_9524,N_5326,N_5261);
and U9525 (N_9525,N_6795,N_4721);
and U9526 (N_9526,N_4534,N_4801);
and U9527 (N_9527,N_6732,N_4778);
xnor U9528 (N_9528,N_4905,N_7312);
nand U9529 (N_9529,N_5162,N_6395);
nand U9530 (N_9530,N_7273,N_6943);
xor U9531 (N_9531,N_6758,N_7793);
or U9532 (N_9532,N_5059,N_4618);
and U9533 (N_9533,N_7393,N_4184);
and U9534 (N_9534,N_7856,N_5220);
nand U9535 (N_9535,N_6966,N_6098);
and U9536 (N_9536,N_6278,N_5955);
or U9537 (N_9537,N_7106,N_4715);
nand U9538 (N_9538,N_7424,N_7319);
xor U9539 (N_9539,N_7133,N_5233);
nor U9540 (N_9540,N_6496,N_6288);
or U9541 (N_9541,N_5638,N_5289);
nand U9542 (N_9542,N_6582,N_7189);
xnor U9543 (N_9543,N_4479,N_4574);
nand U9544 (N_9544,N_5154,N_6619);
nor U9545 (N_9545,N_4784,N_7109);
and U9546 (N_9546,N_4828,N_6669);
and U9547 (N_9547,N_6312,N_7150);
nor U9548 (N_9548,N_6801,N_6635);
and U9549 (N_9549,N_7045,N_5281);
nor U9550 (N_9550,N_6612,N_4502);
and U9551 (N_9551,N_6570,N_6484);
or U9552 (N_9552,N_6534,N_5339);
or U9553 (N_9553,N_4579,N_4948);
nor U9554 (N_9554,N_4206,N_5537);
xnor U9555 (N_9555,N_7727,N_4791);
and U9556 (N_9556,N_4605,N_5057);
or U9557 (N_9557,N_4127,N_7369);
xnor U9558 (N_9558,N_4561,N_7683);
or U9559 (N_9559,N_6366,N_6038);
or U9560 (N_9560,N_4360,N_6033);
nor U9561 (N_9561,N_6096,N_5925);
xnor U9562 (N_9562,N_5185,N_5071);
xor U9563 (N_9563,N_7726,N_4804);
nand U9564 (N_9564,N_5968,N_4875);
nor U9565 (N_9565,N_6293,N_6661);
and U9566 (N_9566,N_4877,N_5291);
nand U9567 (N_9567,N_4780,N_5263);
xnor U9568 (N_9568,N_5853,N_5635);
xnor U9569 (N_9569,N_7840,N_4960);
xor U9570 (N_9570,N_6504,N_5985);
xnor U9571 (N_9571,N_4925,N_6781);
nor U9572 (N_9572,N_6860,N_6763);
nor U9573 (N_9573,N_6767,N_7396);
xor U9574 (N_9574,N_5475,N_4876);
and U9575 (N_9575,N_5514,N_5961);
and U9576 (N_9576,N_5361,N_7675);
xor U9577 (N_9577,N_5806,N_5140);
nand U9578 (N_9578,N_5020,N_6711);
nand U9579 (N_9579,N_5653,N_7013);
nor U9580 (N_9580,N_5759,N_4325);
nor U9581 (N_9581,N_6957,N_6045);
nand U9582 (N_9582,N_4014,N_5730);
nand U9583 (N_9583,N_7036,N_7022);
xor U9584 (N_9584,N_7228,N_6607);
nor U9585 (N_9585,N_5039,N_6397);
nand U9586 (N_9586,N_6238,N_4706);
xor U9587 (N_9587,N_5164,N_5958);
xnor U9588 (N_9588,N_7337,N_6204);
nand U9589 (N_9589,N_5247,N_4746);
nor U9590 (N_9590,N_7288,N_4542);
and U9591 (N_9591,N_7180,N_7781);
and U9592 (N_9592,N_5979,N_5950);
nor U9593 (N_9593,N_5655,N_4362);
and U9594 (N_9594,N_7749,N_4376);
and U9595 (N_9595,N_6652,N_6412);
xor U9596 (N_9596,N_7206,N_5940);
xor U9597 (N_9597,N_4386,N_5101);
nor U9598 (N_9598,N_4955,N_6076);
nand U9599 (N_9599,N_4395,N_5030);
nor U9600 (N_9600,N_5269,N_4998);
nand U9601 (N_9601,N_7783,N_7557);
and U9602 (N_9602,N_7425,N_7864);
or U9603 (N_9603,N_7817,N_4970);
and U9604 (N_9604,N_4037,N_5496);
nand U9605 (N_9605,N_5670,N_5213);
and U9606 (N_9606,N_6861,N_7556);
or U9607 (N_9607,N_6577,N_5928);
nor U9608 (N_9608,N_5417,N_6830);
nor U9609 (N_9609,N_6690,N_6402);
xor U9610 (N_9610,N_4484,N_6182);
nor U9611 (N_9611,N_6507,N_5866);
nor U9612 (N_9612,N_5276,N_7200);
nor U9613 (N_9613,N_4735,N_5282);
nor U9614 (N_9614,N_4028,N_6535);
nand U9615 (N_9615,N_5772,N_6212);
xnor U9616 (N_9616,N_4632,N_6863);
and U9617 (N_9617,N_7254,N_6106);
and U9618 (N_9618,N_5981,N_4737);
or U9619 (N_9619,N_5443,N_7881);
or U9620 (N_9620,N_7703,N_5521);
xor U9621 (N_9621,N_6084,N_7448);
xnor U9622 (N_9622,N_5409,N_7358);
nand U9623 (N_9623,N_5074,N_4483);
xor U9624 (N_9624,N_7219,N_6147);
nor U9625 (N_9625,N_4280,N_6680);
and U9626 (N_9626,N_5719,N_4197);
xnor U9627 (N_9627,N_5893,N_6588);
or U9628 (N_9628,N_4319,N_7552);
and U9629 (N_9629,N_7520,N_7334);
xor U9630 (N_9630,N_5457,N_5049);
nand U9631 (N_9631,N_6111,N_7873);
nand U9632 (N_9632,N_4733,N_6933);
and U9633 (N_9633,N_5640,N_7960);
nor U9634 (N_9634,N_7692,N_4626);
and U9635 (N_9635,N_5109,N_7993);
nor U9636 (N_9636,N_4364,N_4696);
and U9637 (N_9637,N_6600,N_6875);
or U9638 (N_9638,N_6090,N_4075);
or U9639 (N_9639,N_7768,N_6232);
nand U9640 (N_9640,N_5335,N_7941);
and U9641 (N_9641,N_6442,N_5595);
xnor U9642 (N_9642,N_5258,N_5498);
xnor U9643 (N_9643,N_6176,N_6696);
nor U9644 (N_9644,N_6455,N_5338);
or U9645 (N_9645,N_5825,N_6004);
nand U9646 (N_9646,N_5978,N_6249);
xor U9647 (N_9647,N_7091,N_4100);
nand U9648 (N_9648,N_5761,N_6697);
xnor U9649 (N_9649,N_4991,N_5776);
and U9650 (N_9650,N_6254,N_4621);
and U9651 (N_9651,N_5367,N_6485);
or U9652 (N_9652,N_4601,N_6074);
and U9653 (N_9653,N_4752,N_7350);
nor U9654 (N_9654,N_5673,N_5988);
nor U9655 (N_9655,N_5628,N_4958);
or U9656 (N_9656,N_6568,N_4508);
and U9657 (N_9657,N_7778,N_5172);
nand U9658 (N_9658,N_7354,N_4628);
or U9659 (N_9659,N_5823,N_7548);
xnor U9660 (N_9660,N_5766,N_5503);
or U9661 (N_9661,N_4669,N_7823);
and U9662 (N_9662,N_6614,N_7811);
nand U9663 (N_9663,N_4461,N_5956);
and U9664 (N_9664,N_4289,N_7434);
xor U9665 (N_9665,N_7451,N_4615);
nor U9666 (N_9666,N_7240,N_5711);
nand U9667 (N_9667,N_4805,N_5752);
xor U9668 (N_9668,N_5816,N_5442);
nand U9669 (N_9669,N_6310,N_5687);
and U9670 (N_9670,N_7866,N_7554);
and U9671 (N_9671,N_7452,N_4761);
and U9672 (N_9672,N_7867,N_5113);
nand U9673 (N_9673,N_4859,N_6469);
xor U9674 (N_9674,N_6715,N_7108);
and U9675 (N_9675,N_6001,N_6422);
and U9676 (N_9676,N_6871,N_7087);
xor U9677 (N_9677,N_6891,N_4586);
nor U9678 (N_9678,N_4825,N_4937);
nand U9679 (N_9679,N_4813,N_7243);
and U9680 (N_9680,N_5265,N_5682);
or U9681 (N_9681,N_4499,N_7121);
and U9682 (N_9682,N_5649,N_4705);
or U9683 (N_9683,N_5528,N_6687);
nand U9684 (N_9684,N_7512,N_5610);
and U9685 (N_9685,N_7798,N_5221);
nor U9686 (N_9686,N_5674,N_7637);
and U9687 (N_9687,N_6645,N_7103);
nor U9688 (N_9688,N_5085,N_4258);
nand U9689 (N_9689,N_6333,N_4754);
nand U9690 (N_9690,N_7161,N_6946);
xnor U9691 (N_9691,N_5272,N_6519);
nor U9692 (N_9692,N_4231,N_4807);
and U9693 (N_9693,N_4139,N_5104);
nand U9694 (N_9694,N_6925,N_4042);
nand U9695 (N_9695,N_7579,N_7538);
xor U9696 (N_9696,N_4889,N_7698);
or U9697 (N_9697,N_5090,N_7170);
nand U9698 (N_9698,N_5229,N_4647);
or U9699 (N_9699,N_6593,N_6611);
nand U9700 (N_9700,N_7111,N_7570);
xnor U9701 (N_9701,N_7504,N_6930);
and U9702 (N_9702,N_6821,N_7672);
or U9703 (N_9703,N_4339,N_6673);
or U9704 (N_9704,N_6849,N_7833);
nor U9705 (N_9705,N_5378,N_6735);
and U9706 (N_9706,N_7493,N_7898);
and U9707 (N_9707,N_7301,N_4800);
or U9708 (N_9708,N_7061,N_7543);
or U9709 (N_9709,N_7863,N_4512);
and U9710 (N_9710,N_7123,N_5685);
xnor U9711 (N_9711,N_7988,N_7501);
xnor U9712 (N_9712,N_6834,N_4179);
or U9713 (N_9713,N_6436,N_7596);
nor U9714 (N_9714,N_4774,N_6713);
nor U9715 (N_9715,N_5389,N_5522);
nand U9716 (N_9716,N_4145,N_7990);
xnor U9717 (N_9717,N_7006,N_7937);
nor U9718 (N_9718,N_6812,N_5365);
or U9719 (N_9719,N_4641,N_6580);
nor U9720 (N_9720,N_4204,N_4571);
or U9721 (N_9721,N_7942,N_7850);
and U9722 (N_9722,N_6921,N_7660);
and U9723 (N_9723,N_5679,N_4794);
nand U9724 (N_9724,N_4814,N_4050);
or U9725 (N_9725,N_5881,N_7874);
or U9726 (N_9726,N_5299,N_4098);
nand U9727 (N_9727,N_4077,N_5249);
and U9728 (N_9728,N_7758,N_4610);
and U9729 (N_9729,N_6659,N_4293);
and U9730 (N_9730,N_5783,N_5015);
xnor U9731 (N_9731,N_5117,N_4102);
and U9732 (N_9732,N_5596,N_6750);
nor U9733 (N_9733,N_7413,N_6736);
and U9734 (N_9734,N_4658,N_6151);
nor U9735 (N_9735,N_4265,N_7563);
and U9736 (N_9736,N_4138,N_7280);
nor U9737 (N_9737,N_6139,N_4840);
and U9738 (N_9738,N_5061,N_5688);
nand U9739 (N_9739,N_6270,N_5486);
and U9740 (N_9740,N_5639,N_4002);
nand U9741 (N_9741,N_4370,N_5841);
or U9742 (N_9742,N_4352,N_5305);
nor U9743 (N_9743,N_5116,N_4924);
and U9744 (N_9744,N_5695,N_4121);
and U9745 (N_9745,N_7909,N_5459);
nor U9746 (N_9746,N_7412,N_7847);
nand U9747 (N_9747,N_4748,N_6344);
xor U9748 (N_9748,N_5519,N_5942);
nor U9749 (N_9749,N_7093,N_7884);
nor U9750 (N_9750,N_7314,N_7848);
or U9751 (N_9751,N_5609,N_4044);
nand U9752 (N_9752,N_5725,N_7574);
and U9753 (N_9753,N_7211,N_7521);
nor U9754 (N_9754,N_4856,N_5929);
and U9755 (N_9755,N_5896,N_7454);
and U9756 (N_9756,N_7469,N_4459);
or U9757 (N_9757,N_4065,N_7764);
or U9758 (N_9758,N_5742,N_7162);
and U9759 (N_9759,N_6447,N_4664);
and U9760 (N_9760,N_4292,N_5875);
xor U9761 (N_9761,N_7281,N_4436);
nand U9762 (N_9762,N_6423,N_4087);
nor U9763 (N_9763,N_4165,N_5386);
or U9764 (N_9764,N_7043,N_7376);
and U9765 (N_9765,N_6596,N_6431);
and U9766 (N_9766,N_5786,N_5657);
and U9767 (N_9767,N_4978,N_4407);
nand U9768 (N_9768,N_4530,N_5240);
nand U9769 (N_9769,N_5260,N_6536);
or U9770 (N_9770,N_7373,N_7330);
and U9771 (N_9771,N_4168,N_5184);
nand U9772 (N_9772,N_4410,N_5845);
nand U9773 (N_9773,N_4719,N_4504);
or U9774 (N_9774,N_5251,N_6809);
nor U9775 (N_9775,N_6040,N_4865);
or U9776 (N_9776,N_7067,N_6492);
nand U9777 (N_9777,N_6722,N_5738);
or U9778 (N_9778,N_7070,N_4639);
or U9779 (N_9779,N_5275,N_5887);
nand U9780 (N_9780,N_6266,N_7382);
and U9781 (N_9781,N_6602,N_4005);
nand U9782 (N_9782,N_6263,N_6131);
nor U9783 (N_9783,N_5949,N_5480);
nand U9784 (N_9784,N_4527,N_5222);
or U9785 (N_9785,N_4025,N_4788);
nor U9786 (N_9786,N_6655,N_5842);
or U9787 (N_9787,N_5560,N_5573);
nor U9788 (N_9788,N_6816,N_5283);
or U9789 (N_9789,N_6817,N_7114);
nor U9790 (N_9790,N_7342,N_4305);
nor U9791 (N_9791,N_6171,N_6658);
xor U9792 (N_9792,N_4500,N_7716);
or U9793 (N_9793,N_6300,N_4718);
or U9794 (N_9794,N_7120,N_6677);
xnor U9795 (N_9795,N_5416,N_7827);
xnor U9796 (N_9796,N_7634,N_5903);
and U9797 (N_9797,N_6425,N_4854);
xnor U9798 (N_9798,N_7957,N_4537);
nor U9799 (N_9799,N_4283,N_5890);
nor U9800 (N_9800,N_7815,N_5671);
nand U9801 (N_9801,N_5586,N_6199);
and U9802 (N_9802,N_7149,N_5430);
nor U9803 (N_9803,N_5824,N_7253);
nor U9804 (N_9804,N_4901,N_4279);
and U9805 (N_9805,N_7773,N_5621);
and U9806 (N_9806,N_7038,N_6214);
nand U9807 (N_9807,N_5132,N_5518);
nor U9808 (N_9808,N_6480,N_4080);
nand U9809 (N_9809,N_7542,N_4058);
or U9810 (N_9810,N_7858,N_7265);
xor U9811 (N_9811,N_6327,N_6617);
nand U9812 (N_9812,N_5223,N_4787);
nor U9813 (N_9813,N_5741,N_5423);
xnor U9814 (N_9814,N_5904,N_4401);
xnor U9815 (N_9815,N_6912,N_7751);
nand U9816 (N_9816,N_7138,N_5962);
or U9817 (N_9817,N_7462,N_5063);
or U9818 (N_9818,N_4458,N_7088);
nand U9819 (N_9819,N_7307,N_4398);
and U9820 (N_9820,N_7834,N_7391);
and U9821 (N_9821,N_5035,N_7987);
and U9822 (N_9822,N_6926,N_5957);
xor U9823 (N_9823,N_4704,N_5895);
nor U9824 (N_9824,N_7148,N_4802);
or U9825 (N_9825,N_7619,N_7083);
or U9826 (N_9826,N_5992,N_6307);
nand U9827 (N_9827,N_7507,N_7015);
nor U9828 (N_9828,N_4217,N_7841);
or U9829 (N_9829,N_6466,N_7277);
nor U9830 (N_9830,N_6847,N_4032);
or U9831 (N_9831,N_5097,N_4427);
and U9832 (N_9832,N_7107,N_7055);
or U9833 (N_9833,N_4413,N_5726);
xor U9834 (N_9834,N_5765,N_4513);
nor U9835 (N_9835,N_4445,N_7517);
nand U9836 (N_9836,N_7896,N_5739);
nand U9837 (N_9837,N_7575,N_6975);
nand U9838 (N_9838,N_5729,N_4853);
and U9839 (N_9839,N_5774,N_4251);
nand U9840 (N_9840,N_4243,N_7594);
or U9841 (N_9841,N_4594,N_4066);
nand U9842 (N_9842,N_5576,N_7071);
nand U9843 (N_9843,N_4120,N_5424);
and U9844 (N_9844,N_5491,N_6039);
nor U9845 (N_9845,N_4245,N_4072);
and U9846 (N_9846,N_4230,N_6406);
and U9847 (N_9847,N_4070,N_6459);
xnor U9848 (N_9848,N_6163,N_7849);
nor U9849 (N_9849,N_5706,N_5909);
nor U9850 (N_9850,N_5320,N_6029);
or U9851 (N_9851,N_6605,N_6072);
nor U9852 (N_9852,N_5933,N_7380);
or U9853 (N_9853,N_5989,N_6892);
nand U9854 (N_9854,N_5351,N_5801);
xor U9855 (N_9855,N_7131,N_7587);
nor U9856 (N_9856,N_7725,N_5070);
nor U9857 (N_9857,N_7122,N_6609);
nand U9858 (N_9858,N_4338,N_7496);
nand U9859 (N_9859,N_5855,N_4886);
nand U9860 (N_9860,N_6982,N_4021);
or U9861 (N_9861,N_4681,N_4048);
or U9862 (N_9862,N_7246,N_7880);
and U9863 (N_9863,N_5469,N_4208);
nor U9864 (N_9864,N_6815,N_7468);
nand U9865 (N_9865,N_7861,N_6291);
and U9866 (N_9866,N_4808,N_6903);
nand U9867 (N_9867,N_5466,N_5792);
xor U9868 (N_9868,N_7352,N_7141);
nor U9869 (N_9869,N_6112,N_7164);
xor U9870 (N_9870,N_4440,N_5547);
nor U9871 (N_9871,N_7560,N_6211);
xor U9872 (N_9872,N_6391,N_4118);
or U9873 (N_9873,N_7346,N_6332);
nand U9874 (N_9874,N_6320,N_4491);
nor U9875 (N_9875,N_6774,N_6006);
xor U9876 (N_9876,N_6935,N_6502);
xnor U9877 (N_9877,N_6919,N_4337);
xnor U9878 (N_9878,N_5555,N_5594);
nor U9879 (N_9879,N_4592,N_6595);
nand U9880 (N_9880,N_6885,N_7528);
nor U9881 (N_9881,N_5201,N_6043);
nand U9882 (N_9882,N_4585,N_7938);
nor U9883 (N_9883,N_6554,N_4355);
or U9884 (N_9884,N_6144,N_6974);
or U9885 (N_9885,N_5959,N_7657);
or U9886 (N_9886,N_5540,N_7304);
nor U9887 (N_9887,N_5995,N_4313);
nor U9888 (N_9888,N_7064,N_4838);
nor U9889 (N_9889,N_6026,N_4450);
and U9890 (N_9890,N_7029,N_6449);
or U9891 (N_9891,N_5660,N_7483);
and U9892 (N_9892,N_6049,N_5613);
nand U9893 (N_9893,N_6558,N_5936);
nor U9894 (N_9894,N_6741,N_7780);
or U9895 (N_9895,N_5641,N_7711);
nand U9896 (N_9896,N_7400,N_5946);
nor U9897 (N_9897,N_6573,N_5183);
xor U9898 (N_9898,N_7871,N_5775);
nor U9899 (N_9899,N_4603,N_6743);
nand U9900 (N_9900,N_7155,N_5777);
and U9901 (N_9901,N_4668,N_7665);
xnor U9902 (N_9902,N_6884,N_4747);
xor U9903 (N_9903,N_5530,N_7674);
nor U9904 (N_9904,N_4342,N_5002);
nand U9905 (N_9905,N_6567,N_4285);
or U9906 (N_9906,N_5680,N_5665);
nor U9907 (N_9907,N_4128,N_4141);
and U9908 (N_9908,N_7865,N_6579);
xor U9909 (N_9909,N_6194,N_6746);
or U9910 (N_9910,N_5100,N_4514);
and U9911 (N_9911,N_7707,N_4062);
nor U9912 (N_9912,N_5264,N_5643);
xnor U9913 (N_9913,N_7831,N_4894);
and U9914 (N_9914,N_7629,N_4824);
or U9915 (N_9915,N_5485,N_4757);
and U9916 (N_9916,N_6689,N_5349);
nor U9917 (N_9917,N_5278,N_5165);
nor U9918 (N_9918,N_6035,N_5048);
or U9919 (N_9919,N_6698,N_6525);
nand U9920 (N_9920,N_7248,N_4692);
xnor U9921 (N_9921,N_5273,N_4071);
or U9922 (N_9922,N_6433,N_4186);
or U9923 (N_9923,N_5619,N_6539);
nor U9924 (N_9924,N_4822,N_7338);
nand U9925 (N_9925,N_4878,N_4529);
or U9926 (N_9926,N_6313,N_7586);
nor U9927 (N_9927,N_4556,N_6373);
nand U9928 (N_9928,N_4426,N_7356);
and U9929 (N_9929,N_6044,N_6100);
or U9930 (N_9930,N_7271,N_7597);
and U9931 (N_9931,N_5731,N_5474);
and U9932 (N_9932,N_7089,N_7506);
and U9933 (N_9933,N_7487,N_5578);
nand U9934 (N_9934,N_7442,N_7914);
nand U9935 (N_9935,N_6813,N_4569);
nor U9936 (N_9936,N_6213,N_5608);
and U9937 (N_9937,N_5874,N_6247);
nor U9938 (N_9938,N_7449,N_7800);
nor U9939 (N_9939,N_6839,N_7900);
nor U9940 (N_9940,N_5499,N_6104);
xor U9941 (N_9941,N_6099,N_4837);
nor U9942 (N_9942,N_5589,N_6014);
nand U9943 (N_9943,N_6337,N_7470);
xnor U9944 (N_9944,N_4496,N_6623);
nor U9945 (N_9945,N_7569,N_6367);
nor U9946 (N_9946,N_6264,N_6976);
nor U9947 (N_9947,N_6407,N_5218);
nor U9948 (N_9948,N_4347,N_6061);
and U9949 (N_9949,N_7426,N_5171);
or U9950 (N_9950,N_6917,N_5863);
and U9951 (N_9951,N_7389,N_5590);
xnor U9952 (N_9952,N_5124,N_4425);
nand U9953 (N_9953,N_5919,N_7429);
nand U9954 (N_9954,N_6720,N_5501);
and U9955 (N_9955,N_6838,N_5128);
and U9956 (N_9956,N_7826,N_4175);
and U9957 (N_9957,N_5527,N_6031);
or U9958 (N_9958,N_5238,N_4522);
or U9959 (N_9959,N_7492,N_4373);
or U9960 (N_9960,N_4244,N_7229);
or U9961 (N_9961,N_7421,N_5421);
nand U9962 (N_9962,N_6475,N_4252);
nor U9963 (N_9963,N_5740,N_4766);
or U9964 (N_9964,N_7752,N_6103);
xnor U9965 (N_9965,N_6161,N_7323);
nor U9966 (N_9966,N_5705,N_6807);
nand U9967 (N_9967,N_5615,N_6225);
and U9968 (N_9968,N_4584,N_5552);
or U9969 (N_9969,N_4640,N_4432);
or U9970 (N_9970,N_5872,N_4437);
nor U9971 (N_9971,N_4295,N_5876);
or U9972 (N_9972,N_5878,N_4944);
nor U9973 (N_9973,N_6201,N_5831);
or U9974 (N_9974,N_6537,N_4350);
nand U9975 (N_9975,N_5067,N_7503);
or U9976 (N_9976,N_6823,N_4460);
nor U9977 (N_9977,N_4276,N_5369);
or U9978 (N_9978,N_6046,N_6949);
nand U9979 (N_9979,N_4799,N_7465);
nand U9980 (N_9980,N_4873,N_6704);
nor U9981 (N_9981,N_4366,N_7194);
xnor U9982 (N_9982,N_4564,N_7099);
or U9983 (N_9983,N_4543,N_6166);
nand U9984 (N_9984,N_7303,N_5449);
xnor U9985 (N_9985,N_7526,N_4091);
nand U9986 (N_9986,N_4871,N_5304);
or U9987 (N_9987,N_7432,N_6675);
nor U9988 (N_9988,N_4680,N_7838);
nor U9989 (N_9989,N_6200,N_7978);
and U9990 (N_9990,N_5053,N_4358);
and U9991 (N_9991,N_5698,N_4965);
and U9992 (N_9992,N_6920,N_7816);
xnor U9993 (N_9993,N_7404,N_5762);
nand U9994 (N_9994,N_5182,N_4893);
nand U9995 (N_9995,N_7760,N_6399);
and U9996 (N_9996,N_6780,N_4441);
xor U9997 (N_9997,N_7595,N_7607);
nand U9998 (N_9998,N_7644,N_4917);
and U9999 (N_9999,N_5340,N_7222);
xnor U10000 (N_10000,N_6284,N_5157);
nand U10001 (N_10001,N_7215,N_5046);
nand U10002 (N_10002,N_5993,N_4010);
xor U10003 (N_10003,N_6086,N_5701);
nand U10004 (N_10004,N_5105,N_4077);
nand U10005 (N_10005,N_7858,N_5703);
nand U10006 (N_10006,N_6493,N_7961);
nor U10007 (N_10007,N_7854,N_6926);
nor U10008 (N_10008,N_4676,N_5317);
or U10009 (N_10009,N_6506,N_5867);
nor U10010 (N_10010,N_6563,N_6315);
and U10011 (N_10011,N_7088,N_4605);
nand U10012 (N_10012,N_6061,N_4242);
xnor U10013 (N_10013,N_4177,N_6610);
nand U10014 (N_10014,N_5124,N_6778);
nand U10015 (N_10015,N_5499,N_4721);
nand U10016 (N_10016,N_5081,N_7255);
or U10017 (N_10017,N_7179,N_6020);
and U10018 (N_10018,N_5463,N_5485);
nor U10019 (N_10019,N_4541,N_5439);
and U10020 (N_10020,N_6604,N_7704);
nor U10021 (N_10021,N_7809,N_6438);
nor U10022 (N_10022,N_7219,N_6626);
and U10023 (N_10023,N_7166,N_7186);
and U10024 (N_10024,N_4862,N_7012);
nand U10025 (N_10025,N_4815,N_7684);
and U10026 (N_10026,N_4390,N_4400);
nor U10027 (N_10027,N_7245,N_5207);
or U10028 (N_10028,N_7241,N_5794);
nand U10029 (N_10029,N_7191,N_4547);
or U10030 (N_10030,N_4697,N_6672);
xor U10031 (N_10031,N_4924,N_7619);
xnor U10032 (N_10032,N_7507,N_6544);
and U10033 (N_10033,N_6430,N_7025);
nor U10034 (N_10034,N_5678,N_4160);
xor U10035 (N_10035,N_4139,N_6586);
nor U10036 (N_10036,N_4246,N_7707);
xor U10037 (N_10037,N_4280,N_7494);
or U10038 (N_10038,N_7339,N_4126);
and U10039 (N_10039,N_5418,N_6658);
nor U10040 (N_10040,N_6953,N_4995);
nand U10041 (N_10041,N_6860,N_6562);
or U10042 (N_10042,N_4632,N_6458);
nand U10043 (N_10043,N_7584,N_5724);
nand U10044 (N_10044,N_6122,N_4412);
xor U10045 (N_10045,N_4450,N_4958);
and U10046 (N_10046,N_6207,N_7570);
nand U10047 (N_10047,N_4941,N_6848);
xor U10048 (N_10048,N_4242,N_7040);
and U10049 (N_10049,N_7131,N_4354);
xnor U10050 (N_10050,N_5203,N_6408);
or U10051 (N_10051,N_4583,N_6454);
and U10052 (N_10052,N_7918,N_7948);
or U10053 (N_10053,N_7390,N_5452);
nor U10054 (N_10054,N_6415,N_6894);
nand U10055 (N_10055,N_7729,N_5363);
nand U10056 (N_10056,N_4836,N_5903);
nor U10057 (N_10057,N_6983,N_6059);
nand U10058 (N_10058,N_6589,N_5499);
nand U10059 (N_10059,N_6056,N_4134);
nor U10060 (N_10060,N_7002,N_4643);
nor U10061 (N_10061,N_7638,N_5791);
and U10062 (N_10062,N_7177,N_7071);
nor U10063 (N_10063,N_4704,N_6902);
xnor U10064 (N_10064,N_5281,N_4207);
xor U10065 (N_10065,N_7484,N_4411);
and U10066 (N_10066,N_7799,N_7370);
nand U10067 (N_10067,N_6880,N_5551);
xnor U10068 (N_10068,N_7399,N_6184);
or U10069 (N_10069,N_4826,N_5105);
xor U10070 (N_10070,N_4318,N_7644);
xor U10071 (N_10071,N_7875,N_4181);
nor U10072 (N_10072,N_6698,N_6210);
and U10073 (N_10073,N_6594,N_4882);
nor U10074 (N_10074,N_4049,N_5218);
xor U10075 (N_10075,N_7787,N_4169);
nand U10076 (N_10076,N_7611,N_5349);
or U10077 (N_10077,N_6844,N_6839);
xor U10078 (N_10078,N_5846,N_7155);
xor U10079 (N_10079,N_5383,N_4641);
or U10080 (N_10080,N_4802,N_7755);
nand U10081 (N_10081,N_4177,N_5810);
or U10082 (N_10082,N_5098,N_6412);
or U10083 (N_10083,N_5853,N_4768);
or U10084 (N_10084,N_4391,N_7549);
nand U10085 (N_10085,N_7891,N_7668);
and U10086 (N_10086,N_5114,N_7284);
or U10087 (N_10087,N_4292,N_4433);
xnor U10088 (N_10088,N_4118,N_4966);
nor U10089 (N_10089,N_6855,N_4412);
xor U10090 (N_10090,N_4240,N_5460);
or U10091 (N_10091,N_7357,N_4062);
and U10092 (N_10092,N_6948,N_7524);
nor U10093 (N_10093,N_4384,N_7430);
or U10094 (N_10094,N_5144,N_7493);
nand U10095 (N_10095,N_4431,N_5061);
nand U10096 (N_10096,N_4259,N_5379);
nand U10097 (N_10097,N_6878,N_5383);
nor U10098 (N_10098,N_6740,N_5449);
and U10099 (N_10099,N_4457,N_6060);
nand U10100 (N_10100,N_7182,N_7610);
and U10101 (N_10101,N_7630,N_6594);
and U10102 (N_10102,N_4133,N_4438);
nor U10103 (N_10103,N_6196,N_7068);
nor U10104 (N_10104,N_6495,N_5142);
and U10105 (N_10105,N_5767,N_6432);
xnor U10106 (N_10106,N_7067,N_6643);
xnor U10107 (N_10107,N_7484,N_5476);
and U10108 (N_10108,N_4053,N_5816);
nor U10109 (N_10109,N_4898,N_7609);
nor U10110 (N_10110,N_6653,N_7153);
xor U10111 (N_10111,N_7403,N_6169);
xnor U10112 (N_10112,N_7678,N_6711);
xor U10113 (N_10113,N_5264,N_6181);
or U10114 (N_10114,N_4367,N_7168);
and U10115 (N_10115,N_7307,N_7336);
and U10116 (N_10116,N_6327,N_5767);
nand U10117 (N_10117,N_6239,N_6154);
or U10118 (N_10118,N_4678,N_4053);
nand U10119 (N_10119,N_6599,N_7399);
or U10120 (N_10120,N_4795,N_7500);
xnor U10121 (N_10121,N_4396,N_7107);
and U10122 (N_10122,N_6993,N_5597);
and U10123 (N_10123,N_7917,N_7354);
xor U10124 (N_10124,N_6241,N_4794);
or U10125 (N_10125,N_7176,N_7403);
xor U10126 (N_10126,N_4227,N_5457);
or U10127 (N_10127,N_5625,N_7853);
and U10128 (N_10128,N_5854,N_6439);
and U10129 (N_10129,N_5620,N_6812);
nand U10130 (N_10130,N_4243,N_4969);
nand U10131 (N_10131,N_4974,N_7348);
or U10132 (N_10132,N_5692,N_5056);
nor U10133 (N_10133,N_7211,N_4047);
and U10134 (N_10134,N_6153,N_6743);
and U10135 (N_10135,N_6039,N_6605);
nand U10136 (N_10136,N_7111,N_5595);
nor U10137 (N_10137,N_6668,N_7888);
xor U10138 (N_10138,N_5239,N_7405);
xnor U10139 (N_10139,N_7159,N_6104);
xnor U10140 (N_10140,N_7216,N_6318);
and U10141 (N_10141,N_7053,N_7131);
and U10142 (N_10142,N_4239,N_7549);
xnor U10143 (N_10143,N_7344,N_4252);
xnor U10144 (N_10144,N_7254,N_5691);
nand U10145 (N_10145,N_5998,N_5664);
nand U10146 (N_10146,N_4506,N_5349);
or U10147 (N_10147,N_5084,N_4858);
and U10148 (N_10148,N_4107,N_6534);
and U10149 (N_10149,N_5669,N_6929);
and U10150 (N_10150,N_7931,N_5324);
or U10151 (N_10151,N_4567,N_5736);
nor U10152 (N_10152,N_4940,N_5475);
nand U10153 (N_10153,N_4493,N_4051);
nor U10154 (N_10154,N_4065,N_5339);
nor U10155 (N_10155,N_6488,N_6073);
nor U10156 (N_10156,N_7629,N_6133);
nor U10157 (N_10157,N_4327,N_4433);
xor U10158 (N_10158,N_7555,N_7145);
xnor U10159 (N_10159,N_6832,N_4640);
or U10160 (N_10160,N_6523,N_7715);
and U10161 (N_10161,N_4289,N_6092);
or U10162 (N_10162,N_4912,N_4586);
and U10163 (N_10163,N_6264,N_7731);
or U10164 (N_10164,N_7264,N_5779);
nand U10165 (N_10165,N_4219,N_6903);
or U10166 (N_10166,N_5764,N_5519);
or U10167 (N_10167,N_5796,N_5210);
or U10168 (N_10168,N_7816,N_4620);
or U10169 (N_10169,N_6509,N_6204);
and U10170 (N_10170,N_6302,N_5630);
xor U10171 (N_10171,N_5737,N_5272);
xor U10172 (N_10172,N_7959,N_7866);
or U10173 (N_10173,N_4359,N_7613);
or U10174 (N_10174,N_7121,N_4535);
nand U10175 (N_10175,N_5038,N_4785);
xnor U10176 (N_10176,N_4498,N_6787);
xnor U10177 (N_10177,N_5349,N_6961);
nor U10178 (N_10178,N_4379,N_5532);
nor U10179 (N_10179,N_5215,N_7868);
and U10180 (N_10180,N_6233,N_4218);
nand U10181 (N_10181,N_7647,N_6348);
or U10182 (N_10182,N_7862,N_5106);
and U10183 (N_10183,N_6929,N_4370);
and U10184 (N_10184,N_7117,N_5632);
and U10185 (N_10185,N_7113,N_7334);
and U10186 (N_10186,N_5557,N_4738);
xnor U10187 (N_10187,N_7439,N_4378);
and U10188 (N_10188,N_6721,N_7333);
and U10189 (N_10189,N_4606,N_6996);
nand U10190 (N_10190,N_6111,N_7989);
or U10191 (N_10191,N_5030,N_5341);
or U10192 (N_10192,N_5970,N_4502);
or U10193 (N_10193,N_7391,N_5711);
and U10194 (N_10194,N_4436,N_7846);
nand U10195 (N_10195,N_5072,N_4164);
or U10196 (N_10196,N_5133,N_6194);
or U10197 (N_10197,N_6970,N_5903);
nor U10198 (N_10198,N_7461,N_5905);
nor U10199 (N_10199,N_4406,N_6822);
or U10200 (N_10200,N_4787,N_4205);
xor U10201 (N_10201,N_7918,N_6292);
and U10202 (N_10202,N_7496,N_5178);
xor U10203 (N_10203,N_6873,N_6383);
or U10204 (N_10204,N_6938,N_6048);
xnor U10205 (N_10205,N_6096,N_4893);
and U10206 (N_10206,N_6961,N_7674);
or U10207 (N_10207,N_5580,N_4057);
xnor U10208 (N_10208,N_7132,N_5810);
nand U10209 (N_10209,N_4653,N_4170);
xor U10210 (N_10210,N_4652,N_5344);
nor U10211 (N_10211,N_6038,N_4056);
and U10212 (N_10212,N_7856,N_4097);
and U10213 (N_10213,N_7207,N_4579);
and U10214 (N_10214,N_7662,N_4718);
nor U10215 (N_10215,N_6123,N_5494);
nand U10216 (N_10216,N_5945,N_4367);
nor U10217 (N_10217,N_5338,N_4650);
or U10218 (N_10218,N_7319,N_7976);
and U10219 (N_10219,N_5027,N_7593);
or U10220 (N_10220,N_5445,N_7611);
nand U10221 (N_10221,N_6728,N_6009);
nor U10222 (N_10222,N_6425,N_6652);
xnor U10223 (N_10223,N_4518,N_7738);
nand U10224 (N_10224,N_5669,N_5872);
xnor U10225 (N_10225,N_5321,N_5939);
nand U10226 (N_10226,N_5239,N_4381);
and U10227 (N_10227,N_7958,N_7445);
nor U10228 (N_10228,N_7661,N_5929);
or U10229 (N_10229,N_5728,N_5344);
or U10230 (N_10230,N_5352,N_4275);
and U10231 (N_10231,N_6613,N_7020);
and U10232 (N_10232,N_7813,N_6165);
xor U10233 (N_10233,N_5650,N_7738);
xor U10234 (N_10234,N_5787,N_5045);
nand U10235 (N_10235,N_4440,N_6861);
and U10236 (N_10236,N_7021,N_5127);
or U10237 (N_10237,N_5058,N_5915);
and U10238 (N_10238,N_6354,N_6361);
nor U10239 (N_10239,N_7922,N_5686);
or U10240 (N_10240,N_7201,N_5269);
nor U10241 (N_10241,N_6692,N_5651);
xor U10242 (N_10242,N_7524,N_5851);
nor U10243 (N_10243,N_7287,N_5799);
xor U10244 (N_10244,N_6683,N_7016);
and U10245 (N_10245,N_7196,N_4784);
or U10246 (N_10246,N_6756,N_5960);
or U10247 (N_10247,N_6487,N_6495);
xor U10248 (N_10248,N_4896,N_7461);
xnor U10249 (N_10249,N_4343,N_6277);
nor U10250 (N_10250,N_6450,N_7558);
nor U10251 (N_10251,N_5222,N_6272);
xor U10252 (N_10252,N_6106,N_7923);
nor U10253 (N_10253,N_4229,N_7664);
or U10254 (N_10254,N_5787,N_6623);
nor U10255 (N_10255,N_7743,N_5894);
nand U10256 (N_10256,N_5354,N_7706);
nor U10257 (N_10257,N_5585,N_6341);
nand U10258 (N_10258,N_4741,N_5714);
xor U10259 (N_10259,N_7568,N_5580);
or U10260 (N_10260,N_6955,N_7191);
and U10261 (N_10261,N_5568,N_7950);
and U10262 (N_10262,N_5446,N_6100);
xor U10263 (N_10263,N_7827,N_5248);
or U10264 (N_10264,N_6315,N_6736);
nor U10265 (N_10265,N_7409,N_6994);
nand U10266 (N_10266,N_4167,N_4844);
or U10267 (N_10267,N_6239,N_4641);
nand U10268 (N_10268,N_5572,N_7097);
nand U10269 (N_10269,N_7908,N_6524);
nand U10270 (N_10270,N_6492,N_6914);
and U10271 (N_10271,N_6872,N_7343);
nand U10272 (N_10272,N_4366,N_6036);
and U10273 (N_10273,N_7419,N_6205);
nor U10274 (N_10274,N_7499,N_5468);
xnor U10275 (N_10275,N_4741,N_5900);
nor U10276 (N_10276,N_6904,N_7907);
nand U10277 (N_10277,N_6418,N_7938);
and U10278 (N_10278,N_6691,N_6626);
nor U10279 (N_10279,N_6633,N_6734);
xor U10280 (N_10280,N_5818,N_7774);
and U10281 (N_10281,N_6452,N_7271);
and U10282 (N_10282,N_6591,N_7338);
or U10283 (N_10283,N_5563,N_7708);
xor U10284 (N_10284,N_7282,N_6128);
or U10285 (N_10285,N_6724,N_7252);
or U10286 (N_10286,N_7151,N_6495);
and U10287 (N_10287,N_4474,N_7283);
xor U10288 (N_10288,N_4386,N_5221);
xnor U10289 (N_10289,N_7515,N_6231);
xor U10290 (N_10290,N_5635,N_7466);
nand U10291 (N_10291,N_6763,N_6091);
and U10292 (N_10292,N_4852,N_6866);
nor U10293 (N_10293,N_7491,N_5880);
or U10294 (N_10294,N_7445,N_4270);
xor U10295 (N_10295,N_7010,N_6979);
nor U10296 (N_10296,N_6723,N_4612);
nand U10297 (N_10297,N_5287,N_7964);
nand U10298 (N_10298,N_6800,N_5449);
or U10299 (N_10299,N_5862,N_7815);
nor U10300 (N_10300,N_4140,N_5649);
and U10301 (N_10301,N_6480,N_7894);
and U10302 (N_10302,N_7642,N_5945);
or U10303 (N_10303,N_7287,N_5907);
nand U10304 (N_10304,N_5678,N_6995);
nand U10305 (N_10305,N_4207,N_4765);
xnor U10306 (N_10306,N_7337,N_5829);
or U10307 (N_10307,N_5890,N_6214);
nor U10308 (N_10308,N_7147,N_5335);
or U10309 (N_10309,N_4643,N_7470);
nand U10310 (N_10310,N_7328,N_7802);
xor U10311 (N_10311,N_7406,N_5705);
or U10312 (N_10312,N_5982,N_6629);
and U10313 (N_10313,N_7559,N_7837);
and U10314 (N_10314,N_4571,N_4168);
and U10315 (N_10315,N_7791,N_4158);
or U10316 (N_10316,N_4465,N_7360);
nor U10317 (N_10317,N_7076,N_6738);
xnor U10318 (N_10318,N_7977,N_6245);
nor U10319 (N_10319,N_6653,N_4425);
nand U10320 (N_10320,N_6922,N_7970);
and U10321 (N_10321,N_7536,N_6110);
or U10322 (N_10322,N_6063,N_6252);
xnor U10323 (N_10323,N_6808,N_6477);
xnor U10324 (N_10324,N_5456,N_6310);
nor U10325 (N_10325,N_6112,N_4774);
nor U10326 (N_10326,N_5107,N_5290);
or U10327 (N_10327,N_4157,N_5587);
nor U10328 (N_10328,N_4384,N_5162);
nand U10329 (N_10329,N_5809,N_6611);
and U10330 (N_10330,N_5923,N_5737);
xor U10331 (N_10331,N_5514,N_7749);
nor U10332 (N_10332,N_6998,N_7694);
and U10333 (N_10333,N_6317,N_7020);
nor U10334 (N_10334,N_6861,N_5997);
nand U10335 (N_10335,N_7113,N_6876);
nand U10336 (N_10336,N_7022,N_4731);
or U10337 (N_10337,N_5677,N_5487);
xnor U10338 (N_10338,N_7770,N_6599);
and U10339 (N_10339,N_7153,N_5020);
or U10340 (N_10340,N_5902,N_7043);
nand U10341 (N_10341,N_4363,N_4566);
xnor U10342 (N_10342,N_5672,N_4578);
nand U10343 (N_10343,N_4217,N_5705);
or U10344 (N_10344,N_4967,N_5152);
or U10345 (N_10345,N_5408,N_4310);
xor U10346 (N_10346,N_7551,N_5378);
xor U10347 (N_10347,N_7119,N_6596);
nor U10348 (N_10348,N_7831,N_6768);
or U10349 (N_10349,N_4512,N_6476);
or U10350 (N_10350,N_5485,N_4121);
or U10351 (N_10351,N_4211,N_6937);
xor U10352 (N_10352,N_6195,N_5586);
xor U10353 (N_10353,N_6305,N_5612);
nor U10354 (N_10354,N_4262,N_7702);
and U10355 (N_10355,N_4325,N_4367);
and U10356 (N_10356,N_6438,N_4485);
nor U10357 (N_10357,N_6145,N_5545);
nand U10358 (N_10358,N_7669,N_7772);
or U10359 (N_10359,N_6390,N_6363);
or U10360 (N_10360,N_6235,N_4016);
nor U10361 (N_10361,N_6267,N_4233);
or U10362 (N_10362,N_4792,N_4760);
xor U10363 (N_10363,N_4214,N_6902);
or U10364 (N_10364,N_4756,N_6326);
and U10365 (N_10365,N_7776,N_4863);
and U10366 (N_10366,N_7809,N_4817);
or U10367 (N_10367,N_5897,N_7483);
nor U10368 (N_10368,N_4250,N_5807);
xnor U10369 (N_10369,N_4445,N_4192);
nand U10370 (N_10370,N_7678,N_6816);
and U10371 (N_10371,N_6495,N_4888);
nor U10372 (N_10372,N_5507,N_6371);
and U10373 (N_10373,N_6786,N_4754);
and U10374 (N_10374,N_5102,N_4088);
or U10375 (N_10375,N_7161,N_7789);
xor U10376 (N_10376,N_5272,N_6804);
xnor U10377 (N_10377,N_5166,N_5824);
nand U10378 (N_10378,N_7508,N_5354);
xnor U10379 (N_10379,N_4119,N_6566);
or U10380 (N_10380,N_7195,N_4743);
nor U10381 (N_10381,N_6147,N_4714);
nor U10382 (N_10382,N_5330,N_6539);
or U10383 (N_10383,N_6035,N_6998);
nand U10384 (N_10384,N_7349,N_6958);
nand U10385 (N_10385,N_6876,N_6197);
xnor U10386 (N_10386,N_6620,N_6424);
or U10387 (N_10387,N_6163,N_5231);
or U10388 (N_10388,N_6677,N_7479);
xor U10389 (N_10389,N_4288,N_7417);
and U10390 (N_10390,N_4480,N_4963);
and U10391 (N_10391,N_6963,N_4702);
nor U10392 (N_10392,N_6286,N_4301);
nor U10393 (N_10393,N_6518,N_6192);
and U10394 (N_10394,N_4494,N_7560);
or U10395 (N_10395,N_7435,N_5312);
nor U10396 (N_10396,N_5306,N_7041);
or U10397 (N_10397,N_4473,N_5203);
and U10398 (N_10398,N_7417,N_4534);
and U10399 (N_10399,N_6529,N_5514);
nand U10400 (N_10400,N_4271,N_4958);
xor U10401 (N_10401,N_7208,N_7673);
or U10402 (N_10402,N_4498,N_5186);
nand U10403 (N_10403,N_7740,N_6502);
and U10404 (N_10404,N_6322,N_5770);
and U10405 (N_10405,N_4530,N_5867);
nor U10406 (N_10406,N_7558,N_6588);
xnor U10407 (N_10407,N_6845,N_6558);
nand U10408 (N_10408,N_6323,N_6470);
xor U10409 (N_10409,N_5446,N_7379);
nand U10410 (N_10410,N_5125,N_7398);
xor U10411 (N_10411,N_6239,N_6295);
and U10412 (N_10412,N_6720,N_7942);
nand U10413 (N_10413,N_5033,N_6652);
nand U10414 (N_10414,N_4546,N_5486);
xnor U10415 (N_10415,N_5361,N_7468);
nand U10416 (N_10416,N_5451,N_5613);
and U10417 (N_10417,N_7673,N_4371);
and U10418 (N_10418,N_7077,N_7465);
nor U10419 (N_10419,N_4244,N_6090);
nand U10420 (N_10420,N_5053,N_6673);
xor U10421 (N_10421,N_6290,N_5459);
and U10422 (N_10422,N_4255,N_5031);
xor U10423 (N_10423,N_7562,N_7497);
or U10424 (N_10424,N_5514,N_5011);
or U10425 (N_10425,N_6910,N_7213);
nor U10426 (N_10426,N_4751,N_4297);
xor U10427 (N_10427,N_4228,N_5459);
nand U10428 (N_10428,N_7324,N_4719);
nand U10429 (N_10429,N_4235,N_7954);
and U10430 (N_10430,N_4392,N_4672);
xor U10431 (N_10431,N_4515,N_4058);
xor U10432 (N_10432,N_7815,N_4648);
and U10433 (N_10433,N_7228,N_6980);
xnor U10434 (N_10434,N_7381,N_4020);
or U10435 (N_10435,N_7789,N_4429);
and U10436 (N_10436,N_4879,N_4972);
or U10437 (N_10437,N_4536,N_6470);
or U10438 (N_10438,N_5979,N_7405);
xor U10439 (N_10439,N_4349,N_4337);
or U10440 (N_10440,N_4685,N_7029);
xnor U10441 (N_10441,N_5586,N_7679);
or U10442 (N_10442,N_5351,N_4027);
nor U10443 (N_10443,N_4451,N_4538);
nor U10444 (N_10444,N_4205,N_7039);
and U10445 (N_10445,N_4446,N_7467);
and U10446 (N_10446,N_6036,N_6020);
or U10447 (N_10447,N_4265,N_4884);
nor U10448 (N_10448,N_6835,N_6778);
nand U10449 (N_10449,N_6581,N_4983);
nand U10450 (N_10450,N_6080,N_4378);
xnor U10451 (N_10451,N_4928,N_7570);
xnor U10452 (N_10452,N_4897,N_5932);
and U10453 (N_10453,N_6642,N_5543);
xnor U10454 (N_10454,N_7226,N_5137);
nor U10455 (N_10455,N_4257,N_7064);
nor U10456 (N_10456,N_4195,N_5277);
nor U10457 (N_10457,N_4252,N_5289);
nand U10458 (N_10458,N_7676,N_5670);
nand U10459 (N_10459,N_4073,N_5519);
and U10460 (N_10460,N_7363,N_5879);
or U10461 (N_10461,N_5666,N_5066);
xnor U10462 (N_10462,N_4717,N_5299);
nor U10463 (N_10463,N_5569,N_7722);
and U10464 (N_10464,N_4758,N_5778);
or U10465 (N_10465,N_7203,N_4089);
nand U10466 (N_10466,N_5634,N_7059);
and U10467 (N_10467,N_5273,N_7063);
nor U10468 (N_10468,N_4241,N_4182);
or U10469 (N_10469,N_6676,N_4052);
nand U10470 (N_10470,N_7471,N_6647);
and U10471 (N_10471,N_6503,N_6423);
nand U10472 (N_10472,N_5815,N_4554);
or U10473 (N_10473,N_4903,N_6100);
and U10474 (N_10474,N_6147,N_7167);
nand U10475 (N_10475,N_5560,N_7959);
nand U10476 (N_10476,N_4486,N_4981);
or U10477 (N_10477,N_7179,N_6548);
nor U10478 (N_10478,N_6199,N_7822);
and U10479 (N_10479,N_4766,N_7388);
nor U10480 (N_10480,N_5648,N_4928);
and U10481 (N_10481,N_6295,N_5235);
nor U10482 (N_10482,N_4919,N_5943);
xor U10483 (N_10483,N_4167,N_5513);
or U10484 (N_10484,N_5724,N_6678);
xnor U10485 (N_10485,N_6549,N_6613);
or U10486 (N_10486,N_6728,N_5669);
or U10487 (N_10487,N_5080,N_6539);
or U10488 (N_10488,N_6621,N_5405);
or U10489 (N_10489,N_4879,N_4878);
or U10490 (N_10490,N_6716,N_6970);
or U10491 (N_10491,N_4658,N_6119);
or U10492 (N_10492,N_4377,N_5755);
and U10493 (N_10493,N_6339,N_4428);
xnor U10494 (N_10494,N_6812,N_5279);
xor U10495 (N_10495,N_5247,N_4405);
xor U10496 (N_10496,N_5831,N_6204);
nand U10497 (N_10497,N_7764,N_5611);
nor U10498 (N_10498,N_5075,N_6475);
xnor U10499 (N_10499,N_7114,N_5944);
nor U10500 (N_10500,N_6494,N_4453);
and U10501 (N_10501,N_7935,N_7934);
and U10502 (N_10502,N_7750,N_5672);
or U10503 (N_10503,N_6084,N_5811);
xnor U10504 (N_10504,N_6285,N_4108);
or U10505 (N_10505,N_7561,N_4246);
or U10506 (N_10506,N_6851,N_6010);
and U10507 (N_10507,N_4531,N_6595);
nand U10508 (N_10508,N_4731,N_5762);
and U10509 (N_10509,N_4159,N_6775);
nor U10510 (N_10510,N_5152,N_4784);
xnor U10511 (N_10511,N_4378,N_7055);
and U10512 (N_10512,N_4040,N_5093);
or U10513 (N_10513,N_4652,N_6820);
nand U10514 (N_10514,N_5272,N_5424);
nand U10515 (N_10515,N_6617,N_7905);
xor U10516 (N_10516,N_7651,N_4838);
nand U10517 (N_10517,N_4688,N_7516);
xnor U10518 (N_10518,N_4449,N_6895);
xnor U10519 (N_10519,N_4277,N_5608);
nand U10520 (N_10520,N_4260,N_6980);
and U10521 (N_10521,N_7725,N_4893);
nor U10522 (N_10522,N_4493,N_7097);
nor U10523 (N_10523,N_4058,N_5489);
or U10524 (N_10524,N_4430,N_7010);
xnor U10525 (N_10525,N_7624,N_5601);
and U10526 (N_10526,N_5259,N_6251);
or U10527 (N_10527,N_6396,N_5164);
nand U10528 (N_10528,N_6484,N_7173);
or U10529 (N_10529,N_7570,N_5631);
xnor U10530 (N_10530,N_5348,N_5880);
and U10531 (N_10531,N_4104,N_7553);
xnor U10532 (N_10532,N_5653,N_6430);
nand U10533 (N_10533,N_5086,N_6739);
nand U10534 (N_10534,N_4937,N_7413);
or U10535 (N_10535,N_7795,N_6695);
or U10536 (N_10536,N_4246,N_5819);
or U10537 (N_10537,N_7802,N_6964);
nand U10538 (N_10538,N_6972,N_4699);
or U10539 (N_10539,N_5866,N_4312);
or U10540 (N_10540,N_6007,N_5704);
nand U10541 (N_10541,N_5404,N_7346);
or U10542 (N_10542,N_5115,N_7980);
xnor U10543 (N_10543,N_7545,N_7684);
nand U10544 (N_10544,N_6673,N_5561);
xnor U10545 (N_10545,N_7171,N_7591);
xnor U10546 (N_10546,N_7057,N_7243);
nor U10547 (N_10547,N_6573,N_4414);
nor U10548 (N_10548,N_5389,N_6778);
or U10549 (N_10549,N_4246,N_4711);
and U10550 (N_10550,N_5915,N_6332);
xnor U10551 (N_10551,N_7442,N_7714);
nor U10552 (N_10552,N_5013,N_6617);
and U10553 (N_10553,N_4359,N_4846);
and U10554 (N_10554,N_5983,N_6300);
xnor U10555 (N_10555,N_5916,N_4646);
xnor U10556 (N_10556,N_5997,N_5065);
nor U10557 (N_10557,N_6545,N_7013);
nor U10558 (N_10558,N_4995,N_6739);
nand U10559 (N_10559,N_5668,N_4078);
xor U10560 (N_10560,N_4055,N_6350);
or U10561 (N_10561,N_7202,N_4099);
nand U10562 (N_10562,N_7433,N_6560);
or U10563 (N_10563,N_7178,N_4074);
and U10564 (N_10564,N_7379,N_4630);
nor U10565 (N_10565,N_5964,N_4748);
nand U10566 (N_10566,N_5681,N_4217);
xnor U10567 (N_10567,N_5612,N_7383);
or U10568 (N_10568,N_7669,N_6931);
nor U10569 (N_10569,N_5635,N_6901);
nor U10570 (N_10570,N_6005,N_7229);
nand U10571 (N_10571,N_6604,N_4752);
nor U10572 (N_10572,N_7732,N_6766);
nor U10573 (N_10573,N_6948,N_7098);
and U10574 (N_10574,N_4945,N_4508);
or U10575 (N_10575,N_6229,N_7025);
and U10576 (N_10576,N_4415,N_5125);
nand U10577 (N_10577,N_4108,N_5903);
nor U10578 (N_10578,N_6535,N_5924);
and U10579 (N_10579,N_7330,N_5200);
nand U10580 (N_10580,N_7014,N_5168);
xnor U10581 (N_10581,N_6740,N_6754);
nand U10582 (N_10582,N_6067,N_5960);
nand U10583 (N_10583,N_4642,N_7138);
nand U10584 (N_10584,N_7011,N_7575);
nand U10585 (N_10585,N_4702,N_6489);
nand U10586 (N_10586,N_7842,N_6359);
nor U10587 (N_10587,N_6776,N_4714);
xnor U10588 (N_10588,N_7990,N_7699);
or U10589 (N_10589,N_7801,N_7380);
nand U10590 (N_10590,N_7381,N_4874);
xor U10591 (N_10591,N_6159,N_6250);
xnor U10592 (N_10592,N_7509,N_7004);
nand U10593 (N_10593,N_4329,N_6476);
xor U10594 (N_10594,N_6287,N_5579);
nand U10595 (N_10595,N_6402,N_4277);
xnor U10596 (N_10596,N_6951,N_4457);
and U10597 (N_10597,N_4556,N_4836);
nor U10598 (N_10598,N_4299,N_5937);
and U10599 (N_10599,N_6066,N_6211);
and U10600 (N_10600,N_4209,N_5479);
and U10601 (N_10601,N_4072,N_4251);
xnor U10602 (N_10602,N_5014,N_7216);
xnor U10603 (N_10603,N_4275,N_5908);
and U10604 (N_10604,N_7900,N_7383);
nand U10605 (N_10605,N_6006,N_7546);
nand U10606 (N_10606,N_5983,N_5634);
and U10607 (N_10607,N_7442,N_6528);
xor U10608 (N_10608,N_7653,N_6549);
xor U10609 (N_10609,N_7822,N_5181);
xor U10610 (N_10610,N_6781,N_4726);
nand U10611 (N_10611,N_6678,N_7112);
or U10612 (N_10612,N_5306,N_6005);
xor U10613 (N_10613,N_6887,N_6210);
xor U10614 (N_10614,N_6968,N_5175);
nor U10615 (N_10615,N_7246,N_7182);
nor U10616 (N_10616,N_6789,N_5545);
and U10617 (N_10617,N_7188,N_6324);
and U10618 (N_10618,N_7260,N_5886);
xnor U10619 (N_10619,N_6408,N_7826);
nor U10620 (N_10620,N_5651,N_4464);
nor U10621 (N_10621,N_4611,N_7063);
or U10622 (N_10622,N_6027,N_7830);
or U10623 (N_10623,N_7117,N_5277);
nand U10624 (N_10624,N_6702,N_5687);
nor U10625 (N_10625,N_5781,N_6398);
xnor U10626 (N_10626,N_4042,N_5079);
nand U10627 (N_10627,N_6666,N_6689);
and U10628 (N_10628,N_5141,N_4764);
xor U10629 (N_10629,N_7156,N_4552);
and U10630 (N_10630,N_7913,N_7801);
nor U10631 (N_10631,N_4170,N_6812);
and U10632 (N_10632,N_6434,N_6484);
nand U10633 (N_10633,N_4524,N_7127);
and U10634 (N_10634,N_4841,N_5756);
or U10635 (N_10635,N_4138,N_7130);
nor U10636 (N_10636,N_7202,N_5698);
xor U10637 (N_10637,N_6773,N_7927);
nand U10638 (N_10638,N_4818,N_6995);
and U10639 (N_10639,N_5572,N_5746);
nor U10640 (N_10640,N_6760,N_5784);
or U10641 (N_10641,N_6646,N_6704);
nand U10642 (N_10642,N_4872,N_7392);
xnor U10643 (N_10643,N_4492,N_5227);
or U10644 (N_10644,N_5800,N_5580);
nand U10645 (N_10645,N_5508,N_4122);
and U10646 (N_10646,N_7146,N_7617);
xor U10647 (N_10647,N_5343,N_6815);
and U10648 (N_10648,N_5930,N_6275);
xnor U10649 (N_10649,N_7338,N_6368);
or U10650 (N_10650,N_4605,N_4422);
or U10651 (N_10651,N_4140,N_6417);
xor U10652 (N_10652,N_7594,N_6174);
and U10653 (N_10653,N_7044,N_6970);
or U10654 (N_10654,N_6300,N_5124);
xor U10655 (N_10655,N_5325,N_5011);
xor U10656 (N_10656,N_5686,N_7828);
or U10657 (N_10657,N_7502,N_5987);
nor U10658 (N_10658,N_5925,N_7803);
nor U10659 (N_10659,N_7248,N_5658);
or U10660 (N_10660,N_4550,N_6483);
xor U10661 (N_10661,N_5270,N_7611);
and U10662 (N_10662,N_5619,N_5676);
xnor U10663 (N_10663,N_5252,N_6047);
or U10664 (N_10664,N_4369,N_7020);
and U10665 (N_10665,N_4471,N_4662);
nor U10666 (N_10666,N_4266,N_7084);
or U10667 (N_10667,N_6371,N_4588);
and U10668 (N_10668,N_6987,N_4273);
nand U10669 (N_10669,N_5173,N_4861);
nand U10670 (N_10670,N_5192,N_6726);
xnor U10671 (N_10671,N_5202,N_7953);
nor U10672 (N_10672,N_7481,N_4133);
xnor U10673 (N_10673,N_5612,N_7781);
nand U10674 (N_10674,N_7144,N_6049);
and U10675 (N_10675,N_5404,N_7541);
xor U10676 (N_10676,N_4193,N_7585);
xor U10677 (N_10677,N_4766,N_6281);
nand U10678 (N_10678,N_5436,N_5674);
nor U10679 (N_10679,N_7108,N_4729);
xor U10680 (N_10680,N_7688,N_4573);
xnor U10681 (N_10681,N_5401,N_7530);
xnor U10682 (N_10682,N_4711,N_4771);
or U10683 (N_10683,N_7566,N_6908);
nor U10684 (N_10684,N_5843,N_7682);
or U10685 (N_10685,N_7352,N_5432);
and U10686 (N_10686,N_4444,N_4228);
and U10687 (N_10687,N_5750,N_4656);
and U10688 (N_10688,N_5071,N_6012);
or U10689 (N_10689,N_7286,N_4988);
nand U10690 (N_10690,N_7521,N_6993);
xor U10691 (N_10691,N_5013,N_7604);
xor U10692 (N_10692,N_4777,N_5726);
or U10693 (N_10693,N_7192,N_4221);
nand U10694 (N_10694,N_4155,N_6634);
nand U10695 (N_10695,N_6095,N_5169);
nand U10696 (N_10696,N_7449,N_6921);
or U10697 (N_10697,N_7350,N_7875);
or U10698 (N_10698,N_4074,N_4226);
xnor U10699 (N_10699,N_7421,N_6753);
and U10700 (N_10700,N_5629,N_4306);
xor U10701 (N_10701,N_7439,N_4054);
nor U10702 (N_10702,N_5694,N_4420);
nor U10703 (N_10703,N_4089,N_4311);
or U10704 (N_10704,N_5162,N_6152);
xnor U10705 (N_10705,N_5504,N_5063);
or U10706 (N_10706,N_5578,N_5913);
and U10707 (N_10707,N_5524,N_5456);
or U10708 (N_10708,N_5887,N_7723);
nor U10709 (N_10709,N_4460,N_6881);
or U10710 (N_10710,N_4328,N_6863);
and U10711 (N_10711,N_4058,N_5204);
nand U10712 (N_10712,N_5345,N_4236);
nand U10713 (N_10713,N_6634,N_5160);
nor U10714 (N_10714,N_5798,N_5742);
or U10715 (N_10715,N_6291,N_6317);
or U10716 (N_10716,N_4303,N_5922);
nand U10717 (N_10717,N_7330,N_6538);
and U10718 (N_10718,N_5619,N_7493);
or U10719 (N_10719,N_7505,N_4402);
nand U10720 (N_10720,N_5683,N_6700);
nand U10721 (N_10721,N_4816,N_5459);
nor U10722 (N_10722,N_5448,N_7148);
nand U10723 (N_10723,N_5305,N_5337);
or U10724 (N_10724,N_6151,N_7656);
nor U10725 (N_10725,N_6163,N_4273);
and U10726 (N_10726,N_5358,N_6503);
nor U10727 (N_10727,N_7770,N_7954);
nand U10728 (N_10728,N_5579,N_6450);
nor U10729 (N_10729,N_5187,N_4801);
or U10730 (N_10730,N_4716,N_7515);
nor U10731 (N_10731,N_4480,N_6562);
xor U10732 (N_10732,N_4135,N_5474);
nor U10733 (N_10733,N_5029,N_6112);
and U10734 (N_10734,N_5593,N_6323);
or U10735 (N_10735,N_4328,N_5977);
nor U10736 (N_10736,N_4472,N_7588);
xnor U10737 (N_10737,N_5506,N_4517);
and U10738 (N_10738,N_4961,N_7662);
or U10739 (N_10739,N_7529,N_4133);
or U10740 (N_10740,N_6626,N_5625);
nand U10741 (N_10741,N_6624,N_6778);
nand U10742 (N_10742,N_4831,N_4057);
or U10743 (N_10743,N_6909,N_5102);
xor U10744 (N_10744,N_5654,N_7390);
xor U10745 (N_10745,N_7784,N_5732);
xor U10746 (N_10746,N_6624,N_6072);
nand U10747 (N_10747,N_5918,N_7714);
nor U10748 (N_10748,N_5207,N_5317);
or U10749 (N_10749,N_7519,N_4266);
xor U10750 (N_10750,N_7917,N_4280);
nor U10751 (N_10751,N_6210,N_5367);
xor U10752 (N_10752,N_5191,N_7412);
nor U10753 (N_10753,N_7942,N_4210);
xor U10754 (N_10754,N_6067,N_5700);
xor U10755 (N_10755,N_6729,N_6980);
nor U10756 (N_10756,N_5905,N_5295);
or U10757 (N_10757,N_6585,N_5703);
nor U10758 (N_10758,N_4042,N_6443);
or U10759 (N_10759,N_7869,N_4189);
xnor U10760 (N_10760,N_7179,N_6126);
nand U10761 (N_10761,N_7399,N_6622);
nand U10762 (N_10762,N_4125,N_7368);
xor U10763 (N_10763,N_7099,N_7727);
nand U10764 (N_10764,N_5183,N_5792);
xnor U10765 (N_10765,N_4348,N_7271);
xor U10766 (N_10766,N_7467,N_5015);
nand U10767 (N_10767,N_7710,N_7205);
and U10768 (N_10768,N_6532,N_5274);
and U10769 (N_10769,N_5732,N_5187);
xor U10770 (N_10770,N_5358,N_4989);
nor U10771 (N_10771,N_6156,N_5373);
nand U10772 (N_10772,N_6823,N_4826);
nor U10773 (N_10773,N_4127,N_4373);
or U10774 (N_10774,N_7497,N_4473);
or U10775 (N_10775,N_5503,N_6125);
and U10776 (N_10776,N_6191,N_4706);
nor U10777 (N_10777,N_6696,N_7871);
and U10778 (N_10778,N_4087,N_7011);
xnor U10779 (N_10779,N_6135,N_6756);
or U10780 (N_10780,N_7564,N_5053);
nand U10781 (N_10781,N_7905,N_4882);
nand U10782 (N_10782,N_6820,N_5001);
and U10783 (N_10783,N_6069,N_5600);
and U10784 (N_10784,N_6548,N_7759);
nor U10785 (N_10785,N_5849,N_5768);
or U10786 (N_10786,N_4767,N_7384);
xnor U10787 (N_10787,N_6116,N_5100);
xnor U10788 (N_10788,N_5604,N_7078);
or U10789 (N_10789,N_5406,N_4634);
xnor U10790 (N_10790,N_7910,N_4725);
nor U10791 (N_10791,N_4041,N_6611);
or U10792 (N_10792,N_4489,N_6702);
nor U10793 (N_10793,N_4623,N_5382);
or U10794 (N_10794,N_7214,N_5916);
nand U10795 (N_10795,N_7555,N_7962);
and U10796 (N_10796,N_4506,N_5613);
xor U10797 (N_10797,N_5496,N_4730);
or U10798 (N_10798,N_6480,N_6883);
xor U10799 (N_10799,N_4710,N_6994);
and U10800 (N_10800,N_7087,N_6774);
or U10801 (N_10801,N_7653,N_5867);
xor U10802 (N_10802,N_5925,N_7716);
nor U10803 (N_10803,N_4887,N_4077);
nand U10804 (N_10804,N_5834,N_5155);
and U10805 (N_10805,N_5132,N_5613);
and U10806 (N_10806,N_6064,N_5508);
xnor U10807 (N_10807,N_7819,N_6654);
or U10808 (N_10808,N_5403,N_6373);
nor U10809 (N_10809,N_4731,N_6050);
and U10810 (N_10810,N_5653,N_4039);
xnor U10811 (N_10811,N_4193,N_5839);
or U10812 (N_10812,N_6635,N_5211);
nor U10813 (N_10813,N_5270,N_4724);
nor U10814 (N_10814,N_5496,N_5909);
nor U10815 (N_10815,N_4386,N_5450);
nor U10816 (N_10816,N_5203,N_6527);
xnor U10817 (N_10817,N_5728,N_6061);
nand U10818 (N_10818,N_6965,N_5664);
nand U10819 (N_10819,N_6880,N_5440);
nand U10820 (N_10820,N_7644,N_5393);
or U10821 (N_10821,N_7904,N_6168);
nor U10822 (N_10822,N_6362,N_5437);
nand U10823 (N_10823,N_4744,N_5464);
nand U10824 (N_10824,N_5758,N_6195);
nor U10825 (N_10825,N_6195,N_5781);
and U10826 (N_10826,N_5133,N_7887);
and U10827 (N_10827,N_7477,N_6026);
and U10828 (N_10828,N_4417,N_5073);
and U10829 (N_10829,N_4244,N_4769);
nor U10830 (N_10830,N_5202,N_7907);
xor U10831 (N_10831,N_7050,N_6210);
and U10832 (N_10832,N_6334,N_7693);
xnor U10833 (N_10833,N_7763,N_7225);
and U10834 (N_10834,N_5594,N_5959);
nand U10835 (N_10835,N_7492,N_5580);
nor U10836 (N_10836,N_4363,N_5657);
and U10837 (N_10837,N_7364,N_4479);
xor U10838 (N_10838,N_5447,N_7269);
nor U10839 (N_10839,N_7094,N_4698);
or U10840 (N_10840,N_7125,N_7806);
xor U10841 (N_10841,N_6612,N_4005);
nor U10842 (N_10842,N_6480,N_7296);
or U10843 (N_10843,N_7315,N_6544);
and U10844 (N_10844,N_5780,N_4196);
xnor U10845 (N_10845,N_7504,N_6609);
or U10846 (N_10846,N_6721,N_7870);
nand U10847 (N_10847,N_6146,N_4744);
xnor U10848 (N_10848,N_5697,N_7050);
or U10849 (N_10849,N_7297,N_4375);
or U10850 (N_10850,N_6386,N_5317);
and U10851 (N_10851,N_4349,N_7807);
nor U10852 (N_10852,N_6282,N_4566);
nand U10853 (N_10853,N_6833,N_6050);
or U10854 (N_10854,N_7635,N_7757);
xnor U10855 (N_10855,N_5797,N_5770);
xor U10856 (N_10856,N_7714,N_7691);
xnor U10857 (N_10857,N_4653,N_5865);
and U10858 (N_10858,N_5394,N_6923);
xnor U10859 (N_10859,N_6866,N_6790);
or U10860 (N_10860,N_5498,N_6585);
or U10861 (N_10861,N_4591,N_5937);
and U10862 (N_10862,N_7032,N_5121);
and U10863 (N_10863,N_4655,N_4352);
xor U10864 (N_10864,N_6252,N_5300);
xnor U10865 (N_10865,N_7779,N_7567);
nand U10866 (N_10866,N_5822,N_4885);
and U10867 (N_10867,N_6875,N_7002);
xor U10868 (N_10868,N_4421,N_4361);
and U10869 (N_10869,N_6406,N_4341);
or U10870 (N_10870,N_4910,N_6073);
nor U10871 (N_10871,N_4416,N_7306);
nor U10872 (N_10872,N_7221,N_5611);
nor U10873 (N_10873,N_7846,N_6687);
or U10874 (N_10874,N_4703,N_5032);
nor U10875 (N_10875,N_6365,N_6282);
xnor U10876 (N_10876,N_4123,N_4264);
and U10877 (N_10877,N_7495,N_4257);
or U10878 (N_10878,N_6422,N_6909);
nor U10879 (N_10879,N_7352,N_4019);
and U10880 (N_10880,N_5273,N_7957);
nor U10881 (N_10881,N_6324,N_4643);
xor U10882 (N_10882,N_5766,N_4712);
and U10883 (N_10883,N_4146,N_7365);
nor U10884 (N_10884,N_6425,N_6679);
nor U10885 (N_10885,N_4175,N_6702);
nand U10886 (N_10886,N_6527,N_6025);
nor U10887 (N_10887,N_5136,N_7428);
and U10888 (N_10888,N_5130,N_7163);
or U10889 (N_10889,N_4222,N_6552);
xnor U10890 (N_10890,N_4851,N_5031);
xor U10891 (N_10891,N_4628,N_7562);
nor U10892 (N_10892,N_6156,N_7376);
or U10893 (N_10893,N_6835,N_4669);
xnor U10894 (N_10894,N_5332,N_4200);
and U10895 (N_10895,N_7586,N_6873);
nand U10896 (N_10896,N_7161,N_4012);
xor U10897 (N_10897,N_6806,N_5415);
and U10898 (N_10898,N_6758,N_5520);
nor U10899 (N_10899,N_7211,N_7027);
and U10900 (N_10900,N_6901,N_7665);
or U10901 (N_10901,N_6874,N_5347);
nor U10902 (N_10902,N_7981,N_4680);
nand U10903 (N_10903,N_7275,N_4707);
nor U10904 (N_10904,N_5140,N_6321);
and U10905 (N_10905,N_7308,N_5237);
or U10906 (N_10906,N_7811,N_7708);
and U10907 (N_10907,N_5964,N_6090);
and U10908 (N_10908,N_6778,N_4697);
nand U10909 (N_10909,N_5715,N_5363);
xor U10910 (N_10910,N_7810,N_6658);
or U10911 (N_10911,N_6575,N_6166);
xor U10912 (N_10912,N_5418,N_7708);
and U10913 (N_10913,N_7622,N_4910);
and U10914 (N_10914,N_4483,N_4966);
nand U10915 (N_10915,N_7973,N_7727);
nor U10916 (N_10916,N_4301,N_6385);
and U10917 (N_10917,N_7023,N_4372);
and U10918 (N_10918,N_6613,N_5108);
and U10919 (N_10919,N_7525,N_7168);
or U10920 (N_10920,N_5548,N_6675);
or U10921 (N_10921,N_4552,N_5544);
xnor U10922 (N_10922,N_7680,N_4648);
nand U10923 (N_10923,N_7319,N_7669);
or U10924 (N_10924,N_7204,N_5023);
xnor U10925 (N_10925,N_6957,N_7349);
nor U10926 (N_10926,N_4271,N_7488);
nor U10927 (N_10927,N_7559,N_5022);
and U10928 (N_10928,N_6399,N_7126);
or U10929 (N_10929,N_6915,N_4638);
nor U10930 (N_10930,N_7131,N_7651);
xor U10931 (N_10931,N_4724,N_6177);
nor U10932 (N_10932,N_5484,N_7399);
or U10933 (N_10933,N_7087,N_5203);
nor U10934 (N_10934,N_7462,N_4514);
and U10935 (N_10935,N_4025,N_7036);
or U10936 (N_10936,N_4573,N_4496);
or U10937 (N_10937,N_5243,N_4509);
nor U10938 (N_10938,N_5919,N_4663);
and U10939 (N_10939,N_6918,N_7548);
or U10940 (N_10940,N_7295,N_5547);
nor U10941 (N_10941,N_5622,N_4009);
and U10942 (N_10942,N_5966,N_5135);
or U10943 (N_10943,N_5919,N_6149);
or U10944 (N_10944,N_5332,N_6143);
nand U10945 (N_10945,N_4728,N_6640);
nor U10946 (N_10946,N_4174,N_5965);
xor U10947 (N_10947,N_4085,N_4903);
xnor U10948 (N_10948,N_5602,N_7958);
nand U10949 (N_10949,N_7193,N_4448);
xnor U10950 (N_10950,N_4192,N_4631);
and U10951 (N_10951,N_4012,N_6716);
nand U10952 (N_10952,N_4879,N_7054);
or U10953 (N_10953,N_4852,N_6601);
xor U10954 (N_10954,N_6895,N_7900);
or U10955 (N_10955,N_4770,N_5942);
nor U10956 (N_10956,N_6274,N_4978);
nand U10957 (N_10957,N_4331,N_4967);
and U10958 (N_10958,N_5429,N_4527);
nor U10959 (N_10959,N_6513,N_5140);
or U10960 (N_10960,N_6028,N_4994);
and U10961 (N_10961,N_7769,N_6288);
xnor U10962 (N_10962,N_5825,N_4272);
nor U10963 (N_10963,N_4308,N_4879);
nor U10964 (N_10964,N_4300,N_5854);
and U10965 (N_10965,N_4425,N_7278);
and U10966 (N_10966,N_7057,N_4544);
and U10967 (N_10967,N_4958,N_7016);
nor U10968 (N_10968,N_4990,N_5459);
nand U10969 (N_10969,N_5195,N_6567);
xor U10970 (N_10970,N_5381,N_4115);
or U10971 (N_10971,N_4023,N_6594);
nand U10972 (N_10972,N_4208,N_4379);
nand U10973 (N_10973,N_4334,N_5750);
xnor U10974 (N_10974,N_7617,N_5135);
and U10975 (N_10975,N_7549,N_6932);
nor U10976 (N_10976,N_6234,N_6266);
nand U10977 (N_10977,N_5672,N_7118);
or U10978 (N_10978,N_4781,N_4002);
nand U10979 (N_10979,N_7835,N_7722);
xnor U10980 (N_10980,N_7937,N_6103);
nand U10981 (N_10981,N_5522,N_5243);
nand U10982 (N_10982,N_7998,N_4141);
nor U10983 (N_10983,N_7868,N_7748);
and U10984 (N_10984,N_6530,N_4117);
and U10985 (N_10985,N_5832,N_7820);
xor U10986 (N_10986,N_6773,N_4749);
xnor U10987 (N_10987,N_4818,N_4322);
nor U10988 (N_10988,N_6194,N_5297);
or U10989 (N_10989,N_6798,N_4495);
xor U10990 (N_10990,N_4094,N_7369);
nand U10991 (N_10991,N_6177,N_5358);
xnor U10992 (N_10992,N_6394,N_4393);
or U10993 (N_10993,N_4048,N_7713);
or U10994 (N_10994,N_7826,N_4346);
nand U10995 (N_10995,N_4065,N_5306);
and U10996 (N_10996,N_7707,N_5425);
xnor U10997 (N_10997,N_7153,N_6744);
nor U10998 (N_10998,N_7349,N_6557);
and U10999 (N_10999,N_4331,N_7139);
xnor U11000 (N_11000,N_7773,N_6439);
and U11001 (N_11001,N_5437,N_7276);
nor U11002 (N_11002,N_5755,N_4859);
nor U11003 (N_11003,N_6904,N_6173);
or U11004 (N_11004,N_6868,N_6923);
xor U11005 (N_11005,N_5556,N_7762);
or U11006 (N_11006,N_5540,N_4077);
or U11007 (N_11007,N_5386,N_7041);
xnor U11008 (N_11008,N_4210,N_4101);
xor U11009 (N_11009,N_5304,N_4222);
and U11010 (N_11010,N_7860,N_4399);
xor U11011 (N_11011,N_7930,N_7640);
xor U11012 (N_11012,N_7357,N_5360);
or U11013 (N_11013,N_7405,N_4802);
nor U11014 (N_11014,N_6185,N_6134);
or U11015 (N_11015,N_4880,N_5288);
and U11016 (N_11016,N_5323,N_5326);
xnor U11017 (N_11017,N_4151,N_4905);
nor U11018 (N_11018,N_6924,N_5089);
xnor U11019 (N_11019,N_7376,N_4957);
or U11020 (N_11020,N_6564,N_5654);
or U11021 (N_11021,N_6204,N_5807);
nand U11022 (N_11022,N_5184,N_7426);
nor U11023 (N_11023,N_5679,N_7727);
nor U11024 (N_11024,N_5304,N_7128);
or U11025 (N_11025,N_6303,N_5733);
xnor U11026 (N_11026,N_5567,N_6573);
and U11027 (N_11027,N_7225,N_4907);
nor U11028 (N_11028,N_4953,N_6259);
nor U11029 (N_11029,N_6707,N_6098);
or U11030 (N_11030,N_4908,N_5060);
or U11031 (N_11031,N_5223,N_6079);
nor U11032 (N_11032,N_7635,N_7182);
nand U11033 (N_11033,N_5932,N_6343);
or U11034 (N_11034,N_7104,N_6722);
and U11035 (N_11035,N_6485,N_6390);
xor U11036 (N_11036,N_4990,N_7903);
and U11037 (N_11037,N_4264,N_4039);
nand U11038 (N_11038,N_4869,N_5975);
nand U11039 (N_11039,N_5037,N_5268);
xnor U11040 (N_11040,N_5208,N_6700);
nor U11041 (N_11041,N_5431,N_6020);
or U11042 (N_11042,N_4077,N_7854);
nand U11043 (N_11043,N_4050,N_4134);
nand U11044 (N_11044,N_6124,N_6528);
nand U11045 (N_11045,N_7925,N_6070);
or U11046 (N_11046,N_6384,N_7180);
or U11047 (N_11047,N_5658,N_7096);
or U11048 (N_11048,N_7334,N_4911);
and U11049 (N_11049,N_7896,N_5064);
nor U11050 (N_11050,N_4922,N_7656);
and U11051 (N_11051,N_6318,N_4581);
nand U11052 (N_11052,N_7944,N_5462);
nor U11053 (N_11053,N_4977,N_4872);
and U11054 (N_11054,N_5596,N_4789);
nand U11055 (N_11055,N_7730,N_7836);
or U11056 (N_11056,N_6666,N_7135);
nand U11057 (N_11057,N_6622,N_6349);
nand U11058 (N_11058,N_4530,N_4451);
nor U11059 (N_11059,N_7745,N_6688);
xor U11060 (N_11060,N_4645,N_5411);
or U11061 (N_11061,N_6886,N_7517);
xor U11062 (N_11062,N_7299,N_6447);
and U11063 (N_11063,N_5018,N_7386);
nand U11064 (N_11064,N_7664,N_6920);
or U11065 (N_11065,N_7348,N_4360);
and U11066 (N_11066,N_5340,N_7418);
nor U11067 (N_11067,N_7406,N_7518);
nor U11068 (N_11068,N_7007,N_5834);
nand U11069 (N_11069,N_4695,N_4982);
and U11070 (N_11070,N_4925,N_5917);
or U11071 (N_11071,N_4349,N_6192);
nand U11072 (N_11072,N_7392,N_5765);
or U11073 (N_11073,N_5290,N_7530);
xnor U11074 (N_11074,N_5495,N_4509);
and U11075 (N_11075,N_7843,N_6847);
or U11076 (N_11076,N_6243,N_7356);
or U11077 (N_11077,N_6085,N_5312);
or U11078 (N_11078,N_4513,N_5154);
nand U11079 (N_11079,N_5153,N_4235);
nand U11080 (N_11080,N_7746,N_4619);
or U11081 (N_11081,N_5143,N_5066);
or U11082 (N_11082,N_4260,N_6664);
xnor U11083 (N_11083,N_4574,N_7766);
and U11084 (N_11084,N_6957,N_6578);
xnor U11085 (N_11085,N_6747,N_4977);
xor U11086 (N_11086,N_6129,N_7551);
nor U11087 (N_11087,N_7100,N_6277);
or U11088 (N_11088,N_5799,N_7469);
and U11089 (N_11089,N_4623,N_4651);
nand U11090 (N_11090,N_6481,N_4507);
or U11091 (N_11091,N_4195,N_6097);
nor U11092 (N_11092,N_4766,N_7944);
or U11093 (N_11093,N_6983,N_5520);
xnor U11094 (N_11094,N_5831,N_6982);
and U11095 (N_11095,N_4605,N_5367);
xor U11096 (N_11096,N_4911,N_4073);
xor U11097 (N_11097,N_4632,N_4802);
xor U11098 (N_11098,N_6262,N_7140);
nand U11099 (N_11099,N_5719,N_5125);
or U11100 (N_11100,N_6770,N_6278);
nand U11101 (N_11101,N_5299,N_5357);
xor U11102 (N_11102,N_6274,N_4397);
and U11103 (N_11103,N_4294,N_4221);
or U11104 (N_11104,N_6239,N_6937);
nor U11105 (N_11105,N_7149,N_5368);
or U11106 (N_11106,N_4744,N_5243);
xnor U11107 (N_11107,N_6319,N_6455);
nor U11108 (N_11108,N_5845,N_7793);
nor U11109 (N_11109,N_6143,N_7800);
nand U11110 (N_11110,N_6874,N_7805);
nand U11111 (N_11111,N_5271,N_6824);
nand U11112 (N_11112,N_5334,N_6636);
or U11113 (N_11113,N_7411,N_5493);
and U11114 (N_11114,N_4965,N_4450);
xor U11115 (N_11115,N_6197,N_4598);
xor U11116 (N_11116,N_5710,N_7332);
and U11117 (N_11117,N_4684,N_4508);
xnor U11118 (N_11118,N_5659,N_5667);
xnor U11119 (N_11119,N_5502,N_5917);
or U11120 (N_11120,N_5736,N_4298);
nor U11121 (N_11121,N_4506,N_5492);
xnor U11122 (N_11122,N_6502,N_7565);
or U11123 (N_11123,N_4351,N_4498);
or U11124 (N_11124,N_5809,N_7150);
nor U11125 (N_11125,N_7927,N_5877);
xnor U11126 (N_11126,N_4144,N_7446);
or U11127 (N_11127,N_5258,N_5293);
and U11128 (N_11128,N_7080,N_5317);
xor U11129 (N_11129,N_4329,N_7233);
nor U11130 (N_11130,N_5370,N_5693);
nand U11131 (N_11131,N_7878,N_5605);
nand U11132 (N_11132,N_5815,N_7384);
or U11133 (N_11133,N_6811,N_5112);
or U11134 (N_11134,N_7698,N_6993);
and U11135 (N_11135,N_6971,N_7300);
or U11136 (N_11136,N_6381,N_4847);
nand U11137 (N_11137,N_5775,N_6391);
nor U11138 (N_11138,N_7838,N_6645);
nor U11139 (N_11139,N_7090,N_6366);
nor U11140 (N_11140,N_4850,N_7364);
xor U11141 (N_11141,N_6169,N_7898);
and U11142 (N_11142,N_6012,N_6762);
xnor U11143 (N_11143,N_4721,N_5593);
xor U11144 (N_11144,N_7316,N_4981);
xnor U11145 (N_11145,N_7407,N_4745);
nand U11146 (N_11146,N_6317,N_5155);
nand U11147 (N_11147,N_4003,N_4610);
or U11148 (N_11148,N_4519,N_4672);
nand U11149 (N_11149,N_4980,N_7255);
and U11150 (N_11150,N_5127,N_4425);
or U11151 (N_11151,N_5849,N_7750);
nand U11152 (N_11152,N_7941,N_6412);
or U11153 (N_11153,N_6173,N_5984);
and U11154 (N_11154,N_4511,N_4135);
nor U11155 (N_11155,N_7211,N_4543);
nor U11156 (N_11156,N_5913,N_7414);
nand U11157 (N_11157,N_5555,N_7334);
nor U11158 (N_11158,N_4016,N_4652);
and U11159 (N_11159,N_4524,N_7677);
nor U11160 (N_11160,N_4296,N_5480);
xor U11161 (N_11161,N_4594,N_7025);
or U11162 (N_11162,N_5460,N_6202);
and U11163 (N_11163,N_6106,N_4707);
nor U11164 (N_11164,N_6596,N_6394);
and U11165 (N_11165,N_7077,N_5549);
xor U11166 (N_11166,N_7548,N_7901);
nor U11167 (N_11167,N_4755,N_6908);
or U11168 (N_11168,N_7806,N_7269);
nand U11169 (N_11169,N_4271,N_6459);
xnor U11170 (N_11170,N_4055,N_4984);
nor U11171 (N_11171,N_6951,N_7965);
or U11172 (N_11172,N_6621,N_4875);
xnor U11173 (N_11173,N_5631,N_5134);
and U11174 (N_11174,N_5387,N_5147);
or U11175 (N_11175,N_4738,N_4425);
xnor U11176 (N_11176,N_7839,N_7769);
xor U11177 (N_11177,N_5098,N_7809);
nor U11178 (N_11178,N_7358,N_6819);
and U11179 (N_11179,N_4479,N_7461);
xor U11180 (N_11180,N_5794,N_6854);
and U11181 (N_11181,N_4878,N_5604);
xor U11182 (N_11182,N_6655,N_6557);
nor U11183 (N_11183,N_7532,N_5783);
nor U11184 (N_11184,N_7680,N_6198);
or U11185 (N_11185,N_4683,N_5540);
nor U11186 (N_11186,N_7209,N_7244);
xnor U11187 (N_11187,N_5338,N_6330);
nand U11188 (N_11188,N_6485,N_5393);
nand U11189 (N_11189,N_6542,N_7049);
nand U11190 (N_11190,N_7450,N_7794);
or U11191 (N_11191,N_6280,N_6868);
nand U11192 (N_11192,N_7931,N_7445);
nor U11193 (N_11193,N_6397,N_7923);
and U11194 (N_11194,N_6049,N_4986);
xor U11195 (N_11195,N_4387,N_5437);
nor U11196 (N_11196,N_4647,N_4838);
xor U11197 (N_11197,N_4819,N_5694);
nor U11198 (N_11198,N_7989,N_5691);
or U11199 (N_11199,N_4958,N_5567);
or U11200 (N_11200,N_6099,N_7188);
xor U11201 (N_11201,N_7187,N_5488);
nand U11202 (N_11202,N_4457,N_7079);
nor U11203 (N_11203,N_5349,N_7067);
xnor U11204 (N_11204,N_5239,N_4419);
and U11205 (N_11205,N_7886,N_7076);
nor U11206 (N_11206,N_5897,N_7747);
or U11207 (N_11207,N_4644,N_6764);
xor U11208 (N_11208,N_6172,N_7082);
nor U11209 (N_11209,N_7969,N_7822);
or U11210 (N_11210,N_6061,N_4765);
xnor U11211 (N_11211,N_4577,N_7166);
nand U11212 (N_11212,N_4337,N_6140);
or U11213 (N_11213,N_5660,N_5922);
and U11214 (N_11214,N_4021,N_7367);
nor U11215 (N_11215,N_5848,N_5625);
nor U11216 (N_11216,N_7893,N_4932);
and U11217 (N_11217,N_4306,N_7449);
and U11218 (N_11218,N_7324,N_7757);
nor U11219 (N_11219,N_6975,N_7328);
and U11220 (N_11220,N_7381,N_4424);
nor U11221 (N_11221,N_5732,N_6689);
nand U11222 (N_11222,N_5268,N_7533);
nor U11223 (N_11223,N_4172,N_5445);
nor U11224 (N_11224,N_5936,N_6059);
xor U11225 (N_11225,N_4286,N_7084);
nor U11226 (N_11226,N_6573,N_7857);
and U11227 (N_11227,N_4394,N_5996);
or U11228 (N_11228,N_4793,N_4560);
xor U11229 (N_11229,N_4028,N_4066);
nand U11230 (N_11230,N_4523,N_4041);
xor U11231 (N_11231,N_4725,N_4754);
or U11232 (N_11232,N_4719,N_4296);
xor U11233 (N_11233,N_6483,N_7720);
xor U11234 (N_11234,N_7500,N_5667);
nor U11235 (N_11235,N_7592,N_6080);
xnor U11236 (N_11236,N_4786,N_4999);
nor U11237 (N_11237,N_6141,N_4519);
nor U11238 (N_11238,N_6372,N_4745);
nor U11239 (N_11239,N_4041,N_6907);
nand U11240 (N_11240,N_4675,N_4729);
nor U11241 (N_11241,N_6620,N_4809);
and U11242 (N_11242,N_5489,N_6954);
nand U11243 (N_11243,N_5242,N_6073);
nand U11244 (N_11244,N_6286,N_7270);
nand U11245 (N_11245,N_5502,N_4030);
and U11246 (N_11246,N_6979,N_6702);
or U11247 (N_11247,N_4829,N_5206);
nor U11248 (N_11248,N_7746,N_4564);
xnor U11249 (N_11249,N_4578,N_5398);
or U11250 (N_11250,N_4928,N_7787);
nand U11251 (N_11251,N_7613,N_7976);
xor U11252 (N_11252,N_7782,N_7542);
nand U11253 (N_11253,N_4591,N_4128);
xnor U11254 (N_11254,N_6963,N_4337);
or U11255 (N_11255,N_6091,N_6249);
and U11256 (N_11256,N_6515,N_5863);
and U11257 (N_11257,N_5574,N_6570);
or U11258 (N_11258,N_5166,N_5449);
nor U11259 (N_11259,N_4154,N_5589);
xor U11260 (N_11260,N_7367,N_5602);
nor U11261 (N_11261,N_4040,N_5107);
nand U11262 (N_11262,N_6477,N_6738);
nor U11263 (N_11263,N_5541,N_7700);
xor U11264 (N_11264,N_6747,N_7892);
or U11265 (N_11265,N_5122,N_4080);
nand U11266 (N_11266,N_4318,N_5837);
nand U11267 (N_11267,N_5816,N_7848);
nand U11268 (N_11268,N_7769,N_4724);
or U11269 (N_11269,N_6323,N_5102);
or U11270 (N_11270,N_5903,N_7678);
nand U11271 (N_11271,N_5043,N_5184);
nor U11272 (N_11272,N_6309,N_7667);
nor U11273 (N_11273,N_6785,N_6144);
nand U11274 (N_11274,N_4316,N_6850);
xnor U11275 (N_11275,N_6077,N_6938);
or U11276 (N_11276,N_4689,N_6237);
and U11277 (N_11277,N_7751,N_4846);
and U11278 (N_11278,N_7332,N_5004);
nand U11279 (N_11279,N_7200,N_6265);
nand U11280 (N_11280,N_4792,N_4577);
nor U11281 (N_11281,N_7291,N_5077);
and U11282 (N_11282,N_6012,N_7712);
nor U11283 (N_11283,N_5762,N_7525);
and U11284 (N_11284,N_5834,N_4623);
and U11285 (N_11285,N_7148,N_5422);
nor U11286 (N_11286,N_4624,N_5062);
nand U11287 (N_11287,N_6446,N_4974);
xor U11288 (N_11288,N_7715,N_5088);
nor U11289 (N_11289,N_6793,N_5667);
or U11290 (N_11290,N_4133,N_4643);
or U11291 (N_11291,N_5374,N_6812);
nand U11292 (N_11292,N_7910,N_7936);
nor U11293 (N_11293,N_4264,N_7997);
nor U11294 (N_11294,N_5379,N_4209);
xor U11295 (N_11295,N_5162,N_6115);
nand U11296 (N_11296,N_7225,N_7505);
and U11297 (N_11297,N_4445,N_5185);
or U11298 (N_11298,N_4589,N_6776);
and U11299 (N_11299,N_6778,N_5901);
xor U11300 (N_11300,N_5042,N_5386);
or U11301 (N_11301,N_7298,N_5343);
and U11302 (N_11302,N_7904,N_7520);
nor U11303 (N_11303,N_5851,N_6407);
nand U11304 (N_11304,N_5656,N_4799);
xnor U11305 (N_11305,N_7974,N_5914);
or U11306 (N_11306,N_5523,N_4665);
nand U11307 (N_11307,N_7045,N_4242);
xor U11308 (N_11308,N_7761,N_6973);
nor U11309 (N_11309,N_4513,N_5607);
xor U11310 (N_11310,N_7494,N_5812);
nand U11311 (N_11311,N_4157,N_4839);
or U11312 (N_11312,N_7449,N_5985);
or U11313 (N_11313,N_4009,N_5275);
nor U11314 (N_11314,N_4579,N_6703);
nor U11315 (N_11315,N_5213,N_5599);
nand U11316 (N_11316,N_6956,N_4134);
nor U11317 (N_11317,N_7275,N_7082);
or U11318 (N_11318,N_4338,N_5023);
nand U11319 (N_11319,N_6441,N_6814);
nand U11320 (N_11320,N_6181,N_5716);
or U11321 (N_11321,N_7635,N_4611);
and U11322 (N_11322,N_6611,N_6790);
or U11323 (N_11323,N_6873,N_5911);
nor U11324 (N_11324,N_6547,N_7593);
xor U11325 (N_11325,N_5712,N_5150);
or U11326 (N_11326,N_4520,N_6741);
and U11327 (N_11327,N_7445,N_7001);
or U11328 (N_11328,N_6115,N_5733);
or U11329 (N_11329,N_6597,N_7184);
xor U11330 (N_11330,N_5937,N_6271);
or U11331 (N_11331,N_6818,N_5536);
or U11332 (N_11332,N_7514,N_7374);
nor U11333 (N_11333,N_5079,N_7234);
nor U11334 (N_11334,N_6402,N_7840);
and U11335 (N_11335,N_5502,N_6864);
nand U11336 (N_11336,N_6184,N_4598);
or U11337 (N_11337,N_4931,N_5337);
nor U11338 (N_11338,N_7217,N_7674);
nor U11339 (N_11339,N_6845,N_5519);
and U11340 (N_11340,N_7139,N_4100);
and U11341 (N_11341,N_7443,N_7498);
or U11342 (N_11342,N_5534,N_4051);
or U11343 (N_11343,N_6064,N_6792);
xnor U11344 (N_11344,N_5390,N_6365);
or U11345 (N_11345,N_6747,N_4272);
or U11346 (N_11346,N_7150,N_6009);
nand U11347 (N_11347,N_5828,N_5422);
or U11348 (N_11348,N_5427,N_7805);
nor U11349 (N_11349,N_4846,N_4756);
nor U11350 (N_11350,N_7085,N_4891);
or U11351 (N_11351,N_6158,N_7393);
xor U11352 (N_11352,N_6321,N_5821);
xor U11353 (N_11353,N_4270,N_4259);
nand U11354 (N_11354,N_4430,N_4347);
nand U11355 (N_11355,N_7404,N_5396);
nand U11356 (N_11356,N_5478,N_7387);
xnor U11357 (N_11357,N_7097,N_5826);
or U11358 (N_11358,N_6142,N_7190);
xnor U11359 (N_11359,N_6080,N_4745);
nor U11360 (N_11360,N_7919,N_4258);
and U11361 (N_11361,N_5681,N_7519);
nand U11362 (N_11362,N_6867,N_7417);
nor U11363 (N_11363,N_5911,N_4309);
nor U11364 (N_11364,N_6089,N_7400);
xnor U11365 (N_11365,N_4933,N_5753);
nand U11366 (N_11366,N_4871,N_4126);
and U11367 (N_11367,N_6940,N_6984);
xor U11368 (N_11368,N_7050,N_5493);
or U11369 (N_11369,N_6865,N_7520);
and U11370 (N_11370,N_7692,N_7738);
xor U11371 (N_11371,N_4672,N_6419);
xor U11372 (N_11372,N_7837,N_6388);
nor U11373 (N_11373,N_4812,N_6706);
xor U11374 (N_11374,N_4958,N_6387);
or U11375 (N_11375,N_6184,N_5716);
nand U11376 (N_11376,N_7153,N_6991);
or U11377 (N_11377,N_6191,N_6968);
nor U11378 (N_11378,N_5789,N_4003);
or U11379 (N_11379,N_4926,N_6642);
or U11380 (N_11380,N_4697,N_4588);
or U11381 (N_11381,N_6809,N_5742);
nand U11382 (N_11382,N_7576,N_7889);
or U11383 (N_11383,N_4655,N_5871);
or U11384 (N_11384,N_7167,N_7949);
nor U11385 (N_11385,N_5178,N_7308);
or U11386 (N_11386,N_4530,N_5365);
and U11387 (N_11387,N_6842,N_6803);
nand U11388 (N_11388,N_7110,N_6546);
nand U11389 (N_11389,N_4927,N_5808);
and U11390 (N_11390,N_7372,N_5625);
nand U11391 (N_11391,N_4009,N_4800);
nor U11392 (N_11392,N_5196,N_4783);
and U11393 (N_11393,N_5807,N_4383);
or U11394 (N_11394,N_4009,N_5108);
or U11395 (N_11395,N_6810,N_5799);
and U11396 (N_11396,N_4581,N_5988);
and U11397 (N_11397,N_6870,N_6830);
or U11398 (N_11398,N_7168,N_4520);
or U11399 (N_11399,N_6746,N_7608);
nor U11400 (N_11400,N_7781,N_7739);
or U11401 (N_11401,N_6900,N_4410);
nor U11402 (N_11402,N_5651,N_5266);
xor U11403 (N_11403,N_4617,N_5293);
and U11404 (N_11404,N_4307,N_4241);
xnor U11405 (N_11405,N_7068,N_4281);
nand U11406 (N_11406,N_5821,N_7346);
and U11407 (N_11407,N_7642,N_5520);
nor U11408 (N_11408,N_6232,N_5074);
nor U11409 (N_11409,N_7913,N_6611);
nand U11410 (N_11410,N_6835,N_6479);
and U11411 (N_11411,N_7105,N_5102);
nand U11412 (N_11412,N_5776,N_4182);
xnor U11413 (N_11413,N_5147,N_5019);
xnor U11414 (N_11414,N_5558,N_6803);
nand U11415 (N_11415,N_7700,N_7055);
nor U11416 (N_11416,N_6675,N_6194);
and U11417 (N_11417,N_5044,N_7312);
and U11418 (N_11418,N_5090,N_4549);
nor U11419 (N_11419,N_4029,N_4415);
xor U11420 (N_11420,N_5497,N_4523);
and U11421 (N_11421,N_7886,N_7471);
or U11422 (N_11422,N_7103,N_5260);
and U11423 (N_11423,N_6603,N_7574);
or U11424 (N_11424,N_6192,N_7476);
and U11425 (N_11425,N_4963,N_5633);
nand U11426 (N_11426,N_7881,N_7232);
nor U11427 (N_11427,N_6339,N_7720);
or U11428 (N_11428,N_6835,N_7931);
or U11429 (N_11429,N_7127,N_6892);
or U11430 (N_11430,N_5367,N_7926);
nor U11431 (N_11431,N_6192,N_4170);
or U11432 (N_11432,N_5739,N_5875);
or U11433 (N_11433,N_7982,N_4587);
xnor U11434 (N_11434,N_6264,N_7764);
nand U11435 (N_11435,N_5529,N_7517);
xor U11436 (N_11436,N_7874,N_7657);
nor U11437 (N_11437,N_4264,N_6206);
or U11438 (N_11438,N_7372,N_5617);
xor U11439 (N_11439,N_4659,N_7908);
or U11440 (N_11440,N_5387,N_6314);
and U11441 (N_11441,N_7875,N_7313);
nor U11442 (N_11442,N_6674,N_5770);
nor U11443 (N_11443,N_6063,N_6501);
xnor U11444 (N_11444,N_4444,N_4542);
nand U11445 (N_11445,N_7955,N_4691);
or U11446 (N_11446,N_5453,N_4616);
nor U11447 (N_11447,N_4205,N_5058);
xor U11448 (N_11448,N_4700,N_4156);
or U11449 (N_11449,N_4500,N_4527);
xor U11450 (N_11450,N_5890,N_5947);
xor U11451 (N_11451,N_5217,N_7957);
nand U11452 (N_11452,N_6957,N_7315);
or U11453 (N_11453,N_5549,N_5909);
nand U11454 (N_11454,N_7627,N_4459);
nand U11455 (N_11455,N_4635,N_5816);
nor U11456 (N_11456,N_4966,N_6712);
nor U11457 (N_11457,N_4636,N_6871);
nor U11458 (N_11458,N_7823,N_6744);
or U11459 (N_11459,N_7448,N_7244);
or U11460 (N_11460,N_5298,N_7011);
or U11461 (N_11461,N_5504,N_6748);
xnor U11462 (N_11462,N_7748,N_7702);
or U11463 (N_11463,N_5492,N_5304);
and U11464 (N_11464,N_4415,N_4533);
nor U11465 (N_11465,N_4991,N_4113);
or U11466 (N_11466,N_7011,N_4490);
nor U11467 (N_11467,N_6162,N_6990);
nor U11468 (N_11468,N_4672,N_4764);
nor U11469 (N_11469,N_6015,N_7370);
and U11470 (N_11470,N_7294,N_6345);
nor U11471 (N_11471,N_4213,N_5619);
nand U11472 (N_11472,N_5596,N_4708);
nand U11473 (N_11473,N_6078,N_7848);
or U11474 (N_11474,N_4445,N_6707);
xor U11475 (N_11475,N_6066,N_7833);
nand U11476 (N_11476,N_6572,N_7656);
and U11477 (N_11477,N_6121,N_4564);
or U11478 (N_11478,N_4291,N_5394);
nor U11479 (N_11479,N_4434,N_7191);
xnor U11480 (N_11480,N_7671,N_6568);
and U11481 (N_11481,N_6191,N_4622);
nor U11482 (N_11482,N_5347,N_4862);
and U11483 (N_11483,N_7637,N_7295);
nor U11484 (N_11484,N_5673,N_5788);
or U11485 (N_11485,N_6841,N_7707);
or U11486 (N_11486,N_5756,N_5633);
nand U11487 (N_11487,N_7820,N_5267);
nand U11488 (N_11488,N_5665,N_7865);
xnor U11489 (N_11489,N_6965,N_7483);
nand U11490 (N_11490,N_6545,N_6721);
or U11491 (N_11491,N_5520,N_4460);
and U11492 (N_11492,N_4800,N_7879);
and U11493 (N_11493,N_7780,N_7667);
nor U11494 (N_11494,N_5514,N_5315);
nand U11495 (N_11495,N_5552,N_7357);
nand U11496 (N_11496,N_4703,N_5855);
nand U11497 (N_11497,N_4582,N_6426);
or U11498 (N_11498,N_4476,N_6164);
or U11499 (N_11499,N_6412,N_4867);
nand U11500 (N_11500,N_6960,N_5327);
nor U11501 (N_11501,N_7659,N_7291);
nand U11502 (N_11502,N_7631,N_6803);
nor U11503 (N_11503,N_7225,N_6222);
xor U11504 (N_11504,N_5283,N_4071);
nand U11505 (N_11505,N_7786,N_6650);
nor U11506 (N_11506,N_7013,N_6266);
or U11507 (N_11507,N_7860,N_6105);
or U11508 (N_11508,N_6394,N_5902);
nand U11509 (N_11509,N_5043,N_5826);
nor U11510 (N_11510,N_7091,N_5755);
xor U11511 (N_11511,N_4859,N_4674);
or U11512 (N_11512,N_7708,N_6826);
or U11513 (N_11513,N_7910,N_6309);
nand U11514 (N_11514,N_7304,N_6182);
or U11515 (N_11515,N_7179,N_5729);
nand U11516 (N_11516,N_7202,N_4845);
nand U11517 (N_11517,N_6205,N_7393);
nand U11518 (N_11518,N_7712,N_5308);
nor U11519 (N_11519,N_6528,N_6808);
and U11520 (N_11520,N_6033,N_7556);
or U11521 (N_11521,N_5951,N_4889);
or U11522 (N_11522,N_5137,N_7328);
and U11523 (N_11523,N_6607,N_7643);
nand U11524 (N_11524,N_5935,N_5969);
nor U11525 (N_11525,N_5694,N_6939);
xor U11526 (N_11526,N_5533,N_6220);
xnor U11527 (N_11527,N_7905,N_6738);
nand U11528 (N_11528,N_5279,N_7462);
nor U11529 (N_11529,N_6483,N_7060);
nor U11530 (N_11530,N_7217,N_6009);
or U11531 (N_11531,N_5615,N_4598);
and U11532 (N_11532,N_6391,N_6067);
or U11533 (N_11533,N_4089,N_5642);
nand U11534 (N_11534,N_5543,N_5085);
xnor U11535 (N_11535,N_5624,N_6414);
and U11536 (N_11536,N_6331,N_7971);
or U11537 (N_11537,N_4515,N_4975);
or U11538 (N_11538,N_7510,N_6274);
and U11539 (N_11539,N_6647,N_7527);
xnor U11540 (N_11540,N_4371,N_4174);
nor U11541 (N_11541,N_4795,N_7142);
nor U11542 (N_11542,N_5002,N_6478);
or U11543 (N_11543,N_7712,N_5828);
xnor U11544 (N_11544,N_5031,N_5918);
xor U11545 (N_11545,N_5973,N_5383);
xnor U11546 (N_11546,N_6072,N_5127);
and U11547 (N_11547,N_7144,N_5361);
xor U11548 (N_11548,N_4221,N_4401);
nand U11549 (N_11549,N_7985,N_6518);
nand U11550 (N_11550,N_7759,N_6582);
xor U11551 (N_11551,N_4567,N_4389);
nand U11552 (N_11552,N_5103,N_4197);
xnor U11553 (N_11553,N_6177,N_6929);
xnor U11554 (N_11554,N_6568,N_7569);
nor U11555 (N_11555,N_4020,N_4555);
and U11556 (N_11556,N_5516,N_6035);
nor U11557 (N_11557,N_6410,N_5911);
and U11558 (N_11558,N_4031,N_7451);
nand U11559 (N_11559,N_4945,N_4913);
xnor U11560 (N_11560,N_7564,N_4738);
xor U11561 (N_11561,N_6470,N_7797);
and U11562 (N_11562,N_6289,N_7896);
and U11563 (N_11563,N_6383,N_5123);
nor U11564 (N_11564,N_6351,N_5577);
nor U11565 (N_11565,N_7081,N_5825);
nand U11566 (N_11566,N_4734,N_7531);
or U11567 (N_11567,N_7955,N_4312);
nand U11568 (N_11568,N_7634,N_7992);
or U11569 (N_11569,N_5260,N_7733);
nand U11570 (N_11570,N_4644,N_5869);
and U11571 (N_11571,N_4286,N_4685);
nor U11572 (N_11572,N_5973,N_5596);
xor U11573 (N_11573,N_5074,N_6615);
and U11574 (N_11574,N_4086,N_6782);
or U11575 (N_11575,N_7395,N_5207);
or U11576 (N_11576,N_4527,N_4610);
or U11577 (N_11577,N_7194,N_6725);
or U11578 (N_11578,N_6177,N_7455);
nand U11579 (N_11579,N_7814,N_4569);
and U11580 (N_11580,N_6742,N_5828);
xnor U11581 (N_11581,N_5735,N_4761);
nor U11582 (N_11582,N_7528,N_7964);
nor U11583 (N_11583,N_6492,N_6470);
nand U11584 (N_11584,N_5664,N_6178);
nor U11585 (N_11585,N_4260,N_7952);
xor U11586 (N_11586,N_5810,N_4800);
nand U11587 (N_11587,N_7167,N_4295);
nor U11588 (N_11588,N_7840,N_5249);
xor U11589 (N_11589,N_4406,N_6802);
and U11590 (N_11590,N_7504,N_7978);
or U11591 (N_11591,N_5525,N_6450);
or U11592 (N_11592,N_7478,N_6643);
nand U11593 (N_11593,N_4960,N_6680);
nor U11594 (N_11594,N_5365,N_7020);
nor U11595 (N_11595,N_6173,N_6199);
nand U11596 (N_11596,N_4709,N_4894);
xor U11597 (N_11597,N_4706,N_6263);
nand U11598 (N_11598,N_6906,N_6151);
nand U11599 (N_11599,N_6105,N_5904);
xor U11600 (N_11600,N_6049,N_7655);
nor U11601 (N_11601,N_4658,N_5215);
nor U11602 (N_11602,N_4930,N_7525);
nor U11603 (N_11603,N_5513,N_5304);
nand U11604 (N_11604,N_6119,N_6999);
and U11605 (N_11605,N_7671,N_5030);
nor U11606 (N_11606,N_5296,N_6585);
nand U11607 (N_11607,N_4525,N_5121);
or U11608 (N_11608,N_6595,N_4699);
nor U11609 (N_11609,N_6861,N_7607);
and U11610 (N_11610,N_5996,N_5948);
and U11611 (N_11611,N_5246,N_7910);
nor U11612 (N_11612,N_7061,N_4147);
nand U11613 (N_11613,N_5546,N_5677);
nand U11614 (N_11614,N_5279,N_4751);
xor U11615 (N_11615,N_6036,N_6260);
or U11616 (N_11616,N_6236,N_6025);
and U11617 (N_11617,N_5555,N_7279);
nor U11618 (N_11618,N_7143,N_7881);
or U11619 (N_11619,N_6494,N_4659);
nand U11620 (N_11620,N_7699,N_4747);
nor U11621 (N_11621,N_6029,N_4182);
xnor U11622 (N_11622,N_7097,N_6856);
nor U11623 (N_11623,N_7947,N_6231);
nand U11624 (N_11624,N_6172,N_5839);
and U11625 (N_11625,N_5101,N_4351);
nand U11626 (N_11626,N_6207,N_7201);
or U11627 (N_11627,N_5231,N_7030);
or U11628 (N_11628,N_6329,N_5983);
and U11629 (N_11629,N_6129,N_5165);
and U11630 (N_11630,N_7306,N_7866);
and U11631 (N_11631,N_6180,N_7169);
nor U11632 (N_11632,N_5925,N_4848);
nor U11633 (N_11633,N_7186,N_4354);
nand U11634 (N_11634,N_4208,N_6526);
nor U11635 (N_11635,N_6915,N_6234);
nand U11636 (N_11636,N_6835,N_5010);
or U11637 (N_11637,N_7518,N_7904);
nand U11638 (N_11638,N_4387,N_5839);
xor U11639 (N_11639,N_6534,N_6189);
nor U11640 (N_11640,N_6467,N_4255);
and U11641 (N_11641,N_7189,N_7759);
and U11642 (N_11642,N_7178,N_6978);
and U11643 (N_11643,N_7571,N_4493);
nor U11644 (N_11644,N_6597,N_4113);
nand U11645 (N_11645,N_5114,N_7161);
xor U11646 (N_11646,N_4227,N_6052);
nor U11647 (N_11647,N_7616,N_4175);
xnor U11648 (N_11648,N_5139,N_4938);
nor U11649 (N_11649,N_6021,N_7779);
nand U11650 (N_11650,N_5192,N_4172);
or U11651 (N_11651,N_4408,N_4322);
xor U11652 (N_11652,N_4130,N_5397);
and U11653 (N_11653,N_4455,N_4964);
xor U11654 (N_11654,N_6354,N_7090);
nand U11655 (N_11655,N_5742,N_6641);
nor U11656 (N_11656,N_5634,N_4780);
or U11657 (N_11657,N_4780,N_4874);
nor U11658 (N_11658,N_6844,N_6104);
nor U11659 (N_11659,N_5758,N_5700);
or U11660 (N_11660,N_4787,N_6205);
nand U11661 (N_11661,N_5207,N_5731);
and U11662 (N_11662,N_7733,N_7300);
nor U11663 (N_11663,N_6626,N_7098);
or U11664 (N_11664,N_6275,N_6473);
nor U11665 (N_11665,N_6923,N_4909);
nand U11666 (N_11666,N_4102,N_5600);
nand U11667 (N_11667,N_4259,N_6041);
or U11668 (N_11668,N_6802,N_6581);
nor U11669 (N_11669,N_7915,N_6827);
xor U11670 (N_11670,N_5474,N_6168);
and U11671 (N_11671,N_7482,N_5890);
xnor U11672 (N_11672,N_5289,N_5746);
or U11673 (N_11673,N_4268,N_7917);
and U11674 (N_11674,N_7704,N_7495);
nand U11675 (N_11675,N_4714,N_6170);
or U11676 (N_11676,N_7348,N_4310);
nor U11677 (N_11677,N_5642,N_4590);
nand U11678 (N_11678,N_5648,N_5007);
and U11679 (N_11679,N_5162,N_6234);
xnor U11680 (N_11680,N_4152,N_7891);
nand U11681 (N_11681,N_7090,N_4296);
nor U11682 (N_11682,N_4401,N_6828);
or U11683 (N_11683,N_5956,N_4153);
or U11684 (N_11684,N_4002,N_6269);
xor U11685 (N_11685,N_4816,N_4762);
xnor U11686 (N_11686,N_7651,N_7785);
xor U11687 (N_11687,N_5268,N_7041);
nor U11688 (N_11688,N_4475,N_4695);
nor U11689 (N_11689,N_4007,N_7637);
xnor U11690 (N_11690,N_7828,N_5804);
xor U11691 (N_11691,N_5980,N_5682);
nor U11692 (N_11692,N_4339,N_6884);
nor U11693 (N_11693,N_4648,N_5815);
nand U11694 (N_11694,N_5910,N_6898);
xor U11695 (N_11695,N_4438,N_7986);
or U11696 (N_11696,N_7349,N_7438);
nand U11697 (N_11697,N_5704,N_5238);
xor U11698 (N_11698,N_7964,N_5706);
or U11699 (N_11699,N_6501,N_6771);
xor U11700 (N_11700,N_5820,N_6856);
nand U11701 (N_11701,N_5233,N_4303);
xnor U11702 (N_11702,N_7103,N_6874);
nand U11703 (N_11703,N_7413,N_6435);
xnor U11704 (N_11704,N_5418,N_7065);
nor U11705 (N_11705,N_7767,N_4260);
or U11706 (N_11706,N_7559,N_6707);
nand U11707 (N_11707,N_7079,N_5303);
nand U11708 (N_11708,N_6402,N_7045);
xnor U11709 (N_11709,N_7419,N_6700);
nor U11710 (N_11710,N_5415,N_7678);
xnor U11711 (N_11711,N_6001,N_5189);
xnor U11712 (N_11712,N_5688,N_5230);
nand U11713 (N_11713,N_6032,N_4806);
nor U11714 (N_11714,N_6893,N_5490);
nor U11715 (N_11715,N_4578,N_7535);
xor U11716 (N_11716,N_5871,N_6210);
nor U11717 (N_11717,N_6758,N_6224);
or U11718 (N_11718,N_6081,N_4010);
xnor U11719 (N_11719,N_6374,N_7519);
nand U11720 (N_11720,N_7214,N_4692);
xor U11721 (N_11721,N_5610,N_5453);
and U11722 (N_11722,N_6136,N_4754);
nor U11723 (N_11723,N_6828,N_4919);
or U11724 (N_11724,N_6163,N_4120);
xor U11725 (N_11725,N_4045,N_6882);
xnor U11726 (N_11726,N_7585,N_4316);
or U11727 (N_11727,N_6108,N_5828);
or U11728 (N_11728,N_6103,N_6942);
xor U11729 (N_11729,N_6977,N_5922);
and U11730 (N_11730,N_7201,N_5511);
nand U11731 (N_11731,N_5672,N_6817);
or U11732 (N_11732,N_4195,N_4788);
and U11733 (N_11733,N_6506,N_5640);
xor U11734 (N_11734,N_4847,N_4796);
xnor U11735 (N_11735,N_4770,N_5618);
nand U11736 (N_11736,N_5637,N_4365);
xnor U11737 (N_11737,N_7798,N_5181);
or U11738 (N_11738,N_6548,N_7882);
and U11739 (N_11739,N_6951,N_6126);
nand U11740 (N_11740,N_6326,N_7174);
and U11741 (N_11741,N_7594,N_6737);
nand U11742 (N_11742,N_5154,N_5624);
and U11743 (N_11743,N_4784,N_6976);
and U11744 (N_11744,N_5923,N_4633);
or U11745 (N_11745,N_4938,N_6506);
nor U11746 (N_11746,N_7449,N_5761);
nand U11747 (N_11747,N_5946,N_7520);
nand U11748 (N_11748,N_6894,N_6064);
xnor U11749 (N_11749,N_6484,N_7133);
or U11750 (N_11750,N_6143,N_6239);
nand U11751 (N_11751,N_5758,N_7974);
nand U11752 (N_11752,N_6621,N_6594);
nor U11753 (N_11753,N_6973,N_7673);
or U11754 (N_11754,N_4619,N_7583);
xor U11755 (N_11755,N_7000,N_6879);
xor U11756 (N_11756,N_4605,N_4252);
nor U11757 (N_11757,N_4110,N_4168);
xnor U11758 (N_11758,N_5407,N_4883);
nor U11759 (N_11759,N_4474,N_7717);
or U11760 (N_11760,N_6490,N_7997);
nor U11761 (N_11761,N_5443,N_4309);
nand U11762 (N_11762,N_5773,N_6388);
and U11763 (N_11763,N_7546,N_7044);
xor U11764 (N_11764,N_6263,N_5221);
and U11765 (N_11765,N_5343,N_7985);
xnor U11766 (N_11766,N_6795,N_6061);
and U11767 (N_11767,N_4660,N_4079);
or U11768 (N_11768,N_6719,N_6473);
xnor U11769 (N_11769,N_6250,N_4972);
and U11770 (N_11770,N_7290,N_7081);
nor U11771 (N_11771,N_5209,N_4244);
or U11772 (N_11772,N_6060,N_4225);
nor U11773 (N_11773,N_4287,N_6044);
nand U11774 (N_11774,N_6300,N_6920);
or U11775 (N_11775,N_6495,N_6656);
or U11776 (N_11776,N_7391,N_7451);
and U11777 (N_11777,N_5775,N_4045);
or U11778 (N_11778,N_6511,N_7808);
or U11779 (N_11779,N_6499,N_7965);
nor U11780 (N_11780,N_6845,N_5225);
nand U11781 (N_11781,N_7893,N_6109);
and U11782 (N_11782,N_4133,N_7888);
or U11783 (N_11783,N_5846,N_7054);
nand U11784 (N_11784,N_4541,N_7284);
xor U11785 (N_11785,N_6286,N_7123);
and U11786 (N_11786,N_7164,N_7714);
or U11787 (N_11787,N_5577,N_7234);
nor U11788 (N_11788,N_6329,N_5654);
and U11789 (N_11789,N_6885,N_4545);
and U11790 (N_11790,N_7921,N_5977);
nand U11791 (N_11791,N_4488,N_5373);
nor U11792 (N_11792,N_7901,N_6298);
xor U11793 (N_11793,N_5083,N_4957);
nand U11794 (N_11794,N_5893,N_5139);
and U11795 (N_11795,N_6360,N_6918);
or U11796 (N_11796,N_4627,N_7705);
or U11797 (N_11797,N_4064,N_4029);
nand U11798 (N_11798,N_6495,N_6839);
or U11799 (N_11799,N_7083,N_7945);
and U11800 (N_11800,N_6918,N_7770);
or U11801 (N_11801,N_4304,N_4057);
nor U11802 (N_11802,N_4951,N_6296);
nor U11803 (N_11803,N_6742,N_4928);
and U11804 (N_11804,N_6266,N_7349);
or U11805 (N_11805,N_6459,N_4786);
nor U11806 (N_11806,N_4208,N_7638);
nand U11807 (N_11807,N_7477,N_4139);
nor U11808 (N_11808,N_7581,N_4441);
and U11809 (N_11809,N_5205,N_6128);
nand U11810 (N_11810,N_4340,N_5719);
nand U11811 (N_11811,N_4070,N_6530);
nand U11812 (N_11812,N_6947,N_5795);
xor U11813 (N_11813,N_7983,N_6751);
nand U11814 (N_11814,N_7883,N_4005);
or U11815 (N_11815,N_7076,N_4139);
or U11816 (N_11816,N_7184,N_5207);
and U11817 (N_11817,N_4741,N_4059);
and U11818 (N_11818,N_4397,N_5631);
nand U11819 (N_11819,N_6736,N_6940);
xnor U11820 (N_11820,N_4016,N_5041);
or U11821 (N_11821,N_6968,N_5597);
nor U11822 (N_11822,N_7446,N_7548);
nand U11823 (N_11823,N_6242,N_4740);
or U11824 (N_11824,N_4574,N_5795);
or U11825 (N_11825,N_7177,N_6536);
or U11826 (N_11826,N_7298,N_6011);
or U11827 (N_11827,N_6517,N_4752);
xnor U11828 (N_11828,N_7749,N_7576);
nor U11829 (N_11829,N_6984,N_7207);
and U11830 (N_11830,N_4409,N_6738);
nor U11831 (N_11831,N_7830,N_6370);
nor U11832 (N_11832,N_4546,N_7935);
and U11833 (N_11833,N_5486,N_4485);
or U11834 (N_11834,N_6293,N_4898);
or U11835 (N_11835,N_5622,N_7385);
nand U11836 (N_11836,N_6841,N_4521);
nor U11837 (N_11837,N_7936,N_7432);
or U11838 (N_11838,N_6675,N_5095);
and U11839 (N_11839,N_6523,N_5982);
xnor U11840 (N_11840,N_5344,N_4437);
nor U11841 (N_11841,N_7186,N_7562);
or U11842 (N_11842,N_4814,N_4678);
and U11843 (N_11843,N_7725,N_4833);
xor U11844 (N_11844,N_4625,N_5777);
nor U11845 (N_11845,N_5752,N_6671);
nor U11846 (N_11846,N_5838,N_6387);
xnor U11847 (N_11847,N_7867,N_6204);
or U11848 (N_11848,N_4736,N_6226);
and U11849 (N_11849,N_4508,N_6839);
nor U11850 (N_11850,N_7349,N_5168);
nand U11851 (N_11851,N_5693,N_5837);
and U11852 (N_11852,N_5521,N_4767);
xor U11853 (N_11853,N_5020,N_7647);
nand U11854 (N_11854,N_4858,N_5032);
or U11855 (N_11855,N_4413,N_7498);
nor U11856 (N_11856,N_6866,N_7149);
xor U11857 (N_11857,N_7390,N_7767);
or U11858 (N_11858,N_4874,N_7437);
and U11859 (N_11859,N_7734,N_6573);
and U11860 (N_11860,N_6676,N_4527);
or U11861 (N_11861,N_5200,N_6344);
and U11862 (N_11862,N_6763,N_6085);
nand U11863 (N_11863,N_4614,N_6913);
or U11864 (N_11864,N_7286,N_4076);
or U11865 (N_11865,N_4653,N_6181);
or U11866 (N_11866,N_7614,N_5457);
xnor U11867 (N_11867,N_7992,N_5534);
xnor U11868 (N_11868,N_7996,N_4504);
nand U11869 (N_11869,N_6259,N_7073);
nor U11870 (N_11870,N_5090,N_5378);
or U11871 (N_11871,N_5210,N_7070);
or U11872 (N_11872,N_7964,N_4635);
and U11873 (N_11873,N_7972,N_5178);
nor U11874 (N_11874,N_5854,N_5614);
or U11875 (N_11875,N_4941,N_5243);
nor U11876 (N_11876,N_6707,N_6703);
and U11877 (N_11877,N_6519,N_5305);
nor U11878 (N_11878,N_5684,N_7152);
nand U11879 (N_11879,N_4571,N_6453);
and U11880 (N_11880,N_6377,N_5885);
nand U11881 (N_11881,N_6097,N_6458);
nand U11882 (N_11882,N_4905,N_4090);
or U11883 (N_11883,N_7136,N_7076);
nor U11884 (N_11884,N_7157,N_6856);
or U11885 (N_11885,N_4944,N_6539);
nor U11886 (N_11886,N_7303,N_7837);
nor U11887 (N_11887,N_4992,N_6111);
and U11888 (N_11888,N_4223,N_6884);
nor U11889 (N_11889,N_7931,N_6948);
xnor U11890 (N_11890,N_7207,N_7161);
xnor U11891 (N_11891,N_6575,N_7338);
and U11892 (N_11892,N_6515,N_6227);
xor U11893 (N_11893,N_6045,N_5165);
xnor U11894 (N_11894,N_6031,N_6681);
and U11895 (N_11895,N_6923,N_6443);
and U11896 (N_11896,N_6739,N_7618);
and U11897 (N_11897,N_5583,N_4610);
xor U11898 (N_11898,N_5874,N_6579);
nand U11899 (N_11899,N_6108,N_6293);
nand U11900 (N_11900,N_5980,N_4515);
nand U11901 (N_11901,N_4618,N_4417);
xor U11902 (N_11902,N_6673,N_5069);
and U11903 (N_11903,N_5037,N_6043);
or U11904 (N_11904,N_7961,N_4648);
nand U11905 (N_11905,N_5715,N_4000);
xnor U11906 (N_11906,N_5030,N_6038);
and U11907 (N_11907,N_6257,N_5651);
or U11908 (N_11908,N_5570,N_5797);
nor U11909 (N_11909,N_4787,N_7407);
or U11910 (N_11910,N_4452,N_4225);
xor U11911 (N_11911,N_4534,N_5342);
nand U11912 (N_11912,N_6200,N_4283);
or U11913 (N_11913,N_6255,N_6584);
nand U11914 (N_11914,N_4624,N_6743);
nor U11915 (N_11915,N_5370,N_5392);
nor U11916 (N_11916,N_4982,N_4123);
or U11917 (N_11917,N_4928,N_4497);
or U11918 (N_11918,N_4117,N_6613);
or U11919 (N_11919,N_4081,N_6856);
nor U11920 (N_11920,N_6005,N_6090);
nand U11921 (N_11921,N_6070,N_7427);
and U11922 (N_11922,N_7021,N_4393);
nand U11923 (N_11923,N_5994,N_4276);
or U11924 (N_11924,N_5732,N_7003);
nand U11925 (N_11925,N_5680,N_6990);
or U11926 (N_11926,N_7912,N_5612);
and U11927 (N_11927,N_7886,N_7269);
or U11928 (N_11928,N_7184,N_7492);
nand U11929 (N_11929,N_5579,N_6574);
nand U11930 (N_11930,N_4202,N_5909);
and U11931 (N_11931,N_6004,N_6471);
xnor U11932 (N_11932,N_6359,N_5316);
xnor U11933 (N_11933,N_7201,N_7523);
nand U11934 (N_11934,N_5286,N_4389);
and U11935 (N_11935,N_5256,N_6792);
or U11936 (N_11936,N_6867,N_7120);
nor U11937 (N_11937,N_6349,N_7690);
xnor U11938 (N_11938,N_6687,N_7057);
and U11939 (N_11939,N_4889,N_5241);
or U11940 (N_11940,N_5714,N_7749);
and U11941 (N_11941,N_5648,N_7926);
nor U11942 (N_11942,N_5108,N_6770);
or U11943 (N_11943,N_7077,N_5910);
and U11944 (N_11944,N_5123,N_5497);
or U11945 (N_11945,N_6922,N_6108);
and U11946 (N_11946,N_6392,N_5931);
and U11947 (N_11947,N_4962,N_7339);
nand U11948 (N_11948,N_4301,N_4950);
nand U11949 (N_11949,N_5909,N_4316);
nor U11950 (N_11950,N_4200,N_6159);
and U11951 (N_11951,N_6211,N_4775);
nand U11952 (N_11952,N_4541,N_6795);
xnor U11953 (N_11953,N_4628,N_4287);
xor U11954 (N_11954,N_6220,N_7005);
xnor U11955 (N_11955,N_6870,N_7481);
nor U11956 (N_11956,N_4633,N_4035);
nand U11957 (N_11957,N_4461,N_5774);
xor U11958 (N_11958,N_4021,N_5928);
nand U11959 (N_11959,N_7258,N_7993);
or U11960 (N_11960,N_7190,N_6600);
nand U11961 (N_11961,N_7058,N_4259);
nand U11962 (N_11962,N_5632,N_6923);
nor U11963 (N_11963,N_6137,N_6667);
and U11964 (N_11964,N_7015,N_6146);
nor U11965 (N_11965,N_5320,N_5782);
and U11966 (N_11966,N_4200,N_6538);
and U11967 (N_11967,N_7509,N_4169);
or U11968 (N_11968,N_4567,N_6296);
nor U11969 (N_11969,N_7423,N_7868);
nor U11970 (N_11970,N_6073,N_4689);
xor U11971 (N_11971,N_7666,N_6342);
nand U11972 (N_11972,N_4848,N_5566);
nor U11973 (N_11973,N_6070,N_5890);
or U11974 (N_11974,N_5845,N_4748);
and U11975 (N_11975,N_5819,N_7988);
nor U11976 (N_11976,N_6983,N_5647);
xnor U11977 (N_11977,N_4866,N_7994);
xnor U11978 (N_11978,N_5701,N_4435);
or U11979 (N_11979,N_7399,N_7871);
nor U11980 (N_11980,N_6961,N_5106);
xnor U11981 (N_11981,N_7778,N_5839);
and U11982 (N_11982,N_6355,N_5653);
nor U11983 (N_11983,N_5021,N_7871);
nand U11984 (N_11984,N_5652,N_5320);
or U11985 (N_11985,N_7211,N_5879);
nand U11986 (N_11986,N_6649,N_6546);
and U11987 (N_11987,N_4551,N_6746);
xnor U11988 (N_11988,N_4514,N_5108);
and U11989 (N_11989,N_7354,N_4446);
and U11990 (N_11990,N_6162,N_7712);
xnor U11991 (N_11991,N_5722,N_6432);
nand U11992 (N_11992,N_4509,N_6119);
xnor U11993 (N_11993,N_4293,N_7184);
nand U11994 (N_11994,N_4264,N_6874);
or U11995 (N_11995,N_6865,N_4636);
nor U11996 (N_11996,N_6911,N_6074);
xor U11997 (N_11997,N_7722,N_7708);
nor U11998 (N_11998,N_7239,N_6926);
or U11999 (N_11999,N_5752,N_5060);
nor U12000 (N_12000,N_9477,N_8030);
and U12001 (N_12001,N_9911,N_9654);
or U12002 (N_12002,N_8138,N_10808);
nor U12003 (N_12003,N_11446,N_8739);
nand U12004 (N_12004,N_11886,N_9525);
nor U12005 (N_12005,N_8359,N_10352);
nand U12006 (N_12006,N_10804,N_9956);
xnor U12007 (N_12007,N_9532,N_10276);
xnor U12008 (N_12008,N_8533,N_8613);
nor U12009 (N_12009,N_9621,N_10973);
or U12010 (N_12010,N_10245,N_10536);
xor U12011 (N_12011,N_9342,N_10111);
nand U12012 (N_12012,N_9830,N_11475);
xnor U12013 (N_12013,N_10786,N_8783);
xnor U12014 (N_12014,N_10794,N_10697);
and U12015 (N_12015,N_8190,N_9350);
and U12016 (N_12016,N_10300,N_10323);
and U12017 (N_12017,N_8235,N_8049);
and U12018 (N_12018,N_8832,N_10320);
xnor U12019 (N_12019,N_10223,N_11431);
and U12020 (N_12020,N_8699,N_8874);
or U12021 (N_12021,N_8590,N_10458);
and U12022 (N_12022,N_11250,N_10494);
nand U12023 (N_12023,N_11322,N_9708);
xnor U12024 (N_12024,N_9984,N_10184);
and U12025 (N_12025,N_10237,N_9707);
nor U12026 (N_12026,N_10366,N_8773);
and U12027 (N_12027,N_11303,N_10167);
xor U12028 (N_12028,N_10055,N_8144);
or U12029 (N_12029,N_9693,N_10698);
and U12030 (N_12030,N_8503,N_9294);
nor U12031 (N_12031,N_9838,N_8857);
or U12032 (N_12032,N_11672,N_11779);
xor U12033 (N_12033,N_11517,N_10066);
and U12034 (N_12034,N_9127,N_11048);
nor U12035 (N_12035,N_8114,N_9929);
xnor U12036 (N_12036,N_11414,N_8285);
xnor U12037 (N_12037,N_10068,N_9015);
and U12038 (N_12038,N_9107,N_8695);
and U12039 (N_12039,N_11413,N_11149);
nand U12040 (N_12040,N_11704,N_9326);
and U12041 (N_12041,N_10369,N_11646);
and U12042 (N_12042,N_10082,N_9455);
or U12043 (N_12043,N_11123,N_10283);
or U12044 (N_12044,N_10582,N_11072);
and U12045 (N_12045,N_11767,N_9320);
nand U12046 (N_12046,N_8646,N_9121);
or U12047 (N_12047,N_9970,N_9168);
and U12048 (N_12048,N_10307,N_11366);
nor U12049 (N_12049,N_9356,N_10824);
nand U12050 (N_12050,N_10641,N_9202);
nor U12051 (N_12051,N_9579,N_10752);
or U12052 (N_12052,N_11891,N_8703);
or U12053 (N_12053,N_11273,N_9007);
or U12054 (N_12054,N_9146,N_8764);
nand U12055 (N_12055,N_9427,N_8504);
and U12056 (N_12056,N_10972,N_11068);
or U12057 (N_12057,N_10190,N_10810);
and U12058 (N_12058,N_11144,N_9275);
nand U12059 (N_12059,N_8345,N_11329);
or U12060 (N_12060,N_9233,N_8330);
or U12061 (N_12061,N_9059,N_8328);
and U12062 (N_12062,N_10646,N_10478);
nand U12063 (N_12063,N_11998,N_9507);
xor U12064 (N_12064,N_11391,N_11463);
or U12065 (N_12065,N_9804,N_11674);
or U12066 (N_12066,N_10056,N_8928);
or U12067 (N_12067,N_8844,N_10001);
or U12068 (N_12068,N_10971,N_10875);
and U12069 (N_12069,N_11778,N_9623);
nand U12070 (N_12070,N_8333,N_9467);
xor U12071 (N_12071,N_11138,N_8270);
or U12072 (N_12072,N_11980,N_10687);
xor U12073 (N_12073,N_9663,N_9600);
and U12074 (N_12074,N_10654,N_10774);
nor U12075 (N_12075,N_8602,N_11938);
nand U12076 (N_12076,N_8553,N_11612);
nand U12077 (N_12077,N_9296,N_8212);
xnor U12078 (N_12078,N_10628,N_11400);
or U12079 (N_12079,N_10147,N_10756);
and U12080 (N_12080,N_10400,N_8506);
nand U12081 (N_12081,N_8236,N_8472);
and U12082 (N_12082,N_10094,N_10793);
or U12083 (N_12083,N_9229,N_8203);
or U12084 (N_12084,N_11529,N_10685);
nand U12085 (N_12085,N_8195,N_9259);
nand U12086 (N_12086,N_11814,N_9983);
xor U12087 (N_12087,N_11963,N_10541);
xor U12088 (N_12088,N_9496,N_8916);
xnor U12089 (N_12089,N_11701,N_8591);
nor U12090 (N_12090,N_8241,N_11520);
xor U12091 (N_12091,N_9826,N_9158);
nand U12092 (N_12092,N_10806,N_9411);
nor U12093 (N_12093,N_11900,N_10014);
and U12094 (N_12094,N_11757,N_9875);
xnor U12095 (N_12095,N_8932,N_8186);
and U12096 (N_12096,N_9499,N_11683);
nand U12097 (N_12097,N_11765,N_10045);
nor U12098 (N_12098,N_8197,N_10749);
or U12099 (N_12099,N_8470,N_10043);
nor U12100 (N_12100,N_8765,N_10615);
nor U12101 (N_12101,N_10613,N_10269);
or U12102 (N_12102,N_10809,N_11733);
nand U12103 (N_12103,N_9814,N_9057);
nor U12104 (N_12104,N_8015,N_8223);
nand U12105 (N_12105,N_10538,N_11602);
nor U12106 (N_12106,N_10943,N_11562);
nor U12107 (N_12107,N_10069,N_11309);
xor U12108 (N_12108,N_11226,N_11533);
xnor U12109 (N_12109,N_8657,N_8277);
nand U12110 (N_12110,N_10939,N_11164);
xor U12111 (N_12111,N_10290,N_11764);
or U12112 (N_12112,N_8700,N_10493);
xnor U12113 (N_12113,N_8656,N_10181);
xnor U12114 (N_12114,N_9094,N_8122);
xor U12115 (N_12115,N_10399,N_10206);
xnor U12116 (N_12116,N_8670,N_10472);
or U12117 (N_12117,N_9381,N_9246);
nor U12118 (N_12118,N_9243,N_10829);
nor U12119 (N_12119,N_8158,N_9771);
and U12120 (N_12120,N_8774,N_10408);
xor U12121 (N_12121,N_10149,N_9068);
xnor U12122 (N_12122,N_9918,N_11402);
and U12123 (N_12123,N_11357,N_11990);
and U12124 (N_12124,N_11324,N_9919);
nor U12125 (N_12125,N_9188,N_11595);
xor U12126 (N_12126,N_9250,N_11544);
and U12127 (N_12127,N_11023,N_8704);
nor U12128 (N_12128,N_8856,N_9831);
nor U12129 (N_12129,N_11464,N_10643);
xor U12130 (N_12130,N_9644,N_11842);
nand U12131 (N_12131,N_9159,N_9374);
nand U12132 (N_12132,N_11537,N_10311);
nand U12133 (N_12133,N_10508,N_8334);
and U12134 (N_12134,N_10414,N_8685);
and U12135 (N_12135,N_8967,N_10632);
nand U12136 (N_12136,N_8040,N_11394);
xnor U12137 (N_12137,N_8130,N_8389);
or U12138 (N_12138,N_8770,N_8641);
and U12139 (N_12139,N_8425,N_9049);
nor U12140 (N_12140,N_11477,N_10105);
nor U12141 (N_12141,N_11699,N_10688);
and U12142 (N_12142,N_11925,N_8775);
xor U12143 (N_12143,N_9548,N_9536);
xnor U12144 (N_12144,N_9131,N_9828);
xnor U12145 (N_12145,N_11777,N_8527);
and U12146 (N_12146,N_11165,N_8034);
and U12147 (N_12147,N_9797,N_10337);
and U12148 (N_12148,N_8023,N_9030);
xnor U12149 (N_12149,N_9054,N_11540);
nor U12150 (N_12150,N_11791,N_11307);
xnor U12151 (N_12151,N_10821,N_9387);
nand U12152 (N_12152,N_9223,N_9558);
and U12153 (N_12153,N_11830,N_11975);
nand U12154 (N_12154,N_10521,N_8500);
and U12155 (N_12155,N_10452,N_10722);
xnor U12156 (N_12156,N_11272,N_9475);
nand U12157 (N_12157,N_11535,N_9098);
nand U12158 (N_12158,N_9530,N_8315);
xor U12159 (N_12159,N_10898,N_8464);
and U12160 (N_12160,N_9369,N_11241);
nor U12161 (N_12161,N_9907,N_10405);
and U12162 (N_12162,N_8925,N_10780);
nor U12163 (N_12163,N_8202,N_10222);
or U12164 (N_12164,N_11043,N_11255);
nor U12165 (N_12165,N_9994,N_9459);
xnor U12166 (N_12166,N_9000,N_11770);
and U12167 (N_12167,N_10227,N_8970);
xnor U12168 (N_12168,N_8788,N_8038);
and U12169 (N_12169,N_11092,N_11417);
nor U12170 (N_12170,N_11404,N_10189);
and U12171 (N_12171,N_9930,N_11542);
or U12172 (N_12172,N_10463,N_10611);
and U12173 (N_12173,N_11706,N_8213);
xor U12174 (N_12174,N_9478,N_11343);
or U12175 (N_12175,N_11775,N_10371);
nand U12176 (N_12176,N_9314,N_10612);
xor U12177 (N_12177,N_9402,N_8511);
nand U12178 (N_12178,N_8907,N_9239);
xnor U12179 (N_12179,N_10980,N_10107);
nor U12180 (N_12180,N_11368,N_8361);
xnor U12181 (N_12181,N_9864,N_10777);
and U12182 (N_12182,N_10339,N_9563);
nand U12183 (N_12183,N_9572,N_9135);
nand U12184 (N_12184,N_9393,N_11205);
and U12185 (N_12185,N_9965,N_8754);
and U12186 (N_12186,N_11292,N_11982);
nand U12187 (N_12187,N_8892,N_8601);
and U12188 (N_12188,N_9438,N_8674);
and U12189 (N_12189,N_9612,N_9975);
xnor U12190 (N_12190,N_11330,N_8609);
nand U12191 (N_12191,N_8742,N_10140);
or U12192 (N_12192,N_10594,N_8480);
nor U12193 (N_12193,N_9647,N_10090);
nand U12194 (N_12194,N_9792,N_8939);
nor U12195 (N_12195,N_9340,N_11953);
xor U12196 (N_12196,N_11739,N_11481);
nor U12197 (N_12197,N_11689,N_11457);
and U12198 (N_12198,N_8363,N_11182);
or U12199 (N_12199,N_10575,N_8148);
xnor U12200 (N_12200,N_8006,N_8082);
nand U12201 (N_12201,N_11424,N_9473);
or U12202 (N_12202,N_9577,N_11580);
nand U12203 (N_12203,N_9271,N_10555);
nand U12204 (N_12204,N_10755,N_9470);
nand U12205 (N_12205,N_8914,N_11937);
nor U12206 (N_12206,N_10878,N_11768);
and U12207 (N_12207,N_9101,N_10087);
xnor U12208 (N_12208,N_9145,N_8753);
nor U12209 (N_12209,N_10827,N_8465);
nor U12210 (N_12210,N_9784,N_11118);
or U12211 (N_12211,N_11808,N_8991);
xnor U12212 (N_12212,N_8147,N_11628);
and U12213 (N_12213,N_9901,N_11419);
xnor U12214 (N_12214,N_8043,N_8638);
nand U12215 (N_12215,N_8273,N_9443);
xnor U12216 (N_12216,N_10299,N_9856);
nand U12217 (N_12217,N_10424,N_9531);
nand U12218 (N_12218,N_9685,N_8296);
nor U12219 (N_12219,N_11145,N_8721);
or U12220 (N_12220,N_10692,N_9768);
nor U12221 (N_12221,N_11684,N_11895);
and U12222 (N_12222,N_8937,N_10077);
xor U12223 (N_12223,N_8650,N_9781);
nand U12224 (N_12224,N_9916,N_8085);
and U12225 (N_12225,N_8278,N_11676);
and U12226 (N_12226,N_11934,N_10762);
nor U12227 (N_12227,N_8708,N_10266);
nand U12228 (N_12228,N_10250,N_11455);
nor U12229 (N_12229,N_11142,N_11609);
nand U12230 (N_12230,N_9697,N_8749);
nand U12231 (N_12231,N_10433,N_8189);
nor U12232 (N_12232,N_9153,N_11451);
and U12233 (N_12233,N_11390,N_11279);
xor U12234 (N_12234,N_10524,N_11319);
nor U12235 (N_12235,N_11162,N_8099);
nand U12236 (N_12236,N_10434,N_9723);
and U12237 (N_12237,N_8476,N_11723);
xor U12238 (N_12238,N_9026,N_9656);
or U12239 (N_12239,N_9328,N_8672);
xnor U12240 (N_12240,N_11984,N_10955);
and U12241 (N_12241,N_8945,N_9757);
nor U12242 (N_12242,N_8073,N_9086);
and U12243 (N_12243,N_10454,N_11783);
xnor U12244 (N_12244,N_10409,N_8319);
nand U12245 (N_12245,N_9946,N_8522);
nor U12246 (N_12246,N_9292,N_9016);
nor U12247 (N_12247,N_8473,N_8793);
xnor U12248 (N_12248,N_11835,N_10715);
and U12249 (N_12249,N_10159,N_11927);
or U12250 (N_12250,N_8912,N_9075);
nor U12251 (N_12251,N_9509,N_11868);
nand U12252 (N_12252,N_8630,N_10543);
xnor U12253 (N_12253,N_10258,N_8179);
xnor U12254 (N_12254,N_8649,N_10637);
nand U12255 (N_12255,N_10835,N_10221);
nand U12256 (N_12256,N_11751,N_8289);
nor U12257 (N_12257,N_9779,N_9706);
and U12258 (N_12258,N_10681,N_8899);
nand U12259 (N_12259,N_10909,N_10744);
or U12260 (N_12260,N_9542,N_11894);
xor U12261 (N_12261,N_9872,N_8654);
and U12262 (N_12262,N_10616,N_8563);
xnor U12263 (N_12263,N_11734,N_11902);
nor U12264 (N_12264,N_9047,N_8283);
nor U12265 (N_12265,N_9002,N_8012);
xnor U12266 (N_12266,N_9841,N_10492);
nand U12267 (N_12267,N_8255,N_11872);
nor U12268 (N_12268,N_11240,N_11582);
xnor U12269 (N_12269,N_11590,N_9554);
nand U12270 (N_12270,N_11386,N_11572);
and U12271 (N_12271,N_10041,N_9192);
nor U12272 (N_12272,N_11556,N_9187);
nand U12273 (N_12273,N_10818,N_9742);
or U12274 (N_12274,N_11664,N_11642);
and U12275 (N_12275,N_9601,N_9245);
xnor U12276 (N_12276,N_9373,N_9799);
or U12277 (N_12277,N_8702,N_10195);
nand U12278 (N_12278,N_10747,N_8933);
or U12279 (N_12279,N_8083,N_8784);
xor U12280 (N_12280,N_11470,N_8767);
nor U12281 (N_12281,N_10247,N_10280);
nand U12282 (N_12282,N_11126,N_9767);
and U12283 (N_12283,N_8824,N_8370);
nor U12284 (N_12284,N_9576,N_8399);
and U12285 (N_12285,N_8194,N_8575);
xor U12286 (N_12286,N_8528,N_8436);
nand U12287 (N_12287,N_11211,N_9186);
nor U12288 (N_12288,N_10015,N_8410);
and U12289 (N_12289,N_8295,N_10870);
or U12290 (N_12290,N_11379,N_11482);
nand U12291 (N_12291,N_10882,N_10071);
or U12292 (N_12292,N_8926,N_11013);
nand U12293 (N_12293,N_9746,N_8694);
nor U12294 (N_12294,N_8965,N_10095);
xor U12295 (N_12295,N_9898,N_8141);
xor U12296 (N_12296,N_8380,N_9204);
or U12297 (N_12297,N_10378,N_10602);
and U12298 (N_12298,N_11163,N_8176);
nand U12299 (N_12299,N_9801,N_8584);
nor U12300 (N_12300,N_11547,N_11552);
or U12301 (N_12301,N_8438,N_11971);
and U12302 (N_12302,N_8351,N_11685);
nand U12303 (N_12303,N_8080,N_11131);
nand U12304 (N_12304,N_8948,N_8797);
and U12305 (N_12305,N_9604,N_11921);
nor U12306 (N_12306,N_8651,N_10451);
or U12307 (N_12307,N_10481,N_8297);
xor U12308 (N_12308,N_10032,N_9912);
nor U12309 (N_12309,N_10441,N_11452);
or U12310 (N_12310,N_8632,N_10552);
xnor U12311 (N_12311,N_9266,N_9691);
nor U12312 (N_12312,N_9696,N_11541);
or U12313 (N_12313,N_11172,N_9811);
nand U12314 (N_12314,N_9070,N_9191);
and U12315 (N_12315,N_11864,N_8011);
and U12316 (N_12316,N_11978,N_11467);
nand U12317 (N_12317,N_10607,N_9646);
xnor U12318 (N_12318,N_10800,N_8055);
xnor U12319 (N_12319,N_8227,N_9555);
nor U12320 (N_12320,N_8730,N_8863);
or U12321 (N_12321,N_9458,N_9425);
nor U12322 (N_12322,N_11443,N_9931);
xnor U12323 (N_12323,N_9333,N_10178);
xnor U12324 (N_12324,N_8963,N_11784);
nor U12325 (N_12325,N_9991,N_8451);
xor U12326 (N_12326,N_8495,N_9766);
nor U12327 (N_12327,N_9113,N_8725);
and U12328 (N_12328,N_10872,N_8454);
nor U12329 (N_12329,N_11619,N_9439);
nor U12330 (N_12330,N_11857,N_9545);
and U12331 (N_12331,N_11675,N_10830);
and U12332 (N_12332,N_9658,N_10881);
xor U12333 (N_12333,N_9018,N_9743);
nand U12334 (N_12334,N_10557,N_11846);
xnor U12335 (N_12335,N_10765,N_11371);
nand U12336 (N_12336,N_9132,N_10288);
nor U12337 (N_12337,N_10461,N_10631);
or U12338 (N_12338,N_11854,N_10998);
nor U12339 (N_12339,N_8384,N_9943);
and U12340 (N_12340,N_11466,N_10305);
xnor U12341 (N_12341,N_11209,N_8185);
nand U12342 (N_12342,N_10229,N_8004);
nand U12343 (N_12343,N_10207,N_9090);
nand U12344 (N_12344,N_11663,N_9594);
nand U12345 (N_12345,N_10623,N_8393);
or U12346 (N_12346,N_9344,N_10131);
or U12347 (N_12347,N_11640,N_10025);
nand U12348 (N_12348,N_9005,N_9632);
xnor U12349 (N_12349,N_11922,N_9605);
nand U12350 (N_12350,N_10334,N_9974);
or U12351 (N_12351,N_11432,N_11084);
xor U12352 (N_12352,N_11037,N_8002);
and U12353 (N_12353,N_10532,N_10263);
nor U12354 (N_12354,N_8348,N_10328);
nand U12355 (N_12355,N_11603,N_8516);
and U12356 (N_12356,N_9653,N_9861);
or U12357 (N_12357,N_8175,N_10185);
xor U12358 (N_12358,N_9992,N_10338);
nand U12359 (N_12359,N_10460,N_9206);
or U12360 (N_12360,N_9445,N_10315);
or U12361 (N_12361,N_9669,N_11360);
nand U12362 (N_12362,N_8752,N_9041);
nor U12363 (N_12363,N_11096,N_8132);
nor U12364 (N_12364,N_8673,N_10389);
xnor U12365 (N_12365,N_10136,N_9451);
and U12366 (N_12366,N_10439,N_11492);
nand U12367 (N_12367,N_10480,N_8758);
or U12368 (N_12368,N_9392,N_8940);
nand U12369 (N_12369,N_11009,N_9379);
and U12370 (N_12370,N_8645,N_11016);
or U12371 (N_12371,N_10942,N_8806);
nand U12372 (N_12372,N_9407,N_10891);
nor U12373 (N_12373,N_11625,N_11183);
or U12374 (N_12374,N_9595,N_11742);
nor U12375 (N_12375,N_10385,N_8054);
nand U12376 (N_12376,N_10841,N_9009);
or U12377 (N_12377,N_9715,N_10811);
or U12378 (N_12378,N_10767,N_9276);
nor U12379 (N_12379,N_9376,N_9598);
xor U12380 (N_12380,N_10349,N_9520);
or U12381 (N_12381,N_9985,N_9815);
or U12382 (N_12382,N_10781,N_8312);
nand U12383 (N_12383,N_10908,N_8231);
nor U12384 (N_12384,N_10076,N_10255);
xor U12385 (N_12385,N_10495,N_11313);
nor U12386 (N_12386,N_8534,N_9808);
nand U12387 (N_12387,N_8885,N_10825);
nor U12388 (N_12388,N_8184,N_9463);
and U12389 (N_12389,N_8385,N_10332);
or U12390 (N_12390,N_8412,N_9544);
xor U12391 (N_12391,N_11323,N_8072);
nor U12392 (N_12392,N_9888,N_10970);
and U12393 (N_12393,N_11063,N_10547);
nor U12394 (N_12394,N_11066,N_11352);
xnor U12395 (N_12395,N_10108,N_8424);
and U12396 (N_12396,N_10198,N_11245);
nand U12397 (N_12397,N_8403,N_9152);
nand U12398 (N_12398,N_10992,N_11383);
and U12399 (N_12399,N_10587,N_10933);
nor U12400 (N_12400,N_10644,N_9701);
nor U12401 (N_12401,N_8274,N_8572);
nor U12402 (N_12402,N_9747,N_10106);
nand U12403 (N_12403,N_11546,N_9378);
nand U12404 (N_12404,N_11782,N_9065);
and U12405 (N_12405,N_9011,N_10191);
or U12406 (N_12406,N_10924,N_9251);
nor U12407 (N_12407,N_10469,N_11000);
and U12408 (N_12408,N_11363,N_8620);
or U12409 (N_12409,N_8779,N_8124);
and U12410 (N_12410,N_10026,N_10516);
nand U12411 (N_12411,N_11844,N_8787);
nor U12412 (N_12412,N_10626,N_9112);
nand U12413 (N_12413,N_8876,N_8986);
and U12414 (N_12414,N_9692,N_9926);
nor U12415 (N_12415,N_8173,N_8756);
or U12416 (N_12416,N_8057,N_8873);
or U12417 (N_12417,N_9556,N_11416);
xnor U12418 (N_12418,N_10329,N_11244);
xor U12419 (N_12419,N_9236,N_10622);
or U12420 (N_12420,N_10520,N_8120);
and U12421 (N_12421,N_8335,N_11650);
xnor U12422 (N_12422,N_10121,N_11003);
nor U12423 (N_12423,N_8959,N_8938);
or U12424 (N_12424,N_9226,N_10265);
xor U12425 (N_12425,N_9010,N_11662);
or U12426 (N_12426,N_9116,N_11997);
xor U12427 (N_12427,N_10267,N_8008);
xnor U12428 (N_12428,N_8468,N_9966);
nor U12429 (N_12429,N_9960,N_11382);
and U12430 (N_12430,N_8430,N_9321);
xnor U12431 (N_12431,N_8628,N_11461);
or U12432 (N_12432,N_10270,N_10444);
xor U12433 (N_12433,N_10850,N_9834);
xor U12434 (N_12434,N_11175,N_10843);
nand U12435 (N_12435,N_11206,N_10540);
or U12436 (N_12436,N_9104,N_9675);
nor U12437 (N_12437,N_9248,N_8751);
or U12438 (N_12438,N_11132,N_10148);
nand U12439 (N_12439,N_11150,N_8492);
nand U12440 (N_12440,N_11358,N_11333);
nand U12441 (N_12441,N_9428,N_10348);
xnor U12442 (N_12442,N_11690,N_10655);
nand U12443 (N_12443,N_8760,N_8401);
nor U12444 (N_12444,N_8368,N_10736);
and U12445 (N_12445,N_9616,N_8371);
and U12446 (N_12446,N_9031,N_11034);
nand U12447 (N_12447,N_11302,N_10502);
and U12448 (N_12448,N_11201,N_11283);
or U12449 (N_12449,N_10391,N_8096);
nor U12450 (N_12450,N_10930,N_11756);
nor U12451 (N_12451,N_8538,N_8982);
xor U12452 (N_12452,N_11137,N_9606);
nor U12453 (N_12453,N_9882,N_10836);
nand U12454 (N_12454,N_11944,N_9414);
xnor U12455 (N_12455,N_8587,N_10231);
nand U12456 (N_12456,N_11850,N_11881);
xor U12457 (N_12457,N_10138,N_11353);
xnor U12458 (N_12458,N_10062,N_11247);
and U12459 (N_12459,N_11823,N_10497);
and U12460 (N_12460,N_10928,N_10487);
xor U12461 (N_12461,N_11671,N_11010);
or U12462 (N_12462,N_10274,N_11280);
and U12463 (N_12463,N_11729,N_8629);
nor U12464 (N_12464,N_9777,N_9704);
xnor U12465 (N_12465,N_8518,N_8855);
nand U12466 (N_12466,N_11213,N_11061);
xnor U12467 (N_12467,N_8759,N_10426);
nand U12468 (N_12468,N_8485,N_11920);
or U12469 (N_12469,N_8053,N_9357);
nor U12470 (N_12470,N_8160,N_9590);
nor U12471 (N_12471,N_9674,N_10717);
nor U12472 (N_12472,N_9717,N_8137);
xor U12473 (N_12473,N_9114,N_11809);
nor U12474 (N_12474,N_10847,N_9617);
and U12475 (N_12475,N_11418,N_9752);
and U12476 (N_12476,N_10900,N_11833);
or U12477 (N_12477,N_11763,N_10669);
and U12478 (N_12478,N_9263,N_9868);
nor U12479 (N_12479,N_11026,N_10565);
xor U12480 (N_12480,N_8108,N_11393);
and U12481 (N_12481,N_8417,N_10416);
xnor U12482 (N_12482,N_10115,N_8847);
and U12483 (N_12483,N_11566,N_9079);
or U12484 (N_12484,N_8905,N_9137);
or U12485 (N_12485,N_9761,N_10982);
nor U12486 (N_12486,N_10620,N_11698);
and U12487 (N_12487,N_11038,N_10505);
nand U12488 (N_12488,N_8852,N_8551);
or U12489 (N_12489,N_9111,N_9267);
or U12490 (N_12490,N_8092,N_9178);
and U12491 (N_12491,N_10395,N_8955);
xnor U12492 (N_12492,N_8155,N_9535);
or U12493 (N_12493,N_9115,N_9077);
xor U12494 (N_12494,N_11665,N_8068);
nor U12495 (N_12495,N_11267,N_9679);
or U12496 (N_12496,N_9909,N_9798);
nand U12497 (N_12497,N_11011,N_8850);
xnor U12498 (N_12498,N_11204,N_8036);
or U12499 (N_12499,N_10696,N_10008);
or U12500 (N_12500,N_9441,N_9643);
xor U12501 (N_12501,N_11217,N_11306);
and U12502 (N_12502,N_10559,N_11364);
nand U12503 (N_12503,N_8881,N_11233);
and U12504 (N_12504,N_11125,N_9698);
nor U12505 (N_12505,N_8691,N_9652);
or U12506 (N_12506,N_8306,N_8254);
nor U12507 (N_12507,N_10913,N_9769);
and U12508 (N_12508,N_10238,N_8104);
or U12509 (N_12509,N_8688,N_10445);
nand U12510 (N_12510,N_11522,N_10009);
nand U12511 (N_12511,N_11993,N_9958);
nand U12512 (N_12512,N_10914,N_11928);
nor U12513 (N_12513,N_11679,N_8327);
xnor U12514 (N_12514,N_9859,N_10498);
nand U12515 (N_12515,N_10635,N_9687);
nor U12516 (N_12516,N_11696,N_11870);
nand U12517 (N_12517,N_10618,N_9863);
nand U12518 (N_12518,N_8462,N_8118);
or U12519 (N_12519,N_11827,N_8596);
nor U12520 (N_12520,N_8619,N_11472);
or U12521 (N_12521,N_8693,N_9124);
xnor U12522 (N_12522,N_10118,N_9689);
and U12523 (N_12523,N_11780,N_8958);
nor U12524 (N_12524,N_8149,N_10513);
nor U12525 (N_12525,N_11143,N_9963);
nor U12526 (N_12526,N_10172,N_10740);
and U12527 (N_12527,N_11456,N_10325);
nand U12528 (N_12528,N_10394,N_8253);
xnor U12529 (N_12529,N_9227,N_9899);
and U12530 (N_12530,N_9607,N_8031);
nor U12531 (N_12531,N_10336,N_10650);
xnor U12532 (N_12532,N_11715,N_10479);
and U12533 (N_12533,N_9361,N_8887);
or U12534 (N_12534,N_11331,N_8458);
or U12535 (N_12535,N_8561,N_8383);
nand U12536 (N_12536,N_10950,N_11627);
and U12537 (N_12537,N_9222,N_9313);
and U12538 (N_12538,N_8279,N_9497);
xor U12539 (N_12539,N_10868,N_11802);
nand U12540 (N_12540,N_11304,N_11055);
or U12541 (N_12541,N_11995,N_11224);
xor U12542 (N_12542,N_10851,N_9712);
and U12543 (N_12543,N_11519,N_10564);
nand U12544 (N_12544,N_11709,N_10573);
nor U12545 (N_12545,N_8117,N_8557);
and U12546 (N_12546,N_8994,N_9614);
xnor U12547 (N_12547,N_11570,N_8408);
and U12548 (N_12548,N_11600,N_9372);
nand U12549 (N_12549,N_10608,N_10219);
nor U12550 (N_12550,N_10303,N_11258);
nor U12551 (N_12551,N_9209,N_8224);
nor U12552 (N_12552,N_10122,N_9048);
nand U12553 (N_12553,N_10456,N_9613);
nor U12554 (N_12554,N_8187,N_8342);
and U12555 (N_12555,N_11579,N_9422);
nand U12556 (N_12556,N_11766,N_10940);
and U12557 (N_12557,N_8828,N_9396);
and U12558 (N_12558,N_10029,N_10934);
and U12559 (N_12559,N_9329,N_10035);
nor U12560 (N_12560,N_11889,N_10296);
nand U12561 (N_12561,N_11605,N_8623);
and U12562 (N_12562,N_11940,N_10278);
nor U12563 (N_12563,N_8105,N_11238);
and U12564 (N_12564,N_9805,N_10537);
nand U12565 (N_12565,N_8696,N_8299);
xnor U12566 (N_12566,N_11644,N_11342);
and U12567 (N_12567,N_8192,N_11395);
or U12568 (N_12568,N_11356,N_9274);
and U12569 (N_12569,N_10983,N_10096);
or U12570 (N_12570,N_11588,N_10862);
nand U12571 (N_12571,N_9775,N_9920);
nand U12572 (N_12572,N_8125,N_10621);
nand U12573 (N_12573,N_8772,N_10586);
xnor U12574 (N_12574,N_9190,N_9234);
nand U12575 (N_12575,N_9662,N_8210);
xnor U12576 (N_12576,N_10533,N_9793);
and U12577 (N_12577,N_11473,N_8367);
nand U12578 (N_12578,N_9773,N_8512);
xor U12579 (N_12579,N_8890,N_11133);
or U12580 (N_12580,N_11598,N_8448);
nor U12581 (N_12581,N_8423,N_10570);
nand U12582 (N_12582,N_11212,N_11177);
or U12583 (N_12583,N_8726,N_8323);
or U12584 (N_12584,N_9353,N_9363);
nand U12585 (N_12585,N_8428,N_9574);
or U12586 (N_12586,N_9733,N_9491);
and U12587 (N_12587,N_10387,N_8497);
nor U12588 (N_12588,N_8329,N_10944);
and U12589 (N_12589,N_10033,N_11029);
and U12590 (N_12590,N_9889,N_11661);
and U12591 (N_12591,N_9207,N_10874);
xnor U12592 (N_12592,N_10135,N_11067);
nor U12593 (N_12593,N_8801,N_11559);
nor U12594 (N_12594,N_8079,N_11667);
and U12595 (N_12595,N_11405,N_10588);
nand U12596 (N_12596,N_10291,N_10302);
and U12597 (N_12597,N_10584,N_8262);
nor U12598 (N_12598,N_10085,N_9256);
nand U12599 (N_12599,N_8435,N_9599);
and U12600 (N_12600,N_9238,N_9684);
nor U12601 (N_12601,N_8305,N_9624);
and U12602 (N_12602,N_10488,N_8390);
nor U12603 (N_12603,N_11514,N_11959);
xor U12604 (N_12604,N_8156,N_8456);
nand U12605 (N_12605,N_8027,N_11508);
xor U12606 (N_12606,N_11086,N_8833);
xnor U12607 (N_12607,N_11191,N_10163);
nor U12608 (N_12608,N_9748,N_10511);
and U12609 (N_12609,N_11707,N_11019);
xnor U12610 (N_12610,N_11635,N_10817);
xnor U12611 (N_12611,N_10853,N_11490);
nand U12612 (N_12612,N_10335,N_10246);
or U12613 (N_12613,N_11741,N_8415);
or U12614 (N_12614,N_11597,N_8745);
nor U12615 (N_12615,N_9914,N_10088);
nor U12616 (N_12616,N_11750,N_10945);
nor U12617 (N_12617,N_10840,N_9044);
xor U12618 (N_12618,N_10432,N_11274);
and U12619 (N_12619,N_10925,N_8338);
and U12620 (N_12620,N_9833,N_9409);
or U12621 (N_12621,N_10380,N_11896);
or U12622 (N_12622,N_9620,N_8675);
and U12623 (N_12623,N_11392,N_11311);
nor U12624 (N_12624,N_10012,N_10176);
or U12625 (N_12625,N_9050,N_9479);
xor U12626 (N_12626,N_11847,N_8444);
or U12627 (N_12627,N_11560,N_8523);
or U12628 (N_12628,N_8063,N_11745);
nor U12629 (N_12629,N_11495,N_11315);
nand U12630 (N_12630,N_11314,N_10214);
nor U12631 (N_12631,N_9802,N_10504);
or U12632 (N_12632,N_11688,N_8529);
nand U12633 (N_12633,N_11349,N_8232);
xnor U12634 (N_12634,N_10425,N_9330);
and U12635 (N_12635,N_10556,N_11500);
or U12636 (N_12636,N_10218,N_8550);
xor U12637 (N_12637,N_9442,N_10331);
nor U12638 (N_12638,N_11981,N_11972);
and U12639 (N_12639,N_9847,N_11929);
nor U12640 (N_12640,N_11912,N_11115);
nand U12641 (N_12641,N_11090,N_9205);
nand U12642 (N_12642,N_8634,N_10802);
or U12643 (N_12643,N_8103,N_8505);
and U12644 (N_12644,N_8720,N_8123);
and U12645 (N_12645,N_10558,N_11565);
nand U12646 (N_12646,N_9144,N_8349);
nand U12647 (N_12647,N_10730,N_10151);
and U12648 (N_12648,N_11873,N_8067);
nor U12649 (N_12649,N_9118,N_9628);
or U12650 (N_12650,N_9823,N_10298);
nor U12651 (N_12651,N_11269,N_8951);
or U12652 (N_12652,N_8269,N_11636);
nor U12653 (N_12653,N_10053,N_10473);
and U12654 (N_12654,N_10030,N_10897);
nand U12655 (N_12655,N_8616,N_10625);
nand U12656 (N_12656,N_11797,N_9254);
and U12657 (N_12657,N_8286,N_11278);
or U12658 (N_12658,N_10022,N_9857);
xnor U12659 (N_12659,N_9244,N_10061);
xor U12660 (N_12660,N_9588,N_10926);
or U12661 (N_12661,N_9272,N_9462);
or U12662 (N_12662,N_8280,N_8519);
nor U12663 (N_12663,N_9584,N_8019);
xnor U12664 (N_12664,N_9456,N_9786);
or U12665 (N_12665,N_8029,N_11397);
nand U12666 (N_12666,N_8261,N_11151);
nand U12667 (N_12667,N_11248,N_8795);
nor U12668 (N_12668,N_9673,N_9703);
xnor U12669 (N_12669,N_8585,N_9560);
xnor U12670 (N_12670,N_8732,N_8025);
xnor U12671 (N_12671,N_8291,N_11488);
nand U12672 (N_12672,N_9877,N_11321);
nand U12673 (N_12673,N_10049,N_11079);
nor U12674 (N_12674,N_10097,N_11007);
and U12675 (N_12675,N_9288,N_9106);
nor U12676 (N_12676,N_10915,N_9933);
and U12677 (N_12677,N_9928,N_8701);
nor U12678 (N_12678,N_11040,N_11139);
nor U12679 (N_12679,N_9695,N_11948);
xnor U12680 (N_12680,N_9890,N_11532);
and U12681 (N_12681,N_9283,N_8331);
nand U12682 (N_12682,N_11480,N_11285);
nor U12683 (N_12683,N_11989,N_8134);
nor U12684 (N_12684,N_8898,N_8740);
and U12685 (N_12685,N_11649,N_9141);
or U12686 (N_12686,N_10124,N_10719);
or U12687 (N_12687,N_8178,N_9610);
and U12688 (N_12688,N_8757,N_9770);
or U12689 (N_12689,N_10450,N_8169);
nand U12690 (N_12690,N_9690,N_9518);
xor U12691 (N_12691,N_9935,N_10393);
nor U12692 (N_12692,N_9506,N_11262);
xnor U12693 (N_12693,N_10392,N_11259);
or U12694 (N_12694,N_8163,N_10419);
or U12695 (N_12695,N_9894,N_11486);
nor U12696 (N_12696,N_8392,N_10292);
xor U12697 (N_12697,N_10662,N_10718);
and U12698 (N_12698,N_10849,N_9783);
nor U12699 (N_12699,N_9126,N_8239);
nor U12700 (N_12700,N_11773,N_11774);
and U12701 (N_12701,N_11154,N_11824);
and U12702 (N_12702,N_10249,N_9482);
or U12703 (N_12703,N_9138,N_9388);
xor U12704 (N_12704,N_9084,N_10217);
or U12705 (N_12705,N_9170,N_10801);
or U12706 (N_12706,N_9835,N_11437);
and U12707 (N_12707,N_8064,N_11787);
nor U12708 (N_12708,N_11821,N_8976);
and U12709 (N_12709,N_9231,N_8871);
xnor U12710 (N_12710,N_11265,N_8683);
nand U12711 (N_12711,N_9173,N_11398);
xor U12712 (N_12712,N_11915,N_9587);
nand U12713 (N_12713,N_11232,N_8450);
or U12714 (N_12714,N_10407,N_8233);
nand U12715 (N_12715,N_10117,N_9028);
nand U12716 (N_12716,N_10491,N_10403);
or U12717 (N_12717,N_11668,N_8372);
or U12718 (N_12718,N_10462,N_10512);
or U12719 (N_12719,N_10661,N_10578);
nand U12720 (N_12720,N_8711,N_11287);
xnor U12721 (N_12721,N_8265,N_8135);
or U12722 (N_12722,N_10357,N_10368);
nand U12723 (N_12723,N_10466,N_9936);
nand U12724 (N_12724,N_9290,N_9546);
nor U12725 (N_12725,N_8024,N_9568);
or U12726 (N_12726,N_11498,N_8374);
nand U12727 (N_12727,N_9807,N_8562);
and U12728 (N_12728,N_10652,N_8679);
or U12729 (N_12729,N_11851,N_9855);
xnor U12730 (N_12730,N_11173,N_9527);
xor U12731 (N_12731,N_8867,N_9417);
nand U12732 (N_12732,N_9008,N_8091);
xor U12733 (N_12733,N_9371,N_9096);
nand U12734 (N_12734,N_8457,N_9302);
and U12735 (N_12735,N_11613,N_10209);
nor U12736 (N_12736,N_11994,N_9308);
and U12737 (N_12737,N_8215,N_9822);
and U12738 (N_12738,N_9200,N_11062);
xnor U12739 (N_12739,N_10317,N_8493);
nor U12740 (N_12740,N_11337,N_10196);
xnor U12741 (N_12741,N_9678,N_8910);
or U12742 (N_12742,N_9800,N_9884);
or U12743 (N_12743,N_9431,N_11501);
or U12744 (N_12744,N_11008,N_10037);
or U12745 (N_12745,N_8849,N_10899);
nand U12746 (N_12746,N_9354,N_11762);
nand U12747 (N_12747,N_8502,N_11208);
xnor U12748 (N_12748,N_9871,N_9418);
and U12749 (N_12749,N_10969,N_10693);
xnor U12750 (N_12750,N_11070,N_10888);
xnor U12751 (N_12751,N_8248,N_10701);
nand U12752 (N_12752,N_8829,N_9705);
nor U12753 (N_12753,N_9751,N_9921);
nor U12754 (N_12754,N_8094,N_11180);
nor U12755 (N_12755,N_11345,N_11839);
xor U12756 (N_12756,N_10251,N_8478);
and U12757 (N_12757,N_8151,N_10410);
nor U12758 (N_12758,N_8000,N_8843);
or U12759 (N_12759,N_10966,N_10664);
nor U12760 (N_12760,N_11318,N_11387);
and U12761 (N_12761,N_10072,N_8655);
nand U12762 (N_12762,N_10284,N_9977);
and U12763 (N_12763,N_10746,N_9570);
or U12764 (N_12764,N_10984,N_11970);
or U12765 (N_12765,N_9947,N_9967);
xnor U12766 (N_12766,N_9750,N_10074);
and U12767 (N_12767,N_11291,N_9728);
nor U12768 (N_12768,N_11874,N_11999);
nand U12769 (N_12769,N_11469,N_8355);
nor U12770 (N_12770,N_10958,N_9562);
xnor U12771 (N_12771,N_9424,N_8234);
xnor U12772 (N_12772,N_11025,N_8889);
nand U12773 (N_12773,N_8191,N_10860);
xor U12774 (N_12774,N_10485,N_10133);
or U12775 (N_12775,N_10542,N_8337);
or U12776 (N_12776,N_10567,N_9739);
xor U12777 (N_12777,N_10732,N_9323);
nor U12778 (N_12778,N_10880,N_8687);
nor U12779 (N_12779,N_8566,N_9902);
xnor U12780 (N_12780,N_11385,N_8919);
nor U12781 (N_12781,N_10826,N_9163);
and U12782 (N_12782,N_8543,N_11962);
or U12783 (N_12783,N_8044,N_9119);
nand U12784 (N_12784,N_10912,N_11246);
xnor U12785 (N_12785,N_11237,N_10186);
nand U12786 (N_12786,N_8369,N_8126);
and U12787 (N_12787,N_10000,N_9870);
nor U12788 (N_12788,N_8205,N_10630);
xnor U12789 (N_12789,N_8886,N_11430);
nand U12790 (N_12790,N_10002,N_9736);
xnor U12791 (N_12791,N_9869,N_11006);
and U12792 (N_12792,N_9637,N_11071);
nand U12793 (N_12793,N_11648,N_9311);
or U12794 (N_12794,N_9731,N_9430);
nand U12795 (N_12795,N_10893,N_8583);
xnor U12796 (N_12796,N_8437,N_10277);
nand U12797 (N_12797,N_8058,N_10769);
or U12798 (N_12798,N_8736,N_11810);
nand U12799 (N_12799,N_9433,N_9541);
nor U12800 (N_12800,N_9524,N_9021);
xnor U12801 (N_12801,N_11634,N_8113);
and U12802 (N_12802,N_11736,N_10905);
xnor U12803 (N_12803,N_9633,N_8292);
nor U12804 (N_12804,N_11977,N_8592);
xnor U12805 (N_12805,N_9552,N_8924);
xor U12806 (N_12806,N_11786,N_11899);
nor U12807 (N_12807,N_9569,N_11618);
or U12808 (N_12808,N_8486,N_10386);
nand U12809 (N_12809,N_8906,N_9829);
or U12810 (N_12810,N_10931,N_11638);
and U12811 (N_12811,N_8193,N_8983);
xnor U12812 (N_12812,N_9553,N_11687);
and U12813 (N_12813,N_11712,N_9437);
nor U12814 (N_12814,N_10775,N_11629);
and U12815 (N_12815,N_10092,N_11639);
or U12816 (N_12816,N_10995,N_8552);
or U12817 (N_12817,N_11867,N_9180);
nor U12818 (N_12818,N_10728,N_9316);
xnor U12819 (N_12819,N_9299,N_10523);
nand U12820 (N_12820,N_9241,N_9851);
nand U12821 (N_12821,N_9515,N_9547);
nor U12822 (N_12822,N_11624,N_11643);
xor U12823 (N_12823,N_8510,N_10103);
xnor U12824 (N_12824,N_10668,N_9718);
and U12825 (N_12825,N_9726,N_11607);
and U12826 (N_12826,N_8477,N_11035);
nor U12827 (N_12827,N_9908,N_10576);
nor U12828 (N_12828,N_11620,N_8966);
nor U12829 (N_12829,N_9611,N_9686);
and U12830 (N_12830,N_11251,N_8666);
nor U12831 (N_12831,N_8984,N_8242);
nor U12832 (N_12832,N_11943,N_10963);
nor U12833 (N_12833,N_11776,N_10020);
nor U12834 (N_12834,N_10761,N_10848);
or U12835 (N_12835,N_11949,N_8409);
xnor U12836 (N_12836,N_10126,N_9681);
or U12837 (N_12837,N_10128,N_8712);
nor U12838 (N_12838,N_11193,N_11746);
nor U12839 (N_12839,N_8989,N_9940);
xor U12840 (N_12840,N_9203,N_10373);
or U12841 (N_12841,N_8360,N_11983);
nor U12842 (N_12842,N_11192,N_8294);
xor U12843 (N_12843,N_11892,N_8643);
and U12844 (N_12844,N_10601,N_11300);
nand U12845 (N_12845,N_10724,N_11910);
or U12846 (N_12846,N_11339,N_8220);
xnor U12847 (N_12847,N_10411,N_10649);
xor U12848 (N_12848,N_8606,N_10790);
nand U12849 (N_12849,N_8142,N_8501);
nand U12850 (N_12850,N_8625,N_11594);
or U12851 (N_12851,N_9922,N_8766);
xor U12852 (N_12852,N_9795,N_11841);
nor U12853 (N_12853,N_10819,N_11276);
xor U12854 (N_12854,N_9110,N_10065);
and U12855 (N_12855,N_10640,N_8796);
xnor U12856 (N_12856,N_10947,N_8750);
nand U12857 (N_12857,N_11521,N_9523);
and U12858 (N_12858,N_8075,N_9993);
or U12859 (N_12859,N_10318,N_9512);
nand U12860 (N_12860,N_11289,N_10431);
and U12861 (N_12861,N_10951,N_9360);
and U12862 (N_12862,N_11996,N_10663);
and U12863 (N_12863,N_11257,N_8048);
xor U12864 (N_12864,N_8706,N_8257);
and U12865 (N_12865,N_8418,N_9763);
nand U12866 (N_12866,N_10465,N_11991);
xnor U12867 (N_12867,N_10889,N_9957);
nor U12868 (N_12868,N_11719,N_10376);
nor U12869 (N_12869,N_9230,N_8250);
or U12870 (N_12870,N_11124,N_11788);
nand U12871 (N_12871,N_9729,N_8714);
xnor U12872 (N_12872,N_10739,N_9659);
and U12873 (N_12873,N_10771,N_8466);
nor U12874 (N_12874,N_10680,N_10375);
and U12875 (N_12875,N_10721,N_10954);
nand U12876 (N_12876,N_8467,N_11945);
and U12877 (N_12877,N_9608,N_11317);
nor U12878 (N_12878,N_11381,N_8298);
and U12879 (N_12879,N_8259,N_10443);
and U12880 (N_12880,N_9528,N_9117);
nor U12881 (N_12881,N_11158,N_8780);
or U12882 (N_12882,N_9976,N_11713);
and U12883 (N_12883,N_10435,N_10585);
or U12884 (N_12884,N_8047,N_11575);
and U12885 (N_12885,N_8362,N_8482);
xor U12886 (N_12886,N_10200,N_11448);
nand U12887 (N_12887,N_11148,N_8007);
nand U12888 (N_12888,N_10048,N_10202);
or U12889 (N_12889,N_10671,N_10735);
nand U12890 (N_12890,N_8535,N_11057);
and U12891 (N_12891,N_10501,N_11888);
or U12892 (N_12892,N_11680,N_11095);
xor U12893 (N_12893,N_9401,N_8540);
nor U12894 (N_12894,N_9842,N_10627);
or U12895 (N_12895,N_10785,N_8271);
xor U12896 (N_12896,N_11812,N_10795);
nor U12897 (N_12897,N_10146,N_10281);
and U12898 (N_12898,N_10729,N_9095);
nand U12899 (N_12899,N_11449,N_9645);
and U12900 (N_12900,N_9324,N_10743);
or U12901 (N_12901,N_10367,N_8003);
or U12902 (N_12902,N_10114,N_9812);
nor U12903 (N_12903,N_11485,N_9218);
nor U12904 (N_12904,N_9264,N_10877);
or U12905 (N_12905,N_10996,N_8768);
and U12906 (N_12906,N_11103,N_9778);
and U12907 (N_12907,N_9004,N_11286);
or U12908 (N_12908,N_8880,N_11523);
xnor U12909 (N_12909,N_11800,N_9465);
nand U12910 (N_12910,N_8875,N_8314);
and U12911 (N_12911,N_8903,N_11914);
nand U12912 (N_12912,N_8782,N_9897);
xnor U12913 (N_12913,N_8181,N_10589);
nor U12914 (N_12914,N_10346,N_11524);
and U12915 (N_12915,N_11816,N_8032);
nor U12916 (N_12916,N_9959,N_8860);
or U12917 (N_12917,N_8520,N_10057);
or U12918 (N_12918,N_11410,N_10690);
nand U12919 (N_12919,N_10977,N_8814);
or U12920 (N_12920,N_9064,N_9640);
and U12921 (N_12921,N_10506,N_10215);
nor U12922 (N_12922,N_9952,N_10027);
nor U12923 (N_12923,N_8290,N_10442);
nand U12924 (N_12924,N_10321,N_9900);
and U12925 (N_12925,N_11438,N_11178);
xor U12926 (N_12926,N_10170,N_8052);
or U12927 (N_12927,N_8225,N_11326);
or U12928 (N_12928,N_10194,N_8868);
or U12929 (N_12929,N_10179,N_10839);
nor U12930 (N_12930,N_8211,N_8009);
xnor U12931 (N_12931,N_8326,N_9913);
nand U12932 (N_12932,N_11852,N_9759);
and U12933 (N_12933,N_11020,N_10844);
or U12934 (N_12934,N_11753,N_10324);
or U12935 (N_12935,N_10228,N_9150);
xnor U12936 (N_12936,N_10678,N_8204);
xor U12937 (N_12937,N_10295,N_8526);
and U12938 (N_12938,N_11911,N_9082);
and U12939 (N_12939,N_10659,N_9511);
nor U12940 (N_12940,N_9651,N_8954);
nand U12941 (N_12941,N_9154,N_9103);
or U12942 (N_12942,N_11838,N_11725);
nor U12943 (N_12943,N_11036,N_10946);
nand U12944 (N_12944,N_11496,N_8998);
nor U12945 (N_12945,N_11711,N_8805);
and U12946 (N_12946,N_11557,N_8394);
or U12947 (N_12947,N_10957,N_8987);
nor U12948 (N_12948,N_9423,N_9213);
or U12949 (N_12949,N_9033,N_11077);
xnor U12950 (N_12950,N_11433,N_10257);
nand U12951 (N_12951,N_10517,N_9649);
nand U12952 (N_12952,N_8097,N_11181);
nor U12953 (N_12953,N_11435,N_8827);
and U12954 (N_12954,N_8459,N_9140);
nand U12955 (N_12955,N_10018,N_11884);
or U12956 (N_12956,N_9694,N_9184);
xor U12957 (N_12957,N_9351,N_10449);
or U12958 (N_12958,N_10782,N_8174);
or U12959 (N_12959,N_11754,N_9448);
and U12960 (N_12960,N_10593,N_9961);
or U12961 (N_12961,N_11803,N_11235);
xor U12962 (N_12962,N_8001,N_10286);
xnor U12963 (N_12963,N_8631,N_9375);
or U12964 (N_12964,N_9301,N_9210);
xor U12965 (N_12965,N_10546,N_10798);
xor U12966 (N_12966,N_8682,N_10901);
nor U12967 (N_12967,N_9749,N_11506);
and U12968 (N_12968,N_10141,N_8608);
and U12969 (N_12969,N_8816,N_9609);
and U12970 (N_12970,N_10129,N_10210);
xnor U12971 (N_12971,N_10152,N_11128);
xnor U12972 (N_12972,N_11081,N_10051);
or U12973 (N_12973,N_9941,N_8400);
or U12974 (N_12974,N_9099,N_10143);
nor U12975 (N_12975,N_10322,N_9161);
xor U12976 (N_12976,N_11458,N_10748);
or U12977 (N_12977,N_11848,N_11134);
and U12978 (N_12978,N_11024,N_10638);
or U12979 (N_12979,N_9083,N_11316);
nand U12980 (N_12980,N_8028,N_8375);
xnor U12981 (N_12981,N_8943,N_11871);
xor U12982 (N_12982,N_8644,N_10109);
xor U12983 (N_12983,N_9175,N_10047);
and U12984 (N_12984,N_10093,N_9214);
xor U12985 (N_12985,N_8037,N_11856);
or U12986 (N_12986,N_10962,N_10596);
and U12987 (N_12987,N_8406,N_9774);
nor U12988 (N_12988,N_11214,N_10326);
xnor U12989 (N_12989,N_8817,N_9297);
nor U12990 (N_12990,N_11218,N_10656);
xor U12991 (N_12991,N_8115,N_9581);
and U12992 (N_12992,N_11666,N_8432);
xor U12993 (N_12993,N_11799,N_10700);
and U12994 (N_12994,N_11044,N_10686);
or U12995 (N_12995,N_9298,N_8258);
or U12996 (N_12996,N_9592,N_11421);
or U12997 (N_12997,N_11834,N_11335);
nor U12998 (N_12998,N_8810,N_8172);
and U12999 (N_12999,N_10917,N_9307);
nand U13000 (N_13000,N_11608,N_8840);
nand U13001 (N_13001,N_9816,N_11825);
and U13002 (N_13002,N_11908,N_8264);
or U13003 (N_13003,N_9164,N_10279);
xor U13004 (N_13004,N_8396,N_10895);
xnor U13005 (N_13005,N_8309,N_11616);
xor U13006 (N_13006,N_9434,N_11122);
and U13007 (N_13007,N_8206,N_10153);
and U13008 (N_13008,N_10876,N_8786);
nor U13009 (N_13009,N_9199,N_11219);
and U13010 (N_13010,N_10468,N_11906);
xor U13011 (N_13011,N_10903,N_10213);
nand U13012 (N_13012,N_10519,N_9339);
and U13013 (N_13013,N_11534,N_9765);
nor U13014 (N_13014,N_11260,N_9309);
and U13015 (N_13015,N_8975,N_9225);
nand U13016 (N_13016,N_9073,N_9839);
nand U13017 (N_13017,N_10382,N_10787);
or U13018 (N_13018,N_10812,N_8698);
nand U13019 (N_13019,N_10297,N_10127);
xnor U13020 (N_13020,N_9683,N_9760);
nand U13021 (N_13021,N_11747,N_11752);
nor U13022 (N_13022,N_9513,N_8035);
nand U13023 (N_13023,N_11744,N_9785);
nor U13024 (N_13024,N_9636,N_8610);
nor U13025 (N_13025,N_11156,N_9881);
and U13026 (N_13026,N_11186,N_9949);
and U13027 (N_13027,N_8781,N_8710);
nand U13028 (N_13028,N_9969,N_11549);
nor U13029 (N_13029,N_11633,N_8376);
xor U13030 (N_13030,N_9501,N_9072);
and U13031 (N_13031,N_9051,N_9193);
or U13032 (N_13032,N_9183,N_9488);
or U13033 (N_13033,N_11056,N_11021);
and U13034 (N_13034,N_11843,N_9951);
and U13035 (N_13035,N_8733,N_9370);
nor U13036 (N_13036,N_8597,N_10856);
nor U13037 (N_13037,N_8152,N_9661);
nor U13038 (N_13038,N_8252,N_10145);
nand U13039 (N_13039,N_11059,N_8888);
and U13040 (N_13040,N_11798,N_10742);
nor U13041 (N_13041,N_11054,N_11091);
or U13042 (N_13042,N_10600,N_9461);
nor U13043 (N_13043,N_11439,N_8960);
and U13044 (N_13044,N_8626,N_11202);
xor U13045 (N_13045,N_11954,N_11716);
or U13046 (N_13046,N_9516,N_10455);
nor U13047 (N_13047,N_11655,N_9268);
nor U13048 (N_13048,N_11678,N_8378);
or U13049 (N_13049,N_11264,N_11109);
and U13050 (N_13050,N_8441,N_11880);
nand U13051 (N_13051,N_10396,N_10733);
and U13052 (N_13052,N_10551,N_11127);
and U13053 (N_13053,N_8481,N_9171);
nand U13054 (N_13054,N_8969,N_11815);
nor U13055 (N_13055,N_8988,N_10475);
and U13056 (N_13056,N_10175,N_8061);
or U13057 (N_13057,N_8870,N_11530);
or U13058 (N_13058,N_10658,N_11047);
xnor U13059 (N_13059,N_10932,N_11015);
nand U13060 (N_13060,N_8411,N_10916);
nand U13061 (N_13061,N_8111,N_8549);
nor U13062 (N_13062,N_9444,N_9408);
xor U13063 (N_13063,N_11697,N_9917);
and U13064 (N_13064,N_9194,N_11436);
and U13065 (N_13065,N_11907,N_11220);
or U13066 (N_13066,N_10527,N_9362);
nor U13067 (N_13067,N_10549,N_11078);
and U13068 (N_13068,N_9737,N_11119);
xnor U13069 (N_13069,N_9081,N_11076);
xor U13070 (N_13070,N_10884,N_10535);
or U13071 (N_13071,N_11931,N_9130);
xnor U13072 (N_13072,N_11960,N_10694);
nor U13073 (N_13073,N_10791,N_9734);
or U13074 (N_13074,N_8013,N_8153);
and U13075 (N_13075,N_9998,N_8498);
xnor U13076 (N_13076,N_10010,N_10406);
nand U13077 (N_13077,N_10383,N_11822);
and U13078 (N_13078,N_8709,N_8240);
nand U13079 (N_13079,N_9058,N_11083);
xor U13080 (N_13080,N_9810,N_11234);
or U13081 (N_13081,N_9078,N_9450);
nand U13082 (N_13082,N_8662,N_11373);
xor U13083 (N_13083,N_9586,N_11340);
xor U13084 (N_13084,N_9631,N_8728);
or U13085 (N_13085,N_9336,N_11460);
xor U13086 (N_13086,N_10343,N_10873);
nand U13087 (N_13087,N_8183,N_11805);
nand U13088 (N_13088,N_8853,N_10490);
nand U13089 (N_13089,N_8588,N_8373);
nor U13090 (N_13090,N_9756,N_8640);
or U13091 (N_13091,N_10230,N_11869);
and U13092 (N_13092,N_8531,N_11966);
and U13093 (N_13093,N_10017,N_8941);
xor U13094 (N_13094,N_10285,N_11167);
nand U13095 (N_13095,N_10212,N_11445);
and U13096 (N_13096,N_9725,N_11412);
nand U13097 (N_13097,N_9883,N_10773);
nand U13098 (N_13098,N_11577,N_11829);
and U13099 (N_13099,N_9416,N_11189);
nand U13100 (N_13100,N_11793,N_10763);
nor U13101 (N_13101,N_9027,N_8395);
nand U13102 (N_13102,N_8364,N_10471);
nand U13103 (N_13103,N_10470,N_10956);
or U13104 (N_13104,N_8615,N_8066);
or U13105 (N_13105,N_11308,N_11471);
nor U13106 (N_13106,N_11196,N_9221);
xnor U13107 (N_13107,N_10529,N_9794);
nor U13108 (N_13108,N_9968,N_11875);
xnor U13109 (N_13109,N_8266,N_9744);
nor U13110 (N_13110,N_11714,N_9740);
or U13111 (N_13111,N_9738,N_9630);
and U13112 (N_13112,N_10438,N_11299);
nand U13113 (N_13113,N_9366,N_9454);
nor U13114 (N_13114,N_8968,N_8325);
and U13115 (N_13115,N_8354,N_9291);
nor U13116 (N_13116,N_10166,N_9091);
xor U13117 (N_13117,N_8665,N_8559);
nor U13118 (N_13118,N_10714,N_10636);
nand U13119 (N_13119,N_8633,N_9727);
nor U13120 (N_13120,N_8821,N_11263);
xor U13121 (N_13121,N_8322,N_9055);
nor U13122 (N_13122,N_10330,N_11332);
or U13123 (N_13123,N_9216,N_9097);
and U13124 (N_13124,N_11512,N_9886);
nor U13125 (N_13125,N_10130,N_10205);
nor U13126 (N_13126,N_9688,N_11022);
xor U13127 (N_13127,N_9165,N_8690);
or U13128 (N_13128,N_11468,N_11551);
or U13129 (N_13129,N_8116,N_10965);
nand U13130 (N_13130,N_8532,N_9906);
and U13131 (N_13131,N_10474,N_8804);
or U13132 (N_13132,N_11585,N_8536);
nand U13133 (N_13133,N_11926,N_8426);
and U13134 (N_13134,N_11877,N_9827);
or U13135 (N_13135,N_11434,N_9100);
nor U13136 (N_13136,N_9504,N_10289);
xor U13137 (N_13137,N_9128,N_9247);
nand U13138 (N_13138,N_8171,N_10287);
xnor U13139 (N_13139,N_10162,N_9788);
nor U13140 (N_13140,N_10563,N_9755);
xnor U13141 (N_13141,N_11538,N_11720);
and U13142 (N_13142,N_10834,N_8166);
nor U13143 (N_13143,N_9212,N_9279);
or U13144 (N_13144,N_10569,N_9818);
or U13145 (N_13145,N_10164,N_10734);
nor U13146 (N_13146,N_11717,N_8405);
and U13147 (N_13147,N_9848,N_9167);
or U13148 (N_13148,N_11489,N_8546);
nand U13149 (N_13149,N_10499,N_9134);
nor U13150 (N_13150,N_9332,N_8878);
nand U13151 (N_13151,N_8895,N_9665);
or U13152 (N_13152,N_10525,N_9012);
and U13153 (N_13153,N_9088,N_10918);
and U13154 (N_13154,N_8713,N_8599);
xor U13155 (N_13155,N_8776,N_8896);
and U13156 (N_13156,N_10388,N_9120);
nor U13157 (N_13157,N_8717,N_10180);
nand U13158 (N_13158,N_8131,N_8949);
xnor U13159 (N_13159,N_9503,N_11045);
nor U13160 (N_13160,N_11732,N_10080);
xnor U13161 (N_13161,N_8748,N_9677);
xnor U13162 (N_13162,N_8300,N_9550);
nand U13163 (N_13163,N_9874,N_9472);
and U13164 (N_13164,N_11135,N_8017);
or U13165 (N_13165,N_8997,N_10070);
xnor U13166 (N_13166,N_8921,N_10137);
nand U13167 (N_13167,N_8541,N_8724);
nor U13168 (N_13168,N_9162,N_10054);
and U13169 (N_13169,N_9040,N_8636);
nand U13170 (N_13170,N_10838,N_10099);
nand U13171 (N_13171,N_8422,N_10252);
and U13172 (N_13172,N_8214,N_11169);
or U13173 (N_13173,N_8811,N_9745);
nor U13174 (N_13174,N_10768,N_11376);
xor U13175 (N_13175,N_8157,N_8033);
nor U13176 (N_13176,N_9852,N_11227);
nor U13177 (N_13177,N_9466,N_11042);
xor U13178 (N_13178,N_11415,N_11032);
xor U13179 (N_13179,N_11992,N_8517);
or U13180 (N_13180,N_11288,N_11459);
nand U13181 (N_13181,N_10429,N_8946);
or U13182 (N_13182,N_11336,N_9262);
or U13183 (N_13183,N_8127,N_11932);
nor U13184 (N_13184,N_9253,N_8839);
or U13185 (N_13185,N_8579,N_8869);
or U13186 (N_13186,N_10858,N_9850);
nor U13187 (N_13187,N_11536,N_8971);
nand U13188 (N_13188,N_10920,N_10526);
and U13189 (N_13189,N_9741,N_11818);
and U13190 (N_13190,N_9905,N_10272);
and U13191 (N_13191,N_11859,N_8288);
and U13192 (N_13192,N_9300,N_10046);
and U13193 (N_13193,N_10892,N_8207);
and U13194 (N_13194,N_11583,N_11703);
xnor U13195 (N_13195,N_8251,N_8398);
nand U13196 (N_13196,N_11503,N_11049);
and U13197 (N_13197,N_11110,N_11277);
or U13198 (N_13198,N_9405,N_11531);
xor U13199 (N_13199,N_10174,N_10007);
nand U13200 (N_13200,N_8560,N_10606);
and U13201 (N_13201,N_10670,N_9711);
nand U13202 (N_13202,N_10595,N_10896);
nor U13203 (N_13203,N_10590,N_10173);
xor U13204 (N_13204,N_10253,N_11682);
nor U13205 (N_13205,N_11005,N_8580);
and U13206 (N_13206,N_9925,N_8201);
nor U13207 (N_13207,N_11001,N_9987);
nor U13208 (N_13208,N_10852,N_11116);
or U13209 (N_13209,N_10139,N_10225);
or U13210 (N_13210,N_11058,N_9537);
nand U13211 (N_13211,N_10861,N_10822);
and U13212 (N_13212,N_8062,N_11065);
and U13213 (N_13213,N_8452,N_9597);
nand U13214 (N_13214,N_9122,N_9676);
nand U13215 (N_13215,N_9713,N_10792);
xor U13216 (N_13216,N_9618,N_9019);
nor U13217 (N_13217,N_11312,N_11548);
or U13218 (N_13218,N_9182,N_11710);
or U13219 (N_13219,N_9722,N_11632);
nand U13220 (N_13220,N_11772,N_8722);
and U13221 (N_13221,N_11406,N_9394);
or U13222 (N_13222,N_9490,N_9062);
nor U13223 (N_13223,N_8276,N_9006);
and U13224 (N_13224,N_11748,N_10657);
nand U13225 (N_13225,N_9382,N_10060);
or U13226 (N_13226,N_8846,N_10960);
and U13227 (N_13227,N_8820,N_9817);
nand U13228 (N_13228,N_10759,N_10776);
and U13229 (N_13229,N_8014,N_9937);
nand U13230 (N_13230,N_10633,N_8800);
xnor U13231 (N_13231,N_11883,N_9481);
nand U13232 (N_13232,N_10484,N_11039);
xnor U13233 (N_13233,N_8794,N_9108);
or U13234 (N_13234,N_8934,N_11310);
or U13235 (N_13235,N_8514,N_11223);
or U13236 (N_13236,N_8668,N_10313);
nand U13237 (N_13237,N_11652,N_10753);
nor U13238 (N_13238,N_11863,N_8256);
nand U13239 (N_13239,N_9682,N_10036);
nor U13240 (N_13240,N_10929,N_10921);
xor U13241 (N_13241,N_9840,N_10760);
and U13242 (N_13242,N_8447,N_8861);
nand U13243 (N_13243,N_10157,N_10482);
nor U13244 (N_13244,N_9635,N_8407);
or U13245 (N_13245,N_8150,N_8617);
and U13246 (N_13246,N_10098,N_9469);
xnor U13247 (N_13247,N_11589,N_8848);
nand U13248 (N_13248,N_11243,N_10483);
or U13249 (N_13249,N_9347,N_11290);
nand U13250 (N_13250,N_9042,N_11479);
nor U13251 (N_13251,N_8977,N_11354);
and U13252 (N_13252,N_10757,N_8676);
or U13253 (N_13253,N_9714,N_9471);
nor U13254 (N_13254,N_11082,N_11372);
nand U13255 (N_13255,N_8581,N_8387);
nor U13256 (N_13256,N_10101,N_11271);
nor U13257 (N_13257,N_11933,N_9625);
xor U13258 (N_13258,N_10738,N_11951);
nand U13259 (N_13259,N_10005,N_11098);
xor U13260 (N_13260,N_10938,N_10684);
or U13261 (N_13261,N_9580,N_9476);
nor U13262 (N_13262,N_8397,N_8391);
and U13263 (N_13263,N_9322,N_11041);
xnor U13264 (N_13264,N_9910,N_8303);
nor U13265 (N_13265,N_9364,N_10142);
and U13266 (N_13266,N_10241,N_9020);
or U13267 (N_13267,N_10235,N_10496);
xor U13268 (N_13268,N_10233,N_10091);
nand U13269 (N_13269,N_11108,N_10642);
and U13270 (N_13270,N_10997,N_8324);
and U13271 (N_13271,N_8743,N_8648);
or U13272 (N_13272,N_9429,N_10293);
and U13273 (N_13273,N_11155,N_10784);
nand U13274 (N_13274,N_10820,N_9948);
nor U13275 (N_13275,N_10989,N_8603);
nor U13276 (N_13276,N_8209,N_11930);
nor U13277 (N_13277,N_9971,N_10182);
nand U13278 (N_13278,N_11487,N_11901);
nand U13279 (N_13279,N_8789,N_11275);
and U13280 (N_13280,N_11351,N_8463);
and U13281 (N_13281,N_8826,N_8884);
and U13282 (N_13282,N_11604,N_11936);
nand U13283 (N_13283,N_11569,N_10699);
xor U13284 (N_13284,N_8569,N_8909);
or U13285 (N_13285,N_8420,N_11705);
or U13286 (N_13286,N_9934,N_11359);
and U13287 (N_13287,N_8453,N_11592);
xor U13288 (N_13288,N_11231,N_10708);
nor U13289 (N_13289,N_11447,N_8542);
nor U13290 (N_13290,N_10171,N_11917);
xnor U13291 (N_13291,N_9603,N_8109);
nor U13292 (N_13292,N_10224,N_8081);
and U13293 (N_13293,N_11728,N_11104);
nand U13294 (N_13294,N_9999,N_10356);
xor U13295 (N_13295,N_8999,N_11584);
or U13296 (N_13296,N_10799,N_10362);
or U13297 (N_13297,N_9149,N_9289);
and U13298 (N_13298,N_11905,N_9578);
nor U13299 (N_13299,N_9824,N_11653);
nand U13300 (N_13300,N_9281,N_9813);
xor U13301 (N_13301,N_11564,N_10545);
or U13302 (N_13302,N_10204,N_8268);
nor U13303 (N_13303,N_9045,N_11362);
xnor U13304 (N_13304,N_11111,N_11188);
xnor U13305 (N_13305,N_9346,N_11601);
and U13306 (N_13306,N_8978,N_11225);
and U13307 (N_13307,N_8245,N_11429);
and U13308 (N_13308,N_10603,N_8807);
nor U13309 (N_13309,N_9543,N_11550);
or U13310 (N_13310,N_10081,N_10562);
or U13311 (N_13311,N_9061,N_9105);
nand U13312 (N_13312,N_10922,N_11200);
or U13313 (N_13313,N_9721,N_9964);
or U13314 (N_13314,N_10078,N_9355);
and U13315 (N_13315,N_11947,N_8823);
xnor U13316 (N_13316,N_10665,N_8069);
nor U13317 (N_13317,N_10372,N_8935);
nor U13318 (N_13318,N_8228,N_11428);
and U13319 (N_13319,N_10871,N_11422);
or U13320 (N_13320,N_9944,N_8089);
nand U13321 (N_13321,N_10239,N_9046);
and U13322 (N_13322,N_9232,N_8831);
nand U13323 (N_13323,N_11441,N_8041);
and U13324 (N_13324,N_8154,N_11543);
and U13325 (N_13325,N_8950,N_10197);
and U13326 (N_13326,N_9384,N_9571);
nor U13327 (N_13327,N_11369,N_10737);
or U13328 (N_13328,N_11518,N_11505);
nor U13329 (N_13329,N_11187,N_8039);
xnor U13330 (N_13330,N_11578,N_9505);
xnor U13331 (N_13331,N_9338,N_9780);
and U13332 (N_13332,N_8237,N_9821);
or U13333 (N_13333,N_10104,N_9923);
and U13334 (N_13334,N_11567,N_8471);
nand U13335 (N_13335,N_9023,N_11916);
or U13336 (N_13336,N_9627,N_8841);
and U13337 (N_13337,N_11450,N_10720);
and U13338 (N_13338,N_8990,N_11677);
or U13339 (N_13339,N_10581,N_10345);
xor U13340 (N_13340,N_11348,N_8198);
xor U13341 (N_13341,N_11985,N_9265);
nand U13342 (N_13342,N_11555,N_9310);
nand U13343 (N_13343,N_10660,N_11197);
xor U13344 (N_13344,N_9395,N_8353);
nor U13345 (N_13345,N_11849,N_10894);
or U13346 (N_13346,N_8140,N_10598);
nand U13347 (N_13347,N_8167,N_8705);
xor U13348 (N_13348,N_9284,N_8567);
nand U13349 (N_13349,N_9252,N_9325);
nor U13350 (N_13350,N_11721,N_10629);
xor U13351 (N_13351,N_9732,N_11659);
nor U13352 (N_13352,N_10365,N_10309);
or U13353 (N_13353,N_11370,N_8377);
nor U13354 (N_13354,N_9151,N_8678);
xor U13355 (N_13355,N_8897,N_11426);
nor U13356 (N_13356,N_8366,N_9622);
and U13357 (N_13357,N_8738,N_10476);
nand U13358 (N_13358,N_9615,N_9142);
and U13359 (N_13359,N_11708,N_10404);
and U13360 (N_13360,N_10673,N_9489);
nor U13361 (N_13361,N_10006,N_11230);
nand U13362 (N_13362,N_11377,N_11141);
or U13363 (N_13363,N_11813,N_8344);
nor U13364 (N_13364,N_11027,N_9240);
or U13365 (N_13365,N_8347,N_8050);
xnor U13366 (N_13366,N_8020,N_9493);
nand U13367 (N_13367,N_9076,N_10340);
or U13368 (N_13368,N_9038,N_11388);
nor U13369 (N_13369,N_10100,N_9080);
nand U13370 (N_13370,N_9492,N_10039);
or U13371 (N_13371,N_11504,N_10857);
xnor U13372 (N_13372,N_8446,N_11378);
nand U13373 (N_13373,N_9217,N_11804);
and U13374 (N_13374,N_8746,N_8859);
nand U13375 (N_13375,N_11198,N_9887);
nand U13376 (N_13376,N_10789,N_8570);
nand U13377 (N_13377,N_11587,N_8356);
nand U13378 (N_13378,N_10797,N_10342);
and U13379 (N_13379,N_8908,N_8647);
or U13380 (N_13380,N_8545,N_10459);
xor U13381 (N_13381,N_9446,N_9634);
xnor U13382 (N_13382,N_9085,N_9551);
nand U13383 (N_13383,N_11622,N_11669);
or U13384 (N_13384,N_10044,N_10959);
or U13385 (N_13385,N_11657,N_8320);
xor U13386 (N_13386,N_9228,N_10672);
xnor U13387 (N_13387,N_11229,N_10907);
or U13388 (N_13388,N_8791,N_8799);
nor U13389 (N_13389,N_8957,N_8652);
or U13390 (N_13390,N_10347,N_11510);
xnor U13391 (N_13391,N_9220,N_8605);
nor U13392 (N_13392,N_10374,N_10676);
or U13393 (N_13393,N_8221,N_10815);
nor U13394 (N_13394,N_11338,N_10865);
xnor U13395 (N_13395,N_11724,N_8219);
or U13396 (N_13396,N_11320,N_9208);
xor U13397 (N_13397,N_8483,N_9447);
nand U13398 (N_13398,N_10423,N_11107);
or U13399 (N_13399,N_11051,N_10994);
nand U13400 (N_13400,N_8917,N_9657);
and U13401 (N_13401,N_11862,N_10282);
or U13402 (N_13402,N_8267,N_11645);
or U13403 (N_13403,N_10028,N_9426);
or U13404 (N_13404,N_8622,N_9758);
xor U13405 (N_13405,N_9709,N_9102);
and U13406 (N_13406,N_9986,N_8488);
and U13407 (N_13407,N_10467,N_8635);
or U13408 (N_13408,N_8618,N_11117);
and U13409 (N_13409,N_11610,N_11693);
nor U13410 (N_13410,N_8509,N_10859);
or U13411 (N_13411,N_10397,N_11760);
or U13412 (N_13412,N_8381,N_10023);
xor U13413 (N_13413,N_10886,N_10264);
nor U13414 (N_13414,N_9219,N_11615);
and U13415 (N_13415,N_11297,N_9700);
xor U13416 (N_13416,N_9866,N_8316);
nor U13417 (N_13417,N_9619,N_11176);
and U13418 (N_13418,N_11328,N_9596);
or U13419 (N_13419,N_11898,N_9486);
nor U13420 (N_13420,N_9953,N_9825);
nor U13421 (N_13421,N_11252,N_8637);
and U13422 (N_13422,N_9484,N_9564);
nor U13423 (N_13423,N_9915,N_9391);
nor U13424 (N_13424,N_11730,N_9854);
nor U13425 (N_13425,N_10948,N_8106);
or U13426 (N_13426,N_9655,N_11350);
nand U13427 (N_13427,N_10011,N_9380);
and U13428 (N_13428,N_11513,N_9498);
or U13429 (N_13429,N_8272,N_8893);
and U13430 (N_13430,N_11136,N_8042);
or U13431 (N_13431,N_10507,N_8913);
nand U13432 (N_13432,N_9730,N_9129);
xnor U13433 (N_13433,N_11890,N_8060);
xnor U13434 (N_13434,N_10751,N_9837);
or U13435 (N_13435,N_10040,N_8996);
or U13436 (N_13436,N_10079,N_10192);
nor U13437 (N_13437,N_10904,N_10379);
and U13438 (N_13438,N_8936,N_8964);
nor U13439 (N_13439,N_11281,N_11563);
nand U13440 (N_13440,N_9719,N_9037);
xnor U13441 (N_13441,N_11478,N_11491);
nand U13442 (N_13442,N_11631,N_8836);
xor U13443 (N_13443,N_8929,N_11681);
nand U13444 (N_13444,N_9452,N_8494);
nand U13445 (N_13445,N_10344,N_10110);
nor U13446 (N_13446,N_9819,N_8778);
and U13447 (N_13447,N_10863,N_8985);
and U13448 (N_13448,N_8586,N_11964);
or U13449 (N_13449,N_9224,N_11399);
and U13450 (N_13450,N_8798,N_9293);
xnor U13451 (N_13451,N_8301,N_11727);
nand U13452 (N_13452,N_11606,N_8196);
xor U13453 (N_13453,N_10161,N_8658);
nand U13454 (N_13454,N_10981,N_11614);
and U13455 (N_13455,N_9642,N_9593);
nor U13456 (N_13456,N_9521,N_9136);
nor U13457 (N_13457,N_10401,N_8671);
and U13458 (N_13458,N_9583,N_11571);
or U13459 (N_13459,N_10883,N_8574);
nand U13460 (N_13460,N_10923,N_11031);
xnor U13461 (N_13461,N_9680,N_11718);
xor U13462 (N_13462,N_8404,N_11375);
or U13463 (N_13463,N_11185,N_11361);
nor U13464 (N_13464,N_8911,N_9879);
nand U13465 (N_13465,N_11965,N_8247);
and U13466 (N_13466,N_10183,N_11140);
nor U13467 (N_13467,N_10003,N_9013);
or U13468 (N_13468,N_8244,N_8812);
nand U13469 (N_13469,N_9670,N_8145);
nand U13470 (N_13470,N_11018,N_10333);
xor U13471 (N_13471,N_10354,N_8558);
nor U13472 (N_13472,N_8487,N_8056);
xnor U13473 (N_13473,N_8216,N_8792);
nor U13474 (N_13474,N_11179,N_10457);
xor U13475 (N_13475,N_11860,N_9672);
xor U13476 (N_13476,N_10591,N_10885);
and U13477 (N_13477,N_10211,N_9260);
xnor U13478 (N_13478,N_9776,N_10695);
nand U13479 (N_13479,N_9699,N_9043);
nand U13480 (N_13480,N_9412,N_11968);
nor U13481 (N_13481,N_8263,N_8071);
or U13482 (N_13482,N_10350,N_11826);
or U13483 (N_13483,N_10704,N_8226);
nand U13484 (N_13484,N_10592,N_9508);
nor U13485 (N_13485,N_11097,N_10059);
nor U13486 (N_13486,N_10716,N_8737);
or U13487 (N_13487,N_9201,N_11673);
or U13488 (N_13488,N_11014,N_8729);
nor U13489 (N_13489,N_11670,N_8129);
and U13490 (N_13490,N_8872,N_8744);
and U13491 (N_13491,N_8484,N_11658);
and U13492 (N_13492,N_11159,N_11961);
or U13493 (N_13493,N_11174,N_11957);
and U13494 (N_13494,N_8416,N_8419);
nand U13495 (N_13495,N_8762,N_8442);
or U13496 (N_13496,N_11089,N_11596);
nand U13497 (N_13497,N_10814,N_9650);
xor U13498 (N_13498,N_9176,N_10203);
xnor U13499 (N_13499,N_10073,N_8496);
or U13500 (N_13500,N_10788,N_10327);
nor U13501 (N_13501,N_8719,N_9494);
xnor U13502 (N_13502,N_8230,N_9003);
nand U13503 (N_13503,N_10845,N_10534);
and U13504 (N_13504,N_10319,N_8741);
nand U13505 (N_13505,N_8332,N_8735);
and U13506 (N_13506,N_10682,N_10999);
nor U13507 (N_13507,N_11453,N_11950);
nor U13508 (N_13508,N_10273,N_10832);
and U13509 (N_13509,N_9390,N_10553);
and U13510 (N_13510,N_11347,N_9385);
nor U13511 (N_13511,N_8808,N_11101);
and U13512 (N_13512,N_10294,N_10648);
or U13513 (N_13513,N_9724,N_9789);
nor U13514 (N_13514,N_10358,N_11153);
nor U13515 (N_13515,N_9420,N_9242);
or U13516 (N_13516,N_10710,N_9029);
nand U13517 (N_13517,N_11293,N_11974);
and U13518 (N_13518,N_10248,N_8508);
or U13519 (N_13519,N_9352,N_9978);
xnor U13520 (N_13520,N_9367,N_11952);
xor U13521 (N_13521,N_8537,N_8414);
xnor U13522 (N_13522,N_11553,N_8962);
or U13523 (N_13523,N_8834,N_11166);
and U13524 (N_13524,N_10583,N_8095);
and U13525 (N_13525,N_9853,N_11801);
and U13526 (N_13526,N_8065,N_11979);
and U13527 (N_13527,N_10016,N_11969);
or U13528 (N_13528,N_10021,N_10988);
or U13529 (N_13529,N_11796,N_11785);
or U13530 (N_13530,N_8755,N_10911);
or U13531 (N_13531,N_9419,N_9764);
nor U13532 (N_13532,N_9399,N_10990);
or U13533 (N_13533,N_10677,N_11028);
or U13534 (N_13534,N_10653,N_9836);
nor U13535 (N_13535,N_8086,N_9273);
xor U13536 (N_13536,N_9257,N_8084);
and U13537 (N_13537,N_8915,N_8293);
xor U13538 (N_13538,N_9345,N_9123);
and U13539 (N_13539,N_10979,N_11831);
xor U13540 (N_13540,N_8059,N_11294);
and U13541 (N_13541,N_8862,N_10316);
nand U13542 (N_13542,N_8133,N_8594);
and U13543 (N_13543,N_9034,N_10667);
or U13544 (N_13544,N_9782,N_8513);
or U13545 (N_13545,N_9335,N_9849);
and U13546 (N_13546,N_9753,N_10428);
nand U13547 (N_13547,N_10120,N_9997);
xor U13548 (N_13548,N_10539,N_11861);
and U13549 (N_13549,N_10867,N_9480);
nor U13550 (N_13550,N_11865,N_11939);
nand U13551 (N_13551,N_8449,N_10361);
nand U13552 (N_13552,N_11918,N_8624);
and U13553 (N_13553,N_11407,N_10935);
or U13554 (N_13554,N_10050,N_9133);
or U13555 (N_13555,N_10580,N_11837);
nand U13556 (N_13556,N_10042,N_8677);
or U13557 (N_13557,N_8659,N_8490);
nand U13558 (N_13558,N_8771,N_9862);
xnor U13559 (N_13559,N_9791,N_8421);
or U13560 (N_13560,N_8548,N_10725);
or U13561 (N_13561,N_10941,N_11100);
or U13562 (N_13562,N_9716,N_9945);
xnor U13563 (N_13563,N_9710,N_9754);
xnor U13564 (N_13564,N_10617,N_11088);
and U13565 (N_13565,N_11157,N_8170);
and U13566 (N_13566,N_9787,N_11806);
nor U13567 (N_13567,N_10854,N_8653);
or U13568 (N_13568,N_11967,N_9160);
xnor U13569 (N_13569,N_9895,N_9671);
xnor U13570 (N_13570,N_10645,N_8882);
or U13571 (N_13571,N_9510,N_11647);
xor U13572 (N_13572,N_8818,N_8669);
xnor U13573 (N_13573,N_9397,N_11093);
xor U13574 (N_13574,N_11325,N_11526);
nor U13575 (N_13575,N_10967,N_8402);
nor U13576 (N_13576,N_10624,N_9666);
nand U13577 (N_13577,N_11836,N_8769);
nand U13578 (N_13578,N_10351,N_9036);
nand U13579 (N_13579,N_10384,N_8864);
nand U13580 (N_13580,N_11203,N_9457);
nand U13581 (N_13581,N_9533,N_9181);
and U13582 (N_13582,N_10706,N_10116);
or U13583 (N_13583,N_8524,N_11876);
nor U13584 (N_13584,N_8972,N_10634);
or U13585 (N_13585,N_10647,N_11866);
nand U13586 (N_13586,N_9927,N_8455);
and U13587 (N_13587,N_8284,N_11630);
and U13588 (N_13588,N_8614,N_10515);
nor U13589 (N_13589,N_10177,N_10522);
or U13590 (N_13590,N_10674,N_8479);
and U13591 (N_13591,N_8321,N_8539);
or U13592 (N_13592,N_9157,N_9436);
or U13593 (N_13593,N_10418,N_10831);
and U13594 (N_13594,N_11879,N_11792);
and U13595 (N_13595,N_9148,N_8973);
nor U13596 (N_13596,N_10639,N_8851);
xor U13597 (N_13597,N_11017,N_11254);
or U13598 (N_13598,N_8883,N_10864);
or U13599 (N_13599,N_10083,N_11568);
nor U13600 (N_13600,N_10448,N_9304);
nand U13601 (N_13601,N_10805,N_11168);
xnor U13602 (N_13602,N_8627,N_10422);
and U13603 (N_13603,N_8461,N_10440);
nor U13604 (N_13604,N_11740,N_9561);
or U13605 (N_13605,N_11239,N_8555);
nor U13606 (N_13606,N_10813,N_10978);
nand U13607 (N_13607,N_11050,N_9567);
xor U13608 (N_13608,N_8891,N_10421);
nand U13609 (N_13609,N_10731,N_11228);
nor U13610 (N_13610,N_8346,N_11820);
nor U13611 (N_13611,N_10666,N_9143);
nand U13612 (N_13612,N_10243,N_8904);
nand U13613 (N_13613,N_11626,N_11561);
or U13614 (N_13614,N_8489,N_11152);
nor U13615 (N_13615,N_11893,N_10063);
nor U13616 (N_13616,N_11694,N_8838);
xor U13617 (N_13617,N_8078,N_11256);
nor U13618 (N_13618,N_9500,N_8953);
nand U13619 (N_13619,N_9315,N_10796);
xnor U13620 (N_13620,N_11700,N_11988);
nand U13621 (N_13621,N_10711,N_11702);
or U13622 (N_13622,N_9891,N_10464);
or U13623 (N_13623,N_11731,N_11656);
nand U13624 (N_13624,N_11074,N_11073);
or U13625 (N_13625,N_10745,N_8604);
and U13626 (N_13626,N_9464,N_10353);
nand U13627 (N_13627,N_8993,N_10308);
and U13628 (N_13628,N_10102,N_11789);
and U13629 (N_13629,N_11611,N_9502);
nand U13630 (N_13630,N_8822,N_8660);
nand U13631 (N_13631,N_9318,N_9762);
or U13632 (N_13632,N_11242,N_8715);
and U13633 (N_13633,N_9629,N_8182);
xor U13634 (N_13634,N_9282,N_9903);
and U13635 (N_13635,N_9017,N_8931);
or U13636 (N_13636,N_9449,N_11832);
xnor U13637 (N_13637,N_8313,N_11484);
nand U13638 (N_13638,N_8667,N_8815);
or U13639 (N_13639,N_9873,N_11795);
and U13640 (N_13640,N_10651,N_9962);
nand U13641 (N_13641,N_10952,N_10446);
or U13642 (N_13642,N_9526,N_10902);
nor U13643 (N_13643,N_8865,N_10381);
nand U13644 (N_13644,N_9331,N_9796);
nor U13645 (N_13645,N_10689,N_9867);
and U13646 (N_13646,N_9585,N_9844);
and U13647 (N_13647,N_9389,N_10976);
nand U13648 (N_13648,N_9487,N_9772);
or U13649 (N_13649,N_10783,N_9892);
and U13650 (N_13650,N_10772,N_10034);
and U13651 (N_13651,N_10510,N_9052);
nand U13652 (N_13652,N_11004,N_11828);
nor U13653 (N_13653,N_9495,N_8243);
nor U13654 (N_13654,N_9280,N_8222);
nor U13655 (N_13655,N_9024,N_8161);
and U13656 (N_13656,N_8727,N_11454);
nor U13657 (N_13657,N_11261,N_10024);
nor U13658 (N_13658,N_9056,N_8866);
nor U13659 (N_13659,N_9846,N_8854);
nand U13660 (N_13660,N_9093,N_9060);
and U13661 (N_13661,N_8246,N_10169);
and U13662 (N_13662,N_8956,N_11105);
xor U13663 (N_13663,N_10705,N_10486);
xor U13664 (N_13664,N_10208,N_11284);
or U13665 (N_13665,N_8304,N_10723);
xor U13666 (N_13666,N_8302,N_8443);
nor U13667 (N_13667,N_9172,N_9155);
and U13668 (N_13668,N_11976,N_11075);
and U13669 (N_13669,N_11444,N_9474);
nor U13670 (N_13670,N_10236,N_11069);
xor U13671 (N_13671,N_11365,N_10604);
nand U13672 (N_13672,N_10816,N_11334);
and U13673 (N_13673,N_10312,N_9566);
nand U13674 (N_13674,N_8689,N_9483);
nor U13675 (N_13675,N_8282,N_10112);
and U13676 (N_13676,N_9092,N_8088);
nor U13677 (N_13677,N_8894,N_8357);
xnor U13678 (N_13678,N_11195,N_11327);
or U13679 (N_13679,N_8340,N_8107);
xnor U13680 (N_13680,N_11497,N_8260);
nor U13681 (N_13681,N_10125,N_11722);
xor U13682 (N_13682,N_11855,N_10301);
or U13683 (N_13683,N_11737,N_10605);
nand U13684 (N_13684,N_10741,N_11114);
xnor U13685 (N_13685,N_11411,N_11502);
nor U13686 (N_13686,N_10415,N_11758);
nand U13687 (N_13687,N_10833,N_9995);
and U13688 (N_13688,N_9410,N_9074);
or U13689 (N_13689,N_8112,N_9602);
nand U13690 (N_13690,N_10927,N_11794);
or U13691 (N_13691,N_9538,N_11380);
or U13692 (N_13692,N_9358,N_8809);
and U13693 (N_13693,N_8731,N_11060);
or U13694 (N_13694,N_10216,N_8582);
xor U13695 (N_13695,N_11878,N_9540);
or U13696 (N_13696,N_10566,N_9174);
or U13697 (N_13697,N_9924,N_11958);
and U13698 (N_13698,N_9319,N_10614);
nand U13699 (N_13699,N_10412,N_10887);
and U13700 (N_13700,N_9166,N_11617);
xor U13701 (N_13701,N_11085,N_8661);
nand U13702 (N_13702,N_10619,N_8578);
xnor U13703 (N_13703,N_10572,N_11539);
nor U13704 (N_13704,N_8005,N_9843);
or U13705 (N_13705,N_9415,N_11121);
or U13706 (N_13706,N_9198,N_9702);
nand U13707 (N_13707,N_11897,N_8664);
or U13708 (N_13708,N_11858,N_11296);
xnor U13709 (N_13709,N_9125,N_8547);
or U13710 (N_13710,N_8830,N_11170);
xnor U13711 (N_13711,N_10364,N_9249);
xor U13712 (N_13712,N_8521,N_8900);
and U13713 (N_13713,N_10675,N_10550);
nor U13714 (N_13714,N_10154,N_11305);
nand U13715 (N_13715,N_9334,N_8992);
or U13716 (N_13716,N_10709,N_8427);
nand U13717 (N_13717,N_8139,N_9641);
nand U13718 (N_13718,N_11840,N_11735);
nand U13719 (N_13719,N_9845,N_8961);
xor U13720 (N_13720,N_9648,N_11781);
xnor U13721 (N_13721,N_10964,N_8433);
xor U13722 (N_13722,N_11184,N_10413);
or U13723 (N_13723,N_8358,N_8379);
nand U13724 (N_13724,N_9195,N_11986);
nand U13725 (N_13725,N_9285,N_9269);
xnor U13726 (N_13726,N_8159,N_11973);
xnor U13727 (N_13727,N_8576,N_11660);
xor U13728 (N_13728,N_10268,N_10031);
and U13729 (N_13729,N_8093,N_11215);
or U13730 (N_13730,N_8098,N_9932);
nand U13731 (N_13731,N_8995,N_10084);
nor U13732 (N_13732,N_8016,N_9305);
or U13733 (N_13733,N_9790,N_8944);
nor U13734 (N_13734,N_8813,N_9667);
nand U13735 (N_13735,N_8217,N_11807);
nor U13736 (N_13736,N_8128,N_8920);
xnor U13737 (N_13737,N_9559,N_9179);
xnor U13738 (N_13738,N_11845,N_11442);
and U13739 (N_13739,N_9460,N_8275);
nor U13740 (N_13740,N_9809,N_11389);
or U13741 (N_13741,N_11295,N_11409);
nand U13742 (N_13742,N_10314,N_8046);
and U13743 (N_13743,N_11210,N_11956);
xnor U13744 (N_13744,N_11507,N_10341);
and U13745 (N_13745,N_8565,N_9534);
xor U13746 (N_13746,N_10262,N_10968);
and U13747 (N_13747,N_8208,N_10754);
nor U13748 (N_13748,N_9990,N_8386);
xnor U13749 (N_13749,N_10242,N_10310);
nor U13750 (N_13750,N_8287,N_10879);
and U13751 (N_13751,N_10890,N_9156);
and U13752 (N_13752,N_11987,N_10514);
and U13753 (N_13753,N_10987,N_9981);
nand U13754 (N_13754,N_8686,N_11686);
xor U13755 (N_13755,N_10993,N_10226);
and U13756 (N_13756,N_10123,N_10509);
and U13757 (N_13757,N_11819,N_11761);
or U13758 (N_13758,N_9255,N_10919);
and U13759 (N_13759,N_8218,N_11904);
or U13760 (N_13760,N_8249,N_9177);
xor U13761 (N_13761,N_8612,N_11574);
nand U13762 (N_13762,N_10156,N_11341);
nand U13763 (N_13763,N_8101,N_9575);
or U13764 (N_13764,N_8474,N_8499);
nand U13765 (N_13765,N_11955,N_11509);
and U13766 (N_13766,N_10427,N_10187);
xnor U13767 (N_13767,N_11249,N_9261);
nand U13768 (N_13768,N_8952,N_11087);
and U13769 (N_13769,N_9820,N_9287);
xor U13770 (N_13770,N_8238,N_10398);
nor U13771 (N_13771,N_10144,N_8922);
nand U13772 (N_13772,N_9514,N_8980);
nor U13773 (N_13773,N_11474,N_8087);
or U13774 (N_13774,N_8723,N_10554);
or U13775 (N_13775,N_8680,N_10004);
nor U13776 (N_13776,N_8707,N_10766);
nand U13777 (N_13777,N_11207,N_10019);
nand U13778 (N_13778,N_11221,N_11194);
xnor U13779 (N_13779,N_8074,N_8077);
nand U13780 (N_13780,N_8684,N_10430);
xnor U13781 (N_13781,N_8718,N_10702);
and U13782 (N_13782,N_8229,N_10477);
nor U13783 (N_13783,N_9400,N_8593);
nand U13784 (N_13784,N_9557,N_11160);
nor U13785 (N_13785,N_11695,N_11427);
and U13786 (N_13786,N_8979,N_11525);
or U13787 (N_13787,N_11346,N_9197);
and U13788 (N_13788,N_10910,N_10363);
nor U13789 (N_13789,N_10560,N_11909);
and U13790 (N_13790,N_10803,N_10119);
or U13791 (N_13791,N_11270,N_11769);
nand U13792 (N_13792,N_10254,N_11599);
nand U13793 (N_13793,N_8927,N_9453);
nand U13794 (N_13794,N_8440,N_8790);
or U13795 (N_13795,N_10436,N_11515);
or U13796 (N_13796,N_8310,N_11465);
xnor U13797 (N_13797,N_11593,N_8842);
and U13798 (N_13798,N_8308,N_8692);
or U13799 (N_13799,N_10823,N_10691);
nand U13800 (N_13800,N_10975,N_9025);
and U13801 (N_13801,N_11253,N_10158);
or U13802 (N_13802,N_11749,N_8589);
xnor U13803 (N_13803,N_10610,N_9972);
and U13804 (N_13804,N_11423,N_9169);
nor U13805 (N_13805,N_10220,N_9529);
nand U13806 (N_13806,N_11374,N_11494);
or U13807 (N_13807,N_11344,N_8825);
nand U13808 (N_13808,N_10500,N_11113);
or U13809 (N_13809,N_8051,N_8475);
nand U13810 (N_13810,N_10599,N_11528);
nor U13811 (N_13811,N_10067,N_9942);
or U13812 (N_13812,N_11511,N_9950);
xnor U13813 (N_13813,N_10986,N_9988);
xor U13814 (N_13814,N_10075,N_9435);
nor U13815 (N_13815,N_9591,N_8761);
nand U13816 (N_13816,N_8930,N_10370);
nand U13817 (N_13817,N_10244,N_11190);
nand U13818 (N_13818,N_10530,N_11147);
xnor U13819 (N_13819,N_9404,N_11146);
xnor U13820 (N_13820,N_11573,N_10807);
nand U13821 (N_13821,N_9860,N_10306);
and U13822 (N_13822,N_9295,N_10160);
xor U13823 (N_13823,N_10058,N_9626);
and U13824 (N_13824,N_10489,N_9440);
or U13825 (N_13825,N_9880,N_10937);
and U13826 (N_13826,N_8663,N_8902);
nor U13827 (N_13827,N_9582,N_8022);
and U13828 (N_13828,N_11094,N_10275);
and U13829 (N_13829,N_11755,N_8121);
and U13830 (N_13830,N_11401,N_8119);
and U13831 (N_13831,N_9383,N_8595);
xor U13832 (N_13832,N_9896,N_8600);
or U13833 (N_13833,N_11408,N_10360);
nand U13834 (N_13834,N_9377,N_10750);
xnor U13835 (N_13835,N_9337,N_10377);
xnor U13836 (N_13836,N_11516,N_9039);
or U13837 (N_13837,N_11236,N_9365);
nand U13838 (N_13838,N_9001,N_11222);
or U13839 (N_13839,N_8577,N_10726);
xnor U13840 (N_13840,N_8918,N_11924);
nand U13841 (N_13841,N_8777,N_10949);
xor U13842 (N_13842,N_11171,N_9938);
nor U13843 (N_13843,N_10453,N_9359);
nand U13844 (N_13844,N_11853,N_9565);
nor U13845 (N_13845,N_10985,N_10842);
xnor U13846 (N_13846,N_9349,N_9069);
and U13847 (N_13847,N_9996,N_11268);
nor U13848 (N_13848,N_11641,N_9071);
or U13849 (N_13849,N_11499,N_8621);
nor U13850 (N_13850,N_10199,N_8642);
and U13851 (N_13851,N_8352,N_11558);
nand U13852 (N_13852,N_9573,N_9539);
nand U13853 (N_13853,N_9485,N_8568);
xor U13854 (N_13854,N_11440,N_8388);
nand U13855 (N_13855,N_10240,N_8177);
nor U13856 (N_13856,N_8598,N_8439);
or U13857 (N_13857,N_11012,N_10837);
xnor U13858 (N_13858,N_9421,N_8901);
xor U13859 (N_13859,N_10770,N_8802);
nand U13860 (N_13860,N_8382,N_11129);
and U13861 (N_13861,N_10518,N_8045);
nand U13862 (N_13862,N_9403,N_8413);
nor U13863 (N_13863,N_9432,N_9014);
nand U13864 (N_13864,N_10703,N_8835);
xnor U13865 (N_13865,N_9139,N_8318);
nand U13866 (N_13866,N_9885,N_9348);
or U13867 (N_13867,N_11367,N_8317);
nand U13868 (N_13868,N_11654,N_9147);
nand U13869 (N_13869,N_9089,N_8076);
xnor U13870 (N_13870,N_10232,N_10259);
xnor U13871 (N_13871,N_10256,N_8100);
nor U13872 (N_13872,N_8544,N_9638);
or U13873 (N_13873,N_10086,N_8021);
nand U13874 (N_13874,N_11811,N_9306);
and U13875 (N_13875,N_8090,N_8026);
nor U13876 (N_13876,N_10013,N_10869);
and U13877 (N_13877,N_10961,N_11903);
xor U13878 (N_13878,N_10417,N_9517);
nand U13879 (N_13879,N_11266,N_10064);
xor U13880 (N_13880,N_9035,N_9063);
xor U13881 (N_13881,N_9237,N_9979);
or U13882 (N_13882,N_9939,N_9668);
or U13883 (N_13883,N_11033,N_8307);
nand U13884 (N_13884,N_11493,N_8365);
nor U13885 (N_13885,N_10906,N_9893);
xor U13886 (N_13886,N_10568,N_10260);
nor U13887 (N_13887,N_10548,N_10574);
or U13888 (N_13888,N_11425,N_9664);
nand U13889 (N_13889,N_11053,N_10402);
and U13890 (N_13890,N_11355,N_8070);
nand U13891 (N_13891,N_10561,N_8199);
nor U13892 (N_13892,N_8556,N_9087);
or U13893 (N_13893,N_10991,N_9343);
xnor U13894 (N_13894,N_11576,N_10132);
and U13895 (N_13895,N_9904,N_8571);
xnor U13896 (N_13896,N_10577,N_9468);
nor U13897 (N_13897,N_8343,N_10113);
xnor U13898 (N_13898,N_8785,N_9806);
xor U13899 (N_13899,N_8018,N_9735);
nand U13900 (N_13900,N_8525,N_11759);
xor U13901 (N_13901,N_10134,N_11130);
or U13902 (N_13902,N_8942,N_11623);
nand U13903 (N_13903,N_9973,N_8445);
nand U13904 (N_13904,N_10201,N_10355);
and U13905 (N_13905,N_8573,N_10168);
nor U13906 (N_13906,N_8515,N_11554);
and U13907 (N_13907,N_8681,N_8431);
and U13908 (N_13908,N_10437,N_11885);
and U13909 (N_13909,N_9660,N_9522);
and U13910 (N_13910,N_11691,N_11462);
and U13911 (N_13911,N_10758,N_9189);
xor U13912 (N_13912,N_9066,N_9109);
nand U13913 (N_13913,N_11882,N_8877);
and U13914 (N_13914,N_11581,N_11935);
xnor U13915 (N_13915,N_8981,N_11545);
nand U13916 (N_13916,N_8879,N_10234);
and U13917 (N_13917,N_9955,N_10271);
or U13918 (N_13918,N_10531,N_9720);
and U13919 (N_13919,N_11651,N_11946);
nor U13920 (N_13920,N_9022,N_9312);
xnor U13921 (N_13921,N_10828,N_8350);
nor U13922 (N_13922,N_10936,N_9386);
nand U13923 (N_13923,N_8162,N_10713);
nor U13924 (N_13924,N_10683,N_11790);
xor U13925 (N_13925,N_8010,N_11301);
and U13926 (N_13926,N_8845,N_9980);
nand U13927 (N_13927,N_8530,N_8837);
or U13928 (N_13928,N_8341,N_11112);
or U13929 (N_13929,N_10420,N_9286);
or U13930 (N_13930,N_11771,N_9368);
and U13931 (N_13931,N_9258,N_11738);
nand U13932 (N_13932,N_11282,N_10038);
nor U13933 (N_13933,N_9277,N_11046);
and U13934 (N_13934,N_9317,N_9196);
nand U13935 (N_13935,N_11637,N_8491);
or U13936 (N_13936,N_9832,N_9278);
nor U13937 (N_13937,N_10866,N_9865);
and U13938 (N_13938,N_11106,N_8974);
and U13939 (N_13939,N_10447,N_8164);
xnor U13940 (N_13940,N_11527,N_8102);
and U13941 (N_13941,N_11887,N_10778);
or U13942 (N_13942,N_9876,N_10609);
and U13943 (N_13943,N_8180,N_8507);
xor U13944 (N_13944,N_11913,N_10304);
or U13945 (N_13945,N_8200,N_11199);
xnor U13946 (N_13946,N_8311,N_8716);
and U13947 (N_13947,N_9878,N_8639);
or U13948 (N_13948,N_8143,N_11817);
nor U13949 (N_13949,N_8923,N_8554);
xnor U13950 (N_13950,N_10571,N_11420);
nor U13951 (N_13951,N_10193,N_10597);
nor U13952 (N_13952,N_8136,N_9549);
nand U13953 (N_13953,N_8763,N_11030);
nor U13954 (N_13954,N_9803,N_10953);
nand U13955 (N_13955,N_10846,N_9327);
or U13956 (N_13956,N_11396,N_9341);
nor U13957 (N_13957,N_11384,N_10390);
xor U13958 (N_13958,N_8165,N_8611);
nand U13959 (N_13959,N_11216,N_8168);
or U13960 (N_13960,N_11064,N_8697);
xnor U13961 (N_13961,N_9406,N_10707);
nand U13962 (N_13962,N_11586,N_8339);
nand U13963 (N_13963,N_11692,N_11743);
xor U13964 (N_13964,N_9989,N_8947);
or U13965 (N_13965,N_10155,N_11052);
nor U13966 (N_13966,N_8734,N_10855);
nor U13967 (N_13967,N_8281,N_11726);
nand U13968 (N_13968,N_9211,N_11298);
nor U13969 (N_13969,N_11476,N_11120);
nand U13970 (N_13970,N_8803,N_8819);
and U13971 (N_13971,N_8146,N_10052);
xnor U13972 (N_13972,N_11942,N_8858);
nand U13973 (N_13973,N_11941,N_8460);
and U13974 (N_13974,N_10544,N_10188);
xor U13975 (N_13975,N_10579,N_9858);
and U13976 (N_13976,N_11099,N_9982);
nand U13977 (N_13977,N_8434,N_9032);
or U13978 (N_13978,N_8110,N_11591);
or U13979 (N_13979,N_8429,N_9413);
or U13980 (N_13980,N_11080,N_10165);
or U13981 (N_13981,N_9589,N_10727);
nor U13982 (N_13982,N_10712,N_10764);
or U13983 (N_13983,N_9067,N_8607);
nand U13984 (N_13984,N_10359,N_11102);
and U13985 (N_13985,N_8747,N_10261);
nor U13986 (N_13986,N_10503,N_11161);
nand U13987 (N_13987,N_8564,N_9270);
nor U13988 (N_13988,N_10089,N_10679);
and U13989 (N_13989,N_11919,N_11483);
nor U13990 (N_13990,N_11002,N_10974);
and U13991 (N_13991,N_9519,N_9215);
xnor U13992 (N_13992,N_9303,N_9954);
or U13993 (N_13993,N_11621,N_8188);
nor U13994 (N_13994,N_10528,N_9235);
or U13995 (N_13995,N_9398,N_8469);
xnor U13996 (N_13996,N_11403,N_8336);
nand U13997 (N_13997,N_10150,N_9639);
nand U13998 (N_13998,N_9185,N_11923);
nand U13999 (N_13999,N_10779,N_9053);
nand U14000 (N_14000,N_11944,N_11986);
nand U14001 (N_14001,N_9454,N_10284);
and U14002 (N_14002,N_9630,N_11107);
nor U14003 (N_14003,N_10620,N_11372);
or U14004 (N_14004,N_10926,N_9913);
or U14005 (N_14005,N_11353,N_11125);
xor U14006 (N_14006,N_10306,N_8918);
and U14007 (N_14007,N_9353,N_10422);
xor U14008 (N_14008,N_11550,N_8502);
or U14009 (N_14009,N_8301,N_8048);
nor U14010 (N_14010,N_11158,N_11055);
nor U14011 (N_14011,N_8068,N_9745);
or U14012 (N_14012,N_11267,N_8921);
or U14013 (N_14013,N_10464,N_9834);
or U14014 (N_14014,N_10374,N_8965);
and U14015 (N_14015,N_8379,N_9955);
xnor U14016 (N_14016,N_9122,N_9779);
nand U14017 (N_14017,N_9504,N_8207);
or U14018 (N_14018,N_11801,N_11309);
and U14019 (N_14019,N_11237,N_9760);
and U14020 (N_14020,N_11300,N_8517);
and U14021 (N_14021,N_10369,N_8669);
and U14022 (N_14022,N_8168,N_8854);
nand U14023 (N_14023,N_11787,N_9610);
and U14024 (N_14024,N_9858,N_8711);
or U14025 (N_14025,N_9639,N_9183);
and U14026 (N_14026,N_10105,N_8107);
or U14027 (N_14027,N_8810,N_9645);
or U14028 (N_14028,N_8724,N_8243);
and U14029 (N_14029,N_9121,N_10103);
nor U14030 (N_14030,N_10760,N_11551);
or U14031 (N_14031,N_9538,N_10780);
and U14032 (N_14032,N_10359,N_8789);
nor U14033 (N_14033,N_9514,N_8438);
nand U14034 (N_14034,N_9860,N_9544);
nor U14035 (N_14035,N_8667,N_11375);
nand U14036 (N_14036,N_8446,N_10286);
or U14037 (N_14037,N_8526,N_9368);
nand U14038 (N_14038,N_10714,N_10868);
or U14039 (N_14039,N_9635,N_9215);
xnor U14040 (N_14040,N_11110,N_10802);
or U14041 (N_14041,N_11748,N_11011);
nand U14042 (N_14042,N_8139,N_11615);
or U14043 (N_14043,N_11543,N_8085);
xor U14044 (N_14044,N_9199,N_8863);
nor U14045 (N_14045,N_11240,N_8296);
nor U14046 (N_14046,N_10419,N_9539);
and U14047 (N_14047,N_9961,N_10700);
nor U14048 (N_14048,N_9526,N_11605);
or U14049 (N_14049,N_11212,N_10727);
and U14050 (N_14050,N_8244,N_8181);
nor U14051 (N_14051,N_8161,N_8553);
xnor U14052 (N_14052,N_11952,N_11981);
nand U14053 (N_14053,N_9904,N_8503);
nor U14054 (N_14054,N_9661,N_10507);
or U14055 (N_14055,N_8954,N_10745);
and U14056 (N_14056,N_9639,N_9976);
and U14057 (N_14057,N_9314,N_11359);
nor U14058 (N_14058,N_8287,N_8390);
or U14059 (N_14059,N_10671,N_9412);
nor U14060 (N_14060,N_11729,N_8164);
xor U14061 (N_14061,N_8612,N_9760);
xor U14062 (N_14062,N_9337,N_8924);
xor U14063 (N_14063,N_11254,N_8890);
xor U14064 (N_14064,N_9332,N_8837);
nor U14065 (N_14065,N_11578,N_10221);
or U14066 (N_14066,N_9356,N_11446);
nand U14067 (N_14067,N_8628,N_11191);
nor U14068 (N_14068,N_10120,N_11047);
nor U14069 (N_14069,N_8980,N_10152);
nand U14070 (N_14070,N_9036,N_11499);
xnor U14071 (N_14071,N_10671,N_11247);
xnor U14072 (N_14072,N_9880,N_9789);
nand U14073 (N_14073,N_8923,N_11405);
and U14074 (N_14074,N_8320,N_10134);
xor U14075 (N_14075,N_8005,N_8806);
nor U14076 (N_14076,N_9998,N_9959);
or U14077 (N_14077,N_11093,N_11425);
and U14078 (N_14078,N_11936,N_9867);
and U14079 (N_14079,N_11040,N_10430);
nand U14080 (N_14080,N_9000,N_11450);
and U14081 (N_14081,N_8588,N_11345);
and U14082 (N_14082,N_10174,N_11386);
or U14083 (N_14083,N_8904,N_10707);
and U14084 (N_14084,N_10889,N_8076);
nor U14085 (N_14085,N_11385,N_11144);
and U14086 (N_14086,N_10609,N_10053);
or U14087 (N_14087,N_11183,N_8982);
or U14088 (N_14088,N_8966,N_10458);
xor U14089 (N_14089,N_8050,N_9521);
or U14090 (N_14090,N_9112,N_11052);
nand U14091 (N_14091,N_10035,N_9489);
and U14092 (N_14092,N_10985,N_10730);
xnor U14093 (N_14093,N_8255,N_11498);
nor U14094 (N_14094,N_11268,N_8981);
xnor U14095 (N_14095,N_10516,N_11960);
nand U14096 (N_14096,N_9239,N_11339);
nor U14097 (N_14097,N_8502,N_9374);
nor U14098 (N_14098,N_10376,N_9352);
xnor U14099 (N_14099,N_9367,N_11529);
or U14100 (N_14100,N_9142,N_10229);
xor U14101 (N_14101,N_9970,N_8821);
and U14102 (N_14102,N_8625,N_10000);
and U14103 (N_14103,N_10407,N_11548);
or U14104 (N_14104,N_9404,N_10140);
and U14105 (N_14105,N_10053,N_8060);
and U14106 (N_14106,N_10366,N_11110);
xor U14107 (N_14107,N_10827,N_8634);
xor U14108 (N_14108,N_11051,N_10323);
nand U14109 (N_14109,N_11510,N_10773);
or U14110 (N_14110,N_9112,N_9077);
xor U14111 (N_14111,N_8186,N_9415);
xnor U14112 (N_14112,N_8667,N_9065);
nand U14113 (N_14113,N_11784,N_11212);
and U14114 (N_14114,N_11459,N_8295);
nand U14115 (N_14115,N_10087,N_10189);
nor U14116 (N_14116,N_11700,N_11510);
or U14117 (N_14117,N_8177,N_11826);
nor U14118 (N_14118,N_8202,N_8805);
nand U14119 (N_14119,N_11902,N_8874);
nand U14120 (N_14120,N_8767,N_8816);
nor U14121 (N_14121,N_8076,N_10297);
nand U14122 (N_14122,N_8408,N_9687);
nand U14123 (N_14123,N_8136,N_10351);
and U14124 (N_14124,N_10263,N_10845);
nand U14125 (N_14125,N_9430,N_11143);
and U14126 (N_14126,N_8417,N_10785);
nand U14127 (N_14127,N_10964,N_11529);
xnor U14128 (N_14128,N_10682,N_9438);
nand U14129 (N_14129,N_9268,N_9105);
xnor U14130 (N_14130,N_8249,N_9089);
or U14131 (N_14131,N_11668,N_10680);
and U14132 (N_14132,N_11607,N_11326);
or U14133 (N_14133,N_10998,N_11908);
xnor U14134 (N_14134,N_10471,N_8554);
and U14135 (N_14135,N_10265,N_9768);
xnor U14136 (N_14136,N_9322,N_9252);
xnor U14137 (N_14137,N_10342,N_11974);
nand U14138 (N_14138,N_8908,N_11166);
nor U14139 (N_14139,N_10226,N_11092);
xnor U14140 (N_14140,N_9142,N_9309);
nand U14141 (N_14141,N_11270,N_8032);
xor U14142 (N_14142,N_11049,N_8331);
or U14143 (N_14143,N_9719,N_10724);
and U14144 (N_14144,N_8870,N_10774);
nor U14145 (N_14145,N_10240,N_8355);
nor U14146 (N_14146,N_9839,N_10518);
or U14147 (N_14147,N_8600,N_10729);
nor U14148 (N_14148,N_9094,N_10516);
nand U14149 (N_14149,N_10288,N_8311);
or U14150 (N_14150,N_10015,N_9163);
and U14151 (N_14151,N_9202,N_8035);
nor U14152 (N_14152,N_8928,N_10141);
nor U14153 (N_14153,N_10034,N_10757);
nand U14154 (N_14154,N_10680,N_9704);
or U14155 (N_14155,N_9282,N_11317);
xor U14156 (N_14156,N_11687,N_11226);
nor U14157 (N_14157,N_8993,N_9923);
or U14158 (N_14158,N_11766,N_9017);
and U14159 (N_14159,N_9157,N_9912);
and U14160 (N_14160,N_10956,N_9690);
nand U14161 (N_14161,N_9379,N_11849);
nor U14162 (N_14162,N_11003,N_10919);
and U14163 (N_14163,N_10205,N_10887);
xnor U14164 (N_14164,N_11222,N_9358);
and U14165 (N_14165,N_11844,N_8826);
nand U14166 (N_14166,N_10217,N_9719);
or U14167 (N_14167,N_8892,N_8931);
nor U14168 (N_14168,N_9628,N_9205);
nand U14169 (N_14169,N_11742,N_11374);
nand U14170 (N_14170,N_10654,N_9739);
xnor U14171 (N_14171,N_8927,N_8598);
xor U14172 (N_14172,N_11482,N_10262);
nor U14173 (N_14173,N_11087,N_10274);
nand U14174 (N_14174,N_10968,N_10403);
nor U14175 (N_14175,N_11225,N_8696);
or U14176 (N_14176,N_9483,N_8694);
and U14177 (N_14177,N_8406,N_11664);
nor U14178 (N_14178,N_8611,N_8881);
or U14179 (N_14179,N_10983,N_10402);
or U14180 (N_14180,N_8829,N_9947);
nand U14181 (N_14181,N_9920,N_9574);
nor U14182 (N_14182,N_10203,N_9349);
or U14183 (N_14183,N_8182,N_11204);
xnor U14184 (N_14184,N_8634,N_11635);
nor U14185 (N_14185,N_8384,N_11283);
and U14186 (N_14186,N_10638,N_8168);
xor U14187 (N_14187,N_8740,N_9792);
xnor U14188 (N_14188,N_8898,N_11210);
nand U14189 (N_14189,N_9738,N_11804);
nor U14190 (N_14190,N_10854,N_8643);
xnor U14191 (N_14191,N_8318,N_8579);
nor U14192 (N_14192,N_8661,N_9865);
nor U14193 (N_14193,N_10824,N_8848);
nor U14194 (N_14194,N_10361,N_9586);
or U14195 (N_14195,N_8994,N_11142);
nor U14196 (N_14196,N_8270,N_11931);
or U14197 (N_14197,N_8185,N_8462);
xnor U14198 (N_14198,N_11137,N_10846);
xnor U14199 (N_14199,N_8796,N_11240);
and U14200 (N_14200,N_10016,N_9549);
or U14201 (N_14201,N_11661,N_8071);
and U14202 (N_14202,N_8693,N_9608);
xor U14203 (N_14203,N_8670,N_10671);
or U14204 (N_14204,N_8079,N_8433);
nand U14205 (N_14205,N_11222,N_8759);
nor U14206 (N_14206,N_10946,N_9913);
xor U14207 (N_14207,N_11666,N_10371);
or U14208 (N_14208,N_11451,N_11676);
and U14209 (N_14209,N_10082,N_11988);
and U14210 (N_14210,N_8920,N_8342);
xnor U14211 (N_14211,N_9437,N_8612);
and U14212 (N_14212,N_11898,N_10619);
nor U14213 (N_14213,N_10971,N_10101);
nor U14214 (N_14214,N_11526,N_11179);
or U14215 (N_14215,N_11254,N_9703);
nor U14216 (N_14216,N_10796,N_9181);
and U14217 (N_14217,N_10080,N_9539);
or U14218 (N_14218,N_11690,N_8493);
and U14219 (N_14219,N_8294,N_10928);
and U14220 (N_14220,N_10591,N_11360);
and U14221 (N_14221,N_10640,N_10908);
xor U14222 (N_14222,N_9339,N_9648);
nand U14223 (N_14223,N_9785,N_10052);
and U14224 (N_14224,N_9943,N_9098);
and U14225 (N_14225,N_10629,N_11063);
nor U14226 (N_14226,N_10657,N_11698);
xnor U14227 (N_14227,N_8814,N_8257);
or U14228 (N_14228,N_8943,N_9540);
and U14229 (N_14229,N_8315,N_8374);
xor U14230 (N_14230,N_10649,N_10948);
xor U14231 (N_14231,N_8211,N_8852);
nor U14232 (N_14232,N_10231,N_8479);
or U14233 (N_14233,N_8926,N_8108);
nand U14234 (N_14234,N_10616,N_11408);
or U14235 (N_14235,N_10446,N_11352);
nor U14236 (N_14236,N_10484,N_11132);
xnor U14237 (N_14237,N_9975,N_11708);
nand U14238 (N_14238,N_10267,N_9598);
xor U14239 (N_14239,N_10566,N_8314);
nand U14240 (N_14240,N_9064,N_11618);
nor U14241 (N_14241,N_9651,N_8118);
nor U14242 (N_14242,N_8623,N_10517);
nand U14243 (N_14243,N_11554,N_10563);
and U14244 (N_14244,N_11148,N_10777);
xnor U14245 (N_14245,N_9010,N_9112);
nor U14246 (N_14246,N_8866,N_9022);
or U14247 (N_14247,N_9284,N_9755);
or U14248 (N_14248,N_9627,N_9280);
or U14249 (N_14249,N_9918,N_10379);
or U14250 (N_14250,N_11765,N_8503);
nand U14251 (N_14251,N_8606,N_10223);
and U14252 (N_14252,N_9575,N_9970);
and U14253 (N_14253,N_10970,N_11400);
and U14254 (N_14254,N_8619,N_9577);
nor U14255 (N_14255,N_8732,N_9261);
xnor U14256 (N_14256,N_11494,N_9837);
nand U14257 (N_14257,N_11986,N_8228);
and U14258 (N_14258,N_10673,N_10370);
and U14259 (N_14259,N_9821,N_11735);
nand U14260 (N_14260,N_10621,N_9586);
nor U14261 (N_14261,N_11613,N_10449);
or U14262 (N_14262,N_8335,N_9584);
nand U14263 (N_14263,N_8979,N_8022);
or U14264 (N_14264,N_9955,N_11947);
or U14265 (N_14265,N_8888,N_10505);
and U14266 (N_14266,N_10819,N_11176);
and U14267 (N_14267,N_11032,N_11707);
xor U14268 (N_14268,N_9305,N_8169);
and U14269 (N_14269,N_9713,N_11582);
or U14270 (N_14270,N_9101,N_8775);
nand U14271 (N_14271,N_10139,N_9968);
or U14272 (N_14272,N_10429,N_11885);
nor U14273 (N_14273,N_9081,N_9926);
or U14274 (N_14274,N_9130,N_9260);
and U14275 (N_14275,N_10213,N_9277);
and U14276 (N_14276,N_11604,N_10718);
nand U14277 (N_14277,N_8000,N_9131);
or U14278 (N_14278,N_10768,N_8715);
nor U14279 (N_14279,N_10267,N_9685);
nand U14280 (N_14280,N_8829,N_11514);
xor U14281 (N_14281,N_9038,N_9218);
or U14282 (N_14282,N_8334,N_9918);
and U14283 (N_14283,N_9006,N_10138);
nor U14284 (N_14284,N_10478,N_8621);
nand U14285 (N_14285,N_11468,N_9456);
or U14286 (N_14286,N_8144,N_10814);
and U14287 (N_14287,N_10667,N_11673);
and U14288 (N_14288,N_8702,N_10473);
xor U14289 (N_14289,N_9337,N_11129);
xor U14290 (N_14290,N_10963,N_8208);
xor U14291 (N_14291,N_11652,N_11839);
and U14292 (N_14292,N_9231,N_9819);
nor U14293 (N_14293,N_10253,N_9726);
xnor U14294 (N_14294,N_11032,N_11525);
nand U14295 (N_14295,N_10691,N_10722);
and U14296 (N_14296,N_11010,N_9311);
nand U14297 (N_14297,N_11359,N_11527);
nand U14298 (N_14298,N_9784,N_10350);
and U14299 (N_14299,N_11949,N_9821);
nand U14300 (N_14300,N_11806,N_8277);
xnor U14301 (N_14301,N_10878,N_10544);
or U14302 (N_14302,N_10904,N_11121);
xnor U14303 (N_14303,N_11427,N_8756);
nand U14304 (N_14304,N_9928,N_10908);
and U14305 (N_14305,N_8636,N_8107);
or U14306 (N_14306,N_8754,N_11296);
and U14307 (N_14307,N_10750,N_9862);
nor U14308 (N_14308,N_9994,N_9118);
or U14309 (N_14309,N_8153,N_9544);
nor U14310 (N_14310,N_10499,N_9653);
or U14311 (N_14311,N_9951,N_8682);
xor U14312 (N_14312,N_11374,N_9445);
nand U14313 (N_14313,N_11583,N_10270);
or U14314 (N_14314,N_9605,N_9906);
nand U14315 (N_14315,N_11132,N_11330);
xnor U14316 (N_14316,N_9467,N_8591);
xnor U14317 (N_14317,N_10003,N_11145);
nor U14318 (N_14318,N_11526,N_10122);
and U14319 (N_14319,N_11406,N_11982);
xor U14320 (N_14320,N_9111,N_10318);
or U14321 (N_14321,N_8031,N_11455);
xnor U14322 (N_14322,N_8505,N_11163);
xnor U14323 (N_14323,N_8841,N_8904);
xnor U14324 (N_14324,N_11509,N_11063);
xor U14325 (N_14325,N_11498,N_10018);
nor U14326 (N_14326,N_9783,N_10418);
and U14327 (N_14327,N_11163,N_10776);
nand U14328 (N_14328,N_8803,N_11389);
xor U14329 (N_14329,N_11099,N_10795);
xor U14330 (N_14330,N_9442,N_11318);
xnor U14331 (N_14331,N_11437,N_10620);
nand U14332 (N_14332,N_9898,N_9677);
xnor U14333 (N_14333,N_10791,N_10261);
or U14334 (N_14334,N_10883,N_8544);
and U14335 (N_14335,N_10857,N_9338);
xor U14336 (N_14336,N_10992,N_11796);
and U14337 (N_14337,N_10351,N_8147);
nand U14338 (N_14338,N_10051,N_9545);
xor U14339 (N_14339,N_11730,N_9836);
nor U14340 (N_14340,N_9644,N_11247);
nand U14341 (N_14341,N_8614,N_11838);
or U14342 (N_14342,N_11808,N_9472);
nor U14343 (N_14343,N_9676,N_11130);
nor U14344 (N_14344,N_9048,N_11795);
or U14345 (N_14345,N_9837,N_9304);
xnor U14346 (N_14346,N_8070,N_11167);
and U14347 (N_14347,N_8881,N_11258);
nand U14348 (N_14348,N_11828,N_10579);
nor U14349 (N_14349,N_10294,N_10506);
nand U14350 (N_14350,N_10860,N_9341);
xor U14351 (N_14351,N_9334,N_9450);
and U14352 (N_14352,N_11512,N_8741);
nand U14353 (N_14353,N_10791,N_8804);
xnor U14354 (N_14354,N_11653,N_9602);
nor U14355 (N_14355,N_11496,N_11743);
nand U14356 (N_14356,N_10901,N_10312);
nand U14357 (N_14357,N_9587,N_10113);
or U14358 (N_14358,N_11781,N_9629);
or U14359 (N_14359,N_10114,N_11794);
or U14360 (N_14360,N_11606,N_8434);
or U14361 (N_14361,N_10844,N_11807);
nand U14362 (N_14362,N_11947,N_8605);
xor U14363 (N_14363,N_9787,N_9221);
nand U14364 (N_14364,N_9390,N_10944);
and U14365 (N_14365,N_11619,N_9689);
or U14366 (N_14366,N_11268,N_8757);
or U14367 (N_14367,N_11426,N_9771);
xor U14368 (N_14368,N_9299,N_9041);
xnor U14369 (N_14369,N_9000,N_9300);
nor U14370 (N_14370,N_10188,N_8391);
xor U14371 (N_14371,N_11548,N_9887);
nand U14372 (N_14372,N_11331,N_9389);
nor U14373 (N_14373,N_9479,N_10006);
nand U14374 (N_14374,N_9773,N_8117);
and U14375 (N_14375,N_8641,N_9307);
xnor U14376 (N_14376,N_9375,N_9873);
nor U14377 (N_14377,N_10693,N_9177);
nand U14378 (N_14378,N_8129,N_8701);
nor U14379 (N_14379,N_8064,N_9325);
nor U14380 (N_14380,N_11510,N_9492);
or U14381 (N_14381,N_11633,N_9586);
and U14382 (N_14382,N_8923,N_11937);
and U14383 (N_14383,N_9966,N_8434);
nand U14384 (N_14384,N_8212,N_11145);
nor U14385 (N_14385,N_8943,N_11894);
xor U14386 (N_14386,N_10745,N_11868);
xnor U14387 (N_14387,N_9240,N_9810);
xor U14388 (N_14388,N_11145,N_9751);
or U14389 (N_14389,N_10553,N_8775);
nor U14390 (N_14390,N_9825,N_9104);
or U14391 (N_14391,N_10817,N_10809);
xor U14392 (N_14392,N_10709,N_9870);
nor U14393 (N_14393,N_11816,N_9312);
or U14394 (N_14394,N_10956,N_10905);
xor U14395 (N_14395,N_11767,N_11162);
nand U14396 (N_14396,N_9445,N_8078);
nor U14397 (N_14397,N_10793,N_9732);
nand U14398 (N_14398,N_9096,N_10450);
and U14399 (N_14399,N_11849,N_10414);
xor U14400 (N_14400,N_11816,N_10132);
nor U14401 (N_14401,N_10435,N_10733);
or U14402 (N_14402,N_9967,N_10150);
nand U14403 (N_14403,N_10038,N_10512);
nand U14404 (N_14404,N_10209,N_9358);
and U14405 (N_14405,N_10461,N_10850);
or U14406 (N_14406,N_8105,N_9196);
nand U14407 (N_14407,N_11568,N_9621);
nand U14408 (N_14408,N_8978,N_10420);
or U14409 (N_14409,N_9868,N_11720);
nand U14410 (N_14410,N_11991,N_10125);
or U14411 (N_14411,N_11065,N_10587);
nor U14412 (N_14412,N_9662,N_8272);
nand U14413 (N_14413,N_8193,N_11438);
or U14414 (N_14414,N_10838,N_11948);
or U14415 (N_14415,N_11028,N_11881);
nand U14416 (N_14416,N_11673,N_9092);
and U14417 (N_14417,N_11004,N_11852);
xnor U14418 (N_14418,N_8207,N_9568);
xnor U14419 (N_14419,N_11888,N_8485);
nor U14420 (N_14420,N_9244,N_10038);
and U14421 (N_14421,N_9860,N_9589);
and U14422 (N_14422,N_10462,N_10190);
or U14423 (N_14423,N_10219,N_9429);
or U14424 (N_14424,N_10334,N_8714);
or U14425 (N_14425,N_9326,N_9926);
nor U14426 (N_14426,N_10215,N_10185);
or U14427 (N_14427,N_11479,N_10594);
nand U14428 (N_14428,N_11942,N_11850);
nand U14429 (N_14429,N_11166,N_8212);
xor U14430 (N_14430,N_8504,N_10880);
nand U14431 (N_14431,N_11867,N_11921);
nor U14432 (N_14432,N_8913,N_9430);
or U14433 (N_14433,N_9532,N_11898);
and U14434 (N_14434,N_8175,N_9969);
xnor U14435 (N_14435,N_10513,N_11176);
and U14436 (N_14436,N_9309,N_8686);
xnor U14437 (N_14437,N_10529,N_8242);
nor U14438 (N_14438,N_11643,N_8507);
nand U14439 (N_14439,N_9552,N_10573);
nor U14440 (N_14440,N_8647,N_10030);
or U14441 (N_14441,N_8682,N_8565);
and U14442 (N_14442,N_10933,N_10879);
xnor U14443 (N_14443,N_10480,N_9133);
and U14444 (N_14444,N_8584,N_11931);
and U14445 (N_14445,N_8859,N_10477);
nor U14446 (N_14446,N_11061,N_11165);
xnor U14447 (N_14447,N_8704,N_9104);
nor U14448 (N_14448,N_9242,N_11740);
nor U14449 (N_14449,N_8081,N_10119);
nor U14450 (N_14450,N_9622,N_9668);
nor U14451 (N_14451,N_9604,N_8989);
nand U14452 (N_14452,N_8348,N_10556);
nand U14453 (N_14453,N_9571,N_9512);
and U14454 (N_14454,N_11012,N_11896);
xnor U14455 (N_14455,N_10017,N_8678);
nor U14456 (N_14456,N_11466,N_9000);
and U14457 (N_14457,N_8927,N_11698);
nand U14458 (N_14458,N_11271,N_9820);
nor U14459 (N_14459,N_11415,N_8993);
and U14460 (N_14460,N_11895,N_9695);
xor U14461 (N_14461,N_10129,N_10793);
nor U14462 (N_14462,N_9488,N_8361);
nor U14463 (N_14463,N_8580,N_10913);
or U14464 (N_14464,N_8465,N_8043);
and U14465 (N_14465,N_8177,N_9732);
nand U14466 (N_14466,N_9739,N_8293);
nand U14467 (N_14467,N_10846,N_8180);
nor U14468 (N_14468,N_8174,N_11074);
and U14469 (N_14469,N_10038,N_8865);
or U14470 (N_14470,N_8307,N_10613);
nor U14471 (N_14471,N_8562,N_11792);
xnor U14472 (N_14472,N_8757,N_10068);
nor U14473 (N_14473,N_9356,N_8141);
xnor U14474 (N_14474,N_8448,N_11278);
or U14475 (N_14475,N_8557,N_10113);
nor U14476 (N_14476,N_11069,N_9311);
nor U14477 (N_14477,N_10154,N_8854);
xor U14478 (N_14478,N_9755,N_10518);
nand U14479 (N_14479,N_8170,N_8693);
nand U14480 (N_14480,N_11463,N_10886);
nor U14481 (N_14481,N_11443,N_8150);
nand U14482 (N_14482,N_11329,N_8891);
nor U14483 (N_14483,N_10282,N_9248);
and U14484 (N_14484,N_11462,N_8374);
nand U14485 (N_14485,N_9211,N_10398);
xnor U14486 (N_14486,N_11968,N_9278);
and U14487 (N_14487,N_10358,N_10092);
and U14488 (N_14488,N_8746,N_10659);
nor U14489 (N_14489,N_8054,N_8891);
or U14490 (N_14490,N_11232,N_8621);
xnor U14491 (N_14491,N_10317,N_10235);
or U14492 (N_14492,N_9874,N_9002);
or U14493 (N_14493,N_8423,N_9678);
nand U14494 (N_14494,N_8789,N_8323);
nand U14495 (N_14495,N_11903,N_10501);
nor U14496 (N_14496,N_11600,N_11601);
nand U14497 (N_14497,N_8516,N_9509);
nor U14498 (N_14498,N_11730,N_9092);
and U14499 (N_14499,N_11619,N_8778);
nand U14500 (N_14500,N_9198,N_8061);
nand U14501 (N_14501,N_8035,N_8193);
xor U14502 (N_14502,N_9592,N_11497);
and U14503 (N_14503,N_11957,N_10907);
or U14504 (N_14504,N_11655,N_11604);
nand U14505 (N_14505,N_10209,N_8731);
nand U14506 (N_14506,N_9696,N_11399);
xnor U14507 (N_14507,N_11875,N_8006);
or U14508 (N_14508,N_10943,N_11235);
and U14509 (N_14509,N_9971,N_11257);
nand U14510 (N_14510,N_8046,N_11201);
nand U14511 (N_14511,N_10078,N_9867);
or U14512 (N_14512,N_8524,N_11046);
or U14513 (N_14513,N_11854,N_10068);
or U14514 (N_14514,N_8587,N_8880);
xnor U14515 (N_14515,N_8436,N_10875);
or U14516 (N_14516,N_9975,N_11228);
nand U14517 (N_14517,N_10357,N_9101);
nor U14518 (N_14518,N_9529,N_8367);
or U14519 (N_14519,N_10938,N_10706);
nand U14520 (N_14520,N_10831,N_9238);
nor U14521 (N_14521,N_9152,N_10903);
or U14522 (N_14522,N_11658,N_9906);
or U14523 (N_14523,N_10398,N_11270);
nand U14524 (N_14524,N_10128,N_10051);
xnor U14525 (N_14525,N_9506,N_11714);
or U14526 (N_14526,N_11336,N_8351);
and U14527 (N_14527,N_8459,N_10455);
nor U14528 (N_14528,N_8355,N_11277);
xor U14529 (N_14529,N_8381,N_9124);
or U14530 (N_14530,N_8050,N_9539);
xnor U14531 (N_14531,N_10590,N_8439);
nor U14532 (N_14532,N_9986,N_11373);
nor U14533 (N_14533,N_11930,N_10431);
xor U14534 (N_14534,N_10275,N_9474);
nor U14535 (N_14535,N_11809,N_8134);
nor U14536 (N_14536,N_11892,N_10382);
or U14537 (N_14537,N_10556,N_10940);
and U14538 (N_14538,N_9106,N_10270);
xor U14539 (N_14539,N_8887,N_9367);
nand U14540 (N_14540,N_10128,N_9966);
nor U14541 (N_14541,N_11350,N_10278);
or U14542 (N_14542,N_10764,N_8639);
or U14543 (N_14543,N_11242,N_8962);
or U14544 (N_14544,N_11465,N_8325);
and U14545 (N_14545,N_9119,N_10656);
or U14546 (N_14546,N_10089,N_8162);
nor U14547 (N_14547,N_9827,N_10826);
xor U14548 (N_14548,N_10584,N_10409);
nand U14549 (N_14549,N_10623,N_8137);
or U14550 (N_14550,N_11624,N_8017);
and U14551 (N_14551,N_8965,N_10923);
or U14552 (N_14552,N_8780,N_8882);
xor U14553 (N_14553,N_10510,N_9239);
and U14554 (N_14554,N_11307,N_11380);
and U14555 (N_14555,N_11840,N_8090);
nand U14556 (N_14556,N_8629,N_9525);
or U14557 (N_14557,N_8455,N_9744);
and U14558 (N_14558,N_8144,N_11943);
nand U14559 (N_14559,N_9380,N_10603);
nand U14560 (N_14560,N_8526,N_8858);
xor U14561 (N_14561,N_11088,N_10411);
nand U14562 (N_14562,N_11110,N_9989);
xor U14563 (N_14563,N_10986,N_8404);
nand U14564 (N_14564,N_11537,N_10882);
xnor U14565 (N_14565,N_8467,N_9270);
xor U14566 (N_14566,N_8228,N_10492);
nand U14567 (N_14567,N_11913,N_8855);
xor U14568 (N_14568,N_8748,N_11859);
or U14569 (N_14569,N_10351,N_10227);
nand U14570 (N_14570,N_11022,N_11559);
nor U14571 (N_14571,N_10788,N_10509);
nor U14572 (N_14572,N_8593,N_8542);
nor U14573 (N_14573,N_9243,N_11548);
xor U14574 (N_14574,N_8018,N_11342);
and U14575 (N_14575,N_11692,N_9208);
and U14576 (N_14576,N_10543,N_8960);
and U14577 (N_14577,N_9496,N_11993);
nor U14578 (N_14578,N_11640,N_10488);
nand U14579 (N_14579,N_11980,N_9106);
or U14580 (N_14580,N_10848,N_11187);
xor U14581 (N_14581,N_9929,N_9211);
or U14582 (N_14582,N_8932,N_11257);
or U14583 (N_14583,N_11625,N_10920);
nor U14584 (N_14584,N_10265,N_10325);
xnor U14585 (N_14585,N_11327,N_11952);
and U14586 (N_14586,N_11772,N_11130);
nand U14587 (N_14587,N_9541,N_10081);
nor U14588 (N_14588,N_11746,N_9006);
nand U14589 (N_14589,N_10536,N_10303);
or U14590 (N_14590,N_8389,N_11046);
and U14591 (N_14591,N_9865,N_11783);
nand U14592 (N_14592,N_9134,N_9315);
xor U14593 (N_14593,N_9012,N_10794);
nand U14594 (N_14594,N_10653,N_9845);
nand U14595 (N_14595,N_9628,N_9550);
and U14596 (N_14596,N_10506,N_11241);
and U14597 (N_14597,N_10244,N_11598);
or U14598 (N_14598,N_9987,N_10508);
nand U14599 (N_14599,N_10707,N_11276);
nand U14600 (N_14600,N_11488,N_8575);
and U14601 (N_14601,N_10433,N_9184);
xnor U14602 (N_14602,N_9876,N_9745);
xnor U14603 (N_14603,N_10143,N_11498);
or U14604 (N_14604,N_10184,N_9585);
nand U14605 (N_14605,N_8298,N_11319);
nand U14606 (N_14606,N_9526,N_8661);
xnor U14607 (N_14607,N_8093,N_10937);
nand U14608 (N_14608,N_10949,N_11962);
nand U14609 (N_14609,N_8382,N_11592);
and U14610 (N_14610,N_8814,N_10955);
xnor U14611 (N_14611,N_9861,N_8620);
and U14612 (N_14612,N_10060,N_8509);
and U14613 (N_14613,N_11903,N_9911);
or U14614 (N_14614,N_9467,N_11251);
and U14615 (N_14615,N_9623,N_10761);
and U14616 (N_14616,N_8394,N_9017);
nand U14617 (N_14617,N_11892,N_10464);
or U14618 (N_14618,N_9523,N_11143);
or U14619 (N_14619,N_8150,N_10309);
xnor U14620 (N_14620,N_8330,N_10705);
nand U14621 (N_14621,N_8654,N_10350);
or U14622 (N_14622,N_9799,N_9551);
nor U14623 (N_14623,N_8891,N_8111);
xnor U14624 (N_14624,N_8778,N_11761);
nand U14625 (N_14625,N_10481,N_9746);
or U14626 (N_14626,N_10037,N_11611);
xor U14627 (N_14627,N_8533,N_8781);
or U14628 (N_14628,N_9007,N_9133);
nor U14629 (N_14629,N_8668,N_8402);
xor U14630 (N_14630,N_9368,N_9459);
or U14631 (N_14631,N_10653,N_8926);
or U14632 (N_14632,N_11846,N_10025);
nand U14633 (N_14633,N_11474,N_10878);
and U14634 (N_14634,N_10800,N_9968);
nor U14635 (N_14635,N_9503,N_9994);
xor U14636 (N_14636,N_9005,N_11111);
or U14637 (N_14637,N_8358,N_10548);
nand U14638 (N_14638,N_8588,N_11097);
nand U14639 (N_14639,N_9122,N_9169);
and U14640 (N_14640,N_8975,N_8036);
and U14641 (N_14641,N_8960,N_9054);
xor U14642 (N_14642,N_8389,N_8386);
and U14643 (N_14643,N_10606,N_11839);
xor U14644 (N_14644,N_11076,N_9918);
and U14645 (N_14645,N_11231,N_11057);
xor U14646 (N_14646,N_9333,N_11483);
nand U14647 (N_14647,N_8625,N_10281);
nor U14648 (N_14648,N_8736,N_8602);
xor U14649 (N_14649,N_10653,N_10458);
and U14650 (N_14650,N_9926,N_11860);
or U14651 (N_14651,N_9888,N_10895);
nand U14652 (N_14652,N_10103,N_9024);
and U14653 (N_14653,N_10984,N_10788);
or U14654 (N_14654,N_11352,N_8949);
and U14655 (N_14655,N_9637,N_9657);
and U14656 (N_14656,N_9028,N_9202);
or U14657 (N_14657,N_8653,N_8862);
nor U14658 (N_14658,N_8064,N_11184);
nor U14659 (N_14659,N_10118,N_11138);
nor U14660 (N_14660,N_8562,N_9016);
nand U14661 (N_14661,N_9457,N_9172);
nor U14662 (N_14662,N_9993,N_11504);
nor U14663 (N_14663,N_10387,N_8389);
nor U14664 (N_14664,N_10793,N_10564);
xnor U14665 (N_14665,N_9457,N_8500);
nor U14666 (N_14666,N_11180,N_11598);
nor U14667 (N_14667,N_11678,N_11410);
nand U14668 (N_14668,N_8946,N_11039);
xnor U14669 (N_14669,N_10338,N_11206);
nor U14670 (N_14670,N_9909,N_9480);
xnor U14671 (N_14671,N_9460,N_9721);
and U14672 (N_14672,N_8479,N_11360);
nor U14673 (N_14673,N_8297,N_11005);
or U14674 (N_14674,N_9781,N_9209);
or U14675 (N_14675,N_11233,N_9039);
nor U14676 (N_14676,N_11601,N_9994);
xor U14677 (N_14677,N_9333,N_10937);
nand U14678 (N_14678,N_11475,N_9719);
and U14679 (N_14679,N_10797,N_11235);
nand U14680 (N_14680,N_9471,N_9352);
xor U14681 (N_14681,N_10449,N_11050);
xnor U14682 (N_14682,N_10516,N_11380);
nand U14683 (N_14683,N_8174,N_8830);
and U14684 (N_14684,N_10848,N_10177);
and U14685 (N_14685,N_11264,N_11119);
nor U14686 (N_14686,N_11036,N_10010);
or U14687 (N_14687,N_11286,N_9318);
xor U14688 (N_14688,N_8980,N_8265);
and U14689 (N_14689,N_9196,N_11706);
xor U14690 (N_14690,N_8497,N_8794);
and U14691 (N_14691,N_9095,N_10910);
nor U14692 (N_14692,N_9227,N_9780);
or U14693 (N_14693,N_10733,N_11038);
nor U14694 (N_14694,N_10763,N_10930);
and U14695 (N_14695,N_8779,N_11906);
and U14696 (N_14696,N_11026,N_8541);
or U14697 (N_14697,N_9749,N_10523);
xnor U14698 (N_14698,N_8032,N_11162);
nor U14699 (N_14699,N_9156,N_8807);
and U14700 (N_14700,N_9017,N_10975);
nor U14701 (N_14701,N_11270,N_11803);
nor U14702 (N_14702,N_9854,N_10194);
nor U14703 (N_14703,N_10067,N_9261);
and U14704 (N_14704,N_9234,N_8124);
nand U14705 (N_14705,N_9986,N_11702);
nor U14706 (N_14706,N_11252,N_10061);
nand U14707 (N_14707,N_8520,N_9183);
nor U14708 (N_14708,N_9072,N_8352);
nor U14709 (N_14709,N_11193,N_10029);
nand U14710 (N_14710,N_8878,N_8222);
and U14711 (N_14711,N_10766,N_9120);
xor U14712 (N_14712,N_8810,N_11577);
or U14713 (N_14713,N_9181,N_8604);
nand U14714 (N_14714,N_8001,N_8722);
nor U14715 (N_14715,N_10166,N_10989);
xor U14716 (N_14716,N_11125,N_9183);
nor U14717 (N_14717,N_11355,N_11648);
and U14718 (N_14718,N_10223,N_11807);
nor U14719 (N_14719,N_10369,N_10202);
nor U14720 (N_14720,N_8739,N_11639);
and U14721 (N_14721,N_8149,N_9200);
and U14722 (N_14722,N_8884,N_9208);
nand U14723 (N_14723,N_10483,N_9875);
or U14724 (N_14724,N_9953,N_9671);
xnor U14725 (N_14725,N_10036,N_8329);
or U14726 (N_14726,N_9108,N_9405);
nand U14727 (N_14727,N_11627,N_9367);
xnor U14728 (N_14728,N_8484,N_8080);
nand U14729 (N_14729,N_8086,N_8421);
and U14730 (N_14730,N_9901,N_8033);
or U14731 (N_14731,N_9721,N_8533);
nor U14732 (N_14732,N_11562,N_10085);
nor U14733 (N_14733,N_9671,N_11758);
nor U14734 (N_14734,N_11521,N_8581);
nor U14735 (N_14735,N_10680,N_11621);
and U14736 (N_14736,N_10935,N_9002);
nor U14737 (N_14737,N_11070,N_10668);
xnor U14738 (N_14738,N_8106,N_8014);
nand U14739 (N_14739,N_11183,N_10741);
or U14740 (N_14740,N_9249,N_10688);
nand U14741 (N_14741,N_8215,N_9137);
xor U14742 (N_14742,N_10909,N_10264);
xor U14743 (N_14743,N_10771,N_11314);
or U14744 (N_14744,N_11594,N_10634);
or U14745 (N_14745,N_8577,N_9605);
and U14746 (N_14746,N_9547,N_9571);
and U14747 (N_14747,N_8745,N_8170);
and U14748 (N_14748,N_11157,N_9708);
or U14749 (N_14749,N_8769,N_9445);
or U14750 (N_14750,N_9165,N_10241);
nor U14751 (N_14751,N_8637,N_9257);
nor U14752 (N_14752,N_9825,N_10293);
or U14753 (N_14753,N_8941,N_8858);
xor U14754 (N_14754,N_10952,N_11749);
nand U14755 (N_14755,N_11363,N_9810);
nor U14756 (N_14756,N_9392,N_8306);
and U14757 (N_14757,N_11858,N_11329);
xor U14758 (N_14758,N_8687,N_10898);
nor U14759 (N_14759,N_10694,N_8087);
or U14760 (N_14760,N_8562,N_8492);
and U14761 (N_14761,N_8727,N_11487);
and U14762 (N_14762,N_10757,N_10849);
nor U14763 (N_14763,N_8666,N_9469);
or U14764 (N_14764,N_10201,N_9703);
nor U14765 (N_14765,N_8882,N_8732);
nand U14766 (N_14766,N_9503,N_9658);
and U14767 (N_14767,N_9132,N_8803);
or U14768 (N_14768,N_9112,N_11419);
or U14769 (N_14769,N_9954,N_10917);
nor U14770 (N_14770,N_9416,N_9147);
nand U14771 (N_14771,N_10584,N_9033);
nor U14772 (N_14772,N_9157,N_11261);
xnor U14773 (N_14773,N_11505,N_9930);
nor U14774 (N_14774,N_8916,N_8180);
and U14775 (N_14775,N_9762,N_11446);
or U14776 (N_14776,N_11785,N_8909);
nor U14777 (N_14777,N_9248,N_11845);
or U14778 (N_14778,N_11243,N_8888);
or U14779 (N_14779,N_8663,N_11822);
nand U14780 (N_14780,N_10066,N_10930);
and U14781 (N_14781,N_11990,N_9041);
nor U14782 (N_14782,N_9284,N_8926);
xnor U14783 (N_14783,N_9971,N_8941);
xnor U14784 (N_14784,N_11275,N_10567);
xnor U14785 (N_14785,N_8257,N_10431);
nand U14786 (N_14786,N_8770,N_11053);
nor U14787 (N_14787,N_11503,N_8720);
nand U14788 (N_14788,N_9476,N_10165);
xnor U14789 (N_14789,N_8456,N_9284);
nor U14790 (N_14790,N_8482,N_11604);
xnor U14791 (N_14791,N_9583,N_10251);
nand U14792 (N_14792,N_11587,N_9764);
and U14793 (N_14793,N_11738,N_8709);
nor U14794 (N_14794,N_8498,N_10851);
xor U14795 (N_14795,N_8625,N_9444);
xnor U14796 (N_14796,N_10264,N_8619);
xor U14797 (N_14797,N_11350,N_11842);
nand U14798 (N_14798,N_11877,N_9004);
nand U14799 (N_14799,N_10500,N_10338);
nand U14800 (N_14800,N_9708,N_10788);
xnor U14801 (N_14801,N_9790,N_9387);
and U14802 (N_14802,N_9708,N_11464);
or U14803 (N_14803,N_11466,N_8096);
and U14804 (N_14804,N_9147,N_8397);
xor U14805 (N_14805,N_8157,N_8750);
or U14806 (N_14806,N_10680,N_9648);
and U14807 (N_14807,N_11247,N_11957);
xor U14808 (N_14808,N_8613,N_8476);
or U14809 (N_14809,N_9487,N_9504);
or U14810 (N_14810,N_11320,N_8930);
and U14811 (N_14811,N_11124,N_8846);
or U14812 (N_14812,N_9951,N_9618);
nand U14813 (N_14813,N_9932,N_10555);
xor U14814 (N_14814,N_10068,N_9242);
nand U14815 (N_14815,N_11469,N_8783);
xnor U14816 (N_14816,N_10374,N_8907);
and U14817 (N_14817,N_9989,N_9914);
and U14818 (N_14818,N_10557,N_8892);
nand U14819 (N_14819,N_10087,N_8693);
or U14820 (N_14820,N_9866,N_8879);
or U14821 (N_14821,N_9328,N_10160);
or U14822 (N_14822,N_8779,N_9298);
and U14823 (N_14823,N_9704,N_8910);
xor U14824 (N_14824,N_8371,N_8064);
nand U14825 (N_14825,N_11430,N_9788);
nand U14826 (N_14826,N_11293,N_8541);
xnor U14827 (N_14827,N_8784,N_10021);
nand U14828 (N_14828,N_11246,N_10620);
xor U14829 (N_14829,N_9795,N_10328);
xor U14830 (N_14830,N_11170,N_8277);
xnor U14831 (N_14831,N_9772,N_8545);
and U14832 (N_14832,N_11541,N_11745);
and U14833 (N_14833,N_10804,N_9124);
nand U14834 (N_14834,N_8073,N_11645);
nand U14835 (N_14835,N_9937,N_10658);
and U14836 (N_14836,N_8180,N_11138);
nand U14837 (N_14837,N_9045,N_9389);
nor U14838 (N_14838,N_11197,N_10800);
and U14839 (N_14839,N_8337,N_11740);
and U14840 (N_14840,N_11295,N_11851);
or U14841 (N_14841,N_11543,N_10230);
or U14842 (N_14842,N_10766,N_10422);
nand U14843 (N_14843,N_9530,N_9308);
and U14844 (N_14844,N_11038,N_11492);
nor U14845 (N_14845,N_8869,N_9669);
nor U14846 (N_14846,N_8733,N_8038);
or U14847 (N_14847,N_11673,N_11145);
nor U14848 (N_14848,N_10692,N_10346);
or U14849 (N_14849,N_11623,N_8540);
and U14850 (N_14850,N_9588,N_9944);
and U14851 (N_14851,N_9526,N_8922);
xor U14852 (N_14852,N_8627,N_10155);
or U14853 (N_14853,N_10117,N_8255);
or U14854 (N_14854,N_10321,N_11375);
xor U14855 (N_14855,N_11719,N_8252);
nor U14856 (N_14856,N_11212,N_10751);
and U14857 (N_14857,N_8035,N_10520);
and U14858 (N_14858,N_11135,N_9109);
xnor U14859 (N_14859,N_10806,N_10957);
nand U14860 (N_14860,N_8511,N_10033);
nor U14861 (N_14861,N_10657,N_8938);
xor U14862 (N_14862,N_11690,N_10961);
nor U14863 (N_14863,N_8856,N_10127);
nand U14864 (N_14864,N_8434,N_10284);
or U14865 (N_14865,N_9342,N_10916);
xor U14866 (N_14866,N_10793,N_11424);
nand U14867 (N_14867,N_11892,N_11755);
nand U14868 (N_14868,N_9198,N_11969);
nor U14869 (N_14869,N_8058,N_11883);
xnor U14870 (N_14870,N_10848,N_9032);
xor U14871 (N_14871,N_9403,N_8896);
nor U14872 (N_14872,N_11469,N_9339);
or U14873 (N_14873,N_8261,N_9095);
or U14874 (N_14874,N_10432,N_8864);
nor U14875 (N_14875,N_11186,N_9687);
or U14876 (N_14876,N_10960,N_8097);
or U14877 (N_14877,N_8713,N_9916);
or U14878 (N_14878,N_8605,N_10654);
xor U14879 (N_14879,N_10250,N_10267);
xor U14880 (N_14880,N_11206,N_10334);
nor U14881 (N_14881,N_9535,N_10406);
nand U14882 (N_14882,N_8658,N_11127);
nor U14883 (N_14883,N_10387,N_8978);
and U14884 (N_14884,N_10412,N_9047);
nor U14885 (N_14885,N_8498,N_9320);
nor U14886 (N_14886,N_8164,N_9969);
or U14887 (N_14887,N_9793,N_11328);
xor U14888 (N_14888,N_10959,N_9021);
xnor U14889 (N_14889,N_11792,N_10089);
nand U14890 (N_14890,N_10225,N_8458);
xor U14891 (N_14891,N_10605,N_10900);
nand U14892 (N_14892,N_9943,N_10756);
or U14893 (N_14893,N_11135,N_8767);
nor U14894 (N_14894,N_8607,N_8446);
and U14895 (N_14895,N_11424,N_8809);
nand U14896 (N_14896,N_11936,N_10446);
nand U14897 (N_14897,N_10454,N_9186);
and U14898 (N_14898,N_10062,N_11167);
or U14899 (N_14899,N_11545,N_11320);
nor U14900 (N_14900,N_10432,N_11663);
nand U14901 (N_14901,N_8196,N_9792);
nand U14902 (N_14902,N_8701,N_8608);
nand U14903 (N_14903,N_11899,N_8811);
nand U14904 (N_14904,N_8175,N_9098);
nand U14905 (N_14905,N_9647,N_9675);
xor U14906 (N_14906,N_9558,N_10988);
xor U14907 (N_14907,N_10888,N_8186);
nand U14908 (N_14908,N_11458,N_11674);
and U14909 (N_14909,N_11280,N_10937);
nor U14910 (N_14910,N_11315,N_8318);
or U14911 (N_14911,N_11933,N_9767);
xnor U14912 (N_14912,N_8053,N_11336);
or U14913 (N_14913,N_11156,N_8767);
nand U14914 (N_14914,N_8499,N_9040);
and U14915 (N_14915,N_9751,N_10421);
nor U14916 (N_14916,N_9891,N_10741);
or U14917 (N_14917,N_8482,N_11941);
nand U14918 (N_14918,N_9426,N_8732);
xnor U14919 (N_14919,N_11890,N_8510);
and U14920 (N_14920,N_11010,N_11783);
nand U14921 (N_14921,N_10685,N_9447);
or U14922 (N_14922,N_10847,N_11726);
or U14923 (N_14923,N_11650,N_8609);
nor U14924 (N_14924,N_8515,N_9904);
xnor U14925 (N_14925,N_8059,N_8509);
nor U14926 (N_14926,N_10679,N_10568);
xnor U14927 (N_14927,N_11558,N_11678);
xor U14928 (N_14928,N_9887,N_10947);
and U14929 (N_14929,N_11701,N_8559);
nor U14930 (N_14930,N_8044,N_10683);
and U14931 (N_14931,N_11402,N_11485);
nand U14932 (N_14932,N_10974,N_11480);
or U14933 (N_14933,N_9987,N_10494);
or U14934 (N_14934,N_10379,N_9141);
nor U14935 (N_14935,N_10583,N_11114);
nor U14936 (N_14936,N_9346,N_11186);
nand U14937 (N_14937,N_10169,N_8123);
xnor U14938 (N_14938,N_8559,N_11123);
or U14939 (N_14939,N_10123,N_9227);
or U14940 (N_14940,N_11035,N_8177);
and U14941 (N_14941,N_11204,N_8631);
nor U14942 (N_14942,N_8011,N_9837);
or U14943 (N_14943,N_9087,N_11173);
nor U14944 (N_14944,N_8399,N_8027);
nand U14945 (N_14945,N_11642,N_9978);
nand U14946 (N_14946,N_9740,N_9570);
or U14947 (N_14947,N_9421,N_8457);
nand U14948 (N_14948,N_8692,N_8254);
nor U14949 (N_14949,N_11151,N_10986);
xor U14950 (N_14950,N_10000,N_11297);
and U14951 (N_14951,N_9059,N_8520);
or U14952 (N_14952,N_8146,N_9915);
nor U14953 (N_14953,N_10162,N_8952);
nand U14954 (N_14954,N_11347,N_9732);
xnor U14955 (N_14955,N_8495,N_10420);
xnor U14956 (N_14956,N_8380,N_9979);
xor U14957 (N_14957,N_11673,N_9874);
xor U14958 (N_14958,N_11031,N_9085);
and U14959 (N_14959,N_8020,N_9848);
nand U14960 (N_14960,N_9432,N_9166);
or U14961 (N_14961,N_11002,N_8501);
xnor U14962 (N_14962,N_11162,N_11497);
or U14963 (N_14963,N_9909,N_8052);
or U14964 (N_14964,N_9794,N_11315);
xnor U14965 (N_14965,N_11615,N_10707);
or U14966 (N_14966,N_10761,N_10811);
nand U14967 (N_14967,N_10364,N_8386);
and U14968 (N_14968,N_10122,N_11144);
or U14969 (N_14969,N_11296,N_8070);
nand U14970 (N_14970,N_9701,N_8801);
and U14971 (N_14971,N_10025,N_9486);
xor U14972 (N_14972,N_9787,N_11422);
nand U14973 (N_14973,N_11267,N_10704);
nor U14974 (N_14974,N_10966,N_11987);
or U14975 (N_14975,N_8000,N_8148);
xnor U14976 (N_14976,N_10820,N_9349);
or U14977 (N_14977,N_8743,N_10967);
and U14978 (N_14978,N_11288,N_9958);
and U14979 (N_14979,N_9796,N_9576);
nor U14980 (N_14980,N_11083,N_11044);
or U14981 (N_14981,N_10129,N_9746);
or U14982 (N_14982,N_11140,N_11633);
or U14983 (N_14983,N_9752,N_8065);
nand U14984 (N_14984,N_11841,N_9327);
and U14985 (N_14985,N_9762,N_11786);
and U14986 (N_14986,N_9380,N_10211);
nand U14987 (N_14987,N_8957,N_8668);
and U14988 (N_14988,N_10786,N_9066);
xnor U14989 (N_14989,N_8182,N_10882);
nand U14990 (N_14990,N_8750,N_10918);
nand U14991 (N_14991,N_10271,N_9928);
nand U14992 (N_14992,N_10044,N_9301);
and U14993 (N_14993,N_8179,N_11932);
nand U14994 (N_14994,N_10791,N_8888);
or U14995 (N_14995,N_9429,N_8444);
nor U14996 (N_14996,N_8823,N_8205);
nor U14997 (N_14997,N_11093,N_10333);
and U14998 (N_14998,N_11355,N_9984);
xor U14999 (N_14999,N_9586,N_11942);
or U15000 (N_15000,N_11866,N_10793);
or U15001 (N_15001,N_8270,N_11146);
nor U15002 (N_15002,N_8794,N_8186);
or U15003 (N_15003,N_10921,N_9660);
and U15004 (N_15004,N_11488,N_10214);
or U15005 (N_15005,N_11879,N_11615);
or U15006 (N_15006,N_8922,N_10080);
xnor U15007 (N_15007,N_8921,N_8917);
or U15008 (N_15008,N_9528,N_11264);
or U15009 (N_15009,N_10707,N_9009);
and U15010 (N_15010,N_11118,N_8700);
xnor U15011 (N_15011,N_11307,N_11185);
or U15012 (N_15012,N_11611,N_9462);
nand U15013 (N_15013,N_10314,N_10958);
nand U15014 (N_15014,N_10795,N_11667);
nand U15015 (N_15015,N_10066,N_10226);
nor U15016 (N_15016,N_9776,N_10005);
or U15017 (N_15017,N_11542,N_11903);
and U15018 (N_15018,N_10689,N_11307);
nor U15019 (N_15019,N_9489,N_10488);
and U15020 (N_15020,N_9904,N_11621);
nand U15021 (N_15021,N_9758,N_11794);
nand U15022 (N_15022,N_11205,N_8059);
nand U15023 (N_15023,N_8550,N_11262);
xor U15024 (N_15024,N_8869,N_9191);
nor U15025 (N_15025,N_9404,N_9368);
and U15026 (N_15026,N_8552,N_8892);
and U15027 (N_15027,N_10175,N_10267);
and U15028 (N_15028,N_8835,N_9174);
nor U15029 (N_15029,N_11195,N_8083);
and U15030 (N_15030,N_8155,N_11676);
nand U15031 (N_15031,N_10623,N_10090);
nand U15032 (N_15032,N_10879,N_10459);
and U15033 (N_15033,N_9855,N_10142);
nand U15034 (N_15034,N_11663,N_9835);
xnor U15035 (N_15035,N_8752,N_9547);
nor U15036 (N_15036,N_9216,N_8766);
xor U15037 (N_15037,N_9458,N_8481);
and U15038 (N_15038,N_11322,N_8850);
nor U15039 (N_15039,N_9790,N_8831);
and U15040 (N_15040,N_9405,N_9864);
xor U15041 (N_15041,N_11947,N_9235);
or U15042 (N_15042,N_10570,N_11218);
xor U15043 (N_15043,N_11796,N_9619);
and U15044 (N_15044,N_11140,N_11080);
nor U15045 (N_15045,N_9033,N_10604);
nor U15046 (N_15046,N_9954,N_11464);
or U15047 (N_15047,N_10014,N_8169);
xnor U15048 (N_15048,N_11987,N_11475);
xor U15049 (N_15049,N_8606,N_8835);
or U15050 (N_15050,N_11799,N_9169);
and U15051 (N_15051,N_11699,N_8024);
nand U15052 (N_15052,N_8422,N_10838);
or U15053 (N_15053,N_11343,N_9454);
xnor U15054 (N_15054,N_9360,N_8538);
and U15055 (N_15055,N_11985,N_9380);
xnor U15056 (N_15056,N_11229,N_11508);
and U15057 (N_15057,N_8885,N_9673);
nor U15058 (N_15058,N_9327,N_8321);
and U15059 (N_15059,N_8170,N_9851);
and U15060 (N_15060,N_10767,N_9038);
nand U15061 (N_15061,N_11472,N_9306);
or U15062 (N_15062,N_8752,N_8380);
nor U15063 (N_15063,N_11992,N_8515);
and U15064 (N_15064,N_9013,N_10509);
nand U15065 (N_15065,N_9135,N_11740);
and U15066 (N_15066,N_11565,N_9575);
xor U15067 (N_15067,N_8591,N_10443);
nand U15068 (N_15068,N_8136,N_10284);
or U15069 (N_15069,N_9729,N_9668);
or U15070 (N_15070,N_10944,N_11916);
xnor U15071 (N_15071,N_11875,N_9367);
nor U15072 (N_15072,N_8131,N_9933);
nand U15073 (N_15073,N_9114,N_8811);
nor U15074 (N_15074,N_10656,N_8248);
and U15075 (N_15075,N_8229,N_8607);
nor U15076 (N_15076,N_8553,N_11577);
nor U15077 (N_15077,N_9015,N_8216);
and U15078 (N_15078,N_11284,N_9504);
and U15079 (N_15079,N_8649,N_11862);
nor U15080 (N_15080,N_8684,N_11110);
nand U15081 (N_15081,N_10549,N_11835);
or U15082 (N_15082,N_9822,N_9672);
nand U15083 (N_15083,N_8092,N_8771);
nand U15084 (N_15084,N_8494,N_10594);
xor U15085 (N_15085,N_11741,N_9191);
and U15086 (N_15086,N_10804,N_8344);
or U15087 (N_15087,N_8302,N_11733);
xor U15088 (N_15088,N_8071,N_10428);
xnor U15089 (N_15089,N_8919,N_10033);
or U15090 (N_15090,N_10828,N_11672);
xnor U15091 (N_15091,N_8499,N_10078);
nor U15092 (N_15092,N_11116,N_9580);
or U15093 (N_15093,N_8869,N_10174);
and U15094 (N_15094,N_10269,N_10401);
nor U15095 (N_15095,N_9231,N_8301);
nor U15096 (N_15096,N_11533,N_10824);
nor U15097 (N_15097,N_10128,N_11696);
xnor U15098 (N_15098,N_11756,N_8672);
nor U15099 (N_15099,N_9262,N_8494);
nor U15100 (N_15100,N_11701,N_11855);
xnor U15101 (N_15101,N_10449,N_10618);
and U15102 (N_15102,N_9737,N_8654);
or U15103 (N_15103,N_11178,N_11360);
nand U15104 (N_15104,N_10162,N_8688);
xnor U15105 (N_15105,N_8967,N_10197);
and U15106 (N_15106,N_8172,N_9075);
xor U15107 (N_15107,N_9174,N_9554);
or U15108 (N_15108,N_9459,N_8667);
nand U15109 (N_15109,N_11312,N_11594);
or U15110 (N_15110,N_8701,N_9947);
nand U15111 (N_15111,N_9301,N_11044);
xor U15112 (N_15112,N_8265,N_10839);
and U15113 (N_15113,N_9811,N_11939);
or U15114 (N_15114,N_10010,N_9608);
nor U15115 (N_15115,N_10724,N_9143);
nor U15116 (N_15116,N_8707,N_10960);
or U15117 (N_15117,N_10623,N_9179);
nor U15118 (N_15118,N_10849,N_8022);
or U15119 (N_15119,N_9227,N_8565);
nand U15120 (N_15120,N_10182,N_10275);
nor U15121 (N_15121,N_8972,N_11141);
nor U15122 (N_15122,N_11075,N_10032);
nand U15123 (N_15123,N_9072,N_10429);
xnor U15124 (N_15124,N_11897,N_10202);
nand U15125 (N_15125,N_8920,N_11802);
and U15126 (N_15126,N_8051,N_10568);
nor U15127 (N_15127,N_8044,N_8623);
nand U15128 (N_15128,N_8552,N_9584);
or U15129 (N_15129,N_8257,N_11533);
nand U15130 (N_15130,N_8227,N_10434);
and U15131 (N_15131,N_9708,N_11828);
nand U15132 (N_15132,N_10964,N_11878);
nor U15133 (N_15133,N_11073,N_10549);
or U15134 (N_15134,N_10058,N_10896);
and U15135 (N_15135,N_10844,N_11385);
nand U15136 (N_15136,N_10878,N_11579);
nor U15137 (N_15137,N_11203,N_10032);
nor U15138 (N_15138,N_10422,N_10430);
nand U15139 (N_15139,N_10470,N_11089);
and U15140 (N_15140,N_8523,N_10176);
nor U15141 (N_15141,N_11160,N_10813);
nor U15142 (N_15142,N_8479,N_11434);
and U15143 (N_15143,N_11921,N_9299);
and U15144 (N_15144,N_9196,N_8296);
and U15145 (N_15145,N_9972,N_9290);
nor U15146 (N_15146,N_8964,N_9853);
nand U15147 (N_15147,N_11089,N_9142);
or U15148 (N_15148,N_9275,N_11289);
and U15149 (N_15149,N_8730,N_9610);
nand U15150 (N_15150,N_11218,N_10126);
nand U15151 (N_15151,N_10290,N_9956);
xnor U15152 (N_15152,N_11757,N_10967);
nor U15153 (N_15153,N_10201,N_8879);
nand U15154 (N_15154,N_11511,N_8165);
and U15155 (N_15155,N_9532,N_11296);
xnor U15156 (N_15156,N_9933,N_9897);
or U15157 (N_15157,N_11784,N_9898);
and U15158 (N_15158,N_10574,N_8453);
and U15159 (N_15159,N_9364,N_9641);
and U15160 (N_15160,N_8107,N_11535);
and U15161 (N_15161,N_11075,N_10266);
xor U15162 (N_15162,N_8265,N_8900);
or U15163 (N_15163,N_10638,N_8474);
nor U15164 (N_15164,N_11090,N_9914);
and U15165 (N_15165,N_10330,N_9180);
nor U15166 (N_15166,N_10363,N_10354);
nand U15167 (N_15167,N_11355,N_10991);
xnor U15168 (N_15168,N_8802,N_8862);
nor U15169 (N_15169,N_11443,N_9535);
nor U15170 (N_15170,N_10361,N_10864);
nand U15171 (N_15171,N_11052,N_10772);
nand U15172 (N_15172,N_10354,N_10733);
nand U15173 (N_15173,N_8891,N_8632);
xnor U15174 (N_15174,N_11422,N_10204);
nand U15175 (N_15175,N_9023,N_11529);
nand U15176 (N_15176,N_10378,N_9079);
nor U15177 (N_15177,N_9992,N_10955);
nor U15178 (N_15178,N_11307,N_10748);
nor U15179 (N_15179,N_8085,N_10548);
xnor U15180 (N_15180,N_8958,N_10243);
and U15181 (N_15181,N_11493,N_10694);
or U15182 (N_15182,N_8626,N_8177);
nand U15183 (N_15183,N_8632,N_8628);
xor U15184 (N_15184,N_11202,N_9540);
nor U15185 (N_15185,N_10468,N_10502);
nor U15186 (N_15186,N_8281,N_10863);
xor U15187 (N_15187,N_8049,N_11352);
and U15188 (N_15188,N_9521,N_9814);
or U15189 (N_15189,N_11683,N_11165);
nor U15190 (N_15190,N_8212,N_8839);
and U15191 (N_15191,N_8406,N_9812);
nor U15192 (N_15192,N_10037,N_8692);
nand U15193 (N_15193,N_10519,N_8401);
and U15194 (N_15194,N_11894,N_11478);
nand U15195 (N_15195,N_8206,N_9103);
and U15196 (N_15196,N_11332,N_10684);
nor U15197 (N_15197,N_11377,N_10173);
nor U15198 (N_15198,N_10085,N_10634);
xor U15199 (N_15199,N_10819,N_10346);
nand U15200 (N_15200,N_9218,N_10265);
and U15201 (N_15201,N_10181,N_11190);
or U15202 (N_15202,N_9956,N_11517);
or U15203 (N_15203,N_11812,N_11755);
xnor U15204 (N_15204,N_9539,N_9964);
nand U15205 (N_15205,N_11857,N_9869);
and U15206 (N_15206,N_11673,N_9219);
nor U15207 (N_15207,N_8004,N_10061);
and U15208 (N_15208,N_8247,N_10784);
xnor U15209 (N_15209,N_10409,N_11234);
or U15210 (N_15210,N_9756,N_11093);
nand U15211 (N_15211,N_11909,N_10795);
nand U15212 (N_15212,N_10744,N_10520);
and U15213 (N_15213,N_10110,N_11980);
and U15214 (N_15214,N_8237,N_11159);
xor U15215 (N_15215,N_10282,N_11568);
nand U15216 (N_15216,N_8423,N_11729);
or U15217 (N_15217,N_11999,N_9638);
or U15218 (N_15218,N_9085,N_8554);
and U15219 (N_15219,N_8221,N_11148);
xor U15220 (N_15220,N_9080,N_8366);
xor U15221 (N_15221,N_9366,N_9969);
xnor U15222 (N_15222,N_10305,N_8274);
nor U15223 (N_15223,N_11223,N_10744);
nor U15224 (N_15224,N_9719,N_11023);
nand U15225 (N_15225,N_11196,N_11425);
and U15226 (N_15226,N_9588,N_11129);
or U15227 (N_15227,N_11264,N_11221);
or U15228 (N_15228,N_8712,N_10100);
or U15229 (N_15229,N_8989,N_8894);
or U15230 (N_15230,N_8492,N_10982);
and U15231 (N_15231,N_9851,N_9953);
nand U15232 (N_15232,N_11293,N_10101);
nand U15233 (N_15233,N_8168,N_10511);
or U15234 (N_15234,N_10625,N_10359);
and U15235 (N_15235,N_11500,N_8088);
nand U15236 (N_15236,N_8239,N_8260);
nor U15237 (N_15237,N_11755,N_9543);
nor U15238 (N_15238,N_10164,N_9356);
nand U15239 (N_15239,N_9252,N_9414);
nor U15240 (N_15240,N_8440,N_11999);
xor U15241 (N_15241,N_10866,N_9118);
and U15242 (N_15242,N_8108,N_10238);
nand U15243 (N_15243,N_10163,N_11010);
nand U15244 (N_15244,N_8061,N_11664);
nor U15245 (N_15245,N_8525,N_8243);
or U15246 (N_15246,N_8719,N_11885);
or U15247 (N_15247,N_10594,N_11645);
nor U15248 (N_15248,N_8494,N_8291);
or U15249 (N_15249,N_8038,N_8715);
or U15250 (N_15250,N_8496,N_9232);
nand U15251 (N_15251,N_9152,N_10317);
xnor U15252 (N_15252,N_8003,N_9503);
nand U15253 (N_15253,N_11002,N_9026);
nand U15254 (N_15254,N_10024,N_9525);
nand U15255 (N_15255,N_11150,N_8091);
nor U15256 (N_15256,N_11241,N_10778);
and U15257 (N_15257,N_8274,N_9581);
nand U15258 (N_15258,N_9960,N_9990);
or U15259 (N_15259,N_11019,N_8269);
xnor U15260 (N_15260,N_10625,N_9212);
xor U15261 (N_15261,N_11705,N_8798);
or U15262 (N_15262,N_11035,N_10973);
and U15263 (N_15263,N_9642,N_8504);
nor U15264 (N_15264,N_10372,N_9156);
xnor U15265 (N_15265,N_10916,N_9662);
nor U15266 (N_15266,N_11230,N_11027);
xor U15267 (N_15267,N_10837,N_10300);
xor U15268 (N_15268,N_11484,N_8232);
nand U15269 (N_15269,N_8186,N_10838);
nand U15270 (N_15270,N_11496,N_11713);
nand U15271 (N_15271,N_10227,N_8136);
nand U15272 (N_15272,N_11755,N_11692);
and U15273 (N_15273,N_10433,N_10350);
or U15274 (N_15274,N_11502,N_10157);
nor U15275 (N_15275,N_8243,N_10304);
and U15276 (N_15276,N_8918,N_10226);
nand U15277 (N_15277,N_10270,N_11763);
nand U15278 (N_15278,N_9250,N_10679);
nand U15279 (N_15279,N_10073,N_10746);
or U15280 (N_15280,N_11634,N_11803);
nand U15281 (N_15281,N_8220,N_10900);
xor U15282 (N_15282,N_8240,N_11720);
xnor U15283 (N_15283,N_11977,N_8439);
nor U15284 (N_15284,N_9840,N_8284);
and U15285 (N_15285,N_10193,N_11684);
and U15286 (N_15286,N_10854,N_8228);
and U15287 (N_15287,N_8032,N_9633);
or U15288 (N_15288,N_8444,N_10796);
or U15289 (N_15289,N_10447,N_8080);
and U15290 (N_15290,N_10035,N_9463);
or U15291 (N_15291,N_8173,N_8037);
and U15292 (N_15292,N_9511,N_11264);
or U15293 (N_15293,N_11750,N_11851);
or U15294 (N_15294,N_11436,N_10932);
or U15295 (N_15295,N_10076,N_10758);
nor U15296 (N_15296,N_8434,N_9624);
nor U15297 (N_15297,N_10809,N_11148);
or U15298 (N_15298,N_10612,N_8300);
nand U15299 (N_15299,N_10166,N_8379);
xor U15300 (N_15300,N_8945,N_9456);
xnor U15301 (N_15301,N_11537,N_11201);
or U15302 (N_15302,N_11371,N_10649);
xor U15303 (N_15303,N_8483,N_11300);
xnor U15304 (N_15304,N_9131,N_10491);
nor U15305 (N_15305,N_11607,N_11647);
and U15306 (N_15306,N_8623,N_8148);
nor U15307 (N_15307,N_9802,N_11063);
and U15308 (N_15308,N_11389,N_9276);
nor U15309 (N_15309,N_8128,N_11543);
xor U15310 (N_15310,N_8313,N_8202);
xnor U15311 (N_15311,N_10500,N_10348);
and U15312 (N_15312,N_8006,N_10690);
xnor U15313 (N_15313,N_8388,N_9520);
or U15314 (N_15314,N_8136,N_9153);
nand U15315 (N_15315,N_9365,N_8954);
nand U15316 (N_15316,N_10619,N_9245);
nor U15317 (N_15317,N_10958,N_10329);
nor U15318 (N_15318,N_9397,N_10233);
nor U15319 (N_15319,N_11730,N_10568);
and U15320 (N_15320,N_10099,N_8700);
nand U15321 (N_15321,N_10601,N_8361);
xor U15322 (N_15322,N_8419,N_8216);
or U15323 (N_15323,N_9756,N_11835);
or U15324 (N_15324,N_10674,N_11956);
nand U15325 (N_15325,N_8355,N_11453);
nand U15326 (N_15326,N_9260,N_8501);
and U15327 (N_15327,N_11448,N_11234);
nand U15328 (N_15328,N_9817,N_8038);
and U15329 (N_15329,N_8630,N_10272);
or U15330 (N_15330,N_10209,N_11741);
nand U15331 (N_15331,N_11740,N_10673);
nor U15332 (N_15332,N_8684,N_8340);
nand U15333 (N_15333,N_11610,N_9977);
and U15334 (N_15334,N_9924,N_8770);
nor U15335 (N_15335,N_10182,N_8618);
nand U15336 (N_15336,N_11098,N_9913);
or U15337 (N_15337,N_11746,N_8816);
nor U15338 (N_15338,N_10382,N_9766);
nand U15339 (N_15339,N_8084,N_9647);
nand U15340 (N_15340,N_10399,N_10748);
and U15341 (N_15341,N_10780,N_11961);
xnor U15342 (N_15342,N_9477,N_10681);
xnor U15343 (N_15343,N_10408,N_8679);
or U15344 (N_15344,N_8345,N_11752);
nor U15345 (N_15345,N_8540,N_8969);
or U15346 (N_15346,N_9593,N_8977);
nand U15347 (N_15347,N_9851,N_10926);
and U15348 (N_15348,N_9084,N_11354);
and U15349 (N_15349,N_11468,N_8258);
nand U15350 (N_15350,N_10223,N_8239);
xor U15351 (N_15351,N_11282,N_11693);
xor U15352 (N_15352,N_10949,N_10292);
or U15353 (N_15353,N_9575,N_9179);
nor U15354 (N_15354,N_9477,N_11621);
and U15355 (N_15355,N_9039,N_10976);
nor U15356 (N_15356,N_9564,N_8626);
and U15357 (N_15357,N_10922,N_10590);
or U15358 (N_15358,N_9172,N_11180);
nor U15359 (N_15359,N_8306,N_9776);
and U15360 (N_15360,N_11950,N_9934);
or U15361 (N_15361,N_10443,N_8395);
nand U15362 (N_15362,N_11401,N_11586);
or U15363 (N_15363,N_9932,N_10269);
or U15364 (N_15364,N_8269,N_10121);
or U15365 (N_15365,N_8849,N_9864);
nand U15366 (N_15366,N_10997,N_10914);
or U15367 (N_15367,N_11536,N_8173);
nor U15368 (N_15368,N_9085,N_10853);
xor U15369 (N_15369,N_10716,N_8434);
or U15370 (N_15370,N_8772,N_9521);
nor U15371 (N_15371,N_9165,N_11095);
nand U15372 (N_15372,N_9330,N_9400);
xor U15373 (N_15373,N_11588,N_8340);
and U15374 (N_15374,N_11058,N_11033);
or U15375 (N_15375,N_11694,N_11291);
nand U15376 (N_15376,N_11837,N_11135);
nor U15377 (N_15377,N_9979,N_8472);
or U15378 (N_15378,N_11429,N_10089);
or U15379 (N_15379,N_10160,N_8268);
nand U15380 (N_15380,N_11953,N_8818);
xor U15381 (N_15381,N_11785,N_9950);
nand U15382 (N_15382,N_11397,N_10440);
xor U15383 (N_15383,N_11206,N_11092);
xor U15384 (N_15384,N_11738,N_8206);
nor U15385 (N_15385,N_9624,N_11485);
or U15386 (N_15386,N_9370,N_9980);
xor U15387 (N_15387,N_8587,N_11003);
nor U15388 (N_15388,N_10171,N_8559);
and U15389 (N_15389,N_10063,N_8270);
nand U15390 (N_15390,N_11710,N_11841);
nor U15391 (N_15391,N_8693,N_9135);
nor U15392 (N_15392,N_11799,N_11685);
or U15393 (N_15393,N_10744,N_9417);
xor U15394 (N_15394,N_8293,N_10952);
or U15395 (N_15395,N_11252,N_9490);
nand U15396 (N_15396,N_9573,N_11831);
nor U15397 (N_15397,N_8668,N_9203);
xnor U15398 (N_15398,N_10125,N_8198);
and U15399 (N_15399,N_10529,N_11831);
xor U15400 (N_15400,N_8730,N_10637);
nor U15401 (N_15401,N_10814,N_8058);
nand U15402 (N_15402,N_9346,N_9855);
or U15403 (N_15403,N_9208,N_11956);
nor U15404 (N_15404,N_9153,N_10822);
or U15405 (N_15405,N_9074,N_9486);
and U15406 (N_15406,N_11174,N_11667);
or U15407 (N_15407,N_9491,N_11256);
nor U15408 (N_15408,N_8245,N_11890);
or U15409 (N_15409,N_11459,N_9194);
or U15410 (N_15410,N_10932,N_8624);
and U15411 (N_15411,N_10969,N_8190);
or U15412 (N_15412,N_8766,N_11527);
or U15413 (N_15413,N_11025,N_9073);
nor U15414 (N_15414,N_10826,N_11677);
or U15415 (N_15415,N_9319,N_9745);
and U15416 (N_15416,N_8201,N_10591);
xor U15417 (N_15417,N_8303,N_8891);
or U15418 (N_15418,N_9078,N_8943);
nor U15419 (N_15419,N_8273,N_10358);
xor U15420 (N_15420,N_10023,N_9774);
xor U15421 (N_15421,N_10591,N_10259);
nand U15422 (N_15422,N_10890,N_10888);
xor U15423 (N_15423,N_9405,N_9707);
nand U15424 (N_15424,N_10798,N_10940);
nand U15425 (N_15425,N_9654,N_9661);
xor U15426 (N_15426,N_10574,N_8149);
nor U15427 (N_15427,N_8963,N_10207);
nand U15428 (N_15428,N_11118,N_9283);
nand U15429 (N_15429,N_9802,N_11747);
xor U15430 (N_15430,N_11521,N_11551);
or U15431 (N_15431,N_9008,N_9010);
or U15432 (N_15432,N_8065,N_11762);
and U15433 (N_15433,N_9767,N_8011);
nand U15434 (N_15434,N_10772,N_10412);
or U15435 (N_15435,N_8639,N_10736);
nor U15436 (N_15436,N_11115,N_11672);
xnor U15437 (N_15437,N_10630,N_11589);
nand U15438 (N_15438,N_9738,N_9038);
nand U15439 (N_15439,N_10761,N_10411);
nor U15440 (N_15440,N_8940,N_10198);
nand U15441 (N_15441,N_11113,N_11464);
or U15442 (N_15442,N_10780,N_9713);
or U15443 (N_15443,N_9448,N_9962);
xor U15444 (N_15444,N_11110,N_11271);
nand U15445 (N_15445,N_9637,N_11825);
nor U15446 (N_15446,N_11774,N_10512);
nand U15447 (N_15447,N_11583,N_8885);
or U15448 (N_15448,N_8007,N_11643);
or U15449 (N_15449,N_9715,N_9518);
and U15450 (N_15450,N_10430,N_9794);
or U15451 (N_15451,N_8708,N_8399);
and U15452 (N_15452,N_11346,N_9828);
or U15453 (N_15453,N_9996,N_11988);
and U15454 (N_15454,N_11908,N_8973);
and U15455 (N_15455,N_11020,N_9299);
and U15456 (N_15456,N_8522,N_9968);
nand U15457 (N_15457,N_10130,N_10789);
or U15458 (N_15458,N_10047,N_10843);
or U15459 (N_15459,N_8947,N_11606);
xnor U15460 (N_15460,N_10165,N_10654);
or U15461 (N_15461,N_11553,N_10380);
and U15462 (N_15462,N_9876,N_11283);
nor U15463 (N_15463,N_10734,N_10408);
and U15464 (N_15464,N_10658,N_8666);
or U15465 (N_15465,N_8249,N_11541);
xnor U15466 (N_15466,N_10753,N_10817);
nand U15467 (N_15467,N_9246,N_10215);
nand U15468 (N_15468,N_8898,N_8267);
nand U15469 (N_15469,N_9846,N_11261);
and U15470 (N_15470,N_8867,N_11103);
or U15471 (N_15471,N_9908,N_8837);
nor U15472 (N_15472,N_10717,N_11382);
nor U15473 (N_15473,N_11955,N_8344);
xor U15474 (N_15474,N_8793,N_10309);
nor U15475 (N_15475,N_9233,N_8478);
and U15476 (N_15476,N_8265,N_9396);
or U15477 (N_15477,N_10854,N_9043);
xor U15478 (N_15478,N_10438,N_9447);
and U15479 (N_15479,N_11448,N_11473);
nor U15480 (N_15480,N_10367,N_10735);
xnor U15481 (N_15481,N_9764,N_9774);
or U15482 (N_15482,N_10813,N_8828);
nor U15483 (N_15483,N_9923,N_10928);
nor U15484 (N_15484,N_9237,N_8514);
nor U15485 (N_15485,N_8229,N_8970);
or U15486 (N_15486,N_10625,N_9649);
xor U15487 (N_15487,N_11646,N_10277);
xor U15488 (N_15488,N_11338,N_10398);
nor U15489 (N_15489,N_10127,N_10298);
or U15490 (N_15490,N_9557,N_10660);
nand U15491 (N_15491,N_11040,N_9544);
nor U15492 (N_15492,N_11878,N_10506);
and U15493 (N_15493,N_10858,N_9639);
or U15494 (N_15494,N_9763,N_8365);
nor U15495 (N_15495,N_8181,N_8632);
nand U15496 (N_15496,N_11048,N_9112);
nor U15497 (N_15497,N_8272,N_9789);
nor U15498 (N_15498,N_10998,N_11305);
nand U15499 (N_15499,N_11605,N_11471);
nand U15500 (N_15500,N_10104,N_11993);
nor U15501 (N_15501,N_10038,N_9259);
nand U15502 (N_15502,N_8969,N_8485);
nand U15503 (N_15503,N_10514,N_11752);
or U15504 (N_15504,N_11147,N_9028);
nand U15505 (N_15505,N_8660,N_10877);
and U15506 (N_15506,N_11198,N_11039);
nor U15507 (N_15507,N_9575,N_9539);
nor U15508 (N_15508,N_11840,N_9340);
xnor U15509 (N_15509,N_8667,N_10533);
xnor U15510 (N_15510,N_9295,N_9284);
or U15511 (N_15511,N_10524,N_8803);
nand U15512 (N_15512,N_9581,N_8087);
or U15513 (N_15513,N_10262,N_9642);
nand U15514 (N_15514,N_10452,N_10703);
nor U15515 (N_15515,N_11025,N_8566);
nand U15516 (N_15516,N_11385,N_9447);
xor U15517 (N_15517,N_10794,N_10473);
nand U15518 (N_15518,N_11818,N_9631);
nor U15519 (N_15519,N_9983,N_11737);
nand U15520 (N_15520,N_10305,N_11827);
nor U15521 (N_15521,N_9061,N_11305);
and U15522 (N_15522,N_9670,N_11959);
xnor U15523 (N_15523,N_11289,N_8273);
and U15524 (N_15524,N_10965,N_11280);
nor U15525 (N_15525,N_11417,N_10054);
nor U15526 (N_15526,N_8517,N_8327);
nor U15527 (N_15527,N_11576,N_9240);
and U15528 (N_15528,N_11233,N_10480);
nand U15529 (N_15529,N_8085,N_8704);
and U15530 (N_15530,N_8278,N_9743);
nor U15531 (N_15531,N_8647,N_11094);
nand U15532 (N_15532,N_8119,N_10935);
or U15533 (N_15533,N_9312,N_8161);
nor U15534 (N_15534,N_11138,N_9028);
nor U15535 (N_15535,N_10260,N_10096);
xnor U15536 (N_15536,N_11924,N_8380);
nor U15537 (N_15537,N_11193,N_11190);
xnor U15538 (N_15538,N_10392,N_8979);
nand U15539 (N_15539,N_8565,N_8373);
nor U15540 (N_15540,N_11166,N_10930);
nor U15541 (N_15541,N_10715,N_11513);
nor U15542 (N_15542,N_10387,N_8780);
and U15543 (N_15543,N_9919,N_10043);
and U15544 (N_15544,N_8829,N_11331);
nor U15545 (N_15545,N_8976,N_9824);
xnor U15546 (N_15546,N_10668,N_9470);
and U15547 (N_15547,N_9862,N_8118);
or U15548 (N_15548,N_8861,N_11822);
xor U15549 (N_15549,N_10630,N_11149);
nor U15550 (N_15550,N_9333,N_11152);
nor U15551 (N_15551,N_8504,N_8503);
nor U15552 (N_15552,N_8741,N_10200);
nor U15553 (N_15553,N_10782,N_9600);
or U15554 (N_15554,N_11044,N_10011);
and U15555 (N_15555,N_8527,N_10358);
nand U15556 (N_15556,N_10157,N_9566);
nand U15557 (N_15557,N_8052,N_10681);
nor U15558 (N_15558,N_9484,N_11414);
and U15559 (N_15559,N_8384,N_11952);
nor U15560 (N_15560,N_9784,N_11849);
or U15561 (N_15561,N_9262,N_10703);
nor U15562 (N_15562,N_10503,N_11276);
or U15563 (N_15563,N_10121,N_9962);
xnor U15564 (N_15564,N_10695,N_8037);
or U15565 (N_15565,N_9792,N_11122);
or U15566 (N_15566,N_11098,N_10624);
nand U15567 (N_15567,N_9089,N_10919);
nor U15568 (N_15568,N_10986,N_9824);
and U15569 (N_15569,N_10624,N_11135);
or U15570 (N_15570,N_11273,N_11709);
or U15571 (N_15571,N_11034,N_11171);
xor U15572 (N_15572,N_10160,N_10909);
nor U15573 (N_15573,N_11491,N_9395);
nor U15574 (N_15574,N_9848,N_10884);
xnor U15575 (N_15575,N_11546,N_11555);
nor U15576 (N_15576,N_11228,N_9555);
nor U15577 (N_15577,N_8596,N_10989);
nand U15578 (N_15578,N_9968,N_9203);
or U15579 (N_15579,N_8580,N_8432);
xnor U15580 (N_15580,N_8247,N_8403);
or U15581 (N_15581,N_8210,N_10679);
or U15582 (N_15582,N_8984,N_8614);
or U15583 (N_15583,N_8043,N_11693);
nand U15584 (N_15584,N_9213,N_9018);
and U15585 (N_15585,N_11056,N_8996);
and U15586 (N_15586,N_9155,N_10861);
and U15587 (N_15587,N_11491,N_8773);
nand U15588 (N_15588,N_9874,N_8945);
nand U15589 (N_15589,N_8472,N_10904);
or U15590 (N_15590,N_9122,N_8579);
or U15591 (N_15591,N_10055,N_11272);
nor U15592 (N_15592,N_10563,N_10997);
or U15593 (N_15593,N_8489,N_11586);
and U15594 (N_15594,N_9328,N_9303);
nand U15595 (N_15595,N_11828,N_8605);
xor U15596 (N_15596,N_11700,N_8890);
or U15597 (N_15597,N_9965,N_11088);
or U15598 (N_15598,N_9976,N_9529);
xnor U15599 (N_15599,N_8552,N_10912);
xnor U15600 (N_15600,N_8307,N_11316);
xnor U15601 (N_15601,N_8333,N_8620);
nand U15602 (N_15602,N_9143,N_11023);
or U15603 (N_15603,N_11048,N_11440);
nand U15604 (N_15604,N_10059,N_8700);
or U15605 (N_15605,N_9813,N_8213);
nand U15606 (N_15606,N_8079,N_8923);
or U15607 (N_15607,N_9185,N_9399);
and U15608 (N_15608,N_9634,N_11508);
nand U15609 (N_15609,N_10555,N_8583);
or U15610 (N_15610,N_9336,N_11181);
xnor U15611 (N_15611,N_8335,N_8515);
and U15612 (N_15612,N_11364,N_10702);
xnor U15613 (N_15613,N_10685,N_9335);
xor U15614 (N_15614,N_10050,N_9374);
and U15615 (N_15615,N_11494,N_8998);
nand U15616 (N_15616,N_9735,N_11602);
and U15617 (N_15617,N_9833,N_11506);
nor U15618 (N_15618,N_11010,N_9411);
and U15619 (N_15619,N_11200,N_10756);
or U15620 (N_15620,N_9973,N_8864);
or U15621 (N_15621,N_10747,N_10368);
and U15622 (N_15622,N_11428,N_9010);
and U15623 (N_15623,N_11311,N_11843);
xnor U15624 (N_15624,N_11674,N_9206);
or U15625 (N_15625,N_11869,N_8048);
nor U15626 (N_15626,N_9369,N_11300);
and U15627 (N_15627,N_11845,N_11796);
xnor U15628 (N_15628,N_10486,N_11712);
nor U15629 (N_15629,N_11308,N_9363);
nor U15630 (N_15630,N_11985,N_9068);
nand U15631 (N_15631,N_9457,N_9235);
or U15632 (N_15632,N_9864,N_9213);
nor U15633 (N_15633,N_8588,N_9917);
or U15634 (N_15634,N_8399,N_10284);
or U15635 (N_15635,N_9268,N_11021);
nand U15636 (N_15636,N_11299,N_11228);
xnor U15637 (N_15637,N_11208,N_9564);
or U15638 (N_15638,N_8476,N_9761);
or U15639 (N_15639,N_10235,N_11544);
or U15640 (N_15640,N_11997,N_11325);
or U15641 (N_15641,N_11310,N_10743);
xnor U15642 (N_15642,N_11312,N_9880);
or U15643 (N_15643,N_11169,N_11553);
nor U15644 (N_15644,N_8406,N_11651);
or U15645 (N_15645,N_8996,N_9395);
xor U15646 (N_15646,N_9608,N_10078);
nand U15647 (N_15647,N_11933,N_8310);
nand U15648 (N_15648,N_10083,N_10210);
nor U15649 (N_15649,N_8120,N_8455);
xnor U15650 (N_15650,N_8431,N_9125);
and U15651 (N_15651,N_11779,N_11666);
and U15652 (N_15652,N_8700,N_9257);
nand U15653 (N_15653,N_9916,N_11898);
nand U15654 (N_15654,N_8597,N_8443);
nor U15655 (N_15655,N_11850,N_10974);
xnor U15656 (N_15656,N_10528,N_8761);
or U15657 (N_15657,N_10236,N_8741);
xnor U15658 (N_15658,N_8868,N_8000);
nor U15659 (N_15659,N_11655,N_8375);
xnor U15660 (N_15660,N_10498,N_8166);
and U15661 (N_15661,N_9147,N_8269);
xnor U15662 (N_15662,N_10114,N_9132);
nand U15663 (N_15663,N_8334,N_11006);
nor U15664 (N_15664,N_11483,N_10588);
nor U15665 (N_15665,N_10369,N_8502);
nor U15666 (N_15666,N_8832,N_9472);
xnor U15667 (N_15667,N_10800,N_9185);
xnor U15668 (N_15668,N_11411,N_11590);
or U15669 (N_15669,N_11266,N_10869);
nor U15670 (N_15670,N_9079,N_8489);
nand U15671 (N_15671,N_8457,N_8389);
nand U15672 (N_15672,N_11658,N_11767);
nand U15673 (N_15673,N_8777,N_11906);
nand U15674 (N_15674,N_11944,N_8666);
nor U15675 (N_15675,N_10624,N_11310);
nor U15676 (N_15676,N_9867,N_9154);
and U15677 (N_15677,N_10372,N_8970);
and U15678 (N_15678,N_10962,N_10712);
and U15679 (N_15679,N_10611,N_11828);
or U15680 (N_15680,N_9579,N_11873);
and U15681 (N_15681,N_10970,N_10492);
xnor U15682 (N_15682,N_8765,N_11398);
and U15683 (N_15683,N_10736,N_10855);
nand U15684 (N_15684,N_8139,N_10908);
xnor U15685 (N_15685,N_9580,N_8574);
nand U15686 (N_15686,N_11502,N_11565);
and U15687 (N_15687,N_10093,N_8621);
or U15688 (N_15688,N_9179,N_9454);
and U15689 (N_15689,N_8708,N_9540);
and U15690 (N_15690,N_8319,N_8513);
or U15691 (N_15691,N_8555,N_11424);
nor U15692 (N_15692,N_9010,N_10299);
and U15693 (N_15693,N_8994,N_10712);
and U15694 (N_15694,N_11767,N_11114);
nand U15695 (N_15695,N_10008,N_11099);
or U15696 (N_15696,N_10290,N_10857);
nand U15697 (N_15697,N_9677,N_10233);
xor U15698 (N_15698,N_11646,N_9821);
nand U15699 (N_15699,N_8128,N_9779);
nor U15700 (N_15700,N_11030,N_8774);
or U15701 (N_15701,N_9519,N_11636);
xnor U15702 (N_15702,N_10329,N_8909);
xnor U15703 (N_15703,N_11367,N_10145);
nor U15704 (N_15704,N_9266,N_11995);
and U15705 (N_15705,N_9501,N_10890);
and U15706 (N_15706,N_10603,N_9744);
xnor U15707 (N_15707,N_10214,N_10322);
and U15708 (N_15708,N_11876,N_11657);
or U15709 (N_15709,N_9983,N_11719);
and U15710 (N_15710,N_10210,N_10530);
and U15711 (N_15711,N_11536,N_8566);
nor U15712 (N_15712,N_11633,N_9754);
nor U15713 (N_15713,N_11157,N_8101);
nand U15714 (N_15714,N_10893,N_11440);
nand U15715 (N_15715,N_8934,N_11609);
nand U15716 (N_15716,N_9162,N_11710);
nor U15717 (N_15717,N_11885,N_11986);
and U15718 (N_15718,N_9308,N_10072);
nor U15719 (N_15719,N_8786,N_8457);
nor U15720 (N_15720,N_8763,N_8553);
nand U15721 (N_15721,N_9719,N_10931);
and U15722 (N_15722,N_11964,N_8734);
or U15723 (N_15723,N_10252,N_9096);
and U15724 (N_15724,N_9931,N_11169);
or U15725 (N_15725,N_11186,N_9800);
and U15726 (N_15726,N_11403,N_11351);
nor U15727 (N_15727,N_8095,N_11546);
xnor U15728 (N_15728,N_9987,N_10772);
xor U15729 (N_15729,N_8514,N_8591);
nand U15730 (N_15730,N_9892,N_8008);
xnor U15731 (N_15731,N_10198,N_10691);
and U15732 (N_15732,N_10080,N_9770);
nor U15733 (N_15733,N_9191,N_9579);
nand U15734 (N_15734,N_9016,N_11802);
nand U15735 (N_15735,N_10939,N_10132);
or U15736 (N_15736,N_10774,N_8491);
xor U15737 (N_15737,N_8015,N_8469);
nand U15738 (N_15738,N_11527,N_10093);
nor U15739 (N_15739,N_10690,N_11581);
or U15740 (N_15740,N_11481,N_9810);
nand U15741 (N_15741,N_8458,N_10290);
xnor U15742 (N_15742,N_10107,N_10022);
nand U15743 (N_15743,N_11278,N_9197);
nor U15744 (N_15744,N_11724,N_11073);
and U15745 (N_15745,N_10435,N_10770);
nand U15746 (N_15746,N_8623,N_10524);
xnor U15747 (N_15747,N_8523,N_10926);
and U15748 (N_15748,N_9094,N_8111);
xor U15749 (N_15749,N_11631,N_9601);
or U15750 (N_15750,N_10853,N_11759);
xor U15751 (N_15751,N_9727,N_8638);
nor U15752 (N_15752,N_11934,N_8627);
nor U15753 (N_15753,N_8241,N_11868);
nand U15754 (N_15754,N_8941,N_11178);
nor U15755 (N_15755,N_9826,N_10444);
and U15756 (N_15756,N_8662,N_9984);
nor U15757 (N_15757,N_11523,N_8993);
xnor U15758 (N_15758,N_9398,N_9601);
xnor U15759 (N_15759,N_8072,N_11981);
nand U15760 (N_15760,N_10414,N_9999);
or U15761 (N_15761,N_8765,N_11652);
nand U15762 (N_15762,N_10312,N_9816);
and U15763 (N_15763,N_10928,N_11602);
and U15764 (N_15764,N_9266,N_8796);
nor U15765 (N_15765,N_10382,N_9850);
and U15766 (N_15766,N_8034,N_10014);
or U15767 (N_15767,N_11113,N_11249);
xnor U15768 (N_15768,N_11851,N_10006);
nor U15769 (N_15769,N_11098,N_9239);
nor U15770 (N_15770,N_11839,N_9647);
or U15771 (N_15771,N_8643,N_11075);
xor U15772 (N_15772,N_10206,N_10891);
or U15773 (N_15773,N_11913,N_11642);
nand U15774 (N_15774,N_10187,N_10139);
or U15775 (N_15775,N_11488,N_10432);
and U15776 (N_15776,N_11056,N_9965);
and U15777 (N_15777,N_10032,N_9190);
nand U15778 (N_15778,N_11000,N_11811);
xor U15779 (N_15779,N_9270,N_10828);
nor U15780 (N_15780,N_10827,N_8680);
nor U15781 (N_15781,N_9263,N_8414);
and U15782 (N_15782,N_10791,N_9545);
nor U15783 (N_15783,N_8287,N_11002);
xor U15784 (N_15784,N_11720,N_10919);
and U15785 (N_15785,N_9951,N_10735);
and U15786 (N_15786,N_8600,N_10519);
xor U15787 (N_15787,N_9224,N_10254);
nor U15788 (N_15788,N_9286,N_11550);
and U15789 (N_15789,N_10244,N_11686);
nor U15790 (N_15790,N_9447,N_8772);
nor U15791 (N_15791,N_8922,N_9215);
nor U15792 (N_15792,N_8558,N_10953);
xor U15793 (N_15793,N_8693,N_11305);
xor U15794 (N_15794,N_9898,N_9202);
nor U15795 (N_15795,N_8326,N_8903);
nor U15796 (N_15796,N_10825,N_8690);
and U15797 (N_15797,N_8986,N_11620);
nor U15798 (N_15798,N_10261,N_8602);
and U15799 (N_15799,N_8718,N_9655);
and U15800 (N_15800,N_11581,N_11140);
and U15801 (N_15801,N_9757,N_11241);
or U15802 (N_15802,N_8643,N_10666);
nand U15803 (N_15803,N_8082,N_11477);
and U15804 (N_15804,N_8492,N_10064);
nor U15805 (N_15805,N_11568,N_10934);
nand U15806 (N_15806,N_10981,N_8319);
or U15807 (N_15807,N_11415,N_8819);
or U15808 (N_15808,N_8042,N_11420);
xor U15809 (N_15809,N_10338,N_8344);
nor U15810 (N_15810,N_8289,N_10511);
nand U15811 (N_15811,N_11313,N_9649);
nand U15812 (N_15812,N_9193,N_11964);
or U15813 (N_15813,N_9277,N_9534);
nand U15814 (N_15814,N_8903,N_10108);
nor U15815 (N_15815,N_11250,N_8315);
xnor U15816 (N_15816,N_11771,N_11467);
or U15817 (N_15817,N_8644,N_10920);
and U15818 (N_15818,N_10344,N_11429);
and U15819 (N_15819,N_10875,N_11428);
nor U15820 (N_15820,N_10387,N_9281);
nand U15821 (N_15821,N_8324,N_9690);
nor U15822 (N_15822,N_11386,N_8299);
and U15823 (N_15823,N_10834,N_9666);
xnor U15824 (N_15824,N_9791,N_10360);
and U15825 (N_15825,N_8507,N_9272);
nand U15826 (N_15826,N_10686,N_9239);
xnor U15827 (N_15827,N_9372,N_11479);
nor U15828 (N_15828,N_8133,N_11089);
nand U15829 (N_15829,N_10608,N_8145);
nand U15830 (N_15830,N_10460,N_10634);
nand U15831 (N_15831,N_9091,N_8202);
and U15832 (N_15832,N_10103,N_8490);
nor U15833 (N_15833,N_8757,N_9670);
nand U15834 (N_15834,N_10628,N_10018);
xnor U15835 (N_15835,N_9536,N_11622);
nand U15836 (N_15836,N_10057,N_10265);
nor U15837 (N_15837,N_9070,N_8276);
or U15838 (N_15838,N_10061,N_8680);
or U15839 (N_15839,N_8615,N_10966);
nor U15840 (N_15840,N_9432,N_8325);
and U15841 (N_15841,N_11519,N_11078);
xnor U15842 (N_15842,N_11890,N_10866);
nor U15843 (N_15843,N_11582,N_10416);
and U15844 (N_15844,N_10719,N_11835);
and U15845 (N_15845,N_8188,N_8017);
and U15846 (N_15846,N_8497,N_11259);
nor U15847 (N_15847,N_9912,N_11003);
or U15848 (N_15848,N_9114,N_11752);
nand U15849 (N_15849,N_9593,N_8501);
nor U15850 (N_15850,N_10716,N_9552);
nor U15851 (N_15851,N_8269,N_8081);
nand U15852 (N_15852,N_8316,N_11448);
and U15853 (N_15853,N_10495,N_8413);
nor U15854 (N_15854,N_10328,N_11387);
nor U15855 (N_15855,N_9106,N_10079);
xor U15856 (N_15856,N_11778,N_11737);
and U15857 (N_15857,N_11456,N_8138);
nor U15858 (N_15858,N_10305,N_11226);
nand U15859 (N_15859,N_10964,N_8314);
xor U15860 (N_15860,N_8552,N_8810);
nand U15861 (N_15861,N_11988,N_10230);
or U15862 (N_15862,N_10119,N_11184);
and U15863 (N_15863,N_9672,N_8284);
xnor U15864 (N_15864,N_8544,N_9115);
and U15865 (N_15865,N_9640,N_10694);
and U15866 (N_15866,N_8573,N_9191);
xnor U15867 (N_15867,N_9585,N_8657);
and U15868 (N_15868,N_9874,N_9694);
xor U15869 (N_15869,N_10332,N_9453);
nor U15870 (N_15870,N_11457,N_11841);
xor U15871 (N_15871,N_9420,N_11246);
and U15872 (N_15872,N_11442,N_11700);
nor U15873 (N_15873,N_9831,N_11991);
nand U15874 (N_15874,N_11653,N_11665);
xor U15875 (N_15875,N_9032,N_11160);
nor U15876 (N_15876,N_8924,N_11028);
or U15877 (N_15877,N_8175,N_11533);
nor U15878 (N_15878,N_10009,N_8297);
nand U15879 (N_15879,N_8447,N_10401);
xnor U15880 (N_15880,N_8170,N_10850);
xnor U15881 (N_15881,N_11958,N_9337);
xor U15882 (N_15882,N_10071,N_10257);
nor U15883 (N_15883,N_8332,N_11138);
nand U15884 (N_15884,N_10547,N_8097);
nor U15885 (N_15885,N_10689,N_8287);
nor U15886 (N_15886,N_9090,N_9657);
nand U15887 (N_15887,N_8798,N_9399);
nor U15888 (N_15888,N_10135,N_10258);
or U15889 (N_15889,N_8708,N_9890);
nor U15890 (N_15890,N_8448,N_8781);
nand U15891 (N_15891,N_9542,N_11905);
or U15892 (N_15892,N_8800,N_10214);
nor U15893 (N_15893,N_11141,N_8393);
nor U15894 (N_15894,N_10124,N_9746);
nor U15895 (N_15895,N_9468,N_10063);
nand U15896 (N_15896,N_11727,N_11298);
nor U15897 (N_15897,N_8472,N_8524);
nand U15898 (N_15898,N_10428,N_11469);
xor U15899 (N_15899,N_11980,N_10616);
nor U15900 (N_15900,N_9719,N_8680);
xor U15901 (N_15901,N_10589,N_11507);
nor U15902 (N_15902,N_10431,N_10517);
or U15903 (N_15903,N_10892,N_8830);
or U15904 (N_15904,N_10888,N_9847);
nand U15905 (N_15905,N_11594,N_9903);
nand U15906 (N_15906,N_10089,N_10564);
xnor U15907 (N_15907,N_9440,N_9080);
or U15908 (N_15908,N_9956,N_8610);
and U15909 (N_15909,N_9015,N_9482);
xnor U15910 (N_15910,N_8907,N_9478);
or U15911 (N_15911,N_8201,N_8116);
and U15912 (N_15912,N_10295,N_11522);
nand U15913 (N_15913,N_11800,N_9215);
and U15914 (N_15914,N_10692,N_8008);
and U15915 (N_15915,N_11239,N_8432);
nand U15916 (N_15916,N_11037,N_10833);
or U15917 (N_15917,N_10084,N_11486);
nand U15918 (N_15918,N_8218,N_11170);
nand U15919 (N_15919,N_10465,N_10281);
or U15920 (N_15920,N_10634,N_8325);
nor U15921 (N_15921,N_8056,N_9527);
nand U15922 (N_15922,N_8965,N_10225);
xnor U15923 (N_15923,N_11294,N_9878);
or U15924 (N_15924,N_11034,N_11622);
or U15925 (N_15925,N_10478,N_11218);
or U15926 (N_15926,N_9597,N_8999);
or U15927 (N_15927,N_8366,N_11570);
nand U15928 (N_15928,N_9380,N_10679);
nand U15929 (N_15929,N_9651,N_10130);
xnor U15930 (N_15930,N_8127,N_11638);
and U15931 (N_15931,N_10672,N_8325);
nand U15932 (N_15932,N_11029,N_9198);
or U15933 (N_15933,N_10885,N_11658);
and U15934 (N_15934,N_10683,N_9976);
xor U15935 (N_15935,N_11814,N_11170);
nor U15936 (N_15936,N_10204,N_11831);
or U15937 (N_15937,N_9517,N_11165);
nor U15938 (N_15938,N_8220,N_8844);
nor U15939 (N_15939,N_11523,N_10613);
nor U15940 (N_15940,N_8213,N_11782);
or U15941 (N_15941,N_10435,N_9200);
or U15942 (N_15942,N_10909,N_11188);
or U15943 (N_15943,N_11574,N_9932);
or U15944 (N_15944,N_9917,N_9582);
nor U15945 (N_15945,N_11506,N_9333);
nand U15946 (N_15946,N_11709,N_11439);
nand U15947 (N_15947,N_10174,N_10531);
nor U15948 (N_15948,N_11251,N_9692);
or U15949 (N_15949,N_9702,N_9778);
and U15950 (N_15950,N_10172,N_10883);
xor U15951 (N_15951,N_8249,N_9872);
xor U15952 (N_15952,N_9841,N_10429);
xor U15953 (N_15953,N_11873,N_8748);
and U15954 (N_15954,N_8676,N_8931);
xnor U15955 (N_15955,N_11236,N_8636);
xnor U15956 (N_15956,N_10630,N_9031);
xnor U15957 (N_15957,N_11735,N_8924);
nand U15958 (N_15958,N_8719,N_10361);
or U15959 (N_15959,N_10520,N_11977);
xor U15960 (N_15960,N_9670,N_9392);
nand U15961 (N_15961,N_8451,N_11912);
nor U15962 (N_15962,N_11682,N_11704);
nor U15963 (N_15963,N_8419,N_9793);
nor U15964 (N_15964,N_8132,N_11365);
xor U15965 (N_15965,N_11706,N_9673);
or U15966 (N_15966,N_10468,N_11255);
and U15967 (N_15967,N_8383,N_8624);
nor U15968 (N_15968,N_11525,N_9796);
and U15969 (N_15969,N_10615,N_9175);
or U15970 (N_15970,N_8812,N_10695);
or U15971 (N_15971,N_9443,N_8094);
or U15972 (N_15972,N_11387,N_8180);
nor U15973 (N_15973,N_9922,N_11834);
and U15974 (N_15974,N_8553,N_10731);
and U15975 (N_15975,N_10846,N_8386);
nand U15976 (N_15976,N_9558,N_10627);
or U15977 (N_15977,N_10735,N_8813);
nand U15978 (N_15978,N_10696,N_9407);
or U15979 (N_15979,N_10107,N_10650);
and U15980 (N_15980,N_10659,N_10764);
nand U15981 (N_15981,N_8583,N_9103);
or U15982 (N_15982,N_8654,N_9149);
xnor U15983 (N_15983,N_9909,N_9293);
xnor U15984 (N_15984,N_8283,N_8204);
nand U15985 (N_15985,N_9486,N_11866);
nor U15986 (N_15986,N_9358,N_10415);
or U15987 (N_15987,N_8100,N_9444);
nor U15988 (N_15988,N_8478,N_8351);
xnor U15989 (N_15989,N_11646,N_8388);
nor U15990 (N_15990,N_11690,N_10445);
and U15991 (N_15991,N_10077,N_8959);
nand U15992 (N_15992,N_9666,N_8260);
or U15993 (N_15993,N_8907,N_11504);
or U15994 (N_15994,N_9209,N_8717);
and U15995 (N_15995,N_9514,N_8728);
nor U15996 (N_15996,N_9327,N_11548);
or U15997 (N_15997,N_9059,N_11565);
xnor U15998 (N_15998,N_9051,N_11292);
nand U15999 (N_15999,N_11476,N_11143);
and U16000 (N_16000,N_12353,N_12008);
or U16001 (N_16001,N_12885,N_14340);
and U16002 (N_16002,N_14994,N_13185);
nand U16003 (N_16003,N_15229,N_14244);
xor U16004 (N_16004,N_15854,N_13024);
and U16005 (N_16005,N_13714,N_14402);
xnor U16006 (N_16006,N_13134,N_15136);
xnor U16007 (N_16007,N_12970,N_12762);
and U16008 (N_16008,N_13957,N_13085);
or U16009 (N_16009,N_12070,N_14866);
and U16010 (N_16010,N_14650,N_15397);
xor U16011 (N_16011,N_15021,N_15283);
and U16012 (N_16012,N_14441,N_13040);
nand U16013 (N_16013,N_12579,N_13995);
nand U16014 (N_16014,N_14872,N_15577);
nor U16015 (N_16015,N_14660,N_14742);
and U16016 (N_16016,N_12368,N_13842);
or U16017 (N_16017,N_12343,N_14109);
and U16018 (N_16018,N_13022,N_15526);
xor U16019 (N_16019,N_15176,N_14853);
nand U16020 (N_16020,N_13588,N_13694);
and U16021 (N_16021,N_13544,N_12703);
nor U16022 (N_16022,N_12243,N_13121);
xor U16023 (N_16023,N_15152,N_15995);
xnor U16024 (N_16024,N_15870,N_15572);
or U16025 (N_16025,N_13920,N_13294);
and U16026 (N_16026,N_15431,N_15480);
nand U16027 (N_16027,N_13048,N_15120);
xnor U16028 (N_16028,N_15316,N_13013);
nor U16029 (N_16029,N_13530,N_14465);
nor U16030 (N_16030,N_12352,N_12534);
nor U16031 (N_16031,N_12587,N_14270);
nand U16032 (N_16032,N_14501,N_12817);
or U16033 (N_16033,N_14392,N_13667);
nor U16034 (N_16034,N_12381,N_15616);
and U16035 (N_16035,N_15991,N_15511);
or U16036 (N_16036,N_13865,N_14530);
xnor U16037 (N_16037,N_13400,N_12224);
and U16038 (N_16038,N_12073,N_12672);
nor U16039 (N_16039,N_14488,N_12053);
or U16040 (N_16040,N_13913,N_12125);
or U16041 (N_16041,N_13613,N_14096);
nor U16042 (N_16042,N_13642,N_15073);
nor U16043 (N_16043,N_15805,N_15005);
nor U16044 (N_16044,N_12198,N_14374);
and U16045 (N_16045,N_13467,N_14756);
and U16046 (N_16046,N_15971,N_15571);
xor U16047 (N_16047,N_13368,N_14970);
and U16048 (N_16048,N_15844,N_12079);
or U16049 (N_16049,N_12895,N_12725);
xor U16050 (N_16050,N_13149,N_15398);
and U16051 (N_16051,N_15912,N_15948);
and U16052 (N_16052,N_15936,N_15047);
nor U16053 (N_16053,N_12156,N_13743);
nor U16054 (N_16054,N_13883,N_12188);
and U16055 (N_16055,N_13100,N_12950);
nor U16056 (N_16056,N_14304,N_14191);
nand U16057 (N_16057,N_13718,N_13773);
and U16058 (N_16058,N_12033,N_15284);
and U16059 (N_16059,N_15430,N_13150);
nand U16060 (N_16060,N_13073,N_13732);
and U16061 (N_16061,N_12722,N_15892);
nor U16062 (N_16062,N_14318,N_13833);
and U16063 (N_16063,N_12558,N_15019);
xor U16064 (N_16064,N_15534,N_12177);
and U16065 (N_16065,N_14447,N_15461);
nor U16066 (N_16066,N_13123,N_13501);
and U16067 (N_16067,N_13899,N_12525);
nand U16068 (N_16068,N_15924,N_13386);
nor U16069 (N_16069,N_15445,N_13958);
xnor U16070 (N_16070,N_15230,N_14512);
and U16071 (N_16071,N_15824,N_15233);
nor U16072 (N_16072,N_14997,N_15266);
xnor U16073 (N_16073,N_12076,N_13515);
nor U16074 (N_16074,N_14554,N_14375);
nand U16075 (N_16075,N_15313,N_15906);
or U16076 (N_16076,N_14503,N_14438);
and U16077 (N_16077,N_12876,N_12946);
or U16078 (N_16078,N_13479,N_15338);
or U16079 (N_16079,N_12975,N_14863);
nand U16080 (N_16080,N_14239,N_12218);
nand U16081 (N_16081,N_13117,N_12489);
nand U16082 (N_16082,N_13858,N_12691);
or U16083 (N_16083,N_15486,N_15950);
or U16084 (N_16084,N_12604,N_13120);
xnor U16085 (N_16085,N_13715,N_15840);
and U16086 (N_16086,N_12554,N_15408);
xor U16087 (N_16087,N_15662,N_15603);
nand U16088 (N_16088,N_14701,N_15114);
xor U16089 (N_16089,N_14149,N_15389);
nand U16090 (N_16090,N_12333,N_12466);
nor U16091 (N_16091,N_15267,N_12618);
or U16092 (N_16092,N_12591,N_15838);
or U16093 (N_16093,N_13115,N_12824);
or U16094 (N_16094,N_14666,N_14152);
nand U16095 (N_16095,N_15998,N_12108);
nor U16096 (N_16096,N_15282,N_13397);
and U16097 (N_16097,N_13829,N_14996);
nor U16098 (N_16098,N_15436,N_15591);
nor U16099 (N_16099,N_14398,N_15209);
nor U16100 (N_16100,N_15368,N_13455);
nor U16101 (N_16101,N_15165,N_12918);
or U16102 (N_16102,N_14927,N_12136);
and U16103 (N_16103,N_15367,N_12199);
and U16104 (N_16104,N_13051,N_15260);
or U16105 (N_16105,N_13355,N_15063);
and U16106 (N_16106,N_13894,N_12271);
nand U16107 (N_16107,N_15192,N_13512);
nand U16108 (N_16108,N_12134,N_15202);
xnor U16109 (N_16109,N_14037,N_14845);
or U16110 (N_16110,N_13432,N_12509);
and U16111 (N_16111,N_14928,N_14547);
xnor U16112 (N_16112,N_14552,N_15536);
nor U16113 (N_16113,N_15538,N_13648);
nand U16114 (N_16114,N_14124,N_15288);
and U16115 (N_16115,N_12653,N_13314);
or U16116 (N_16116,N_12606,N_12598);
or U16117 (N_16117,N_15098,N_15334);
xnor U16118 (N_16118,N_14510,N_14117);
xnor U16119 (N_16119,N_12801,N_12818);
xor U16120 (N_16120,N_14179,N_13356);
nor U16121 (N_16121,N_15447,N_12195);
or U16122 (N_16122,N_12699,N_15708);
or U16123 (N_16123,N_14542,N_15037);
and U16124 (N_16124,N_14361,N_14906);
xor U16125 (N_16125,N_13377,N_13623);
xor U16126 (N_16126,N_12892,N_14017);
and U16127 (N_16127,N_12384,N_12086);
and U16128 (N_16128,N_13854,N_15099);
nor U16129 (N_16129,N_12293,N_13569);
and U16130 (N_16130,N_15032,N_12315);
and U16131 (N_16131,N_12344,N_14550);
or U16132 (N_16132,N_14185,N_13280);
nand U16133 (N_16133,N_15531,N_15770);
and U16134 (N_16134,N_15747,N_13337);
nor U16135 (N_16135,N_15295,N_12562);
or U16136 (N_16136,N_13358,N_13929);
nor U16137 (N_16137,N_13802,N_14540);
and U16138 (N_16138,N_12663,N_14269);
or U16139 (N_16139,N_12694,N_15236);
and U16140 (N_16140,N_15419,N_15305);
and U16141 (N_16141,N_12305,N_15935);
and U16142 (N_16142,N_14704,N_12580);
xor U16143 (N_16143,N_15058,N_12059);
nand U16144 (N_16144,N_12664,N_14246);
or U16145 (N_16145,N_15406,N_15157);
nor U16146 (N_16146,N_13202,N_14846);
nor U16147 (N_16147,N_13195,N_13582);
nand U16148 (N_16148,N_12072,N_13635);
xor U16149 (N_16149,N_12875,N_12584);
nand U16150 (N_16150,N_15756,N_12361);
nand U16151 (N_16151,N_14339,N_12786);
xor U16152 (N_16152,N_13559,N_12829);
and U16153 (N_16153,N_13166,N_13662);
nand U16154 (N_16154,N_14453,N_14710);
xnor U16155 (N_16155,N_13978,N_14468);
or U16156 (N_16156,N_15638,N_12407);
nand U16157 (N_16157,N_14090,N_15439);
or U16158 (N_16158,N_13430,N_12874);
and U16159 (N_16159,N_13934,N_12994);
nor U16160 (N_16160,N_14831,N_12097);
xor U16161 (N_16161,N_12901,N_14781);
and U16162 (N_16162,N_15877,N_15018);
and U16163 (N_16163,N_14966,N_12415);
or U16164 (N_16164,N_13989,N_14419);
nand U16165 (N_16165,N_15641,N_15886);
or U16166 (N_16166,N_14598,N_15839);
nand U16167 (N_16167,N_12745,N_15088);
and U16168 (N_16168,N_12328,N_13423);
nand U16169 (N_16169,N_12091,N_14450);
xor U16170 (N_16170,N_12440,N_13379);
or U16171 (N_16171,N_15787,N_12268);
nand U16172 (N_16172,N_14178,N_12822);
and U16173 (N_16173,N_12768,N_12375);
nor U16174 (N_16174,N_12567,N_13099);
nand U16175 (N_16175,N_12074,N_13760);
and U16176 (N_16176,N_15799,N_12288);
xor U16177 (N_16177,N_14797,N_14665);
nor U16178 (N_16178,N_15469,N_12118);
nand U16179 (N_16179,N_14847,N_12700);
nor U16180 (N_16180,N_14218,N_15275);
xor U16181 (N_16181,N_14464,N_13719);
nor U16182 (N_16182,N_13058,N_13384);
or U16183 (N_16183,N_13723,N_15949);
nor U16184 (N_16184,N_13414,N_14230);
and U16185 (N_16185,N_12056,N_15961);
or U16186 (N_16186,N_12971,N_12696);
or U16187 (N_16187,N_15567,N_12850);
xnor U16188 (N_16188,N_12258,N_15685);
and U16189 (N_16189,N_12411,N_14689);
or U16190 (N_16190,N_12521,N_15816);
nor U16191 (N_16191,N_15774,N_12139);
xnor U16192 (N_16192,N_15198,N_14058);
nand U16193 (N_16193,N_14187,N_12294);
or U16194 (N_16194,N_12857,N_12323);
or U16195 (N_16195,N_13987,N_13381);
nor U16196 (N_16196,N_14955,N_14657);
nand U16197 (N_16197,N_14403,N_12330);
and U16198 (N_16198,N_13407,N_13390);
xor U16199 (N_16199,N_13518,N_14785);
and U16200 (N_16200,N_12648,N_13440);
and U16201 (N_16201,N_14110,N_15166);
nand U16202 (N_16202,N_12940,N_15328);
or U16203 (N_16203,N_13371,N_12427);
xnor U16204 (N_16204,N_12755,N_14265);
and U16205 (N_16205,N_14097,N_12668);
or U16206 (N_16206,N_14498,N_13704);
xor U16207 (N_16207,N_13054,N_15235);
nor U16208 (N_16208,N_15179,N_13770);
nor U16209 (N_16209,N_12821,N_13272);
xnor U16210 (N_16210,N_14770,N_14293);
and U16211 (N_16211,N_14841,N_13266);
nor U16212 (N_16212,N_12853,N_15186);
nand U16213 (N_16213,N_13889,N_13522);
nor U16214 (N_16214,N_14676,N_12608);
nor U16215 (N_16215,N_13462,N_14896);
nor U16216 (N_16216,N_13468,N_14482);
nor U16217 (N_16217,N_12710,N_13309);
or U16218 (N_16218,N_14354,N_12383);
xor U16219 (N_16219,N_14491,N_13447);
nand U16220 (N_16220,N_14397,N_12930);
nand U16221 (N_16221,N_15897,N_15080);
or U16222 (N_16222,N_12684,N_14733);
xor U16223 (N_16223,N_15772,N_12563);
nor U16224 (N_16224,N_12171,N_13621);
and U16225 (N_16225,N_13338,N_12708);
nand U16226 (N_16226,N_15773,N_12005);
nor U16227 (N_16227,N_15505,N_13313);
nor U16228 (N_16228,N_15702,N_12476);
nand U16229 (N_16229,N_14119,N_12908);
nor U16230 (N_16230,N_14065,N_15304);
nand U16231 (N_16231,N_13466,N_15395);
xnor U16232 (N_16232,N_14203,N_15277);
or U16233 (N_16233,N_15119,N_14237);
nand U16234 (N_16234,N_12119,N_14753);
and U16235 (N_16235,N_15732,N_12651);
xnor U16236 (N_16236,N_13231,N_15183);
or U16237 (N_16237,N_13464,N_12233);
or U16238 (N_16238,N_12530,N_15864);
or U16239 (N_16239,N_12779,N_14363);
xor U16240 (N_16240,N_13869,N_13822);
and U16241 (N_16241,N_15409,N_13816);
nor U16242 (N_16242,N_14437,N_15300);
or U16243 (N_16243,N_12756,N_13157);
nand U16244 (N_16244,N_14977,N_13700);
or U16245 (N_16245,N_14499,N_12767);
and U16246 (N_16246,N_15366,N_13003);
and U16247 (N_16247,N_12715,N_12823);
nand U16248 (N_16248,N_15975,N_12403);
and U16249 (N_16249,N_14556,N_15970);
nand U16250 (N_16250,N_15240,N_13665);
nand U16251 (N_16251,N_12652,N_12929);
nor U16252 (N_16252,N_15418,N_12917);
or U16253 (N_16253,N_14856,N_15880);
nor U16254 (N_16254,N_12670,N_12388);
nor U16255 (N_16255,N_15540,N_14036);
and U16256 (N_16256,N_14974,N_15992);
nand U16257 (N_16257,N_13758,N_14003);
nor U16258 (N_16258,N_13285,N_14091);
or U16259 (N_16259,N_15028,N_12448);
xor U16260 (N_16260,N_15384,N_13302);
xnor U16261 (N_16261,N_12002,N_15990);
or U16262 (N_16262,N_14806,N_13260);
nor U16263 (N_16263,N_15330,N_12054);
xnor U16264 (N_16264,N_15673,N_15716);
nand U16265 (N_16265,N_14212,N_13244);
nand U16266 (N_16266,N_14247,N_13975);
and U16267 (N_16267,N_13373,N_14634);
xnor U16268 (N_16268,N_15843,N_13109);
nor U16269 (N_16269,N_13441,N_15051);
nor U16270 (N_16270,N_12522,N_14406);
xor U16271 (N_16271,N_12796,N_13871);
and U16272 (N_16272,N_15889,N_14000);
and U16273 (N_16273,N_14712,N_14999);
or U16274 (N_16274,N_13875,N_15666);
or U16275 (N_16275,N_12758,N_13809);
nand U16276 (N_16276,N_15561,N_13259);
or U16277 (N_16277,N_14102,N_14139);
and U16278 (N_16278,N_14131,N_15378);
and U16279 (N_16279,N_13904,N_15095);
and U16280 (N_16280,N_15132,N_12748);
xnor U16281 (N_16281,N_15464,N_13394);
or U16282 (N_16282,N_14400,N_15713);
nand U16283 (N_16283,N_15331,N_14422);
xnor U16284 (N_16284,N_12516,N_12341);
nand U16285 (N_16285,N_14772,N_14059);
or U16286 (N_16286,N_14953,N_15512);
xor U16287 (N_16287,N_15256,N_12492);
nand U16288 (N_16288,N_15144,N_14624);
xnor U16289 (N_16289,N_14854,N_14415);
and U16290 (N_16290,N_12182,N_14355);
nor U16291 (N_16291,N_12355,N_15882);
xor U16292 (N_16292,N_14352,N_13145);
or U16293 (N_16293,N_13230,N_15108);
xnor U16294 (N_16294,N_12678,N_13977);
nor U16295 (N_16295,N_12458,N_15812);
or U16296 (N_16296,N_12257,N_12799);
or U16297 (N_16297,N_12791,N_13108);
nor U16298 (N_16298,N_13726,N_13248);
xnor U16299 (N_16299,N_12012,N_12193);
nor U16300 (N_16300,N_12178,N_15627);
nor U16301 (N_16301,N_15423,N_14683);
nand U16302 (N_16302,N_12813,N_15011);
xor U16303 (N_16303,N_15215,N_15309);
or U16304 (N_16304,N_12465,N_12172);
nand U16305 (N_16305,N_13321,N_13878);
nor U16306 (N_16306,N_15609,N_15312);
and U16307 (N_16307,N_13520,N_14696);
nor U16308 (N_16308,N_14641,N_14595);
nand U16309 (N_16309,N_13264,N_14381);
or U16310 (N_16310,N_15696,N_13766);
nand U16311 (N_16311,N_14539,N_13942);
nand U16312 (N_16312,N_14262,N_13328);
and U16313 (N_16313,N_15689,N_13255);
nand U16314 (N_16314,N_14489,N_12366);
nand U16315 (N_16315,N_15670,N_15604);
nand U16316 (N_16316,N_12106,N_13892);
nor U16317 (N_16317,N_14055,N_14266);
or U16318 (N_16318,N_15014,N_15139);
and U16319 (N_16319,N_15218,N_14168);
or U16320 (N_16320,N_12599,N_12933);
nor U16321 (N_16321,N_13086,N_15510);
nor U16322 (N_16322,N_14093,N_14827);
and U16323 (N_16323,N_13208,N_12236);
or U16324 (N_16324,N_14703,N_13278);
nor U16325 (N_16325,N_15224,N_15869);
nand U16326 (N_16326,N_15329,N_12246);
xor U16327 (N_16327,N_13606,N_15954);
xor U16328 (N_16328,N_13141,N_12825);
nand U16329 (N_16329,N_15078,N_13031);
nor U16330 (N_16330,N_15010,N_14479);
or U16331 (N_16331,N_15811,N_14599);
nor U16332 (N_16332,N_14444,N_14006);
nand U16333 (N_16333,N_14148,N_15050);
or U16334 (N_16334,N_15668,N_15858);
or U16335 (N_16335,N_15117,N_14534);
nor U16336 (N_16336,N_14757,N_15895);
nor U16337 (N_16337,N_13311,N_13985);
and U16338 (N_16338,N_15500,N_12621);
and U16339 (N_16339,N_12784,N_15519);
xor U16340 (N_16340,N_13463,N_14027);
xor U16341 (N_16341,N_13933,N_12723);
nand U16342 (N_16342,N_12637,N_13542);
and U16343 (N_16343,N_15593,N_12124);
xnor U16344 (N_16344,N_12882,N_14682);
xor U16345 (N_16345,N_13495,N_12986);
and U16346 (N_16346,N_12515,N_12367);
nor U16347 (N_16347,N_13791,N_12585);
or U16348 (N_16348,N_13018,N_14279);
or U16349 (N_16349,N_12300,N_15477);
and U16350 (N_16350,N_14462,N_14805);
xnor U16351 (N_16351,N_12661,N_12350);
or U16352 (N_16352,N_13902,N_14909);
or U16353 (N_16353,N_12497,N_13428);
xor U16354 (N_16354,N_13615,N_15167);
or U16355 (N_16355,N_15530,N_12261);
or U16356 (N_16356,N_13731,N_12886);
xor U16357 (N_16357,N_14649,N_13935);
nand U16358 (N_16358,N_15891,N_14399);
and U16359 (N_16359,N_12281,N_14116);
and U16360 (N_16360,N_13725,N_12701);
and U16361 (N_16361,N_12457,N_15034);
nand U16362 (N_16362,N_14790,N_13911);
xor U16363 (N_16363,N_14362,N_12311);
nand U16364 (N_16364,N_14946,N_15172);
nand U16365 (N_16365,N_15273,N_14427);
nor U16366 (N_16366,N_12265,N_15694);
xnor U16367 (N_16367,N_15046,N_13292);
xor U16368 (N_16368,N_14622,N_14591);
xnor U16369 (N_16369,N_14586,N_13061);
or U16370 (N_16370,N_13560,N_13763);
or U16371 (N_16371,N_14308,N_14963);
nor U16372 (N_16372,N_15589,N_15210);
nand U16373 (N_16373,N_13660,N_14069);
nor U16374 (N_16374,N_13793,N_14889);
nand U16375 (N_16375,N_13133,N_13222);
nand U16376 (N_16376,N_12410,N_12613);
or U16377 (N_16377,N_13136,N_15346);
nand U16378 (N_16378,N_12656,N_13070);
and U16379 (N_16379,N_12215,N_12868);
or U16380 (N_16380,N_14025,N_15463);
xor U16381 (N_16381,N_14186,N_13474);
nand U16382 (N_16382,N_15428,N_15524);
xor U16383 (N_16383,N_12339,N_13749);
nor U16384 (N_16384,N_12942,N_13567);
and U16385 (N_16385,N_13531,N_14233);
nand U16386 (N_16386,N_13279,N_15056);
and U16387 (N_16387,N_13068,N_13446);
nor U16388 (N_16388,N_14633,N_15322);
xor U16389 (N_16389,N_13701,N_13064);
or U16390 (N_16390,N_13286,N_12467);
and U16391 (N_16391,N_13385,N_13658);
and U16392 (N_16392,N_15590,N_12903);
nor U16393 (N_16393,N_15084,N_15916);
nor U16394 (N_16394,N_15135,N_13893);
and U16395 (N_16395,N_14680,N_15247);
nor U16396 (N_16396,N_14394,N_14226);
xnor U16397 (N_16397,N_12095,N_13653);
nand U16398 (N_16398,N_15932,N_13059);
or U16399 (N_16399,N_13383,N_13333);
nor U16400 (N_16400,N_13691,N_12285);
or U16401 (N_16401,N_13299,N_12815);
xor U16402 (N_16402,N_12027,N_14458);
xor U16403 (N_16403,N_13805,N_12941);
nand U16404 (N_16404,N_13332,N_12751);
or U16405 (N_16405,N_14151,N_15111);
xnor U16406 (N_16406,N_14229,N_15009);
and U16407 (N_16407,N_14796,N_15803);
nand U16408 (N_16408,N_15741,N_12235);
or U16409 (N_16409,N_14820,N_14714);
nor U16410 (N_16410,N_13674,N_15206);
xor U16411 (N_16411,N_13004,N_13154);
nand U16412 (N_16412,N_13702,N_13449);
or U16413 (N_16413,N_13663,N_12332);
or U16414 (N_16414,N_12210,N_15197);
nor U16415 (N_16415,N_15353,N_15899);
nand U16416 (N_16416,N_12782,N_12640);
nand U16417 (N_16417,N_12504,N_15944);
or U16418 (N_16418,N_15044,N_13834);
nor U16419 (N_16419,N_14261,N_14267);
or U16420 (N_16420,N_14925,N_12342);
nand U16421 (N_16421,N_13547,N_14662);
or U16422 (N_16422,N_13056,N_13739);
and U16423 (N_16423,N_12559,N_15289);
and U16424 (N_16424,N_13459,N_13354);
xnor U16425 (N_16425,N_13494,N_13376);
and U16426 (N_16426,N_14305,N_14879);
xor U16427 (N_16427,N_14968,N_14590);
and U16428 (N_16428,N_13538,N_12989);
xnor U16429 (N_16429,N_15613,N_15679);
nand U16430 (N_16430,N_12889,N_13951);
or U16431 (N_16431,N_15675,N_12316);
nand U16432 (N_16432,N_15837,N_12928);
and U16433 (N_16433,N_13968,N_15714);
nor U16434 (N_16434,N_13574,N_13888);
or U16435 (N_16435,N_15261,N_12286);
xor U16436 (N_16436,N_15940,N_14720);
and U16437 (N_16437,N_14604,N_12183);
or U16438 (N_16438,N_13523,N_13110);
nand U16439 (N_16439,N_14158,N_15810);
nand U16440 (N_16440,N_12800,N_14306);
nor U16441 (N_16441,N_12911,N_13028);
and U16442 (N_16442,N_14645,N_13856);
and U16443 (N_16443,N_14926,N_13444);
xnor U16444 (N_16444,N_15660,N_14013);
nor U16445 (N_16445,N_13083,N_15631);
nand U16446 (N_16446,N_15158,N_15146);
nor U16447 (N_16447,N_12371,N_13810);
nand U16448 (N_16448,N_15987,N_15758);
xnor U16449 (N_16449,N_15630,N_12159);
nor U16450 (N_16450,N_15841,N_12926);
and U16451 (N_16451,N_15115,N_14615);
nand U16452 (N_16452,N_13839,N_12804);
nand U16453 (N_16453,N_13025,N_14442);
and U16454 (N_16454,N_13140,N_15496);
or U16455 (N_16455,N_14047,N_12409);
nand U16456 (N_16456,N_13063,N_14834);
nor U16457 (N_16457,N_12965,N_13291);
xnor U16458 (N_16458,N_13215,N_15792);
xnor U16459 (N_16459,N_12287,N_13610);
and U16460 (N_16460,N_13811,N_15548);
or U16461 (N_16461,N_14002,N_15988);
nand U16462 (N_16462,N_15997,N_15217);
nand U16463 (N_16463,N_12843,N_14448);
xnor U16464 (N_16464,N_12148,N_13909);
nand U16465 (N_16465,N_15790,N_13919);
or U16466 (N_16466,N_13795,N_12014);
xor U16467 (N_16467,N_13669,N_14976);
or U16468 (N_16468,N_12860,N_14627);
xnor U16469 (N_16469,N_14580,N_14723);
or U16470 (N_16470,N_14287,N_15610);
xnor U16471 (N_16471,N_15723,N_15251);
nand U16472 (N_16472,N_13378,N_13896);
xor U16473 (N_16473,N_15434,N_13183);
nand U16474 (N_16474,N_15101,N_14739);
nand U16475 (N_16475,N_13190,N_13818);
nor U16476 (N_16476,N_13347,N_15539);
xor U16477 (N_16477,N_12690,N_13263);
nor U16478 (N_16478,N_13918,N_12960);
or U16479 (N_16479,N_12772,N_13456);
or U16480 (N_16480,N_15162,N_12162);
and U16481 (N_16481,N_15581,N_15458);
xnor U16482 (N_16482,N_12060,N_15293);
or U16483 (N_16483,N_15110,N_12792);
nor U16484 (N_16484,N_12277,N_14470);
and U16485 (N_16485,N_15624,N_14609);
or U16486 (N_16486,N_13369,N_15865);
or U16487 (N_16487,N_15253,N_12623);
or U16488 (N_16488,N_15559,N_13832);
xor U16489 (N_16489,N_14873,N_14243);
xnor U16490 (N_16490,N_13881,N_12249);
nand U16491 (N_16491,N_13779,N_12679);
or U16492 (N_16492,N_14920,N_13057);
nand U16493 (N_16493,N_13119,N_12998);
xor U16494 (N_16494,N_14326,N_14077);
or U16495 (N_16495,N_15355,N_12961);
nor U16496 (N_16496,N_12462,N_15986);
nand U16497 (N_16497,N_14080,N_15842);
nor U16498 (N_16498,N_15023,N_12577);
and U16499 (N_16499,N_13074,N_13014);
and U16500 (N_16500,N_13817,N_14012);
or U16501 (N_16501,N_14804,N_15007);
xor U16502 (N_16502,N_14589,N_15543);
and U16503 (N_16503,N_12816,N_14718);
or U16504 (N_16504,N_15913,N_13483);
or U16505 (N_16505,N_12044,N_12673);
nor U16506 (N_16506,N_12416,N_14848);
and U16507 (N_16507,N_13304,N_15683);
xor U16508 (N_16508,N_13605,N_15290);
nand U16509 (N_16509,N_13053,N_15254);
nand U16510 (N_16510,N_13603,N_15658);
and U16511 (N_16511,N_15347,N_12113);
nor U16512 (N_16512,N_13290,N_15545);
xnor U16513 (N_16513,N_13664,N_14278);
xor U16514 (N_16514,N_15065,N_12262);
nand U16515 (N_16515,N_12533,N_13124);
nor U16516 (N_16516,N_12956,N_13688);
and U16517 (N_16517,N_12081,N_15821);
nor U16518 (N_16518,N_15532,N_13265);
nand U16519 (N_16519,N_15746,N_14115);
nand U16520 (N_16520,N_14323,N_14505);
or U16521 (N_16521,N_12676,N_12603);
nand U16522 (N_16522,N_14257,N_13079);
xor U16523 (N_16523,N_15719,N_15762);
nand U16524 (N_16524,N_13245,N_14802);
nor U16525 (N_16525,N_12806,N_12031);
or U16526 (N_16526,N_13710,N_12518);
nor U16527 (N_16527,N_15466,N_12234);
or U16528 (N_16528,N_13803,N_13307);
xnor U16529 (N_16529,N_14685,N_14019);
or U16530 (N_16530,N_13938,N_14310);
xor U16531 (N_16531,N_13046,N_15893);
xor U16532 (N_16532,N_12055,N_15653);
nor U16533 (N_16533,N_12098,N_14169);
and U16534 (N_16534,N_15327,N_15173);
and U16535 (N_16535,N_13966,N_15381);
and U16536 (N_16536,N_13607,N_12298);
nand U16537 (N_16537,N_12213,N_15957);
xnor U16538 (N_16538,N_15760,N_13326);
nand U16539 (N_16539,N_14107,N_13203);
or U16540 (N_16540,N_15703,N_13790);
and U16541 (N_16541,N_13257,N_15831);
xor U16542 (N_16542,N_14843,N_15885);
or U16543 (N_16543,N_13585,N_15040);
nor U16544 (N_16544,N_14502,N_13194);
xor U16545 (N_16545,N_12968,N_14205);
nor U16546 (N_16546,N_15123,N_13116);
and U16547 (N_16547,N_15029,N_12879);
nor U16548 (N_16548,N_14150,N_15493);
or U16549 (N_16549,N_12921,N_15319);
or U16550 (N_16550,N_13076,N_15659);
nor U16551 (N_16551,N_15876,N_14652);
and U16552 (N_16552,N_12789,N_15061);
nand U16553 (N_16553,N_14993,N_12483);
xor U16554 (N_16554,N_12514,N_13216);
and U16555 (N_16555,N_13550,N_12369);
and U16556 (N_16556,N_14648,N_12292);
nand U16557 (N_16557,N_14504,N_14838);
nor U16558 (N_16558,N_15748,N_14619);
nor U16559 (N_16559,N_12844,N_14516);
xor U16560 (N_16560,N_15444,N_12493);
xor U16561 (N_16561,N_13780,N_13755);
nand U16562 (N_16562,N_15623,N_13912);
nor U16563 (N_16563,N_13421,N_13860);
nand U16564 (N_16564,N_13946,N_13861);
or U16565 (N_16565,N_15194,N_15656);
and U16566 (N_16566,N_12276,N_15490);
nor U16567 (N_16567,N_15981,N_12624);
or U16568 (N_16568,N_13857,N_15925);
and U16569 (N_16569,N_14803,N_12225);
xnor U16570 (N_16570,N_13435,N_13939);
nand U16571 (N_16571,N_12571,N_15107);
nor U16572 (N_16572,N_12834,N_15953);
nand U16573 (N_16573,N_14771,N_14252);
or U16574 (N_16574,N_15506,N_14023);
nand U16575 (N_16575,N_15104,N_15291);
and U16576 (N_16576,N_15270,N_14043);
or U16577 (N_16577,N_14030,N_14792);
and U16578 (N_16578,N_12163,N_14851);
and U16579 (N_16579,N_14837,N_15875);
nand U16580 (N_16580,N_15642,N_15449);
or U16581 (N_16581,N_14517,N_12160);
and U16582 (N_16582,N_15298,N_12593);
nor U16583 (N_16583,N_12541,N_14167);
nand U16584 (N_16584,N_15456,N_13370);
and U16585 (N_16585,N_14035,N_12473);
nand U16586 (N_16586,N_13983,N_12158);
xnor U16587 (N_16587,N_14668,N_14923);
xnor U16588 (N_16588,N_12902,N_15006);
and U16589 (N_16589,N_12045,N_12977);
xor U16590 (N_16590,N_15048,N_14021);
and U16591 (N_16591,N_13312,N_13774);
xor U16592 (N_16592,N_12220,N_12574);
and U16593 (N_16593,N_15231,N_14018);
and U16594 (N_16594,N_12740,N_12855);
and U16595 (N_16595,N_12006,N_15898);
nand U16596 (N_16596,N_14690,N_12151);
xnor U16597 (N_16597,N_14568,N_14708);
or U16598 (N_16598,N_12283,N_14067);
and U16599 (N_16599,N_12094,N_15438);
nor U16600 (N_16600,N_14232,N_12650);
and U16601 (N_16601,N_13554,N_12726);
and U16602 (N_16602,N_12349,N_12404);
nor U16603 (N_16603,N_14014,N_15580);
or U16604 (N_16604,N_15872,N_14794);
xnor U16605 (N_16605,N_12093,N_14307);
or U16606 (N_16606,N_14766,N_14199);
xor U16607 (N_16607,N_15622,N_15252);
xor U16608 (N_16608,N_13233,N_14902);
nand U16609 (N_16609,N_13593,N_14529);
xor U16610 (N_16610,N_14748,N_12496);
nand U16611 (N_16611,N_12972,N_13672);
nor U16612 (N_16612,N_14587,N_13747);
nand U16613 (N_16613,N_14639,N_12677);
or U16614 (N_16614,N_13961,N_14533);
nand U16615 (N_16615,N_14338,N_12702);
xor U16616 (N_16616,N_13557,N_12190);
or U16617 (N_16617,N_15663,N_13454);
nor U16618 (N_16618,N_15945,N_12635);
nand U16619 (N_16619,N_14424,N_14180);
or U16620 (N_16620,N_15678,N_12142);
nor U16621 (N_16621,N_12067,N_14088);
xnor U16622 (N_16622,N_13325,N_14776);
or U16623 (N_16623,N_13690,N_12746);
and U16624 (N_16624,N_12455,N_15361);
and U16625 (N_16625,N_14862,N_12395);
xor U16626 (N_16626,N_13717,N_12589);
xnor U16627 (N_16627,N_14022,N_14209);
nor U16628 (N_16628,N_15153,N_15620);
and U16629 (N_16629,N_13158,N_14024);
xnor U16630 (N_16630,N_12301,N_13301);
nor U16631 (N_16631,N_14563,N_13005);
and U16632 (N_16632,N_14969,N_12475);
xnor U16633 (N_16633,N_14425,N_15314);
xnor U16634 (N_16634,N_13507,N_15190);
xnor U16635 (N_16635,N_14057,N_13009);
xor U16636 (N_16636,N_14258,N_12413);
and U16637 (N_16637,N_15615,N_15798);
and U16638 (N_16638,N_14176,N_13722);
and U16639 (N_16639,N_12869,N_13931);
or U16640 (N_16640,N_12254,N_12126);
xnor U16641 (N_16641,N_13778,N_13794);
nand U16642 (N_16642,N_13139,N_14749);
or U16643 (N_16643,N_13887,N_14864);
nor U16644 (N_16644,N_14919,N_13424);
xnor U16645 (N_16645,N_13587,N_15090);
or U16646 (N_16646,N_13960,N_12753);
xor U16647 (N_16647,N_13884,N_15460);
nor U16648 (N_16648,N_14317,N_15794);
nor U16649 (N_16649,N_15301,N_15829);
nor U16650 (N_16650,N_12370,N_14369);
nor U16651 (N_16651,N_15244,N_15122);
nand U16652 (N_16652,N_12805,N_12485);
nor U16653 (N_16653,N_15765,N_12472);
nand U16654 (N_16654,N_14432,N_13066);
nand U16655 (N_16655,N_15727,N_13409);
or U16656 (N_16656,N_13306,N_15720);
nor U16657 (N_16657,N_13534,N_14454);
or U16658 (N_16658,N_14998,N_12057);
nand U16659 (N_16659,N_14320,N_14941);
nor U16660 (N_16660,N_12891,N_12004);
xor U16661 (N_16661,N_13580,N_15287);
nor U16662 (N_16662,N_12750,N_14957);
xnor U16663 (N_16663,N_15618,N_13695);
nand U16664 (N_16664,N_13982,N_12322);
or U16665 (N_16665,N_15008,N_12205);
nand U16666 (N_16666,N_15751,N_15067);
and U16667 (N_16667,N_15391,N_12147);
xor U16668 (N_16668,N_15086,N_14347);
or U16669 (N_16669,N_14135,N_15931);
nor U16670 (N_16670,N_12847,N_12674);
or U16671 (N_16671,N_13235,N_15672);
nand U16672 (N_16672,N_15734,N_14223);
xor U16673 (N_16673,N_14121,N_13238);
and U16674 (N_16674,N_15478,N_15412);
nand U16675 (N_16675,N_15781,N_13482);
xnor U16676 (N_16676,N_14647,N_12709);
or U16677 (N_16677,N_15776,N_14576);
nor U16678 (N_16678,N_12038,N_14947);
nand U16679 (N_16679,N_13687,N_13093);
or U16680 (N_16680,N_14282,N_15045);
nor U16681 (N_16681,N_14612,N_13652);
or U16682 (N_16682,N_14490,N_12295);
or U16683 (N_16683,N_15585,N_13303);
or U16684 (N_16684,N_15424,N_15116);
and U16685 (N_16685,N_15066,N_13532);
and U16686 (N_16686,N_15487,N_15553);
or U16687 (N_16687,N_12477,N_14930);
nand U16688 (N_16688,N_14691,N_12146);
nor U16689 (N_16689,N_13436,N_14086);
nor U16690 (N_16690,N_12436,N_15222);
nor U16691 (N_16691,N_14915,N_14737);
nand U16692 (N_16692,N_14706,N_12837);
xnor U16693 (N_16693,N_15292,N_14274);
nand U16694 (N_16694,N_12498,N_14351);
and U16695 (N_16695,N_13282,N_15507);
nor U16696 (N_16696,N_15131,N_15213);
nor U16697 (N_16697,N_13496,N_15557);
nand U16698 (N_16698,N_12110,N_15271);
nand U16699 (N_16699,N_15126,N_14108);
nand U16700 (N_16700,N_13437,N_12351);
xnor U16701 (N_16701,N_13840,N_13492);
nand U16702 (N_16702,N_15907,N_15207);
xor U16703 (N_16703,N_14520,N_14190);
nand U16704 (N_16704,N_12382,N_13801);
xnor U16705 (N_16705,N_13253,N_12536);
nand U16706 (N_16706,N_14493,N_13693);
or U16707 (N_16707,N_14894,N_14137);
nor U16708 (N_16708,N_13320,N_14082);
xnor U16709 (N_16709,N_14521,N_12270);
xnor U16710 (N_16710,N_14087,N_15910);
and U16711 (N_16711,N_13284,N_12164);
xnor U16712 (N_16712,N_15100,N_12675);
and U16713 (N_16713,N_12446,N_15320);
xor U16714 (N_16714,N_13508,N_12916);
nor U16715 (N_16715,N_14601,N_15234);
and U16716 (N_16716,N_15411,N_14852);
and U16717 (N_16717,N_13965,N_14773);
or U16718 (N_16718,N_13457,N_14962);
nand U16719 (N_16719,N_15308,N_15667);
or U16720 (N_16720,N_15817,N_12811);
and U16721 (N_16721,N_15306,N_15909);
or U16722 (N_16722,N_14054,N_13679);
or U16723 (N_16723,N_14536,N_14207);
xor U16724 (N_16724,N_15878,N_15711);
or U16725 (N_16725,N_14545,N_14675);
nor U16726 (N_16726,N_14477,N_13087);
and U16727 (N_16727,N_13570,N_12447);
and U16728 (N_16728,N_14420,N_12775);
and U16729 (N_16729,N_13289,N_14687);
xor U16730 (N_16730,N_15494,N_13706);
nand U16731 (N_16731,N_12468,N_13830);
nor U16732 (N_16732,N_15203,N_14967);
nand U16733 (N_16733,N_15332,N_15392);
and U16734 (N_16734,N_13346,N_12569);
or U16735 (N_16735,N_13173,N_15951);
and U16736 (N_16736,N_14284,N_15709);
or U16737 (N_16737,N_15285,N_12396);
xor U16738 (N_16738,N_12154,N_12399);
nand U16739 (N_16739,N_12766,N_14417);
or U16740 (N_16740,N_15212,N_12572);
nor U16741 (N_16741,N_14163,N_14544);
and U16742 (N_16742,N_14200,N_13042);
xnor U16743 (N_16743,N_15985,N_13258);
nor U16744 (N_16744,N_13470,N_12348);
or U16745 (N_16745,N_13072,N_15016);
or U16746 (N_16746,N_12947,N_12445);
nand U16747 (N_16747,N_13969,N_13350);
and U16748 (N_16748,N_13552,N_13877);
and U16749 (N_16749,N_13944,N_12226);
nor U16750 (N_16750,N_15654,N_12115);
nand U16751 (N_16751,N_14485,N_12963);
and U16752 (N_16752,N_14328,N_12765);
nor U16753 (N_16753,N_15228,N_15164);
and U16754 (N_16754,N_14800,N_12841);
nor U16755 (N_16755,N_15763,N_15200);
or U16756 (N_16756,N_12386,N_15518);
and U16757 (N_16757,N_13419,N_14779);
xor U16758 (N_16758,N_15362,N_12630);
nor U16759 (N_16759,N_15509,N_13172);
and U16760 (N_16760,N_13748,N_14578);
and U16761 (N_16761,N_14588,N_14898);
nor U16762 (N_16762,N_15983,N_14745);
nand U16763 (N_16763,N_14122,N_15470);
nor U16764 (N_16764,N_15551,N_14309);
or U16765 (N_16765,N_14874,N_12944);
xnor U16766 (N_16766,N_14958,N_14154);
nand U16767 (N_16767,N_15879,N_15745);
nor U16768 (N_16768,N_15900,N_14858);
xor U16769 (N_16769,N_13012,N_13019);
xnor U16770 (N_16770,N_12508,N_14812);
or U16771 (N_16771,N_13431,N_13410);
and U16772 (N_16772,N_13819,N_14216);
and U16773 (N_16773,N_15360,N_14337);
or U16774 (N_16774,N_15182,N_12075);
and U16775 (N_16775,N_14421,N_15853);
xor U16776 (N_16776,N_15335,N_12683);
and U16777 (N_16777,N_13214,N_15962);
or U16778 (N_16778,N_15705,N_12241);
nand U16779 (N_16779,N_13254,N_14564);
and U16780 (N_16780,N_14106,N_14064);
xor U16781 (N_16781,N_13319,N_13655);
and U16782 (N_16782,N_13143,N_12145);
or U16783 (N_16783,N_12264,N_13078);
xor U16784 (N_16784,N_15015,N_15674);
xnor U16785 (N_16785,N_12555,N_14694);
nor U16786 (N_16786,N_13848,N_13392);
xor U16787 (N_16787,N_14786,N_14961);
nand U16788 (N_16788,N_14911,N_13427);
or U16789 (N_16789,N_12284,N_15833);
and U16790 (N_16790,N_13647,N_13786);
nor U16791 (N_16791,N_15278,N_13993);
nand U16792 (N_16792,N_12763,N_12718);
nand U16793 (N_16793,N_15697,N_13555);
nand U16794 (N_16794,N_15783,N_13298);
xor U16795 (N_16795,N_14699,N_15919);
or U16796 (N_16796,N_15138,N_15396);
and U16797 (N_16797,N_12432,N_15451);
nand U16798 (N_16798,N_15946,N_13275);
or U16799 (N_16799,N_12469,N_12169);
nor U16800 (N_16800,N_14903,N_12185);
nand U16801 (N_16801,N_13955,N_14071);
nand U16802 (N_16802,N_14395,N_13399);
and U16803 (N_16803,N_14570,N_13497);
and U16804 (N_16804,N_12870,N_12187);
nor U16805 (N_16805,N_12423,N_13439);
and U16806 (N_16806,N_15527,N_12417);
nor U16807 (N_16807,N_14260,N_12007);
xnor U16808 (N_16808,N_13973,N_12966);
nand U16809 (N_16809,N_15168,N_13756);
nor U16810 (N_16810,N_14202,N_14740);
nor U16811 (N_16811,N_15036,N_13262);
and U16812 (N_16812,N_15415,N_13426);
xor U16813 (N_16813,N_12564,N_12083);
xor U16814 (N_16814,N_14656,N_14005);
nor U16815 (N_16815,N_15606,N_12320);
or U16816 (N_16816,N_15219,N_14184);
or U16817 (N_16817,N_15485,N_14522);
xor U16818 (N_16818,N_12704,N_13742);
nor U16819 (N_16819,N_13006,N_13448);
xor U16820 (N_16820,N_14644,N_12736);
and U16821 (N_16821,N_12009,N_12744);
nor U16822 (N_16822,N_13741,N_13945);
xnor U16823 (N_16823,N_14881,N_12336);
nor U16824 (N_16824,N_12540,N_13095);
or U16825 (N_16825,N_15169,N_14312);
and U16826 (N_16826,N_13572,N_12949);
xnor U16827 (N_16827,N_13475,N_12588);
nor U16828 (N_16828,N_15602,N_12480);
xor U16829 (N_16829,N_13198,N_15038);
nand U16830 (N_16830,N_13901,N_13082);
and U16831 (N_16831,N_12638,N_14938);
nor U16832 (N_16832,N_14661,N_13102);
or U16833 (N_16833,N_12781,N_14618);
or U16834 (N_16834,N_13781,N_12317);
nand U16835 (N_16835,N_12737,N_13281);
or U16836 (N_16836,N_13148,N_14007);
xnor U16837 (N_16837,N_13408,N_15068);
or U16838 (N_16838,N_12337,N_13972);
and U16839 (N_16839,N_14754,N_14888);
or U16840 (N_16840,N_13513,N_15976);
or U16841 (N_16841,N_14952,N_13484);
xnor U16842 (N_16842,N_12307,N_14342);
nand U16843 (N_16843,N_14893,N_14391);
and U16844 (N_16844,N_12102,N_12513);
xor U16845 (N_16845,N_12985,N_13703);
and U16846 (N_16846,N_14145,N_14288);
or U16847 (N_16847,N_15646,N_12747);
or U16848 (N_16848,N_15307,N_15339);
and U16849 (N_16849,N_15750,N_13016);
nor U16850 (N_16850,N_14788,N_14053);
and U16851 (N_16851,N_14551,N_12065);
xor U16852 (N_16852,N_13699,N_12743);
and U16853 (N_16853,N_12798,N_14377);
nand U16854 (N_16854,N_15416,N_13608);
or U16855 (N_16855,N_15420,N_12122);
nand U16856 (N_16856,N_15908,N_12063);
xor U16857 (N_16857,N_14204,N_15106);
xnor U16858 (N_16858,N_12887,N_13535);
and U16859 (N_16859,N_14743,N_12302);
nor U16860 (N_16860,N_15550,N_12991);
nor U16861 (N_16861,N_13730,N_13573);
and U16862 (N_16862,N_12017,N_15502);
nor U16863 (N_16863,N_13826,N_14281);
or U16864 (N_16864,N_15280,N_12976);
nand U16865 (N_16865,N_15417,N_14965);
nand U16866 (N_16866,N_12354,N_13796);
or U16867 (N_16867,N_14440,N_14231);
and U16868 (N_16868,N_13249,N_12062);
and U16869 (N_16869,N_15542,N_13502);
nor U16870 (N_16870,N_13372,N_15243);
xnor U16871 (N_16871,N_14433,N_12627);
or U16872 (N_16872,N_13673,N_14144);
and U16873 (N_16873,N_14365,N_12141);
xor U16874 (N_16874,N_13242,N_14388);
xnor U16875 (N_16875,N_15795,N_13943);
or U16876 (N_16876,N_15246,N_15634);
nand U16877 (N_16877,N_12312,N_14378);
nor U16878 (N_16878,N_13698,N_14412);
nor U16879 (N_16879,N_14728,N_15026);
or U16880 (N_16880,N_14734,N_12529);
or U16881 (N_16881,N_12052,N_15105);
and U16882 (N_16882,N_14861,N_12556);
and U16883 (N_16883,N_15124,N_12551);
or U16884 (N_16884,N_13052,N_14343);
nand U16885 (N_16885,N_14253,N_13949);
xnor U16886 (N_16886,N_12208,N_15302);
and U16887 (N_16887,N_12897,N_13343);
or U16888 (N_16888,N_15161,N_14292);
nor U16889 (N_16889,N_14404,N_13953);
and U16890 (N_16890,N_14584,N_13970);
nand U16891 (N_16891,N_14747,N_13753);
xor U16892 (N_16892,N_14767,N_15354);
or U16893 (N_16893,N_13736,N_15484);
nand U16894 (N_16894,N_14042,N_14759);
xor U16895 (N_16895,N_12617,N_15814);
and U16896 (N_16896,N_14789,N_13994);
xor U16897 (N_16897,N_15737,N_14330);
nand U16898 (N_16898,N_14133,N_14436);
or U16899 (N_16899,N_15888,N_15994);
and U16900 (N_16900,N_12430,N_14638);
nand U16901 (N_16901,N_15797,N_13828);
xnor U16902 (N_16902,N_14611,N_12269);
or U16903 (N_16903,N_12741,N_12244);
xnor U16904 (N_16904,N_12168,N_13914);
nand U16905 (N_16905,N_12223,N_12914);
and U16906 (N_16906,N_14494,N_15686);
nand U16907 (N_16907,N_12222,N_15226);
and U16908 (N_16908,N_13937,N_12955);
and U16909 (N_16909,N_14143,N_13420);
nand U16910 (N_16910,N_12573,N_14559);
or U16911 (N_16911,N_15586,N_12978);
or U16912 (N_16912,N_14016,N_13287);
xor U16913 (N_16913,N_14142,N_12935);
nand U16914 (N_16914,N_15272,N_15442);
and U16915 (N_16915,N_12849,N_14836);
and U16916 (N_16916,N_14700,N_14637);
and U16917 (N_16917,N_12616,N_14248);
nand U16918 (N_16918,N_13541,N_15094);
nor U16919 (N_16919,N_12654,N_15850);
nor U16920 (N_16920,N_14428,N_15856);
nor U16921 (N_16921,N_15789,N_12379);
nand U16922 (N_16922,N_14020,N_15255);
nor U16923 (N_16923,N_12420,N_14555);
nand U16924 (N_16924,N_14060,N_14217);
nand U16925 (N_16925,N_12230,N_15757);
or U16926 (N_16926,N_14914,N_12575);
nand U16927 (N_16927,N_13962,N_13917);
nand U16928 (N_16928,N_13524,N_12852);
or U16929 (N_16929,N_12819,N_13161);
nor U16930 (N_16930,N_12019,N_13517);
nor U16931 (N_16931,N_14850,N_12490);
xor U16932 (N_16932,N_14954,N_15941);
nor U16933 (N_16933,N_12561,N_12641);
nor U16934 (N_16934,N_12071,N_15429);
and U16935 (N_16935,N_15363,N_12439);
or U16936 (N_16936,N_14722,N_15488);
xnor U16937 (N_16937,N_14138,N_13241);
and U16938 (N_16938,N_12380,N_13429);
and U16939 (N_16939,N_15237,N_14617);
nor U16940 (N_16940,N_12769,N_13992);
xnor U16941 (N_16941,N_13374,N_13191);
nand U16942 (N_16942,N_14943,N_14942);
nor U16943 (N_16943,N_14583,N_12401);
and U16944 (N_16944,N_14868,N_12152);
nand U16945 (N_16945,N_14807,N_13077);
xnor U16946 (N_16946,N_15569,N_15834);
and U16947 (N_16947,N_13243,N_14684);
nor U16948 (N_16948,N_13310,N_12010);
and U16949 (N_16949,N_13800,N_14473);
xor U16950 (N_16950,N_15150,N_13178);
or U16951 (N_16951,N_13352,N_14670);
or U16952 (N_16952,N_14242,N_14113);
and U16953 (N_16953,N_12738,N_15421);
or U16954 (N_16954,N_12626,N_12565);
and U16955 (N_16955,N_14443,N_12808);
nand U16956 (N_16956,N_14758,N_13256);
and U16957 (N_16957,N_12250,N_15820);
xnor U16958 (N_16958,N_13458,N_13065);
nand U16959 (N_16959,N_13434,N_14198);
nand U16960 (N_16960,N_13020,N_13478);
nor U16961 (N_16961,N_12165,N_13160);
and U16962 (N_16962,N_12391,N_15547);
nor U16963 (N_16963,N_15873,N_13631);
nand U16964 (N_16964,N_12121,N_15584);
xor U16965 (N_16965,N_15448,N_13976);
nor U16966 (N_16966,N_13015,N_14945);
nor U16967 (N_16967,N_12697,N_14172);
and U16968 (N_16968,N_13638,N_14840);
nand U16969 (N_16969,N_14917,N_15336);
xnor U16970 (N_16970,N_12280,N_14594);
and U16971 (N_16971,N_12325,N_15823);
xor U16972 (N_16972,N_14775,N_13422);
nor U16973 (N_16973,N_14674,N_12948);
xor U16974 (N_16974,N_13611,N_13654);
nand U16975 (N_16975,N_14311,N_13798);
and U16976 (N_16976,N_14509,N_14183);
and U16977 (N_16977,N_12717,N_12049);
or U16978 (N_16978,N_15845,N_14877);
or U16979 (N_16979,N_15516,N_15755);
xor U16980 (N_16980,N_12132,N_15939);
nand U16981 (N_16981,N_14089,N_12449);
xnor U16982 (N_16982,N_14129,N_15118);
and U16983 (N_16983,N_12068,N_13936);
xor U16984 (N_16984,N_15785,N_13081);
xnor U16985 (N_16985,N_12842,N_15453);
or U16986 (N_16986,N_14461,N_13490);
nor U16987 (N_16987,N_13342,N_14860);
nand U16988 (N_16988,N_15147,N_15684);
nand U16989 (N_16989,N_14177,N_13080);
xor U16990 (N_16990,N_12080,N_14719);
or U16991 (N_16991,N_15343,N_14950);
and U16992 (N_16992,N_14574,N_12456);
and U16993 (N_16993,N_14396,N_15039);
xor U16994 (N_16994,N_15357,N_13831);
or U16995 (N_16995,N_14672,N_12324);
nand U16996 (N_16996,N_13271,N_13980);
or U16997 (N_16997,N_13846,N_14655);
and U16998 (N_16998,N_14062,N_15340);
xor U16999 (N_16999,N_15759,N_15087);
nor U17000 (N_17000,N_15582,N_13637);
or U17001 (N_17001,N_14164,N_15156);
and U17002 (N_17002,N_13910,N_15724);
nor U17003 (N_17003,N_13711,N_15082);
nand U17004 (N_17004,N_12705,N_14907);
or U17005 (N_17005,N_13090,N_14449);
xnor U17006 (N_17006,N_13131,N_13011);
nor U17007 (N_17007,N_14418,N_14809);
nor U17008 (N_17008,N_15049,N_15220);
nand U17009 (N_17009,N_12867,N_15242);
xnor U17010 (N_17010,N_12934,N_13996);
nor U17011 (N_17011,N_15376,N_14197);
or U17012 (N_17012,N_13329,N_13576);
or U17013 (N_17013,N_14808,N_12107);
or U17014 (N_17014,N_12752,N_15491);
and U17015 (N_17015,N_12035,N_12827);
or U17016 (N_17016,N_13874,N_13783);
or U17017 (N_17017,N_12785,N_14211);
or U17018 (N_17018,N_12778,N_15374);
nor U17019 (N_17019,N_14075,N_15768);
xnor U17020 (N_17020,N_13097,N_15199);
or U17021 (N_17021,N_12306,N_12900);
nor U17022 (N_17022,N_15894,N_12039);
xor U17023 (N_17023,N_14935,N_14986);
nor U17024 (N_17024,N_12266,N_15508);
nand U17025 (N_17025,N_12506,N_15195);
nor U17026 (N_17026,N_15426,N_13824);
nand U17027 (N_17027,N_15558,N_13873);
nor U17028 (N_17028,N_15661,N_13979);
or U17029 (N_17029,N_15079,N_15657);
nor U17030 (N_17030,N_13504,N_14916);
or U17031 (N_17031,N_12064,N_15556);
nand U17032 (N_17032,N_14175,N_12299);
xor U17033 (N_17033,N_14289,N_15070);
nor U17034 (N_17034,N_14389,N_13764);
and U17035 (N_17035,N_14426,N_14810);
nor U17036 (N_17036,N_14567,N_12100);
and U17037 (N_17037,N_15607,N_12474);
nand U17038 (N_17038,N_15276,N_15140);
nand U17039 (N_17039,N_12742,N_15546);
nand U17040 (N_17040,N_12610,N_15977);
or U17041 (N_17041,N_15454,N_12338);
or U17042 (N_17042,N_15379,N_13784);
nor U17043 (N_17043,N_12969,N_12992);
or U17044 (N_17044,N_15151,N_15514);
nand U17045 (N_17045,N_13232,N_14585);
or U17046 (N_17046,N_14553,N_12219);
xnor U17047 (N_17047,N_12832,N_13964);
nand U17048 (N_17048,N_15563,N_14751);
xor U17049 (N_17049,N_14538,N_14524);
and U17050 (N_17050,N_12026,N_15721);
nor U17051 (N_17051,N_14476,N_13196);
xnor U17052 (N_17052,N_15250,N_14671);
nand U17053 (N_17053,N_14153,N_13359);
and U17054 (N_17054,N_14865,N_13661);
nor U17055 (N_17055,N_13096,N_15440);
or U17056 (N_17056,N_12092,N_15232);
xor U17057 (N_17057,N_15482,N_14681);
or U17058 (N_17058,N_13526,N_13349);
xor U17059 (N_17059,N_14677,N_15964);
nor U17060 (N_17060,N_12863,N_15523);
xnor U17061 (N_17061,N_12927,N_14471);
or U17062 (N_17062,N_12291,N_14192);
nor U17063 (N_17063,N_13418,N_12443);
nor U17064 (N_17064,N_13624,N_13225);
and U17065 (N_17065,N_12595,N_15722);
xor U17066 (N_17066,N_13708,N_14275);
and U17067 (N_17067,N_13199,N_12030);
and U17068 (N_17068,N_14379,N_12932);
nand U17069 (N_17069,N_15002,N_14980);
nor U17070 (N_17070,N_14577,N_13201);
xnor U17071 (N_17071,N_15807,N_14372);
and U17072 (N_17072,N_12716,N_12362);
nand U17073 (N_17073,N_13126,N_15625);
nand U17074 (N_17074,N_13709,N_15826);
xnor U17075 (N_17075,N_13098,N_15403);
nand U17076 (N_17076,N_15171,N_13923);
nor U17077 (N_17077,N_12340,N_15390);
xor U17078 (N_17078,N_14201,N_13806);
and U17079 (N_17079,N_12428,N_15069);
nor U17080 (N_17080,N_14349,N_14582);
xor U17081 (N_17081,N_14414,N_14161);
nor U17082 (N_17082,N_13641,N_12500);
and U17083 (N_17083,N_12922,N_12000);
xor U17084 (N_17084,N_15268,N_13029);
nand U17085 (N_17085,N_14359,N_13941);
nand U17086 (N_17086,N_12120,N_14813);
xor U17087 (N_17087,N_12658,N_14407);
and U17088 (N_17088,N_12633,N_13277);
nor U17089 (N_17089,N_14382,N_15955);
and U17090 (N_17090,N_13240,N_15433);
nor U17091 (N_17091,N_12061,N_12890);
or U17092 (N_17092,N_13616,N_15788);
xor U17093 (N_17093,N_12597,N_13525);
nand U17094 (N_17094,N_12713,N_12688);
nor U17095 (N_17095,N_13362,N_12795);
nor U17096 (N_17096,N_14688,N_14206);
nor U17097 (N_17097,N_13948,N_13537);
nor U17098 (N_17098,N_12231,N_14039);
nor U17099 (N_17099,N_13592,N_15052);
xnor U17100 (N_17100,N_12247,N_14483);
and U17101 (N_17101,N_13404,N_13453);
and U17102 (N_17102,N_12576,N_12273);
nand U17103 (N_17103,N_15597,N_15863);
and U17104 (N_17104,N_13239,N_13597);
nor U17105 (N_17105,N_14034,N_13991);
nand U17106 (N_17106,N_14913,N_15178);
nor U17107 (N_17107,N_13577,N_13112);
nor U17108 (N_17108,N_13602,N_13175);
xnor U17109 (N_17109,N_15993,N_12487);
xor U17110 (N_17110,N_13039,N_12943);
and U17111 (N_17111,N_15800,N_13395);
nand U17112 (N_17112,N_13598,N_13211);
nor U17113 (N_17113,N_14387,N_12180);
or U17114 (N_17114,N_14667,N_14259);
or U17115 (N_17115,N_13859,N_15972);
xnor U17116 (N_17116,N_12634,N_12255);
xor U17117 (N_17117,N_14795,N_12858);
or U17118 (N_17118,N_13405,N_13744);
nand U17119 (N_17119,N_13628,N_12279);
xnor U17120 (N_17120,N_12450,N_13599);
nand U17121 (N_17121,N_13252,N_12550);
nor U17122 (N_17122,N_13075,N_12954);
nor U17123 (N_17123,N_15761,N_12984);
xnor U17124 (N_17124,N_14518,N_14887);
xnor U17125 (N_17125,N_15871,N_15942);
and U17126 (N_17126,N_12278,N_14931);
nor U17127 (N_17127,N_15103,N_12217);
nand U17128 (N_17128,N_13300,N_13297);
nor U17129 (N_17129,N_12601,N_13835);
xor U17130 (N_17130,N_12774,N_15109);
and U17131 (N_17131,N_12309,N_15515);
or U17132 (N_17132,N_15216,N_15404);
nand U17133 (N_17133,N_13843,N_15819);
nor U17134 (N_17134,N_14768,N_14451);
and U17135 (N_17135,N_15145,N_14782);
nor U17136 (N_17136,N_12910,N_13044);
xor U17137 (N_17137,N_14038,N_14487);
nor U17138 (N_17138,N_13967,N_12609);
xor U17139 (N_17139,N_15849,N_14083);
xnor U17140 (N_17140,N_15752,N_12032);
nor U17141 (N_17141,N_14240,N_13481);
nand U17142 (N_17142,N_12771,N_15555);
nand U17143 (N_17143,N_15241,N_15093);
nand U17144 (N_17144,N_13156,N_13036);
nor U17145 (N_17145,N_14348,N_14046);
nand U17146 (N_17146,N_12711,N_13591);
nand U17147 (N_17147,N_13761,N_12200);
nand U17148 (N_17148,N_13047,N_14707);
and U17149 (N_17149,N_14249,N_14975);
nor U17150 (N_17150,N_14173,N_13844);
and U17151 (N_17151,N_13209,N_13754);
nand U17152 (N_17152,N_14610,N_15874);
nand U17153 (N_17153,N_13533,N_14826);
xnor U17154 (N_17154,N_15369,N_15933);
xnor U17155 (N_17155,N_15462,N_14651);
nand U17156 (N_17156,N_12041,N_12400);
nor U17157 (N_17157,N_15188,N_12568);
xnor U17158 (N_17158,N_12862,N_12345);
and U17159 (N_17159,N_14673,N_12783);
nand U17160 (N_17160,N_13344,N_12482);
and U17161 (N_17161,N_12528,N_14822);
and U17162 (N_17162,N_14679,N_14384);
or U17163 (N_17163,N_15552,N_15030);
or U17164 (N_17164,N_13493,N_14245);
nor U17165 (N_17165,N_14608,N_15884);
xor U17166 (N_17166,N_12442,N_12374);
nor U17167 (N_17167,N_13155,N_13105);
and U17168 (N_17168,N_14463,N_15092);
nor U17169 (N_17169,N_13144,N_15651);
or U17170 (N_17170,N_15857,N_13412);
or U17171 (N_17171,N_13094,N_13627);
and U17172 (N_17172,N_14910,N_12888);
or U17173 (N_17173,N_13170,N_15326);
or U17174 (N_17174,N_13382,N_15958);
nor U17175 (N_17175,N_13229,N_12835);
xor U17176 (N_17176,N_14761,N_12873);
and U17177 (N_17177,N_13389,N_13879);
and U17178 (N_17178,N_12043,N_14078);
or U17179 (N_17179,N_13506,N_13757);
nand U17180 (N_17180,N_14322,N_14213);
or U17181 (N_17181,N_13510,N_14940);
nand U17182 (N_17182,N_15533,N_15321);
nor U17183 (N_17183,N_14162,N_12175);
nor U17184 (N_17184,N_14350,N_12602);
xor U17185 (N_17185,N_15521,N_13162);
and U17186 (N_17186,N_15341,N_14760);
nor U17187 (N_17187,N_13391,N_12631);
and U17188 (N_17188,N_14074,N_14932);
nand U17189 (N_17189,N_15503,N_15350);
or U17190 (N_17190,N_14335,N_12773);
xnor U17191 (N_17191,N_15201,N_15902);
and U17192 (N_17192,N_15959,N_12952);
nor U17193 (N_17193,N_14193,N_14070);
and U17194 (N_17194,N_13128,N_14746);
and U17195 (N_17195,N_15690,N_15614);
or U17196 (N_17196,N_13581,N_14959);
xor U17197 (N_17197,N_14778,N_12544);
or U17198 (N_17198,N_12174,N_14897);
nand U17199 (N_17199,N_13002,N_13188);
xnor U17200 (N_17200,N_15053,N_13590);
nor U17201 (N_17201,N_12828,N_13807);
xor U17202 (N_17202,N_13954,N_12050);
or U17203 (N_17203,N_15564,N_14621);
and U17204 (N_17204,N_13649,N_12793);
nand U17205 (N_17205,N_14857,N_12803);
and U17206 (N_17206,N_12685,N_13101);
and U17207 (N_17207,N_12957,N_12191);
xor U17208 (N_17208,N_14295,N_12505);
xnor U17209 (N_17209,N_15035,N_15359);
or U17210 (N_17210,N_12760,N_12547);
and U17211 (N_17211,N_13841,N_13341);
or U17212 (N_17212,N_14480,N_13584);
and U17213 (N_17213,N_14466,N_12581);
nand U17214 (N_17214,N_15223,N_13519);
nor U17215 (N_17215,N_12464,N_14044);
xor U17216 (N_17216,N_15373,N_14899);
nand U17217 (N_17217,N_15643,N_12150);
xor U17218 (N_17218,N_15042,N_12461);
xnor U17219 (N_17219,N_13646,N_12069);
nand U17220 (N_17220,N_15476,N_13035);
and U17221 (N_17221,N_12419,N_15479);
nor U17222 (N_17222,N_14455,N_14255);
nand U17223 (N_17223,N_15628,N_14640);
and U17224 (N_17224,N_15380,N_13049);
and U17225 (N_17225,N_12552,N_13771);
xnor U17226 (N_17226,N_14401,N_14068);
nand U17227 (N_17227,N_13692,N_13644);
xnor U17228 (N_17228,N_14603,N_13351);
nand U17229 (N_17229,N_12131,N_14951);
and U17230 (N_17230,N_15358,N_12964);
nand U17231 (N_17231,N_14824,N_15137);
xor U17232 (N_17232,N_12628,N_15655);
nand U17233 (N_17233,N_14511,N_13619);
nand U17234 (N_17234,N_13629,N_14048);
xor U17235 (N_17235,N_15808,N_14755);
or U17236 (N_17236,N_12256,N_12729);
or U17237 (N_17237,N_14405,N_15801);
and U17238 (N_17238,N_15324,N_12211);
nand U17239 (N_17239,N_13836,N_14890);
nand U17240 (N_17240,N_15780,N_12308);
nand U17241 (N_17241,N_13733,N_13707);
nor U17242 (N_17242,N_15474,N_15155);
or U17243 (N_17243,N_15648,N_12542);
nor U17244 (N_17244,N_14170,N_14390);
xor U17245 (N_17245,N_15599,N_13027);
and U17246 (N_17246,N_14219,N_14383);
nand U17247 (N_17247,N_12754,N_12170);
xor U17248 (N_17248,N_14299,N_15513);
and U17249 (N_17249,N_13062,N_15883);
nor U17250 (N_17250,N_15573,N_15520);
or U17251 (N_17251,N_15860,N_12296);
xor U17252 (N_17252,N_14869,N_12221);
or U17253 (N_17253,N_12953,N_14225);
or U17254 (N_17254,N_14527,N_14429);
xnor U17255 (N_17255,N_15859,N_15937);
or U17256 (N_17256,N_12503,N_12356);
and U17257 (N_17257,N_12993,N_14084);
xnor U17258 (N_17258,N_13293,N_12357);
or U17259 (N_17259,N_13334,N_14315);
or U17260 (N_17260,N_13656,N_12155);
xnor U17261 (N_17261,N_15387,N_13527);
xnor U17262 (N_17262,N_13568,N_14762);
xor U17263 (N_17263,N_13738,N_15617);
nor U17264 (N_17264,N_12659,N_15160);
nor U17265 (N_17265,N_15130,N_15184);
xor U17266 (N_17266,N_12667,N_12734);
or U17267 (N_17267,N_13472,N_12437);
or U17268 (N_17268,N_13451,N_13033);
or U17269 (N_17269,N_12334,N_13107);
nand U17270 (N_17270,N_14052,N_15225);
xor U17271 (N_17271,N_12905,N_14605);
nor U17272 (N_17272,N_14344,N_12128);
nand U17273 (N_17273,N_12636,N_15471);
or U17274 (N_17274,N_15127,N_15060);
nor U17275 (N_17275,N_13804,N_13130);
and U17276 (N_17276,N_12216,N_14467);
xor U17277 (N_17277,N_12105,N_15337);
nand U17278 (N_17278,N_14606,N_15296);
nor U17279 (N_17279,N_12421,N_14815);
nand U17280 (N_17280,N_14486,N_12649);
or U17281 (N_17281,N_15437,N_15929);
xnor U17282 (N_17282,N_12112,N_13473);
nand U17283 (N_17283,N_15921,N_14010);
nand U17284 (N_17284,N_13825,N_15731);
xor U17285 (N_17285,N_14987,N_13106);
or U17286 (N_17286,N_13768,N_13189);
nor U17287 (N_17287,N_15544,N_13600);
and U17288 (N_17288,N_13163,N_13797);
xnor U17289 (N_17289,N_15205,N_15177);
xnor U17290 (N_17290,N_12066,N_14985);
or U17291 (N_17291,N_13135,N_15890);
xor U17292 (N_17292,N_13565,N_12470);
nor U17293 (N_17293,N_13247,N_13925);
or U17294 (N_17294,N_12179,N_13268);
nand U17295 (N_17295,N_13926,N_15041);
xor U17296 (N_17296,N_13963,N_12625);
nor U17297 (N_17297,N_15459,N_12424);
nand U17298 (N_17298,N_13633,N_12687);
or U17299 (N_17299,N_12116,N_12084);
or U17300 (N_17300,N_13476,N_12517);
xor U17301 (N_17301,N_15730,N_13388);
or U17302 (N_17302,N_14787,N_15149);
or U17303 (N_17303,N_13882,N_14286);
xnor U17304 (N_17304,N_13589,N_15989);
nor U17305 (N_17305,N_15640,N_15923);
nand U17306 (N_17306,N_13452,N_15855);
nand U17307 (N_17307,N_12881,N_15645);
xor U17308 (N_17308,N_12245,N_14844);
or U17309 (N_17309,N_15264,N_14876);
nor U17310 (N_17310,N_13799,N_12088);
and U17311 (N_17311,N_12491,N_13713);
nand U17312 (N_17312,N_13413,N_15851);
nor U17313 (N_17313,N_15154,N_15649);
nand U17314 (N_17314,N_12251,N_12732);
nor U17315 (N_17315,N_14581,N_12864);
and U17316 (N_17316,N_13177,N_15483);
nand U17317 (N_17317,N_12695,N_12866);
nand U17318 (N_17318,N_14294,N_12662);
xor U17319 (N_17319,N_15349,N_15407);
or U17320 (N_17320,N_12526,N_12089);
nor U17321 (N_17321,N_13549,N_14686);
nand U17322 (N_17322,N_14136,N_13032);
or U17323 (N_17323,N_12201,N_15938);
nor U17324 (N_17324,N_15501,N_14575);
or U17325 (N_17325,N_12877,N_14801);
nor U17326 (N_17326,N_14327,N_13630);
nor U17327 (N_17327,N_12706,N_13626);
nor U17328 (N_17328,N_12924,N_15382);
and U17329 (N_17329,N_14702,N_13720);
xnor U17330 (N_17330,N_14602,N_13677);
nand U17331 (N_17331,N_15033,N_14885);
nor U17332 (N_17332,N_13505,N_15128);
nand U17333 (N_17333,N_14525,N_13974);
nand U17334 (N_17334,N_13445,N_13411);
xnor U17335 (N_17335,N_14892,N_13200);
and U17336 (N_17336,N_14408,N_15239);
nor U17337 (N_17337,N_12728,N_12435);
and U17338 (N_17338,N_13571,N_14004);
nor U17339 (N_17339,N_12721,N_14819);
xnor U17340 (N_17340,N_14120,N_12846);
nor U17341 (N_17341,N_13317,N_12013);
nor U17342 (N_17342,N_15450,N_15262);
nor U17343 (N_17343,N_13489,N_14264);
nor U17344 (N_17344,N_15861,N_13705);
or U17345 (N_17345,N_13366,N_12167);
nor U17346 (N_17346,N_12967,N_14368);
nor U17347 (N_17347,N_15583,N_12883);
and U17348 (N_17348,N_12981,N_15779);
or U17349 (N_17349,N_12714,N_14596);
and U17350 (N_17350,N_13151,N_12532);
or U17351 (N_17351,N_14921,N_13528);
xor U17352 (N_17352,N_12021,N_12974);
and U17353 (N_17353,N_12520,N_12951);
or U17354 (N_17354,N_14492,N_15669);
xnor U17355 (N_17355,N_15435,N_15973);
or U17356 (N_17356,N_13168,N_15457);
nand U17357 (N_17357,N_15728,N_15952);
nand U17358 (N_17358,N_14416,N_12712);
nor U17359 (N_17359,N_13529,N_14535);
nand U17360 (N_17360,N_13792,N_14313);
or U17361 (N_17361,N_15681,N_13330);
and U17362 (N_17362,N_12620,N_15286);
and U17363 (N_17363,N_12945,N_12390);
nor U17364 (N_17364,N_14283,N_12749);
xnor U17365 (N_17365,N_14385,N_14469);
nand U17366 (N_17366,N_14981,N_12788);
or U17367 (N_17367,N_13169,N_13380);
and U17368 (N_17368,N_15960,N_12479);
nor U17369 (N_17369,N_14280,N_15492);
nand U17370 (N_17370,N_15978,N_13539);
or U17371 (N_17371,N_13487,N_15142);
xor U17372 (N_17372,N_13220,N_12898);
nand U17373 (N_17373,N_12878,N_14112);
nand U17374 (N_17374,N_14769,N_14777);
xor U17375 (N_17375,N_14642,N_14445);
nand U17376 (N_17376,N_15809,N_12425);
or U17377 (N_17377,N_12318,N_15356);
xnor U17378 (N_17378,N_15980,N_15969);
nand U17379 (N_17379,N_12511,N_12939);
xor U17380 (N_17380,N_14726,N_14565);
nor U17381 (N_17381,N_13900,N_15535);
nand U17382 (N_17382,N_14157,N_14519);
or U17383 (N_17383,N_15180,N_15465);
or U17384 (N_17384,N_15413,N_13762);
or U17385 (N_17385,N_12826,N_15281);
or U17386 (N_17386,N_14663,N_13561);
xnor U17387 (N_17387,N_13498,N_13928);
nand U17388 (N_17388,N_13553,N_12310);
or U17389 (N_17389,N_15560,N_13682);
xor U17390 (N_17390,N_14984,N_14964);
nand U17391 (N_17391,N_15725,N_15928);
nor U17392 (N_17392,N_14548,N_15733);
nand U17393 (N_17393,N_14346,N_13551);
or U17394 (N_17394,N_14870,N_14049);
and U17395 (N_17395,N_12720,N_13226);
nor U17396 (N_17396,N_14592,N_12962);
or U17397 (N_17397,N_13192,N_12321);
nand U17398 (N_17398,N_12189,N_14526);
or U17399 (N_17399,N_15963,N_12166);
nand U17400 (N_17400,N_15600,N_12260);
nor U17401 (N_17401,N_12707,N_13678);
and U17402 (N_17402,N_13906,N_13091);
nand U17403 (N_17403,N_14228,N_12655);
nand U17404 (N_17404,N_15739,N_14571);
nand U17405 (N_17405,N_12724,N_13251);
and U17406 (N_17406,N_14285,N_15914);
and U17407 (N_17407,N_15652,N_12909);
and U17408 (N_17408,N_13227,N_15299);
nand U17409 (N_17409,N_14654,N_14331);
or U17410 (N_17410,N_13092,N_14832);
xnor U17411 (N_17411,N_15204,N_14227);
nand U17412 (N_17412,N_13668,N_15031);
nor U17413 (N_17413,N_15664,N_15749);
nor U17414 (N_17414,N_13375,N_15371);
nor U17415 (N_17415,N_14716,N_15704);
nand U17416 (N_17416,N_12327,N_15771);
xor U17417 (N_17417,N_12036,N_13586);
or U17418 (N_17418,N_12988,N_15796);
nand U17419 (N_17419,N_14357,N_14236);
or U17420 (N_17420,N_13684,N_14001);
or U17421 (N_17421,N_13815,N_14628);
nor U17422 (N_17422,N_14949,N_15806);
nand U17423 (N_17423,N_14936,N_13625);
and U17424 (N_17424,N_14345,N_15815);
nand U17425 (N_17425,N_14156,N_15394);
or U17426 (N_17426,N_13721,N_12906);
xor U17427 (N_17427,N_15742,N_13812);
nor U17428 (N_17428,N_12378,N_12214);
nor U17429 (N_17429,N_13043,N_13336);
xnor U17430 (N_17430,N_12184,N_13315);
xor U17431 (N_17431,N_15141,N_14367);
nand U17432 (N_17432,N_12326,N_12077);
or U17433 (N_17433,N_15982,N_13323);
or U17434 (N_17434,N_15566,N_13863);
nand U17435 (N_17435,N_14659,N_12037);
and U17436 (N_17436,N_14353,N_15113);
nand U17437 (N_17437,N_14741,N_13981);
and U17438 (N_17438,N_13088,N_12194);
xor U17439 (N_17439,N_15813,N_13988);
xor U17440 (N_17440,N_12471,N_15791);
or U17441 (N_17441,N_14456,N_12546);
and U17442 (N_17442,N_13516,N_13008);
nor U17443 (N_17443,N_14558,N_14623);
or U17444 (N_17444,N_15133,N_14324);
xor U17445 (N_17445,N_13821,N_13886);
and U17446 (N_17446,N_12983,N_12831);
and U17447 (N_17447,N_15024,N_15081);
nor U17448 (N_17448,N_15377,N_12501);
nand U17449 (N_17449,N_12431,N_12402);
nand U17450 (N_17450,N_12358,N_13167);
xor U17451 (N_17451,N_13234,N_12149);
and U17452 (N_17452,N_15102,N_12347);
xor U17453 (N_17453,N_13401,N_12232);
xnor U17454 (N_17454,N_15375,N_15588);
and U17455 (N_17455,N_12586,N_14298);
nor U17456 (N_17456,N_15517,N_15984);
or U17457 (N_17457,N_15637,N_12733);
and U17458 (N_17458,N_14948,N_15825);
nand U17459 (N_17459,N_15621,N_15579);
or U17460 (N_17460,N_13675,N_15441);
xnor U17461 (N_17461,N_13728,N_15592);
or U17462 (N_17462,N_12143,N_14515);
or U17463 (N_17463,N_15020,N_12412);
and U17464 (N_17464,N_15608,N_13417);
and U17465 (N_17465,N_14114,N_15400);
xnor U17466 (N_17466,N_13138,N_12524);
and U17467 (N_17467,N_15832,N_14513);
or U17468 (N_17468,N_12931,N_12809);
nand U17469 (N_17469,N_15074,N_15904);
nand U17470 (N_17470,N_12359,N_12303);
xor U17471 (N_17471,N_14410,N_14105);
nand U17472 (N_17472,N_12204,N_14234);
nand U17473 (N_17473,N_14371,N_14924);
or U17474 (N_17474,N_15896,N_13206);
xnor U17475 (N_17475,N_13870,N_13069);
xor U17476 (N_17476,N_14692,N_14995);
nor U17477 (N_17477,N_12594,N_14496);
and U17478 (N_17478,N_12274,N_14562);
or U17479 (N_17479,N_13324,N_15001);
or U17480 (N_17480,N_14056,N_12459);
nand U17481 (N_17481,N_12376,N_15249);
xnor U17482 (N_17482,N_15000,N_13480);
or U17483 (N_17483,N_14884,N_15769);
nand U17484 (N_17484,N_15947,N_12657);
nand U17485 (N_17485,N_14823,N_14336);
nand U17486 (N_17486,N_14956,N_13142);
or U17487 (N_17487,N_14978,N_14625);
and U17488 (N_17488,N_13485,N_15767);
xor U17489 (N_17489,N_13880,N_14829);
and U17490 (N_17490,N_15943,N_13111);
nand U17491 (N_17491,N_13276,N_15729);
xor U17492 (N_17492,N_13514,N_13639);
and U17493 (N_17493,N_12512,N_15818);
nand U17494 (N_17494,N_12660,N_12639);
nor U17495 (N_17495,N_12919,N_15279);
nor U17496 (N_17496,N_14155,N_15633);
nor U17497 (N_17497,N_13556,N_13897);
or U17498 (N_17498,N_13387,N_14597);
and U17499 (N_17499,N_13898,N_15934);
and U17500 (N_17500,N_14439,N_12510);
and U17501 (N_17501,N_14973,N_15071);
or U17502 (N_17502,N_12196,N_14717);
nand U17503 (N_17503,N_15159,N_14041);
and U17504 (N_17504,N_12228,N_13643);
nor U17505 (N_17505,N_14210,N_15351);
nand U17506 (N_17506,N_14991,N_13997);
or U17507 (N_17507,N_12936,N_13433);
xor U17508 (N_17508,N_15263,N_13885);
nand U17509 (N_17509,N_13971,N_13712);
nor U17510 (N_17510,N_12346,N_13037);
or U17511 (N_17511,N_15782,N_12363);
nand U17512 (N_17512,N_13907,N_12085);
or U17513 (N_17513,N_12408,N_14140);
and U17514 (N_17514,N_15181,N_14334);
or U17515 (N_17515,N_12915,N_12777);
or U17516 (N_17516,N_15786,N_15710);
xnor U17517 (N_17517,N_15422,N_15075);
xnor U17518 (N_17518,N_14653,N_12814);
nand U17519 (N_17519,N_13845,N_14664);
xnor U17520 (N_17520,N_13813,N_15446);
or U17521 (N_17521,N_15650,N_12761);
nand U17522 (N_17522,N_14573,N_13503);
nand U17523 (N_17523,N_14905,N_15852);
xor U17524 (N_17524,N_12980,N_15753);
nand U17525 (N_17525,N_15866,N_14174);
nor U17526 (N_17526,N_15352,N_15027);
xnor U17527 (N_17527,N_15915,N_13636);
nor U17528 (N_17528,N_13578,N_13659);
nand U17529 (N_17529,N_14393,N_13159);
or U17530 (N_17530,N_12313,N_15405);
or U17531 (N_17531,N_14697,N_12871);
xor U17532 (N_17532,N_14992,N_12133);
nor U17533 (N_17533,N_12666,N_12488);
xnor U17534 (N_17534,N_12790,N_14904);
nand U17535 (N_17535,N_13363,N_12289);
xor U17536 (N_17536,N_13127,N_14103);
xor U17537 (N_17537,N_15903,N_14871);
or U17538 (N_17538,N_12463,N_15576);
nand U17539 (N_17539,N_14166,N_15383);
nor U17540 (N_17540,N_14630,N_14215);
xor U17541 (N_17541,N_15017,N_15549);
nand U17542 (N_17542,N_14263,N_14072);
and U17543 (N_17543,N_13890,N_15294);
and U17544 (N_17544,N_13308,N_15594);
nor U17545 (N_17545,N_13751,N_13217);
or U17546 (N_17546,N_12698,N_12797);
nor U17547 (N_17547,N_14631,N_12611);
and U17548 (N_17548,N_14933,N_14181);
nor U17549 (N_17549,N_12499,N_14459);
nor U17550 (N_17550,N_15979,N_15699);
nor U17551 (N_17551,N_15297,N_12240);
and U17552 (N_17552,N_14744,N_13345);
or U17553 (N_17553,N_12140,N_13984);
nor U17554 (N_17554,N_12523,N_15055);
nand U17555 (N_17555,N_12820,N_14329);
and U17556 (N_17556,N_15125,N_13916);
or U17557 (N_17557,N_14735,N_13060);
or U17558 (N_17558,N_13267,N_13396);
xor U17559 (N_17559,N_14646,N_12377);
nor U17560 (N_17560,N_13847,N_15682);
and U17561 (N_17561,N_14031,N_13041);
and U17562 (N_17562,N_14901,N_14549);
or U17563 (N_17563,N_14481,N_14238);
or U17564 (N_17564,N_13067,N_14818);
and U17565 (N_17565,N_14989,N_15967);
nand U17566 (N_17566,N_15208,N_15974);
nor U17567 (N_17567,N_13787,N_14763);
and U17568 (N_17568,N_13734,N_13488);
and U17569 (N_17569,N_15905,N_12048);
nand U17570 (N_17570,N_14918,N_13339);
nor U17571 (N_17571,N_12907,N_14214);
and U17572 (N_17572,N_14126,N_13634);
nand U17573 (N_17573,N_13536,N_12111);
nand U17574 (N_17574,N_15802,N_14332);
xnor U17575 (N_17575,N_12859,N_14709);
or U17576 (N_17576,N_12838,N_14099);
nor U17577 (N_17577,N_13186,N_12787);
or U17578 (N_17578,N_12290,N_13566);
and U17579 (N_17579,N_13775,N_14423);
nor U17580 (N_17580,N_12925,N_13769);
nand U17581 (N_17581,N_13952,N_13361);
and U17582 (N_17582,N_15345,N_12642);
and U17583 (N_17583,N_15766,N_14886);
xor U17584 (N_17584,N_15775,N_13724);
xor U17585 (N_17585,N_15868,N_14732);
nand U17586 (N_17586,N_13104,N_15570);
xor U17587 (N_17587,N_14095,N_12114);
or U17588 (N_17588,N_14695,N_13558);
nor U17589 (N_17589,N_14051,N_12872);
or U17590 (N_17590,N_13563,N_12647);
xnor U17591 (N_17591,N_12839,N_12494);
xor U17592 (N_17592,N_14291,N_13986);
xnor U17593 (N_17593,N_14579,N_13165);
nor U17594 (N_17594,N_14254,N_14127);
nor U17595 (N_17595,N_14146,N_13348);
or U17596 (N_17596,N_15386,N_12028);
xor U17597 (N_17597,N_13545,N_14495);
nor U17598 (N_17598,N_14960,N_14616);
or U17599 (N_17599,N_15013,N_15846);
nand U17600 (N_17600,N_13864,N_12212);
xnor U17601 (N_17601,N_14821,N_14982);
nor U17602 (N_17602,N_12087,N_15175);
and U17603 (N_17603,N_12253,N_12548);
or U17604 (N_17604,N_12912,N_14061);
nand U17605 (N_17605,N_14358,N_12040);
and U17606 (N_17606,N_15784,N_15163);
nand U17607 (N_17607,N_15717,N_15927);
and U17608 (N_17608,N_13670,N_13283);
nor U17609 (N_17609,N_14111,N_13789);
nand U17610 (N_17610,N_15498,N_15043);
nor U17611 (N_17611,N_12263,N_15887);
nand U17612 (N_17612,N_13823,N_13746);
or U17613 (N_17613,N_12719,N_15695);
nor U17614 (N_17614,N_15265,N_13450);
or U17615 (N_17615,N_15830,N_14944);
or U17616 (N_17616,N_12138,N_15691);
and U17617 (N_17617,N_12392,N_14273);
and U17618 (N_17618,N_12051,N_14658);
and U17619 (N_17619,N_15735,N_12123);
nor U17620 (N_17620,N_13940,N_13500);
nand U17621 (N_17621,N_14572,N_14188);
nor U17622 (N_17622,N_15059,N_13164);
and U17623 (N_17623,N_14882,N_13543);
or U17624 (N_17624,N_12209,N_14875);
or U17625 (N_17625,N_15568,N_13132);
and U17626 (N_17626,N_15248,N_15636);
nor U17627 (N_17627,N_14983,N_12206);
nor U17628 (N_17628,N_15687,N_14370);
xnor U17629 (N_17629,N_13210,N_12802);
nor U17630 (N_17630,N_14277,N_14132);
or U17631 (N_17631,N_12387,N_12144);
nor U17632 (N_17632,N_15054,N_14040);
nand U17633 (N_17633,N_14460,N_14409);
or U17634 (N_17634,N_15671,N_14045);
nor U17635 (N_17635,N_13460,N_15999);
nor U17636 (N_17636,N_12537,N_15676);
or U17637 (N_17637,N_12003,N_15410);
nand U17638 (N_17638,N_15743,N_12203);
nand U17639 (N_17639,N_14032,N_13393);
or U17640 (N_17640,N_12426,N_15259);
or U17641 (N_17641,N_12854,N_15452);
xnor U17642 (N_17642,N_15647,N_12973);
nand U17643 (N_17643,N_12810,N_14125);
nand U17644 (N_17644,N_12938,N_13327);
xor U17645 (N_17645,N_12937,N_12757);
or U17646 (N_17646,N_15966,N_13038);
and U17647 (N_17647,N_14507,N_15311);
xor U17648 (N_17648,N_12680,N_15835);
or U17649 (N_17649,N_13666,N_15578);
and U17650 (N_17650,N_15333,N_12275);
and U17651 (N_17651,N_15700,N_15274);
or U17652 (N_17652,N_13891,N_14325);
nor U17653 (N_17653,N_14929,N_13224);
nand U17654 (N_17654,N_14430,N_13017);
nor U17655 (N_17655,N_13686,N_13609);
nand U17656 (N_17656,N_14828,N_13221);
and U17657 (N_17657,N_13905,N_14251);
xnor U17658 (N_17658,N_12329,N_14835);
nand U17659 (N_17659,N_12692,N_15701);
and U17660 (N_17660,N_12181,N_12414);
or U17661 (N_17661,N_14891,N_13270);
xor U17662 (N_17662,N_14321,N_12686);
or U17663 (N_17663,N_14290,N_15497);
or U17664 (N_17664,N_15097,N_13179);
xor U17665 (N_17665,N_14731,N_14523);
xor U17666 (N_17666,N_13583,N_12671);
nor U17667 (N_17667,N_12365,N_15468);
xnor U17668 (N_17668,N_12023,N_15414);
or U17669 (N_17669,N_14736,N_14614);
nand U17670 (N_17670,N_12693,N_13402);
or U17671 (N_17671,N_14130,N_13007);
nor U17672 (N_17672,N_15740,N_12776);
and U17673 (N_17673,N_14271,N_14883);
nand U17674 (N_17674,N_14380,N_13657);
xor U17675 (N_17675,N_12644,N_13486);
nand U17676 (N_17676,N_15170,N_12535);
or U17677 (N_17677,N_13295,N_12130);
nand U17678 (N_17678,N_13903,N_14431);
nor U17679 (N_17679,N_15004,N_14600);
xor U17680 (N_17680,N_12047,N_13146);
nor U17681 (N_17681,N_12096,N_15303);
nand U17682 (N_17682,N_14319,N_13921);
nor U17683 (N_17683,N_13425,N_15587);
and U17684 (N_17684,N_15930,N_13765);
or U17685 (N_17685,N_15385,N_14333);
xor U17686 (N_17686,N_12632,N_12157);
nor U17687 (N_17687,N_12364,N_13956);
nor U17688 (N_17688,N_15881,N_12135);
nor U17689 (N_17689,N_15601,N_12893);
or U17690 (N_17690,N_13596,N_12999);
or U17691 (N_17691,N_13685,N_13228);
xnor U17692 (N_17692,N_13564,N_14301);
xor U17693 (N_17693,N_13612,N_15827);
and U17694 (N_17694,N_14194,N_12899);
or U17695 (N_17695,N_13113,N_12539);
nor U17696 (N_17696,N_15777,N_14303);
nor U17697 (N_17697,N_15495,N_14452);
or U17698 (N_17698,N_13614,N_12669);
nor U17699 (N_17699,N_13316,N_12229);
and U17700 (N_17700,N_13862,N_15121);
xor U17701 (N_17701,N_15342,N_12979);
nand U17702 (N_17702,N_15754,N_12109);
and U17703 (N_17703,N_12304,N_13772);
or U17704 (N_17704,N_14085,N_12481);
xor U17705 (N_17705,N_12619,N_14607);
nand U17706 (N_17706,N_14546,N_15189);
nor U17707 (N_17707,N_14752,N_12101);
and U17708 (N_17708,N_13808,N_13000);
and U17709 (N_17709,N_12197,N_13676);
or U17710 (N_17710,N_12997,N_12607);
and U17711 (N_17711,N_13360,N_12836);
and U17712 (N_17712,N_14593,N_14478);
or U17713 (N_17713,N_13050,N_14566);
xnor U17714 (N_17714,N_15922,N_14798);
or U17715 (N_17715,N_12605,N_14557);
and U17716 (N_17716,N_13999,N_14715);
and U17717 (N_17717,N_13604,N_12995);
nor U17718 (N_17718,N_15402,N_14241);
nor U17719 (N_17719,N_13153,N_15804);
nor U17720 (N_17720,N_13322,N_13895);
nor U17721 (N_17721,N_15245,N_12643);
nand U17722 (N_17722,N_15965,N_15718);
nand U17723 (N_17723,N_14134,N_12373);
nor U17724 (N_17724,N_12406,N_14972);
xnor U17725 (N_17725,N_14356,N_13837);
and U17726 (N_17726,N_13876,N_12560);
nand U17727 (N_17727,N_14101,N_13204);
xor U17728 (N_17728,N_15688,N_12453);
or U17729 (N_17729,N_15611,N_15096);
xnor U17730 (N_17730,N_15901,N_13908);
or U17731 (N_17731,N_15425,N_12011);
nor U17732 (N_17732,N_12495,N_13415);
xnor U17733 (N_17733,N_15238,N_14939);
or U17734 (N_17734,N_15698,N_15193);
and U17735 (N_17735,N_13782,N_15393);
xor U17736 (N_17736,N_13915,N_13010);
or U17737 (N_17737,N_14297,N_13727);
nor U17738 (N_17738,N_15525,N_14765);
nand U17739 (N_17739,N_14009,N_13171);
nor U17740 (N_17740,N_12078,N_15148);
and U17741 (N_17741,N_12527,N_13750);
or U17742 (N_17742,N_12982,N_12845);
nand U17743 (N_17743,N_13814,N_14620);
and U17744 (N_17744,N_15227,N_15083);
xnor U17745 (N_17745,N_13403,N_13187);
and U17746 (N_17746,N_15918,N_15529);
nand U17747 (N_17747,N_14411,N_14066);
xnor U17748 (N_17748,N_15793,N_12557);
nand U17749 (N_17749,N_14366,N_15012);
or U17750 (N_17750,N_12018,N_13318);
nor U17751 (N_17751,N_12025,N_12385);
nand U17752 (N_17752,N_14880,N_12029);
or U17753 (N_17753,N_14435,N_15715);
nand U17754 (N_17754,N_13250,N_15712);
nand U17755 (N_17755,N_12001,N_14839);
nand U17756 (N_17756,N_12622,N_13034);
nor U17757 (N_17757,N_15911,N_12259);
or U17758 (N_17758,N_13180,N_12959);
and U17759 (N_17759,N_13406,N_12807);
nand U17760 (N_17760,N_12848,N_12996);
xor U17761 (N_17761,N_12227,N_15370);
xor U17762 (N_17762,N_12582,N_13236);
nor U17763 (N_17763,N_13205,N_15057);
nand U17764 (N_17764,N_14678,N_13021);
and U17765 (N_17765,N_15143,N_12770);
nor U17766 (N_17766,N_12764,N_15364);
nor U17767 (N_17767,N_12681,N_15596);
nand U17768 (N_17768,N_14937,N_14693);
or U17769 (N_17769,N_12237,N_14222);
or U17770 (N_17770,N_12833,N_14705);
nand U17771 (N_17771,N_12252,N_14457);
nand U17772 (N_17772,N_15076,N_14922);
or U17773 (N_17773,N_13594,N_13745);
xnor U17774 (N_17774,N_13927,N_13465);
nand U17775 (N_17775,N_14118,N_14302);
nor U17776 (N_17776,N_13071,N_15214);
and U17777 (N_17777,N_15632,N_12238);
nor U17778 (N_17778,N_14235,N_15022);
nand U17779 (N_17779,N_13932,N_13767);
and U17780 (N_17780,N_15562,N_12104);
xor U17781 (N_17781,N_13867,N_15574);
nand U17782 (N_17782,N_13219,N_15612);
nor U17783 (N_17783,N_12583,N_13548);
nand U17784 (N_17784,N_13562,N_13471);
or U17785 (N_17785,N_12486,N_14830);
nor U17786 (N_17786,N_14833,N_13777);
or U17787 (N_17787,N_14123,N_14472);
xor U17788 (N_17788,N_13990,N_13129);
xor U17789 (N_17789,N_12856,N_14094);
nor U17790 (N_17790,N_14272,N_13030);
xnor U17791 (N_17791,N_12433,N_14780);
nor U17792 (N_17792,N_15504,N_15848);
nand U17793 (N_17793,N_12015,N_13595);
nor U17794 (N_17794,N_14500,N_14698);
or U17795 (N_17795,N_15427,N_13193);
or U17796 (N_17796,N_12538,N_13274);
and U17797 (N_17797,N_13511,N_15639);
nand U17798 (N_17798,N_14934,N_14855);
and U17799 (N_17799,N_13357,N_12046);
nand U17800 (N_17800,N_12082,N_15003);
and U17801 (N_17801,N_14063,N_13601);
nand U17802 (N_17802,N_12207,N_15554);
nand U17803 (N_17803,N_12502,N_14250);
nor U17804 (N_17804,N_12880,N_12830);
nor U17805 (N_17805,N_15085,N_14076);
nand U17806 (N_17806,N_12507,N_14475);
or U17807 (N_17807,N_14912,N_13855);
nor U17808 (N_17808,N_13103,N_13924);
or U17809 (N_17809,N_12331,N_14613);
xnor U17810 (N_17810,N_14171,N_14195);
nand U17811 (N_17811,N_14636,N_15062);
nor U17812 (N_17812,N_13579,N_13650);
nor U17813 (N_17813,N_15707,N_12739);
nand U17814 (N_17814,N_13853,N_13026);
xnor U17815 (N_17815,N_14908,N_14224);
xor U17816 (N_17816,N_13340,N_14842);
or U17817 (N_17817,N_14541,N_15134);
xor U17818 (N_17818,N_14081,N_14543);
or U17819 (N_17819,N_14011,N_15635);
nand U17820 (N_17820,N_12600,N_13575);
or U17821 (N_17821,N_15481,N_13546);
nand U17822 (N_17822,N_15764,N_14859);
and U17823 (N_17823,N_13118,N_13438);
and U17824 (N_17824,N_14220,N_14713);
and U17825 (N_17825,N_13122,N_13645);
nand U17826 (N_17826,N_12058,N_13335);
nor U17827 (N_17827,N_12689,N_14971);
or U17828 (N_17828,N_15828,N_14104);
or U17829 (N_17829,N_12117,N_14814);
nand U17830 (N_17830,N_12016,N_13947);
nand U17831 (N_17831,N_14783,N_14979);
nor U17832 (N_17832,N_15323,N_15692);
nand U17833 (N_17833,N_15187,N_13785);
or U17834 (N_17834,N_12451,N_14711);
xnor U17835 (N_17835,N_15072,N_13866);
nor U17836 (N_17836,N_14730,N_15522);
nor U17837 (N_17837,N_12460,N_12840);
and U17838 (N_17838,N_12267,N_12202);
nand U17839 (N_17839,N_13683,N_14314);
or U17840 (N_17840,N_13651,N_14268);
and U17841 (N_17841,N_12990,N_13288);
or U17842 (N_17842,N_13620,N_13617);
nand U17843 (N_17843,N_12896,N_12543);
and U17844 (N_17844,N_14221,N_13237);
or U17845 (N_17845,N_14165,N_15221);
or U17846 (N_17846,N_12444,N_13759);
and U17847 (N_17847,N_13207,N_12034);
xor U17848 (N_17848,N_15064,N_13443);
or U17849 (N_17849,N_15926,N_14050);
xnor U17850 (N_17850,N_12153,N_14159);
or U17851 (N_17851,N_14569,N_14373);
and U17852 (N_17852,N_14816,N_12248);
or U17853 (N_17853,N_15091,N_14196);
xnor U17854 (N_17854,N_14508,N_12441);
nor U17855 (N_17855,N_14561,N_15475);
nor U17856 (N_17856,N_14791,N_13174);
xor U17857 (N_17857,N_14727,N_15399);
nand U17858 (N_17858,N_12612,N_15619);
or U17859 (N_17859,N_12780,N_12590);
xnor U17860 (N_17860,N_12389,N_12894);
nor U17861 (N_17861,N_13084,N_14015);
xnor U17862 (N_17862,N_15598,N_13152);
and U17863 (N_17863,N_15956,N_14528);
nand U17864 (N_17864,N_12730,N_14256);
or U17865 (N_17865,N_12549,N_15318);
nor U17866 (N_17866,N_13296,N_15317);
nor U17867 (N_17867,N_14784,N_13364);
or U17868 (N_17868,N_15473,N_13729);
nor U17869 (N_17869,N_13184,N_13125);
and U17870 (N_17870,N_12629,N_15455);
nand U17871 (N_17871,N_15917,N_15401);
nand U17872 (N_17872,N_15269,N_15372);
nor U17873 (N_17873,N_12405,N_15191);
xnor U17874 (N_17874,N_13680,N_15575);
nor U17875 (N_17875,N_15822,N_13181);
and U17876 (N_17876,N_12987,N_13959);
nor U17877 (N_17877,N_13850,N_12020);
and U17878 (N_17878,N_13367,N_12794);
nand U17879 (N_17879,N_14643,N_13632);
nand U17880 (N_17880,N_12434,N_13023);
nor U17881 (N_17881,N_15089,N_13261);
xor U17882 (N_17882,N_12137,N_12319);
xnor U17883 (N_17883,N_15541,N_14497);
nor U17884 (N_17884,N_15325,N_12592);
xnor U17885 (N_17885,N_15025,N_14514);
or U17886 (N_17886,N_12129,N_15862);
xnor U17887 (N_17887,N_14029,N_14632);
nor U17888 (N_17888,N_13137,N_13499);
or U17889 (N_17889,N_12920,N_15344);
nand U17890 (N_17890,N_13618,N_12958);
xor U17891 (N_17891,N_13622,N_14028);
or U17892 (N_17892,N_12360,N_12103);
or U17893 (N_17893,N_12161,N_13218);
or U17894 (N_17894,N_12727,N_14738);
and U17895 (N_17895,N_14988,N_15211);
or U17896 (N_17896,N_13246,N_12394);
and U17897 (N_17897,N_15077,N_12478);
nor U17898 (N_17898,N_15706,N_15185);
and U17899 (N_17899,N_15736,N_14532);
and U17900 (N_17900,N_15626,N_13477);
nor U17901 (N_17901,N_13640,N_12186);
and U17902 (N_17902,N_14878,N_14079);
nor U17903 (N_17903,N_13469,N_12127);
nand U17904 (N_17904,N_14276,N_14316);
nor U17905 (N_17905,N_15443,N_12884);
nand U17906 (N_17906,N_12042,N_14160);
or U17907 (N_17907,N_13740,N_15996);
or U17908 (N_17908,N_14189,N_15467);
xnor U17909 (N_17909,N_15836,N_12904);
xnor U17910 (N_17910,N_12314,N_12297);
nand U17911 (N_17911,N_12022,N_14629);
xnor U17912 (N_17912,N_12665,N_12531);
nor U17913 (N_17913,N_12438,N_12519);
xor U17914 (N_17914,N_14506,N_13922);
nand U17915 (N_17915,N_12176,N_14300);
xnor U17916 (N_17916,N_13681,N_12393);
nand U17917 (N_17917,N_15677,N_14817);
nand U17918 (N_17918,N_15257,N_15744);
xnor U17919 (N_17919,N_12173,N_12372);
and U17920 (N_17920,N_15968,N_12759);
nand U17921 (N_17921,N_15258,N_12099);
nand U17922 (N_17922,N_15605,N_12646);
nor U17923 (N_17923,N_15310,N_15196);
or U17924 (N_17924,N_12596,N_15315);
xor U17925 (N_17925,N_13089,N_13147);
nor U17926 (N_17926,N_12545,N_12272);
xnor U17927 (N_17927,N_14793,N_13820);
and U17928 (N_17928,N_15629,N_14026);
nand U17929 (N_17929,N_13716,N_14811);
nor U17930 (N_17930,N_14296,N_13872);
or U17931 (N_17931,N_15644,N_14182);
nand U17932 (N_17932,N_14990,N_12398);
nor U17933 (N_17933,N_13197,N_12397);
nor U17934 (N_17934,N_15565,N_13689);
xnor U17935 (N_17935,N_14208,N_15472);
or U17936 (N_17936,N_13696,N_12566);
and U17937 (N_17937,N_15595,N_13305);
nand U17938 (N_17938,N_14474,N_14376);
xor U17939 (N_17939,N_12861,N_13509);
nor U17940 (N_17940,N_14669,N_14626);
or U17941 (N_17941,N_14098,N_14092);
nor U17942 (N_17942,N_13223,N_15129);
and U17943 (N_17943,N_13752,N_14725);
nand U17944 (N_17944,N_14100,N_12645);
nor U17945 (N_17945,N_14774,N_12682);
xor U17946 (N_17946,N_15726,N_12335);
nor U17947 (N_17947,N_12429,N_13114);
nand U17948 (N_17948,N_14900,N_14128);
nand U17949 (N_17949,N_14386,N_14724);
xor U17950 (N_17950,N_14033,N_15348);
and U17951 (N_17951,N_13868,N_12454);
and U17952 (N_17952,N_13851,N_12452);
nand U17953 (N_17953,N_15680,N_12192);
nand U17954 (N_17954,N_13331,N_14750);
nand U17955 (N_17955,N_12812,N_13269);
or U17956 (N_17956,N_12614,N_12570);
nand U17957 (N_17957,N_13416,N_15693);
xnor U17958 (N_17958,N_15489,N_13182);
nand U17959 (N_17959,N_15174,N_15847);
nor U17960 (N_17960,N_13697,N_13521);
or U17961 (N_17961,N_14531,N_12553);
and U17962 (N_17962,N_15867,N_15738);
xor U17963 (N_17963,N_12913,N_13827);
xnor U17964 (N_17964,N_14008,N_12090);
xor U17965 (N_17965,N_12865,N_13998);
nor U17966 (N_17966,N_14825,N_13365);
nand U17967 (N_17967,N_15665,N_14537);
nand U17968 (N_17968,N_14341,N_14434);
nor U17969 (N_17969,N_15920,N_14141);
or U17970 (N_17970,N_13353,N_13776);
nand U17971 (N_17971,N_12615,N_12024);
and U17972 (N_17972,N_15778,N_13491);
xnor U17973 (N_17973,N_13737,N_13045);
or U17974 (N_17974,N_14073,N_14560);
xnor U17975 (N_17975,N_14147,N_13671);
nand U17976 (N_17976,N_14895,N_15388);
nor U17977 (N_17977,N_13212,N_14849);
nand U17978 (N_17978,N_12731,N_13055);
nand U17979 (N_17979,N_13930,N_12851);
and U17980 (N_17980,N_12578,N_12735);
nor U17981 (N_17981,N_13273,N_14799);
nand U17982 (N_17982,N_15528,N_14721);
nor U17983 (N_17983,N_14635,N_14413);
nand U17984 (N_17984,N_13001,N_15499);
nand U17985 (N_17985,N_15112,N_12282);
xnor U17986 (N_17986,N_15432,N_13838);
nor U17987 (N_17987,N_14764,N_12923);
or U17988 (N_17988,N_13398,N_14446);
or U17989 (N_17989,N_13950,N_12418);
nor U17990 (N_17990,N_13735,N_13849);
xor U17991 (N_17991,N_13442,N_13852);
nand U17992 (N_17992,N_13788,N_12422);
nand U17993 (N_17993,N_13461,N_13213);
nor U17994 (N_17994,N_14867,N_14484);
and U17995 (N_17995,N_12242,N_13176);
xor U17996 (N_17996,N_14729,N_15537);
or U17997 (N_17997,N_14360,N_14364);
xor U17998 (N_17998,N_13540,N_12484);
and U17999 (N_17999,N_15365,N_12239);
nand U18000 (N_18000,N_15145,N_13725);
xor U18001 (N_18001,N_15749,N_13246);
or U18002 (N_18002,N_15044,N_13967);
and U18003 (N_18003,N_15281,N_14651);
nor U18004 (N_18004,N_12371,N_12243);
and U18005 (N_18005,N_12210,N_15741);
xnor U18006 (N_18006,N_15576,N_12629);
nor U18007 (N_18007,N_15419,N_13072);
nor U18008 (N_18008,N_12707,N_15187);
and U18009 (N_18009,N_15971,N_12201);
nor U18010 (N_18010,N_15473,N_12910);
xor U18011 (N_18011,N_12810,N_15972);
and U18012 (N_18012,N_12130,N_12219);
nand U18013 (N_18013,N_12127,N_12914);
xor U18014 (N_18014,N_13477,N_15536);
nand U18015 (N_18015,N_15562,N_13014);
or U18016 (N_18016,N_15414,N_12216);
xnor U18017 (N_18017,N_12392,N_13792);
nand U18018 (N_18018,N_15110,N_12513);
xnor U18019 (N_18019,N_15743,N_15837);
xnor U18020 (N_18020,N_13932,N_15117);
nand U18021 (N_18021,N_15804,N_14724);
and U18022 (N_18022,N_13035,N_13546);
xor U18023 (N_18023,N_15388,N_15425);
and U18024 (N_18024,N_14034,N_15776);
xnor U18025 (N_18025,N_13183,N_15300);
nand U18026 (N_18026,N_15712,N_15546);
xnor U18027 (N_18027,N_12126,N_14184);
nand U18028 (N_18028,N_14856,N_13423);
and U18029 (N_18029,N_13372,N_12367);
xnor U18030 (N_18030,N_12854,N_12128);
nand U18031 (N_18031,N_14722,N_14918);
xnor U18032 (N_18032,N_14594,N_13936);
nand U18033 (N_18033,N_14518,N_12425);
nand U18034 (N_18034,N_15993,N_13799);
nor U18035 (N_18035,N_12109,N_13209);
and U18036 (N_18036,N_15597,N_12581);
and U18037 (N_18037,N_13178,N_13050);
nand U18038 (N_18038,N_12484,N_15989);
nor U18039 (N_18039,N_13553,N_15267);
nor U18040 (N_18040,N_15244,N_15238);
nor U18041 (N_18041,N_12316,N_12442);
and U18042 (N_18042,N_12625,N_13120);
xnor U18043 (N_18043,N_15251,N_12764);
nor U18044 (N_18044,N_14341,N_13865);
and U18045 (N_18045,N_14354,N_15953);
xor U18046 (N_18046,N_14203,N_15981);
or U18047 (N_18047,N_13019,N_14811);
nand U18048 (N_18048,N_12998,N_14135);
xor U18049 (N_18049,N_14577,N_13017);
nor U18050 (N_18050,N_14012,N_12719);
nor U18051 (N_18051,N_14955,N_14517);
nand U18052 (N_18052,N_12135,N_13296);
xor U18053 (N_18053,N_14806,N_14196);
and U18054 (N_18054,N_12282,N_12237);
nand U18055 (N_18055,N_14100,N_13577);
or U18056 (N_18056,N_12755,N_12911);
nand U18057 (N_18057,N_15145,N_12215);
nor U18058 (N_18058,N_12645,N_13148);
nand U18059 (N_18059,N_12727,N_15685);
nand U18060 (N_18060,N_15536,N_15072);
or U18061 (N_18061,N_15460,N_14499);
and U18062 (N_18062,N_14568,N_12394);
and U18063 (N_18063,N_12235,N_14025);
xor U18064 (N_18064,N_12875,N_14693);
and U18065 (N_18065,N_12972,N_14754);
and U18066 (N_18066,N_13054,N_12739);
or U18067 (N_18067,N_13032,N_12490);
or U18068 (N_18068,N_13729,N_14359);
nand U18069 (N_18069,N_13287,N_14481);
xor U18070 (N_18070,N_14670,N_15100);
xor U18071 (N_18071,N_15693,N_14237);
or U18072 (N_18072,N_13979,N_15898);
or U18073 (N_18073,N_13214,N_12058);
or U18074 (N_18074,N_15979,N_12998);
or U18075 (N_18075,N_13339,N_14909);
nor U18076 (N_18076,N_14499,N_12596);
or U18077 (N_18077,N_12441,N_13100);
nor U18078 (N_18078,N_15034,N_14528);
or U18079 (N_18079,N_13376,N_13089);
xor U18080 (N_18080,N_15849,N_13093);
xnor U18081 (N_18081,N_13360,N_15249);
or U18082 (N_18082,N_12540,N_13403);
xnor U18083 (N_18083,N_13232,N_12934);
xor U18084 (N_18084,N_12040,N_14490);
and U18085 (N_18085,N_14718,N_15483);
or U18086 (N_18086,N_12653,N_14380);
and U18087 (N_18087,N_13356,N_12841);
nor U18088 (N_18088,N_14396,N_14232);
nor U18089 (N_18089,N_12195,N_15751);
nor U18090 (N_18090,N_14445,N_13810);
xor U18091 (N_18091,N_13979,N_12866);
and U18092 (N_18092,N_12969,N_14224);
nor U18093 (N_18093,N_13361,N_15022);
xnor U18094 (N_18094,N_12459,N_15425);
and U18095 (N_18095,N_12943,N_14841);
or U18096 (N_18096,N_15201,N_13679);
and U18097 (N_18097,N_12847,N_14633);
nor U18098 (N_18098,N_14902,N_14033);
xor U18099 (N_18099,N_15787,N_15888);
xnor U18100 (N_18100,N_12050,N_14665);
and U18101 (N_18101,N_13439,N_15463);
xor U18102 (N_18102,N_15924,N_14003);
or U18103 (N_18103,N_13379,N_12870);
nand U18104 (N_18104,N_13159,N_14044);
xnor U18105 (N_18105,N_13061,N_13428);
nor U18106 (N_18106,N_12878,N_12536);
nor U18107 (N_18107,N_12932,N_14578);
nor U18108 (N_18108,N_13394,N_14215);
nor U18109 (N_18109,N_15840,N_13501);
xnor U18110 (N_18110,N_15552,N_14233);
or U18111 (N_18111,N_12281,N_13471);
xnor U18112 (N_18112,N_12018,N_14102);
nand U18113 (N_18113,N_15439,N_13606);
nor U18114 (N_18114,N_15734,N_15053);
xor U18115 (N_18115,N_14345,N_14663);
xor U18116 (N_18116,N_12907,N_12374);
and U18117 (N_18117,N_13469,N_14578);
or U18118 (N_18118,N_12214,N_13142);
nand U18119 (N_18119,N_13529,N_15885);
or U18120 (N_18120,N_13261,N_14214);
nor U18121 (N_18121,N_12176,N_12842);
xor U18122 (N_18122,N_13771,N_12410);
xnor U18123 (N_18123,N_12208,N_13962);
or U18124 (N_18124,N_15490,N_15463);
nor U18125 (N_18125,N_14911,N_12450);
nor U18126 (N_18126,N_15675,N_14836);
and U18127 (N_18127,N_15308,N_15098);
and U18128 (N_18128,N_14853,N_12138);
and U18129 (N_18129,N_13420,N_13162);
or U18130 (N_18130,N_13282,N_12745);
nor U18131 (N_18131,N_15994,N_14332);
nor U18132 (N_18132,N_14605,N_14700);
nand U18133 (N_18133,N_12021,N_14254);
or U18134 (N_18134,N_15122,N_15914);
nor U18135 (N_18135,N_13578,N_15328);
nor U18136 (N_18136,N_13727,N_14956);
nand U18137 (N_18137,N_15649,N_12709);
nand U18138 (N_18138,N_13285,N_15271);
nor U18139 (N_18139,N_13778,N_14486);
and U18140 (N_18140,N_14575,N_13941);
xor U18141 (N_18141,N_15690,N_12343);
nor U18142 (N_18142,N_15789,N_12378);
xor U18143 (N_18143,N_12830,N_14337);
xor U18144 (N_18144,N_15671,N_15113);
nand U18145 (N_18145,N_14986,N_12691);
xor U18146 (N_18146,N_13029,N_12079);
and U18147 (N_18147,N_14134,N_13373);
and U18148 (N_18148,N_12529,N_12992);
and U18149 (N_18149,N_12772,N_12018);
and U18150 (N_18150,N_15245,N_12114);
or U18151 (N_18151,N_13130,N_12650);
or U18152 (N_18152,N_15835,N_13928);
and U18153 (N_18153,N_13085,N_14298);
nor U18154 (N_18154,N_14475,N_15919);
or U18155 (N_18155,N_13762,N_13741);
or U18156 (N_18156,N_13910,N_13434);
nand U18157 (N_18157,N_14710,N_14821);
nor U18158 (N_18158,N_15576,N_15277);
xnor U18159 (N_18159,N_13838,N_14580);
nor U18160 (N_18160,N_12158,N_13339);
nor U18161 (N_18161,N_14787,N_13769);
and U18162 (N_18162,N_15122,N_14438);
xor U18163 (N_18163,N_13545,N_14421);
or U18164 (N_18164,N_13859,N_13512);
nor U18165 (N_18165,N_15652,N_15082);
nor U18166 (N_18166,N_12959,N_12361);
or U18167 (N_18167,N_13026,N_12636);
nor U18168 (N_18168,N_14484,N_12502);
xor U18169 (N_18169,N_14899,N_13890);
and U18170 (N_18170,N_12298,N_13694);
or U18171 (N_18171,N_15914,N_12834);
xor U18172 (N_18172,N_14611,N_15816);
nor U18173 (N_18173,N_13059,N_14210);
and U18174 (N_18174,N_14473,N_14475);
nand U18175 (N_18175,N_14719,N_12491);
and U18176 (N_18176,N_15592,N_12728);
xnor U18177 (N_18177,N_13727,N_12104);
nor U18178 (N_18178,N_15215,N_15314);
xor U18179 (N_18179,N_15093,N_12408);
xnor U18180 (N_18180,N_13021,N_15270);
or U18181 (N_18181,N_15707,N_15678);
and U18182 (N_18182,N_14727,N_13901);
and U18183 (N_18183,N_14289,N_12771);
xnor U18184 (N_18184,N_13419,N_13845);
and U18185 (N_18185,N_15375,N_14175);
nor U18186 (N_18186,N_13454,N_15503);
and U18187 (N_18187,N_13121,N_14691);
and U18188 (N_18188,N_14205,N_13220);
nand U18189 (N_18189,N_12821,N_15284);
and U18190 (N_18190,N_14498,N_13488);
nor U18191 (N_18191,N_13601,N_14630);
nor U18192 (N_18192,N_13839,N_12498);
and U18193 (N_18193,N_13113,N_12813);
and U18194 (N_18194,N_12199,N_15222);
and U18195 (N_18195,N_14109,N_12278);
nand U18196 (N_18196,N_15055,N_12581);
xnor U18197 (N_18197,N_15834,N_15378);
or U18198 (N_18198,N_12501,N_12288);
xor U18199 (N_18199,N_13271,N_14088);
and U18200 (N_18200,N_14923,N_12538);
xor U18201 (N_18201,N_13667,N_14597);
and U18202 (N_18202,N_12404,N_13957);
and U18203 (N_18203,N_14122,N_12228);
or U18204 (N_18204,N_12767,N_13099);
nand U18205 (N_18205,N_15110,N_13490);
xnor U18206 (N_18206,N_13968,N_12792);
or U18207 (N_18207,N_12061,N_12463);
nand U18208 (N_18208,N_12850,N_12483);
xnor U18209 (N_18209,N_14100,N_13386);
and U18210 (N_18210,N_13778,N_13618);
nor U18211 (N_18211,N_15491,N_12524);
xnor U18212 (N_18212,N_13134,N_15542);
and U18213 (N_18213,N_15736,N_12192);
xnor U18214 (N_18214,N_14305,N_12252);
and U18215 (N_18215,N_14504,N_13139);
or U18216 (N_18216,N_15895,N_13252);
and U18217 (N_18217,N_14757,N_13622);
nand U18218 (N_18218,N_14944,N_12445);
and U18219 (N_18219,N_14434,N_14898);
xor U18220 (N_18220,N_14394,N_14066);
xor U18221 (N_18221,N_14106,N_13377);
nor U18222 (N_18222,N_12966,N_14775);
nor U18223 (N_18223,N_15798,N_14936);
nand U18224 (N_18224,N_14179,N_14751);
xnor U18225 (N_18225,N_14288,N_15814);
or U18226 (N_18226,N_14830,N_13671);
nand U18227 (N_18227,N_15581,N_12086);
nand U18228 (N_18228,N_12803,N_13930);
and U18229 (N_18229,N_15654,N_14665);
nand U18230 (N_18230,N_14914,N_13034);
or U18231 (N_18231,N_12809,N_13435);
xor U18232 (N_18232,N_12974,N_12836);
and U18233 (N_18233,N_14428,N_14489);
or U18234 (N_18234,N_14174,N_12160);
and U18235 (N_18235,N_13081,N_15214);
and U18236 (N_18236,N_12139,N_13317);
xor U18237 (N_18237,N_12246,N_15789);
nor U18238 (N_18238,N_12376,N_15378);
nor U18239 (N_18239,N_13635,N_13691);
and U18240 (N_18240,N_13275,N_15959);
or U18241 (N_18241,N_13270,N_13873);
and U18242 (N_18242,N_13232,N_14746);
nor U18243 (N_18243,N_13775,N_14948);
or U18244 (N_18244,N_13829,N_14529);
or U18245 (N_18245,N_13637,N_12614);
nand U18246 (N_18246,N_15313,N_15869);
nor U18247 (N_18247,N_12689,N_15986);
and U18248 (N_18248,N_15011,N_14056);
nor U18249 (N_18249,N_15130,N_15822);
nand U18250 (N_18250,N_14266,N_15338);
or U18251 (N_18251,N_15418,N_13604);
or U18252 (N_18252,N_14933,N_15227);
xnor U18253 (N_18253,N_15607,N_12510);
or U18254 (N_18254,N_15110,N_15927);
or U18255 (N_18255,N_13670,N_12491);
and U18256 (N_18256,N_13042,N_14229);
or U18257 (N_18257,N_12109,N_12668);
or U18258 (N_18258,N_12979,N_14158);
and U18259 (N_18259,N_14803,N_14705);
nor U18260 (N_18260,N_12227,N_14798);
nand U18261 (N_18261,N_15449,N_12332);
nor U18262 (N_18262,N_14493,N_12031);
or U18263 (N_18263,N_12828,N_15837);
xor U18264 (N_18264,N_12076,N_13764);
xnor U18265 (N_18265,N_12559,N_15240);
xnor U18266 (N_18266,N_15907,N_12519);
xor U18267 (N_18267,N_13031,N_15905);
xor U18268 (N_18268,N_12663,N_12755);
nor U18269 (N_18269,N_15517,N_12083);
xor U18270 (N_18270,N_13641,N_13338);
xnor U18271 (N_18271,N_12799,N_14797);
xnor U18272 (N_18272,N_15168,N_14429);
and U18273 (N_18273,N_15583,N_14409);
or U18274 (N_18274,N_12898,N_13760);
nand U18275 (N_18275,N_12915,N_15969);
xor U18276 (N_18276,N_15320,N_15732);
xnor U18277 (N_18277,N_13506,N_15034);
nor U18278 (N_18278,N_15271,N_14963);
xor U18279 (N_18279,N_12067,N_13790);
nand U18280 (N_18280,N_15508,N_14506);
or U18281 (N_18281,N_13018,N_12982);
xor U18282 (N_18282,N_13741,N_14383);
nor U18283 (N_18283,N_13499,N_15710);
and U18284 (N_18284,N_13624,N_12695);
nand U18285 (N_18285,N_14107,N_12763);
or U18286 (N_18286,N_15819,N_14828);
and U18287 (N_18287,N_13081,N_14833);
nor U18288 (N_18288,N_12818,N_14880);
nand U18289 (N_18289,N_12024,N_15285);
nor U18290 (N_18290,N_13197,N_15931);
nand U18291 (N_18291,N_15237,N_15950);
or U18292 (N_18292,N_14748,N_12865);
nand U18293 (N_18293,N_15336,N_15909);
nand U18294 (N_18294,N_14052,N_13993);
nor U18295 (N_18295,N_12851,N_15584);
or U18296 (N_18296,N_13245,N_15079);
nand U18297 (N_18297,N_15451,N_13135);
and U18298 (N_18298,N_15726,N_14188);
xor U18299 (N_18299,N_12711,N_12960);
and U18300 (N_18300,N_13644,N_13959);
or U18301 (N_18301,N_14770,N_15700);
xor U18302 (N_18302,N_14014,N_13906);
nand U18303 (N_18303,N_12111,N_13359);
or U18304 (N_18304,N_15526,N_13758);
nand U18305 (N_18305,N_13772,N_15283);
and U18306 (N_18306,N_12714,N_15229);
and U18307 (N_18307,N_15416,N_14049);
nor U18308 (N_18308,N_15678,N_14268);
nor U18309 (N_18309,N_13558,N_12275);
or U18310 (N_18310,N_13755,N_14040);
nand U18311 (N_18311,N_12735,N_14711);
nand U18312 (N_18312,N_15378,N_14591);
or U18313 (N_18313,N_15721,N_15297);
or U18314 (N_18314,N_15578,N_14626);
and U18315 (N_18315,N_14044,N_14116);
nor U18316 (N_18316,N_14323,N_12114);
xor U18317 (N_18317,N_12484,N_12475);
xor U18318 (N_18318,N_15623,N_12320);
xnor U18319 (N_18319,N_12109,N_14622);
or U18320 (N_18320,N_13162,N_14664);
nand U18321 (N_18321,N_12495,N_15727);
nand U18322 (N_18322,N_13817,N_13039);
and U18323 (N_18323,N_12537,N_13827);
nor U18324 (N_18324,N_13569,N_15283);
and U18325 (N_18325,N_15102,N_15136);
and U18326 (N_18326,N_12586,N_15798);
or U18327 (N_18327,N_12107,N_13657);
and U18328 (N_18328,N_13913,N_15916);
nor U18329 (N_18329,N_14734,N_13860);
nor U18330 (N_18330,N_12139,N_14359);
nand U18331 (N_18331,N_15151,N_12393);
nor U18332 (N_18332,N_12698,N_13985);
nor U18333 (N_18333,N_15544,N_13276);
nand U18334 (N_18334,N_14707,N_15948);
xor U18335 (N_18335,N_12631,N_12167);
nand U18336 (N_18336,N_14534,N_12015);
nor U18337 (N_18337,N_14018,N_14474);
or U18338 (N_18338,N_15303,N_14803);
xor U18339 (N_18339,N_15740,N_13763);
nand U18340 (N_18340,N_15663,N_15125);
or U18341 (N_18341,N_12345,N_13581);
or U18342 (N_18342,N_12565,N_15148);
and U18343 (N_18343,N_14179,N_15685);
and U18344 (N_18344,N_15123,N_14879);
or U18345 (N_18345,N_13531,N_14990);
and U18346 (N_18346,N_13164,N_12007);
xnor U18347 (N_18347,N_15564,N_15129);
and U18348 (N_18348,N_14359,N_13207);
xor U18349 (N_18349,N_15395,N_13045);
xnor U18350 (N_18350,N_13472,N_15585);
or U18351 (N_18351,N_12014,N_13529);
nand U18352 (N_18352,N_14245,N_14942);
nand U18353 (N_18353,N_13524,N_15970);
and U18354 (N_18354,N_13264,N_12497);
nor U18355 (N_18355,N_13290,N_14762);
or U18356 (N_18356,N_13790,N_14592);
nand U18357 (N_18357,N_12013,N_13098);
nand U18358 (N_18358,N_12973,N_12672);
and U18359 (N_18359,N_14808,N_15071);
nand U18360 (N_18360,N_15224,N_13800);
and U18361 (N_18361,N_12771,N_12253);
or U18362 (N_18362,N_14502,N_13763);
nor U18363 (N_18363,N_13500,N_13351);
and U18364 (N_18364,N_14978,N_14948);
nand U18365 (N_18365,N_15024,N_13543);
nor U18366 (N_18366,N_12723,N_12013);
nor U18367 (N_18367,N_14963,N_15014);
nor U18368 (N_18368,N_12409,N_15276);
or U18369 (N_18369,N_13345,N_12603);
nor U18370 (N_18370,N_15796,N_12414);
xnor U18371 (N_18371,N_14903,N_12061);
nor U18372 (N_18372,N_12294,N_14977);
or U18373 (N_18373,N_13893,N_15695);
and U18374 (N_18374,N_14955,N_14136);
and U18375 (N_18375,N_13921,N_12339);
nor U18376 (N_18376,N_12658,N_12299);
or U18377 (N_18377,N_15096,N_14423);
nand U18378 (N_18378,N_13232,N_14446);
xnor U18379 (N_18379,N_14400,N_13054);
nand U18380 (N_18380,N_15418,N_14521);
and U18381 (N_18381,N_14373,N_13109);
nor U18382 (N_18382,N_14501,N_12504);
and U18383 (N_18383,N_15864,N_15515);
xnor U18384 (N_18384,N_14027,N_13402);
or U18385 (N_18385,N_14785,N_13871);
xor U18386 (N_18386,N_13768,N_13001);
xnor U18387 (N_18387,N_14185,N_13818);
nand U18388 (N_18388,N_12782,N_14152);
xnor U18389 (N_18389,N_12223,N_14548);
or U18390 (N_18390,N_15818,N_12886);
nor U18391 (N_18391,N_15798,N_12316);
xor U18392 (N_18392,N_12163,N_13505);
nand U18393 (N_18393,N_12914,N_12121);
xor U18394 (N_18394,N_15470,N_15085);
nor U18395 (N_18395,N_13471,N_13654);
or U18396 (N_18396,N_14448,N_14554);
nor U18397 (N_18397,N_15508,N_12070);
nand U18398 (N_18398,N_14871,N_12877);
nor U18399 (N_18399,N_13854,N_12929);
nand U18400 (N_18400,N_13952,N_13176);
nand U18401 (N_18401,N_13524,N_13636);
and U18402 (N_18402,N_15556,N_13857);
nand U18403 (N_18403,N_13945,N_14980);
or U18404 (N_18404,N_14566,N_15495);
nor U18405 (N_18405,N_13820,N_14057);
nor U18406 (N_18406,N_12154,N_14645);
nand U18407 (N_18407,N_14169,N_15022);
and U18408 (N_18408,N_12508,N_15768);
and U18409 (N_18409,N_14684,N_13150);
or U18410 (N_18410,N_15808,N_12097);
xnor U18411 (N_18411,N_14864,N_15558);
nand U18412 (N_18412,N_12215,N_14643);
xor U18413 (N_18413,N_12342,N_13415);
or U18414 (N_18414,N_14467,N_15626);
or U18415 (N_18415,N_13191,N_12439);
nor U18416 (N_18416,N_13683,N_13871);
nor U18417 (N_18417,N_13549,N_13040);
xnor U18418 (N_18418,N_14333,N_14785);
nor U18419 (N_18419,N_15024,N_14819);
xor U18420 (N_18420,N_12393,N_13462);
and U18421 (N_18421,N_15961,N_12079);
or U18422 (N_18422,N_14891,N_14000);
nor U18423 (N_18423,N_15975,N_15970);
nand U18424 (N_18424,N_15337,N_14548);
nor U18425 (N_18425,N_15341,N_12686);
nand U18426 (N_18426,N_15209,N_14944);
or U18427 (N_18427,N_12278,N_14402);
nor U18428 (N_18428,N_13995,N_14784);
and U18429 (N_18429,N_12437,N_12949);
nand U18430 (N_18430,N_14325,N_12618);
and U18431 (N_18431,N_13082,N_13415);
nor U18432 (N_18432,N_12699,N_15320);
or U18433 (N_18433,N_14199,N_14179);
xor U18434 (N_18434,N_13359,N_15370);
nand U18435 (N_18435,N_13095,N_14263);
and U18436 (N_18436,N_15607,N_14207);
xor U18437 (N_18437,N_12197,N_12945);
xnor U18438 (N_18438,N_14258,N_15932);
xnor U18439 (N_18439,N_12999,N_14396);
or U18440 (N_18440,N_14046,N_12352);
nor U18441 (N_18441,N_14710,N_14415);
nor U18442 (N_18442,N_15189,N_13094);
nand U18443 (N_18443,N_15413,N_15147);
xor U18444 (N_18444,N_14378,N_12574);
nand U18445 (N_18445,N_12709,N_13315);
and U18446 (N_18446,N_15319,N_13441);
xor U18447 (N_18447,N_12675,N_15551);
xnor U18448 (N_18448,N_14923,N_13025);
nand U18449 (N_18449,N_15131,N_14558);
or U18450 (N_18450,N_13216,N_15232);
or U18451 (N_18451,N_14298,N_14856);
and U18452 (N_18452,N_13168,N_13917);
xnor U18453 (N_18453,N_13523,N_13740);
and U18454 (N_18454,N_12568,N_12054);
or U18455 (N_18455,N_14751,N_14043);
and U18456 (N_18456,N_15470,N_14573);
xor U18457 (N_18457,N_15379,N_13460);
and U18458 (N_18458,N_13465,N_14759);
xnor U18459 (N_18459,N_14201,N_13992);
nand U18460 (N_18460,N_14431,N_13213);
and U18461 (N_18461,N_14725,N_15712);
nand U18462 (N_18462,N_12910,N_12100);
nand U18463 (N_18463,N_13733,N_15744);
or U18464 (N_18464,N_14590,N_14615);
xnor U18465 (N_18465,N_12698,N_14659);
and U18466 (N_18466,N_12434,N_14260);
or U18467 (N_18467,N_12931,N_12836);
nor U18468 (N_18468,N_13464,N_13466);
nand U18469 (N_18469,N_15888,N_13640);
and U18470 (N_18470,N_13467,N_13140);
xnor U18471 (N_18471,N_14344,N_13276);
nand U18472 (N_18472,N_12598,N_15067);
nor U18473 (N_18473,N_14067,N_13725);
or U18474 (N_18474,N_14055,N_12055);
nand U18475 (N_18475,N_13131,N_13175);
xnor U18476 (N_18476,N_14888,N_14736);
xor U18477 (N_18477,N_15712,N_13834);
and U18478 (N_18478,N_12102,N_12129);
xnor U18479 (N_18479,N_13786,N_13338);
nand U18480 (N_18480,N_14303,N_12074);
and U18481 (N_18481,N_14971,N_12467);
xor U18482 (N_18482,N_12725,N_15917);
and U18483 (N_18483,N_14879,N_12419);
xnor U18484 (N_18484,N_14456,N_15204);
nor U18485 (N_18485,N_13112,N_12052);
or U18486 (N_18486,N_12798,N_15689);
or U18487 (N_18487,N_14472,N_15483);
nor U18488 (N_18488,N_13534,N_12463);
nor U18489 (N_18489,N_14486,N_15998);
nand U18490 (N_18490,N_13316,N_14350);
and U18491 (N_18491,N_13547,N_13364);
nor U18492 (N_18492,N_12064,N_14678);
or U18493 (N_18493,N_13358,N_13475);
nand U18494 (N_18494,N_12827,N_14493);
nand U18495 (N_18495,N_12635,N_14383);
or U18496 (N_18496,N_14102,N_13298);
and U18497 (N_18497,N_12925,N_13678);
and U18498 (N_18498,N_12943,N_13286);
nor U18499 (N_18499,N_15494,N_13226);
nor U18500 (N_18500,N_12106,N_15778);
xor U18501 (N_18501,N_15117,N_15345);
nor U18502 (N_18502,N_13634,N_14224);
and U18503 (N_18503,N_15897,N_12940);
or U18504 (N_18504,N_13735,N_14554);
nand U18505 (N_18505,N_14137,N_14974);
and U18506 (N_18506,N_14540,N_15168);
or U18507 (N_18507,N_13395,N_13882);
or U18508 (N_18508,N_14493,N_13391);
xnor U18509 (N_18509,N_15573,N_15287);
xnor U18510 (N_18510,N_13472,N_14725);
and U18511 (N_18511,N_14592,N_12612);
xor U18512 (N_18512,N_12572,N_12996);
xnor U18513 (N_18513,N_15635,N_14136);
nand U18514 (N_18514,N_13150,N_15527);
or U18515 (N_18515,N_14706,N_15322);
and U18516 (N_18516,N_12946,N_15256);
or U18517 (N_18517,N_12715,N_14143);
and U18518 (N_18518,N_14047,N_13102);
and U18519 (N_18519,N_15608,N_13830);
or U18520 (N_18520,N_15847,N_12010);
and U18521 (N_18521,N_13131,N_15928);
and U18522 (N_18522,N_15948,N_12556);
xor U18523 (N_18523,N_12995,N_14661);
xnor U18524 (N_18524,N_15849,N_13233);
and U18525 (N_18525,N_12202,N_12104);
nand U18526 (N_18526,N_14159,N_14893);
nand U18527 (N_18527,N_14027,N_14549);
nor U18528 (N_18528,N_15873,N_15855);
or U18529 (N_18529,N_12054,N_15500);
nor U18530 (N_18530,N_12712,N_13218);
or U18531 (N_18531,N_12999,N_14330);
and U18532 (N_18532,N_15080,N_12839);
nand U18533 (N_18533,N_15033,N_12017);
or U18534 (N_18534,N_12306,N_14068);
and U18535 (N_18535,N_14734,N_14244);
or U18536 (N_18536,N_12879,N_13995);
and U18537 (N_18537,N_14878,N_14101);
nand U18538 (N_18538,N_12600,N_12306);
nand U18539 (N_18539,N_13513,N_14117);
nand U18540 (N_18540,N_14678,N_15497);
xnor U18541 (N_18541,N_15018,N_15310);
or U18542 (N_18542,N_14552,N_13970);
xor U18543 (N_18543,N_12568,N_14185);
nor U18544 (N_18544,N_15969,N_13345);
or U18545 (N_18545,N_13673,N_12456);
xor U18546 (N_18546,N_14195,N_12675);
nor U18547 (N_18547,N_15968,N_12691);
nand U18548 (N_18548,N_15891,N_12418);
or U18549 (N_18549,N_12783,N_15803);
nand U18550 (N_18550,N_14847,N_15533);
nand U18551 (N_18551,N_14633,N_15431);
nor U18552 (N_18552,N_13420,N_12767);
nand U18553 (N_18553,N_13281,N_12532);
xnor U18554 (N_18554,N_13843,N_14033);
nor U18555 (N_18555,N_14972,N_12143);
and U18556 (N_18556,N_15177,N_13442);
nand U18557 (N_18557,N_15172,N_14830);
or U18558 (N_18558,N_14231,N_15940);
or U18559 (N_18559,N_14669,N_15229);
nor U18560 (N_18560,N_15220,N_12262);
and U18561 (N_18561,N_13184,N_15617);
and U18562 (N_18562,N_15810,N_15938);
xor U18563 (N_18563,N_14520,N_12554);
nand U18564 (N_18564,N_14321,N_12847);
and U18565 (N_18565,N_13408,N_13633);
and U18566 (N_18566,N_15046,N_13453);
and U18567 (N_18567,N_14445,N_12180);
and U18568 (N_18568,N_14703,N_14253);
nor U18569 (N_18569,N_12672,N_14885);
and U18570 (N_18570,N_12501,N_12970);
nor U18571 (N_18571,N_15124,N_12650);
and U18572 (N_18572,N_12935,N_13613);
or U18573 (N_18573,N_13996,N_13142);
and U18574 (N_18574,N_14061,N_12421);
nand U18575 (N_18575,N_15904,N_14530);
xnor U18576 (N_18576,N_15585,N_13626);
or U18577 (N_18577,N_14193,N_13748);
nand U18578 (N_18578,N_14821,N_15061);
or U18579 (N_18579,N_15476,N_14643);
xor U18580 (N_18580,N_15675,N_15763);
nand U18581 (N_18581,N_13684,N_12223);
nor U18582 (N_18582,N_14885,N_14170);
nor U18583 (N_18583,N_12345,N_14194);
and U18584 (N_18584,N_13901,N_15818);
nand U18585 (N_18585,N_12151,N_13482);
nor U18586 (N_18586,N_14279,N_12823);
nand U18587 (N_18587,N_15388,N_14091);
xnor U18588 (N_18588,N_12647,N_12992);
and U18589 (N_18589,N_15730,N_14846);
xor U18590 (N_18590,N_12202,N_12458);
nor U18591 (N_18591,N_12555,N_15201);
and U18592 (N_18592,N_15405,N_12645);
and U18593 (N_18593,N_14191,N_14173);
nor U18594 (N_18594,N_14743,N_12360);
xnor U18595 (N_18595,N_14720,N_14050);
xnor U18596 (N_18596,N_15147,N_15954);
and U18597 (N_18597,N_14984,N_13503);
xor U18598 (N_18598,N_14339,N_15113);
and U18599 (N_18599,N_13450,N_14666);
or U18600 (N_18600,N_13176,N_14450);
and U18601 (N_18601,N_14000,N_14146);
nor U18602 (N_18602,N_13903,N_13936);
nand U18603 (N_18603,N_14889,N_14692);
xnor U18604 (N_18604,N_14579,N_13346);
nand U18605 (N_18605,N_13984,N_15302);
nor U18606 (N_18606,N_14639,N_15970);
nor U18607 (N_18607,N_13743,N_13492);
and U18608 (N_18608,N_13758,N_12832);
or U18609 (N_18609,N_12950,N_12791);
xor U18610 (N_18610,N_14265,N_13248);
nor U18611 (N_18611,N_14886,N_12638);
and U18612 (N_18612,N_13392,N_14086);
or U18613 (N_18613,N_12512,N_12517);
nor U18614 (N_18614,N_13758,N_15000);
nor U18615 (N_18615,N_15205,N_12689);
nand U18616 (N_18616,N_15034,N_14921);
nor U18617 (N_18617,N_15006,N_15044);
and U18618 (N_18618,N_15670,N_14613);
and U18619 (N_18619,N_14010,N_13882);
nor U18620 (N_18620,N_13780,N_12009);
nor U18621 (N_18621,N_14567,N_12324);
nand U18622 (N_18622,N_14371,N_12420);
and U18623 (N_18623,N_15066,N_12148);
or U18624 (N_18624,N_13734,N_14776);
nand U18625 (N_18625,N_13725,N_15773);
or U18626 (N_18626,N_13638,N_14275);
nand U18627 (N_18627,N_13679,N_12060);
xnor U18628 (N_18628,N_12891,N_12516);
nor U18629 (N_18629,N_15911,N_15738);
and U18630 (N_18630,N_15073,N_15458);
nor U18631 (N_18631,N_15067,N_14343);
or U18632 (N_18632,N_14320,N_12152);
and U18633 (N_18633,N_15026,N_13939);
xor U18634 (N_18634,N_15368,N_12683);
and U18635 (N_18635,N_12611,N_15788);
nand U18636 (N_18636,N_12837,N_14353);
and U18637 (N_18637,N_14864,N_14993);
nor U18638 (N_18638,N_13498,N_12301);
and U18639 (N_18639,N_13847,N_15256);
nor U18640 (N_18640,N_15832,N_12906);
xor U18641 (N_18641,N_13810,N_14167);
nand U18642 (N_18642,N_15037,N_12014);
xor U18643 (N_18643,N_14922,N_14732);
nand U18644 (N_18644,N_13984,N_12479);
xnor U18645 (N_18645,N_14366,N_13860);
nor U18646 (N_18646,N_14154,N_12457);
nor U18647 (N_18647,N_12355,N_12950);
and U18648 (N_18648,N_12919,N_15526);
or U18649 (N_18649,N_14777,N_12205);
xor U18650 (N_18650,N_12505,N_14111);
and U18651 (N_18651,N_14229,N_13855);
nand U18652 (N_18652,N_13110,N_14639);
and U18653 (N_18653,N_12443,N_15195);
nor U18654 (N_18654,N_13090,N_15663);
nor U18655 (N_18655,N_13491,N_12940);
or U18656 (N_18656,N_13180,N_13905);
nand U18657 (N_18657,N_14689,N_15366);
nor U18658 (N_18658,N_13157,N_15534);
xnor U18659 (N_18659,N_14527,N_12650);
and U18660 (N_18660,N_14251,N_14101);
and U18661 (N_18661,N_15152,N_12877);
nand U18662 (N_18662,N_15750,N_15500);
and U18663 (N_18663,N_12096,N_12672);
nor U18664 (N_18664,N_13333,N_15987);
or U18665 (N_18665,N_14385,N_12171);
or U18666 (N_18666,N_13570,N_13779);
and U18667 (N_18667,N_13836,N_13016);
nand U18668 (N_18668,N_13851,N_14151);
xor U18669 (N_18669,N_12211,N_13727);
nor U18670 (N_18670,N_12128,N_15250);
nand U18671 (N_18671,N_13260,N_15782);
or U18672 (N_18672,N_14081,N_14137);
xnor U18673 (N_18673,N_15637,N_12880);
and U18674 (N_18674,N_13540,N_13156);
xor U18675 (N_18675,N_12295,N_15971);
nor U18676 (N_18676,N_15584,N_12578);
and U18677 (N_18677,N_15421,N_14187);
and U18678 (N_18678,N_13354,N_12703);
and U18679 (N_18679,N_13697,N_14637);
nand U18680 (N_18680,N_12730,N_12150);
nand U18681 (N_18681,N_13225,N_12027);
nor U18682 (N_18682,N_13404,N_15537);
and U18683 (N_18683,N_14201,N_12672);
or U18684 (N_18684,N_13827,N_15846);
and U18685 (N_18685,N_14578,N_14895);
and U18686 (N_18686,N_12979,N_13796);
xor U18687 (N_18687,N_14962,N_13251);
or U18688 (N_18688,N_12842,N_14480);
nand U18689 (N_18689,N_14790,N_14201);
nand U18690 (N_18690,N_13423,N_12437);
nor U18691 (N_18691,N_12437,N_14725);
nor U18692 (N_18692,N_13759,N_15554);
and U18693 (N_18693,N_13526,N_13127);
and U18694 (N_18694,N_15828,N_12906);
nand U18695 (N_18695,N_14291,N_15888);
xor U18696 (N_18696,N_13589,N_14989);
nor U18697 (N_18697,N_12042,N_13331);
and U18698 (N_18698,N_13391,N_15709);
nor U18699 (N_18699,N_13164,N_12249);
and U18700 (N_18700,N_13646,N_14368);
and U18701 (N_18701,N_15243,N_13087);
xnor U18702 (N_18702,N_12841,N_14181);
nand U18703 (N_18703,N_13793,N_12813);
xor U18704 (N_18704,N_12186,N_15667);
and U18705 (N_18705,N_14518,N_14756);
xnor U18706 (N_18706,N_14055,N_15282);
nand U18707 (N_18707,N_14247,N_15938);
and U18708 (N_18708,N_12970,N_13278);
and U18709 (N_18709,N_12044,N_13710);
or U18710 (N_18710,N_12891,N_12302);
or U18711 (N_18711,N_14745,N_14390);
nand U18712 (N_18712,N_12589,N_12434);
and U18713 (N_18713,N_15827,N_13479);
nand U18714 (N_18714,N_12127,N_12077);
nor U18715 (N_18715,N_14989,N_13487);
or U18716 (N_18716,N_12812,N_14519);
nand U18717 (N_18717,N_12933,N_13211);
or U18718 (N_18718,N_14949,N_14489);
nor U18719 (N_18719,N_12140,N_12670);
or U18720 (N_18720,N_13476,N_13190);
and U18721 (N_18721,N_14300,N_13965);
and U18722 (N_18722,N_13004,N_14284);
nand U18723 (N_18723,N_14133,N_15193);
and U18724 (N_18724,N_14236,N_12309);
xor U18725 (N_18725,N_13685,N_14083);
xnor U18726 (N_18726,N_14625,N_13345);
xnor U18727 (N_18727,N_15168,N_12345);
nor U18728 (N_18728,N_14229,N_14342);
nand U18729 (N_18729,N_15329,N_12713);
and U18730 (N_18730,N_14284,N_14121);
and U18731 (N_18731,N_14545,N_15059);
and U18732 (N_18732,N_14391,N_13374);
nand U18733 (N_18733,N_13982,N_14844);
nor U18734 (N_18734,N_12470,N_15624);
xnor U18735 (N_18735,N_12103,N_13937);
or U18736 (N_18736,N_15259,N_15914);
nand U18737 (N_18737,N_12960,N_15650);
nand U18738 (N_18738,N_14535,N_13372);
nor U18739 (N_18739,N_15583,N_15152);
and U18740 (N_18740,N_15441,N_15869);
or U18741 (N_18741,N_12511,N_13868);
nand U18742 (N_18742,N_13063,N_15512);
and U18743 (N_18743,N_14685,N_15041);
and U18744 (N_18744,N_12863,N_15329);
or U18745 (N_18745,N_14471,N_13052);
nor U18746 (N_18746,N_12868,N_13811);
nand U18747 (N_18747,N_13838,N_15871);
or U18748 (N_18748,N_14970,N_14608);
nand U18749 (N_18749,N_13985,N_15313);
nand U18750 (N_18750,N_15957,N_13185);
or U18751 (N_18751,N_15690,N_13081);
xor U18752 (N_18752,N_15846,N_12225);
xor U18753 (N_18753,N_12793,N_12787);
or U18754 (N_18754,N_15326,N_14017);
xnor U18755 (N_18755,N_15318,N_15053);
nand U18756 (N_18756,N_15805,N_14887);
and U18757 (N_18757,N_13885,N_12003);
xnor U18758 (N_18758,N_12032,N_15936);
or U18759 (N_18759,N_15988,N_14030);
or U18760 (N_18760,N_14405,N_15966);
nand U18761 (N_18761,N_14685,N_14930);
nor U18762 (N_18762,N_12099,N_15693);
or U18763 (N_18763,N_15092,N_13516);
and U18764 (N_18764,N_14226,N_14662);
xor U18765 (N_18765,N_15089,N_14006);
and U18766 (N_18766,N_13331,N_15665);
or U18767 (N_18767,N_14351,N_15799);
nor U18768 (N_18768,N_12174,N_12069);
nand U18769 (N_18769,N_12302,N_15528);
nand U18770 (N_18770,N_14539,N_15366);
nor U18771 (N_18771,N_13123,N_13006);
and U18772 (N_18772,N_12311,N_14207);
or U18773 (N_18773,N_12296,N_13985);
xnor U18774 (N_18774,N_13929,N_13260);
or U18775 (N_18775,N_15991,N_15538);
and U18776 (N_18776,N_13081,N_15727);
xor U18777 (N_18777,N_12306,N_15823);
nand U18778 (N_18778,N_13066,N_14204);
or U18779 (N_18779,N_15846,N_15989);
xnor U18780 (N_18780,N_15852,N_15676);
xor U18781 (N_18781,N_12290,N_12143);
nor U18782 (N_18782,N_14377,N_12714);
xor U18783 (N_18783,N_12973,N_15267);
or U18784 (N_18784,N_13402,N_14039);
nand U18785 (N_18785,N_14202,N_15152);
and U18786 (N_18786,N_12534,N_15538);
nor U18787 (N_18787,N_13648,N_13429);
or U18788 (N_18788,N_14550,N_15391);
or U18789 (N_18789,N_13830,N_12316);
xnor U18790 (N_18790,N_14387,N_15033);
xor U18791 (N_18791,N_15775,N_15506);
or U18792 (N_18792,N_14534,N_13695);
xnor U18793 (N_18793,N_13767,N_14579);
nor U18794 (N_18794,N_12562,N_14589);
nor U18795 (N_18795,N_15006,N_15067);
or U18796 (N_18796,N_14901,N_14755);
nand U18797 (N_18797,N_13042,N_12874);
nor U18798 (N_18798,N_14810,N_13088);
xor U18799 (N_18799,N_14250,N_14292);
nor U18800 (N_18800,N_12939,N_12057);
or U18801 (N_18801,N_12923,N_13754);
nor U18802 (N_18802,N_12601,N_15934);
and U18803 (N_18803,N_14498,N_13123);
nand U18804 (N_18804,N_14859,N_12518);
nand U18805 (N_18805,N_15542,N_13818);
nor U18806 (N_18806,N_12658,N_13314);
xor U18807 (N_18807,N_13509,N_12130);
and U18808 (N_18808,N_14592,N_12370);
and U18809 (N_18809,N_14521,N_15849);
nor U18810 (N_18810,N_14165,N_15571);
or U18811 (N_18811,N_12980,N_13622);
nand U18812 (N_18812,N_13241,N_15107);
and U18813 (N_18813,N_12594,N_12544);
nand U18814 (N_18814,N_15139,N_13426);
or U18815 (N_18815,N_12594,N_14458);
xor U18816 (N_18816,N_12922,N_15731);
xor U18817 (N_18817,N_14742,N_13818);
nand U18818 (N_18818,N_15946,N_12150);
nor U18819 (N_18819,N_13150,N_12895);
and U18820 (N_18820,N_14718,N_13437);
xnor U18821 (N_18821,N_12954,N_12123);
nand U18822 (N_18822,N_15862,N_12559);
nor U18823 (N_18823,N_14794,N_15148);
nor U18824 (N_18824,N_14827,N_14554);
or U18825 (N_18825,N_13281,N_15408);
or U18826 (N_18826,N_14386,N_14634);
and U18827 (N_18827,N_13552,N_13171);
and U18828 (N_18828,N_15030,N_15709);
or U18829 (N_18829,N_15650,N_12508);
and U18830 (N_18830,N_14436,N_13769);
xnor U18831 (N_18831,N_15533,N_13119);
nand U18832 (N_18832,N_15252,N_12570);
and U18833 (N_18833,N_14884,N_12323);
xnor U18834 (N_18834,N_13177,N_12136);
and U18835 (N_18835,N_13218,N_13145);
xnor U18836 (N_18836,N_13966,N_13567);
xnor U18837 (N_18837,N_13566,N_13555);
nand U18838 (N_18838,N_15589,N_15708);
or U18839 (N_18839,N_14790,N_13185);
nand U18840 (N_18840,N_14638,N_14565);
and U18841 (N_18841,N_13053,N_13064);
xor U18842 (N_18842,N_12499,N_15956);
xnor U18843 (N_18843,N_15059,N_12792);
nor U18844 (N_18844,N_13339,N_12762);
xor U18845 (N_18845,N_15091,N_14759);
or U18846 (N_18846,N_13660,N_13928);
xor U18847 (N_18847,N_13119,N_12392);
or U18848 (N_18848,N_14268,N_12524);
or U18849 (N_18849,N_13503,N_15010);
and U18850 (N_18850,N_14280,N_15087);
xnor U18851 (N_18851,N_15615,N_15266);
xnor U18852 (N_18852,N_13273,N_12307);
nand U18853 (N_18853,N_12782,N_14819);
nand U18854 (N_18854,N_14105,N_15285);
nand U18855 (N_18855,N_14206,N_12648);
xor U18856 (N_18856,N_13031,N_12493);
xor U18857 (N_18857,N_14330,N_13802);
xnor U18858 (N_18858,N_13346,N_13392);
and U18859 (N_18859,N_14867,N_13103);
and U18860 (N_18860,N_13513,N_14100);
or U18861 (N_18861,N_12997,N_14757);
xnor U18862 (N_18862,N_12811,N_14777);
nor U18863 (N_18863,N_12053,N_12520);
or U18864 (N_18864,N_14593,N_15642);
xnor U18865 (N_18865,N_13360,N_14052);
and U18866 (N_18866,N_12323,N_15904);
and U18867 (N_18867,N_13025,N_15938);
nor U18868 (N_18868,N_12223,N_13848);
nand U18869 (N_18869,N_14451,N_14105);
and U18870 (N_18870,N_13196,N_15913);
nor U18871 (N_18871,N_15833,N_14544);
and U18872 (N_18872,N_14813,N_13167);
nor U18873 (N_18873,N_15258,N_12944);
nand U18874 (N_18874,N_14566,N_14692);
nand U18875 (N_18875,N_15406,N_14140);
and U18876 (N_18876,N_12381,N_12659);
nand U18877 (N_18877,N_14980,N_15517);
or U18878 (N_18878,N_12514,N_13371);
nor U18879 (N_18879,N_12409,N_13117);
xor U18880 (N_18880,N_15018,N_13680);
xor U18881 (N_18881,N_14766,N_12121);
nor U18882 (N_18882,N_14790,N_12124);
nand U18883 (N_18883,N_14879,N_13387);
xnor U18884 (N_18884,N_15171,N_14510);
nand U18885 (N_18885,N_14211,N_15726);
or U18886 (N_18886,N_15263,N_14159);
nor U18887 (N_18887,N_12411,N_14473);
nor U18888 (N_18888,N_13990,N_12681);
xnor U18889 (N_18889,N_12088,N_15155);
and U18890 (N_18890,N_15581,N_15970);
nand U18891 (N_18891,N_12610,N_14795);
or U18892 (N_18892,N_15376,N_15719);
xor U18893 (N_18893,N_15456,N_13519);
xnor U18894 (N_18894,N_12086,N_14136);
nor U18895 (N_18895,N_12431,N_12562);
xor U18896 (N_18896,N_14112,N_13593);
or U18897 (N_18897,N_15346,N_14171);
and U18898 (N_18898,N_14652,N_12363);
and U18899 (N_18899,N_14945,N_15553);
nor U18900 (N_18900,N_14471,N_13375);
xnor U18901 (N_18901,N_14440,N_15676);
and U18902 (N_18902,N_14505,N_15833);
or U18903 (N_18903,N_15549,N_14946);
xor U18904 (N_18904,N_12923,N_14355);
or U18905 (N_18905,N_12452,N_15419);
or U18906 (N_18906,N_12152,N_12059);
or U18907 (N_18907,N_12310,N_13728);
xnor U18908 (N_18908,N_14580,N_12978);
nand U18909 (N_18909,N_14426,N_13060);
or U18910 (N_18910,N_12408,N_14799);
nor U18911 (N_18911,N_12423,N_12501);
xor U18912 (N_18912,N_12528,N_13382);
xor U18913 (N_18913,N_12512,N_12357);
xnor U18914 (N_18914,N_15191,N_14860);
and U18915 (N_18915,N_12025,N_13132);
nor U18916 (N_18916,N_14791,N_15702);
nand U18917 (N_18917,N_13235,N_12471);
nand U18918 (N_18918,N_14320,N_13814);
xnor U18919 (N_18919,N_13010,N_12027);
or U18920 (N_18920,N_12083,N_14978);
nand U18921 (N_18921,N_13740,N_12468);
and U18922 (N_18922,N_14589,N_12227);
or U18923 (N_18923,N_13053,N_15049);
and U18924 (N_18924,N_14444,N_13328);
nand U18925 (N_18925,N_13380,N_15577);
nor U18926 (N_18926,N_13135,N_15801);
and U18927 (N_18927,N_15343,N_12294);
or U18928 (N_18928,N_15913,N_14382);
xor U18929 (N_18929,N_14462,N_13285);
and U18930 (N_18930,N_12703,N_13046);
nor U18931 (N_18931,N_14418,N_15593);
or U18932 (N_18932,N_12746,N_13279);
or U18933 (N_18933,N_12578,N_12548);
or U18934 (N_18934,N_13382,N_14655);
nor U18935 (N_18935,N_15165,N_14436);
and U18936 (N_18936,N_15797,N_13923);
nor U18937 (N_18937,N_14954,N_15053);
nor U18938 (N_18938,N_14924,N_12097);
xor U18939 (N_18939,N_13205,N_15521);
and U18940 (N_18940,N_15624,N_13963);
and U18941 (N_18941,N_13207,N_12217);
or U18942 (N_18942,N_15143,N_13938);
nand U18943 (N_18943,N_15726,N_14517);
or U18944 (N_18944,N_13357,N_13762);
xor U18945 (N_18945,N_15296,N_12183);
xnor U18946 (N_18946,N_12890,N_14331);
nor U18947 (N_18947,N_14978,N_14191);
nand U18948 (N_18948,N_15378,N_13467);
xor U18949 (N_18949,N_15984,N_14888);
nor U18950 (N_18950,N_15011,N_14058);
nor U18951 (N_18951,N_15938,N_13493);
and U18952 (N_18952,N_15528,N_13961);
or U18953 (N_18953,N_13659,N_14045);
nor U18954 (N_18954,N_14694,N_12829);
nor U18955 (N_18955,N_13510,N_15759);
and U18956 (N_18956,N_14488,N_12858);
or U18957 (N_18957,N_13518,N_15402);
nand U18958 (N_18958,N_13925,N_15442);
xor U18959 (N_18959,N_15655,N_13288);
nor U18960 (N_18960,N_12791,N_15370);
or U18961 (N_18961,N_13834,N_12384);
nor U18962 (N_18962,N_14381,N_12520);
and U18963 (N_18963,N_13793,N_14496);
nor U18964 (N_18964,N_15119,N_14304);
xnor U18965 (N_18965,N_13412,N_13152);
or U18966 (N_18966,N_15717,N_13651);
xor U18967 (N_18967,N_12800,N_14839);
nor U18968 (N_18968,N_15902,N_14839);
nand U18969 (N_18969,N_15882,N_15043);
and U18970 (N_18970,N_14511,N_12437);
or U18971 (N_18971,N_15477,N_12654);
xor U18972 (N_18972,N_14062,N_13448);
xnor U18973 (N_18973,N_13461,N_13055);
or U18974 (N_18974,N_15531,N_12627);
and U18975 (N_18975,N_13082,N_12897);
or U18976 (N_18976,N_13968,N_13329);
or U18977 (N_18977,N_14969,N_12805);
or U18978 (N_18978,N_15476,N_12366);
nor U18979 (N_18979,N_13888,N_12107);
or U18980 (N_18980,N_14416,N_14621);
or U18981 (N_18981,N_15030,N_14342);
xnor U18982 (N_18982,N_15047,N_12055);
nand U18983 (N_18983,N_12463,N_15942);
nor U18984 (N_18984,N_12004,N_13002);
and U18985 (N_18985,N_15262,N_15455);
nor U18986 (N_18986,N_12756,N_13497);
nor U18987 (N_18987,N_14145,N_12135);
nor U18988 (N_18988,N_15223,N_14337);
or U18989 (N_18989,N_12114,N_14762);
xnor U18990 (N_18990,N_12434,N_13120);
nand U18991 (N_18991,N_12472,N_12275);
or U18992 (N_18992,N_15706,N_12520);
nand U18993 (N_18993,N_13669,N_13052);
nor U18994 (N_18994,N_15249,N_13746);
nor U18995 (N_18995,N_13345,N_15248);
nand U18996 (N_18996,N_12497,N_13894);
nor U18997 (N_18997,N_12146,N_13111);
and U18998 (N_18998,N_12014,N_12567);
and U18999 (N_18999,N_15329,N_14378);
nor U19000 (N_19000,N_14695,N_15114);
nand U19001 (N_19001,N_15333,N_15077);
xnor U19002 (N_19002,N_14972,N_14598);
nand U19003 (N_19003,N_12046,N_14709);
nand U19004 (N_19004,N_15655,N_14374);
xor U19005 (N_19005,N_15870,N_14272);
and U19006 (N_19006,N_13036,N_15905);
nand U19007 (N_19007,N_12578,N_14529);
nand U19008 (N_19008,N_13157,N_13228);
xor U19009 (N_19009,N_13102,N_15455);
nor U19010 (N_19010,N_15452,N_15611);
xnor U19011 (N_19011,N_14988,N_13516);
and U19012 (N_19012,N_14991,N_14214);
and U19013 (N_19013,N_15210,N_15023);
or U19014 (N_19014,N_13924,N_13262);
xor U19015 (N_19015,N_14026,N_12755);
nand U19016 (N_19016,N_12621,N_13587);
or U19017 (N_19017,N_15678,N_12793);
xnor U19018 (N_19018,N_13594,N_14568);
or U19019 (N_19019,N_12282,N_12027);
nor U19020 (N_19020,N_14285,N_15437);
or U19021 (N_19021,N_12057,N_13990);
xnor U19022 (N_19022,N_15124,N_14091);
nand U19023 (N_19023,N_14436,N_15328);
nand U19024 (N_19024,N_14991,N_14892);
nand U19025 (N_19025,N_13091,N_13116);
and U19026 (N_19026,N_15561,N_14051);
nand U19027 (N_19027,N_13657,N_13783);
or U19028 (N_19028,N_12521,N_14402);
or U19029 (N_19029,N_12159,N_13579);
nand U19030 (N_19030,N_13143,N_15358);
nand U19031 (N_19031,N_13946,N_12073);
nand U19032 (N_19032,N_13731,N_15401);
and U19033 (N_19033,N_15154,N_14770);
nor U19034 (N_19034,N_13041,N_15353);
nor U19035 (N_19035,N_13559,N_15181);
xor U19036 (N_19036,N_13491,N_13639);
nand U19037 (N_19037,N_14832,N_13037);
nor U19038 (N_19038,N_15774,N_14820);
xnor U19039 (N_19039,N_12055,N_13595);
or U19040 (N_19040,N_15820,N_13191);
and U19041 (N_19041,N_14362,N_15799);
and U19042 (N_19042,N_13640,N_15048);
nor U19043 (N_19043,N_13541,N_12477);
xor U19044 (N_19044,N_13965,N_14061);
nand U19045 (N_19045,N_13192,N_15733);
nand U19046 (N_19046,N_14081,N_14282);
nor U19047 (N_19047,N_12243,N_13319);
or U19048 (N_19048,N_12180,N_14862);
nor U19049 (N_19049,N_12862,N_14795);
xor U19050 (N_19050,N_12468,N_12129);
or U19051 (N_19051,N_12663,N_15988);
or U19052 (N_19052,N_14249,N_15766);
xor U19053 (N_19053,N_15548,N_14017);
nand U19054 (N_19054,N_15140,N_14555);
nor U19055 (N_19055,N_14983,N_12724);
and U19056 (N_19056,N_12236,N_14040);
xor U19057 (N_19057,N_13313,N_12328);
and U19058 (N_19058,N_14068,N_15249);
nor U19059 (N_19059,N_14899,N_13400);
and U19060 (N_19060,N_13378,N_13844);
and U19061 (N_19061,N_13669,N_12337);
xor U19062 (N_19062,N_14255,N_13650);
nor U19063 (N_19063,N_13630,N_13541);
xnor U19064 (N_19064,N_12256,N_15682);
xnor U19065 (N_19065,N_13228,N_14955);
nor U19066 (N_19066,N_14510,N_15326);
nor U19067 (N_19067,N_14851,N_13667);
and U19068 (N_19068,N_14041,N_12960);
or U19069 (N_19069,N_15393,N_13665);
or U19070 (N_19070,N_15231,N_15379);
nor U19071 (N_19071,N_14170,N_12809);
or U19072 (N_19072,N_13210,N_13288);
and U19073 (N_19073,N_12201,N_14952);
nor U19074 (N_19074,N_14208,N_15308);
nand U19075 (N_19075,N_14289,N_14900);
and U19076 (N_19076,N_13179,N_13281);
and U19077 (N_19077,N_13000,N_13186);
nor U19078 (N_19078,N_15735,N_13052);
xnor U19079 (N_19079,N_15696,N_13281);
nor U19080 (N_19080,N_14184,N_12465);
nor U19081 (N_19081,N_13551,N_14810);
nand U19082 (N_19082,N_15800,N_12477);
or U19083 (N_19083,N_15690,N_12719);
xor U19084 (N_19084,N_14341,N_12895);
nor U19085 (N_19085,N_14937,N_15684);
xnor U19086 (N_19086,N_14635,N_15976);
and U19087 (N_19087,N_14160,N_13778);
nand U19088 (N_19088,N_13058,N_15786);
and U19089 (N_19089,N_15389,N_14571);
xor U19090 (N_19090,N_14186,N_14677);
nand U19091 (N_19091,N_15298,N_12884);
nand U19092 (N_19092,N_13384,N_15453);
nor U19093 (N_19093,N_13163,N_15100);
or U19094 (N_19094,N_15227,N_13055);
nand U19095 (N_19095,N_15559,N_13527);
nand U19096 (N_19096,N_13874,N_14666);
and U19097 (N_19097,N_13161,N_12528);
or U19098 (N_19098,N_15274,N_15642);
xor U19099 (N_19099,N_14219,N_14591);
xnor U19100 (N_19100,N_14566,N_15320);
nor U19101 (N_19101,N_13800,N_12748);
nand U19102 (N_19102,N_12477,N_14787);
nand U19103 (N_19103,N_12976,N_15731);
or U19104 (N_19104,N_13690,N_15834);
nand U19105 (N_19105,N_14930,N_14710);
xnor U19106 (N_19106,N_14652,N_12838);
and U19107 (N_19107,N_15679,N_13251);
and U19108 (N_19108,N_14167,N_14784);
nand U19109 (N_19109,N_15628,N_13211);
nor U19110 (N_19110,N_12998,N_15193);
and U19111 (N_19111,N_14530,N_14227);
xor U19112 (N_19112,N_13964,N_15699);
xnor U19113 (N_19113,N_14331,N_13060);
xor U19114 (N_19114,N_14634,N_13840);
or U19115 (N_19115,N_14592,N_12808);
nor U19116 (N_19116,N_13610,N_15791);
and U19117 (N_19117,N_14855,N_12460);
nor U19118 (N_19118,N_15044,N_13355);
nand U19119 (N_19119,N_14069,N_13609);
and U19120 (N_19120,N_14502,N_15802);
and U19121 (N_19121,N_12860,N_14597);
nor U19122 (N_19122,N_14384,N_12745);
and U19123 (N_19123,N_12036,N_15456);
xnor U19124 (N_19124,N_15734,N_15483);
and U19125 (N_19125,N_12261,N_12661);
nand U19126 (N_19126,N_12482,N_12453);
nand U19127 (N_19127,N_13332,N_14614);
nand U19128 (N_19128,N_13492,N_13236);
xnor U19129 (N_19129,N_13165,N_14139);
nand U19130 (N_19130,N_12896,N_13625);
and U19131 (N_19131,N_13782,N_12839);
or U19132 (N_19132,N_15907,N_13971);
nand U19133 (N_19133,N_14881,N_12261);
nand U19134 (N_19134,N_14791,N_15283);
xnor U19135 (N_19135,N_14652,N_12392);
nor U19136 (N_19136,N_12526,N_15361);
and U19137 (N_19137,N_15523,N_13787);
nor U19138 (N_19138,N_15178,N_15497);
nor U19139 (N_19139,N_15677,N_12935);
nor U19140 (N_19140,N_13987,N_15914);
xnor U19141 (N_19141,N_12256,N_15566);
nor U19142 (N_19142,N_12023,N_13854);
nor U19143 (N_19143,N_14047,N_12794);
xnor U19144 (N_19144,N_13267,N_12811);
xnor U19145 (N_19145,N_13987,N_12319);
xor U19146 (N_19146,N_15884,N_14457);
and U19147 (N_19147,N_15806,N_13525);
nor U19148 (N_19148,N_13655,N_15846);
or U19149 (N_19149,N_12432,N_13172);
nand U19150 (N_19150,N_12480,N_15746);
nor U19151 (N_19151,N_14510,N_12841);
nand U19152 (N_19152,N_14837,N_13485);
xor U19153 (N_19153,N_14522,N_12840);
nand U19154 (N_19154,N_14076,N_13250);
xor U19155 (N_19155,N_15422,N_15932);
and U19156 (N_19156,N_14415,N_12171);
xnor U19157 (N_19157,N_13499,N_12483);
nand U19158 (N_19158,N_13446,N_14661);
nor U19159 (N_19159,N_13261,N_13525);
and U19160 (N_19160,N_13299,N_13736);
and U19161 (N_19161,N_12091,N_14777);
xor U19162 (N_19162,N_13439,N_13201);
xor U19163 (N_19163,N_14626,N_13950);
nand U19164 (N_19164,N_12146,N_14681);
and U19165 (N_19165,N_12504,N_15000);
or U19166 (N_19166,N_12604,N_13892);
or U19167 (N_19167,N_15988,N_15646);
nor U19168 (N_19168,N_14284,N_13306);
or U19169 (N_19169,N_13662,N_12672);
or U19170 (N_19170,N_14870,N_14245);
xor U19171 (N_19171,N_13911,N_13361);
nand U19172 (N_19172,N_13321,N_14771);
or U19173 (N_19173,N_15169,N_14803);
xnor U19174 (N_19174,N_13837,N_14749);
and U19175 (N_19175,N_14849,N_12078);
or U19176 (N_19176,N_15809,N_12437);
nand U19177 (N_19177,N_13726,N_12043);
xor U19178 (N_19178,N_14326,N_12589);
nor U19179 (N_19179,N_15187,N_15235);
nand U19180 (N_19180,N_15697,N_15690);
nor U19181 (N_19181,N_15844,N_14858);
or U19182 (N_19182,N_15473,N_13400);
nand U19183 (N_19183,N_15364,N_12648);
and U19184 (N_19184,N_15311,N_13854);
or U19185 (N_19185,N_15854,N_13139);
nor U19186 (N_19186,N_12718,N_13323);
nor U19187 (N_19187,N_15456,N_13340);
and U19188 (N_19188,N_15340,N_12629);
or U19189 (N_19189,N_14130,N_12369);
xor U19190 (N_19190,N_14271,N_14590);
xor U19191 (N_19191,N_14450,N_15871);
nor U19192 (N_19192,N_12675,N_13073);
or U19193 (N_19193,N_15745,N_12060);
or U19194 (N_19194,N_12255,N_14957);
or U19195 (N_19195,N_12158,N_14536);
nor U19196 (N_19196,N_12141,N_14614);
or U19197 (N_19197,N_15948,N_12492);
or U19198 (N_19198,N_15950,N_15807);
nor U19199 (N_19199,N_14257,N_14615);
nand U19200 (N_19200,N_15353,N_15476);
nand U19201 (N_19201,N_13111,N_14920);
nor U19202 (N_19202,N_14379,N_13248);
or U19203 (N_19203,N_14486,N_12299);
and U19204 (N_19204,N_14168,N_15682);
nand U19205 (N_19205,N_12365,N_13880);
xnor U19206 (N_19206,N_14410,N_12821);
nand U19207 (N_19207,N_14495,N_12184);
nor U19208 (N_19208,N_12286,N_13705);
nand U19209 (N_19209,N_15383,N_14832);
nand U19210 (N_19210,N_13336,N_15480);
nand U19211 (N_19211,N_12851,N_15483);
or U19212 (N_19212,N_13058,N_15325);
and U19213 (N_19213,N_13194,N_12902);
and U19214 (N_19214,N_15759,N_13130);
xor U19215 (N_19215,N_13180,N_12663);
nor U19216 (N_19216,N_12332,N_14536);
nor U19217 (N_19217,N_13080,N_12779);
or U19218 (N_19218,N_14068,N_15171);
or U19219 (N_19219,N_13275,N_13481);
nand U19220 (N_19220,N_12939,N_14682);
nand U19221 (N_19221,N_13449,N_12289);
or U19222 (N_19222,N_15787,N_14767);
xnor U19223 (N_19223,N_13700,N_13651);
xor U19224 (N_19224,N_12145,N_15873);
xor U19225 (N_19225,N_13425,N_14818);
or U19226 (N_19226,N_15379,N_15774);
or U19227 (N_19227,N_12631,N_12438);
or U19228 (N_19228,N_13802,N_14695);
and U19229 (N_19229,N_12240,N_13581);
xor U19230 (N_19230,N_15717,N_13454);
and U19231 (N_19231,N_15484,N_12618);
nor U19232 (N_19232,N_15645,N_15208);
nor U19233 (N_19233,N_12615,N_13199);
xnor U19234 (N_19234,N_15610,N_13524);
xnor U19235 (N_19235,N_13824,N_15701);
nand U19236 (N_19236,N_15820,N_15867);
nor U19237 (N_19237,N_14697,N_15513);
nand U19238 (N_19238,N_12976,N_13844);
nor U19239 (N_19239,N_12454,N_13553);
or U19240 (N_19240,N_12512,N_13382);
nand U19241 (N_19241,N_12623,N_15706);
nand U19242 (N_19242,N_15559,N_14704);
nor U19243 (N_19243,N_15184,N_14700);
nor U19244 (N_19244,N_14358,N_12851);
or U19245 (N_19245,N_13985,N_15303);
nand U19246 (N_19246,N_15593,N_12666);
nand U19247 (N_19247,N_13501,N_14932);
xnor U19248 (N_19248,N_13492,N_12698);
and U19249 (N_19249,N_12674,N_14603);
or U19250 (N_19250,N_14380,N_14660);
xor U19251 (N_19251,N_12615,N_12297);
nand U19252 (N_19252,N_14934,N_13184);
nor U19253 (N_19253,N_13886,N_12066);
nand U19254 (N_19254,N_13770,N_12433);
or U19255 (N_19255,N_12557,N_12703);
or U19256 (N_19256,N_14193,N_12115);
xor U19257 (N_19257,N_12148,N_13936);
nand U19258 (N_19258,N_13796,N_12427);
nor U19259 (N_19259,N_15754,N_12609);
xnor U19260 (N_19260,N_14953,N_15159);
or U19261 (N_19261,N_13082,N_12915);
and U19262 (N_19262,N_13112,N_13612);
nand U19263 (N_19263,N_15748,N_14675);
and U19264 (N_19264,N_15450,N_15257);
and U19265 (N_19265,N_12196,N_14289);
xor U19266 (N_19266,N_12214,N_13621);
or U19267 (N_19267,N_15448,N_14280);
nand U19268 (N_19268,N_13796,N_15557);
nand U19269 (N_19269,N_12756,N_15356);
nand U19270 (N_19270,N_14737,N_13327);
and U19271 (N_19271,N_14084,N_13413);
xnor U19272 (N_19272,N_13456,N_14785);
and U19273 (N_19273,N_14794,N_15363);
xnor U19274 (N_19274,N_12803,N_12092);
and U19275 (N_19275,N_15116,N_15850);
nand U19276 (N_19276,N_14496,N_15356);
nor U19277 (N_19277,N_12913,N_12076);
or U19278 (N_19278,N_13927,N_14056);
xnor U19279 (N_19279,N_14780,N_12864);
and U19280 (N_19280,N_14875,N_14732);
or U19281 (N_19281,N_12214,N_14323);
and U19282 (N_19282,N_13136,N_13846);
and U19283 (N_19283,N_13692,N_15969);
or U19284 (N_19284,N_13047,N_12999);
or U19285 (N_19285,N_13041,N_13162);
nor U19286 (N_19286,N_13558,N_14353);
or U19287 (N_19287,N_13138,N_15925);
or U19288 (N_19288,N_12659,N_13480);
and U19289 (N_19289,N_15047,N_14018);
nor U19290 (N_19290,N_14541,N_13501);
or U19291 (N_19291,N_14531,N_14423);
or U19292 (N_19292,N_15222,N_12094);
nor U19293 (N_19293,N_12201,N_14823);
nor U19294 (N_19294,N_14412,N_13279);
or U19295 (N_19295,N_14234,N_12528);
or U19296 (N_19296,N_15936,N_15206);
xnor U19297 (N_19297,N_12583,N_13384);
or U19298 (N_19298,N_14236,N_12397);
nand U19299 (N_19299,N_13174,N_12258);
or U19300 (N_19300,N_12222,N_14043);
or U19301 (N_19301,N_15655,N_15264);
xnor U19302 (N_19302,N_13540,N_15289);
xor U19303 (N_19303,N_14838,N_13527);
and U19304 (N_19304,N_13355,N_14134);
or U19305 (N_19305,N_15224,N_15189);
or U19306 (N_19306,N_12974,N_12431);
nand U19307 (N_19307,N_14596,N_13520);
and U19308 (N_19308,N_12468,N_13349);
xnor U19309 (N_19309,N_15030,N_15009);
nand U19310 (N_19310,N_13595,N_14016);
nor U19311 (N_19311,N_12934,N_13411);
xnor U19312 (N_19312,N_12359,N_15269);
and U19313 (N_19313,N_13634,N_12121);
or U19314 (N_19314,N_12756,N_12079);
nand U19315 (N_19315,N_13417,N_14096);
nand U19316 (N_19316,N_12459,N_15066);
or U19317 (N_19317,N_14953,N_13398);
and U19318 (N_19318,N_13398,N_13554);
nor U19319 (N_19319,N_13122,N_12355);
xnor U19320 (N_19320,N_13000,N_12598);
nor U19321 (N_19321,N_14091,N_14126);
or U19322 (N_19322,N_13655,N_12777);
xnor U19323 (N_19323,N_15938,N_12281);
nand U19324 (N_19324,N_12804,N_13686);
and U19325 (N_19325,N_15442,N_12915);
nand U19326 (N_19326,N_12874,N_12986);
nor U19327 (N_19327,N_14954,N_12240);
nor U19328 (N_19328,N_13067,N_15387);
or U19329 (N_19329,N_14511,N_12199);
nor U19330 (N_19330,N_12949,N_12305);
nand U19331 (N_19331,N_15830,N_13940);
nor U19332 (N_19332,N_14301,N_13600);
nor U19333 (N_19333,N_12176,N_15437);
or U19334 (N_19334,N_13398,N_14042);
and U19335 (N_19335,N_15167,N_15479);
xnor U19336 (N_19336,N_12264,N_13340);
xor U19337 (N_19337,N_12458,N_14756);
and U19338 (N_19338,N_15875,N_14551);
or U19339 (N_19339,N_13631,N_12233);
nor U19340 (N_19340,N_14203,N_14763);
nand U19341 (N_19341,N_13055,N_13564);
xor U19342 (N_19342,N_12964,N_12828);
or U19343 (N_19343,N_12976,N_15072);
xnor U19344 (N_19344,N_13991,N_15460);
nand U19345 (N_19345,N_12167,N_13864);
xor U19346 (N_19346,N_13123,N_12751);
and U19347 (N_19347,N_14079,N_12395);
nor U19348 (N_19348,N_15082,N_12054);
and U19349 (N_19349,N_15306,N_13328);
or U19350 (N_19350,N_15828,N_13125);
or U19351 (N_19351,N_15830,N_14197);
and U19352 (N_19352,N_15147,N_15555);
xnor U19353 (N_19353,N_13857,N_13153);
nand U19354 (N_19354,N_12872,N_15278);
or U19355 (N_19355,N_14812,N_15752);
and U19356 (N_19356,N_15134,N_15830);
nor U19357 (N_19357,N_12520,N_12467);
nor U19358 (N_19358,N_12399,N_13685);
nor U19359 (N_19359,N_12878,N_12748);
nor U19360 (N_19360,N_12830,N_14369);
nor U19361 (N_19361,N_12952,N_14473);
or U19362 (N_19362,N_14417,N_13599);
and U19363 (N_19363,N_15801,N_13477);
nand U19364 (N_19364,N_12190,N_14318);
nand U19365 (N_19365,N_13456,N_14675);
and U19366 (N_19366,N_13734,N_12705);
nand U19367 (N_19367,N_13591,N_12434);
nand U19368 (N_19368,N_15675,N_12813);
and U19369 (N_19369,N_14800,N_12619);
nand U19370 (N_19370,N_14494,N_13365);
nand U19371 (N_19371,N_15359,N_12425);
nand U19372 (N_19372,N_14778,N_13374);
nor U19373 (N_19373,N_13208,N_13897);
nor U19374 (N_19374,N_14106,N_12442);
or U19375 (N_19375,N_15327,N_12534);
or U19376 (N_19376,N_12249,N_14618);
xor U19377 (N_19377,N_12582,N_12530);
nand U19378 (N_19378,N_12379,N_13683);
and U19379 (N_19379,N_13861,N_12577);
xnor U19380 (N_19380,N_12554,N_14141);
nand U19381 (N_19381,N_14729,N_13404);
or U19382 (N_19382,N_15588,N_14940);
xor U19383 (N_19383,N_12791,N_15919);
or U19384 (N_19384,N_14024,N_13958);
and U19385 (N_19385,N_12994,N_13386);
nor U19386 (N_19386,N_14177,N_15420);
xnor U19387 (N_19387,N_13168,N_13262);
and U19388 (N_19388,N_14299,N_12366);
or U19389 (N_19389,N_14504,N_12045);
nor U19390 (N_19390,N_14787,N_12125);
xor U19391 (N_19391,N_14101,N_12212);
nand U19392 (N_19392,N_13352,N_12052);
nand U19393 (N_19393,N_12445,N_12710);
and U19394 (N_19394,N_14554,N_12640);
xor U19395 (N_19395,N_15283,N_13713);
nand U19396 (N_19396,N_13002,N_12160);
and U19397 (N_19397,N_13142,N_13492);
xnor U19398 (N_19398,N_15646,N_15109);
xor U19399 (N_19399,N_15756,N_13253);
nor U19400 (N_19400,N_14158,N_12094);
nand U19401 (N_19401,N_13086,N_12140);
and U19402 (N_19402,N_14178,N_13625);
xnor U19403 (N_19403,N_15744,N_14545);
nor U19404 (N_19404,N_15116,N_13932);
xnor U19405 (N_19405,N_15657,N_15797);
xor U19406 (N_19406,N_12808,N_14181);
xor U19407 (N_19407,N_14534,N_13652);
nor U19408 (N_19408,N_14294,N_13427);
nor U19409 (N_19409,N_12952,N_14474);
and U19410 (N_19410,N_15015,N_15124);
and U19411 (N_19411,N_13846,N_14628);
and U19412 (N_19412,N_13512,N_12892);
and U19413 (N_19413,N_14668,N_14885);
xor U19414 (N_19414,N_13205,N_12884);
xnor U19415 (N_19415,N_14817,N_15165);
nand U19416 (N_19416,N_12215,N_15310);
or U19417 (N_19417,N_15519,N_15050);
nand U19418 (N_19418,N_13356,N_15149);
or U19419 (N_19419,N_12537,N_12084);
or U19420 (N_19420,N_14137,N_13943);
or U19421 (N_19421,N_14390,N_15715);
nor U19422 (N_19422,N_14734,N_15143);
or U19423 (N_19423,N_12761,N_15801);
xnor U19424 (N_19424,N_12459,N_13309);
or U19425 (N_19425,N_13732,N_14261);
nand U19426 (N_19426,N_15062,N_12765);
or U19427 (N_19427,N_12294,N_13990);
xor U19428 (N_19428,N_15566,N_13837);
and U19429 (N_19429,N_14336,N_14164);
nand U19430 (N_19430,N_13844,N_12353);
nand U19431 (N_19431,N_13199,N_15941);
nand U19432 (N_19432,N_13120,N_15675);
nor U19433 (N_19433,N_14086,N_13396);
nand U19434 (N_19434,N_15441,N_12038);
xnor U19435 (N_19435,N_13573,N_12867);
xnor U19436 (N_19436,N_15038,N_12091);
and U19437 (N_19437,N_14127,N_14662);
and U19438 (N_19438,N_13602,N_13893);
or U19439 (N_19439,N_12625,N_14498);
or U19440 (N_19440,N_12853,N_13646);
xnor U19441 (N_19441,N_13531,N_14342);
or U19442 (N_19442,N_15700,N_12773);
and U19443 (N_19443,N_14535,N_12780);
and U19444 (N_19444,N_14214,N_15951);
nor U19445 (N_19445,N_12429,N_13141);
xor U19446 (N_19446,N_13410,N_13151);
nand U19447 (N_19447,N_15507,N_14805);
xnor U19448 (N_19448,N_15481,N_12028);
nand U19449 (N_19449,N_12651,N_13362);
and U19450 (N_19450,N_14338,N_13922);
nor U19451 (N_19451,N_12726,N_12454);
and U19452 (N_19452,N_12296,N_15926);
nor U19453 (N_19453,N_14100,N_12523);
nand U19454 (N_19454,N_14176,N_14080);
or U19455 (N_19455,N_12168,N_13933);
nand U19456 (N_19456,N_13227,N_12388);
xor U19457 (N_19457,N_13771,N_13221);
xor U19458 (N_19458,N_12665,N_12152);
or U19459 (N_19459,N_13803,N_14620);
nand U19460 (N_19460,N_12573,N_12018);
nor U19461 (N_19461,N_15618,N_15218);
nand U19462 (N_19462,N_12086,N_14483);
nand U19463 (N_19463,N_13854,N_12831);
nor U19464 (N_19464,N_13805,N_14087);
and U19465 (N_19465,N_13977,N_12089);
and U19466 (N_19466,N_15249,N_14477);
or U19467 (N_19467,N_15101,N_15232);
and U19468 (N_19468,N_15237,N_14607);
xnor U19469 (N_19469,N_15414,N_12611);
or U19470 (N_19470,N_13710,N_13397);
and U19471 (N_19471,N_12486,N_13510);
and U19472 (N_19472,N_15744,N_14858);
xnor U19473 (N_19473,N_12956,N_14638);
xor U19474 (N_19474,N_14867,N_15265);
or U19475 (N_19475,N_14033,N_15820);
or U19476 (N_19476,N_13758,N_13827);
nor U19477 (N_19477,N_14163,N_12760);
nand U19478 (N_19478,N_15576,N_13835);
and U19479 (N_19479,N_13239,N_12575);
xnor U19480 (N_19480,N_13728,N_14481);
nor U19481 (N_19481,N_13772,N_15120);
or U19482 (N_19482,N_13013,N_13737);
xnor U19483 (N_19483,N_12742,N_13383);
or U19484 (N_19484,N_13839,N_12552);
or U19485 (N_19485,N_14342,N_15949);
nand U19486 (N_19486,N_12031,N_13473);
nand U19487 (N_19487,N_15188,N_14096);
or U19488 (N_19488,N_12513,N_13939);
and U19489 (N_19489,N_12356,N_12539);
nor U19490 (N_19490,N_12566,N_13228);
xnor U19491 (N_19491,N_13475,N_12894);
nor U19492 (N_19492,N_12864,N_14192);
or U19493 (N_19493,N_15875,N_14768);
xor U19494 (N_19494,N_14597,N_13270);
and U19495 (N_19495,N_14427,N_13773);
and U19496 (N_19496,N_12666,N_13519);
and U19497 (N_19497,N_12210,N_14460);
nand U19498 (N_19498,N_14985,N_14313);
nor U19499 (N_19499,N_15522,N_13134);
xnor U19500 (N_19500,N_12845,N_15698);
nand U19501 (N_19501,N_12313,N_15249);
or U19502 (N_19502,N_15088,N_15501);
or U19503 (N_19503,N_12034,N_14548);
nand U19504 (N_19504,N_15761,N_13257);
or U19505 (N_19505,N_12045,N_13302);
nor U19506 (N_19506,N_13358,N_15545);
or U19507 (N_19507,N_13694,N_14965);
nor U19508 (N_19508,N_13169,N_14613);
nor U19509 (N_19509,N_12459,N_14549);
nor U19510 (N_19510,N_14149,N_14865);
nand U19511 (N_19511,N_15161,N_13624);
xnor U19512 (N_19512,N_14671,N_12320);
nor U19513 (N_19513,N_12475,N_13447);
nor U19514 (N_19514,N_12000,N_12234);
and U19515 (N_19515,N_15830,N_12177);
nor U19516 (N_19516,N_12101,N_13321);
nor U19517 (N_19517,N_15451,N_12761);
nand U19518 (N_19518,N_14748,N_12671);
nand U19519 (N_19519,N_12743,N_15076);
and U19520 (N_19520,N_15677,N_12446);
nand U19521 (N_19521,N_14477,N_15519);
nor U19522 (N_19522,N_12634,N_14735);
xnor U19523 (N_19523,N_15426,N_14945);
nand U19524 (N_19524,N_14627,N_12947);
nand U19525 (N_19525,N_14066,N_14960);
and U19526 (N_19526,N_12798,N_13961);
xnor U19527 (N_19527,N_12758,N_12521);
nor U19528 (N_19528,N_14664,N_13285);
xnor U19529 (N_19529,N_12886,N_13319);
nor U19530 (N_19530,N_12577,N_13611);
xnor U19531 (N_19531,N_15094,N_14384);
nor U19532 (N_19532,N_14300,N_15363);
nand U19533 (N_19533,N_13640,N_12562);
xor U19534 (N_19534,N_14612,N_15224);
or U19535 (N_19535,N_15960,N_12932);
xnor U19536 (N_19536,N_13845,N_12585);
nand U19537 (N_19537,N_13759,N_14970);
and U19538 (N_19538,N_14024,N_14244);
nor U19539 (N_19539,N_12903,N_15726);
nand U19540 (N_19540,N_12040,N_13408);
nor U19541 (N_19541,N_13233,N_14214);
nand U19542 (N_19542,N_14914,N_15682);
nand U19543 (N_19543,N_15427,N_15859);
and U19544 (N_19544,N_14649,N_12467);
and U19545 (N_19545,N_12379,N_13592);
nand U19546 (N_19546,N_12569,N_12907);
xor U19547 (N_19547,N_13703,N_15109);
xor U19548 (N_19548,N_15789,N_12089);
xnor U19549 (N_19549,N_12882,N_14279);
nor U19550 (N_19550,N_15830,N_12374);
or U19551 (N_19551,N_13855,N_12949);
and U19552 (N_19552,N_12110,N_12907);
or U19553 (N_19553,N_15490,N_15054);
xor U19554 (N_19554,N_14145,N_12520);
xnor U19555 (N_19555,N_12695,N_14810);
or U19556 (N_19556,N_15020,N_12858);
or U19557 (N_19557,N_15837,N_12495);
nand U19558 (N_19558,N_14193,N_14242);
nand U19559 (N_19559,N_15861,N_13114);
nand U19560 (N_19560,N_12695,N_13559);
nand U19561 (N_19561,N_14919,N_14957);
xor U19562 (N_19562,N_15469,N_12780);
nand U19563 (N_19563,N_13563,N_14193);
or U19564 (N_19564,N_15598,N_12799);
and U19565 (N_19565,N_13492,N_13146);
xor U19566 (N_19566,N_13434,N_13348);
nand U19567 (N_19567,N_14115,N_13700);
nand U19568 (N_19568,N_14708,N_14083);
nand U19569 (N_19569,N_15231,N_13196);
nor U19570 (N_19570,N_14849,N_13984);
nor U19571 (N_19571,N_14233,N_13374);
xnor U19572 (N_19572,N_13313,N_15169);
and U19573 (N_19573,N_14437,N_13708);
and U19574 (N_19574,N_13533,N_12318);
or U19575 (N_19575,N_15443,N_14147);
and U19576 (N_19576,N_14084,N_12269);
xor U19577 (N_19577,N_13870,N_12972);
nor U19578 (N_19578,N_12506,N_12545);
and U19579 (N_19579,N_14945,N_15370);
xnor U19580 (N_19580,N_13553,N_13615);
nand U19581 (N_19581,N_14106,N_15617);
and U19582 (N_19582,N_15012,N_15712);
nand U19583 (N_19583,N_15477,N_14480);
nand U19584 (N_19584,N_12191,N_12608);
nand U19585 (N_19585,N_15320,N_14726);
nor U19586 (N_19586,N_13156,N_12523);
nor U19587 (N_19587,N_12221,N_14173);
nor U19588 (N_19588,N_12624,N_13062);
and U19589 (N_19589,N_13917,N_13610);
or U19590 (N_19590,N_13888,N_12805);
or U19591 (N_19591,N_14937,N_14833);
xor U19592 (N_19592,N_12665,N_14318);
nor U19593 (N_19593,N_13515,N_13368);
nor U19594 (N_19594,N_14998,N_14159);
nand U19595 (N_19595,N_15756,N_15007);
xor U19596 (N_19596,N_15651,N_14118);
nand U19597 (N_19597,N_15065,N_13482);
xor U19598 (N_19598,N_12142,N_13975);
nor U19599 (N_19599,N_14681,N_14097);
xnor U19600 (N_19600,N_12092,N_15990);
or U19601 (N_19601,N_14783,N_14966);
nand U19602 (N_19602,N_12910,N_13621);
or U19603 (N_19603,N_12919,N_13844);
xnor U19604 (N_19604,N_15531,N_14055);
xnor U19605 (N_19605,N_14930,N_13426);
nor U19606 (N_19606,N_12059,N_15302);
nand U19607 (N_19607,N_14860,N_13366);
xnor U19608 (N_19608,N_12941,N_13959);
nor U19609 (N_19609,N_14712,N_15276);
nand U19610 (N_19610,N_14079,N_12051);
nor U19611 (N_19611,N_14220,N_12493);
nor U19612 (N_19612,N_15896,N_14492);
xnor U19613 (N_19613,N_14163,N_15719);
nor U19614 (N_19614,N_12645,N_13670);
and U19615 (N_19615,N_13412,N_14325);
and U19616 (N_19616,N_15757,N_14058);
nor U19617 (N_19617,N_15618,N_14915);
xor U19618 (N_19618,N_15085,N_13701);
xor U19619 (N_19619,N_15958,N_14795);
and U19620 (N_19620,N_13686,N_15796);
or U19621 (N_19621,N_15821,N_14397);
or U19622 (N_19622,N_13918,N_13470);
nand U19623 (N_19623,N_12226,N_12714);
nor U19624 (N_19624,N_15785,N_13959);
nor U19625 (N_19625,N_15530,N_12267);
and U19626 (N_19626,N_12855,N_14968);
nand U19627 (N_19627,N_14117,N_12980);
xor U19628 (N_19628,N_14906,N_14865);
nand U19629 (N_19629,N_14442,N_15778);
and U19630 (N_19630,N_15580,N_13552);
and U19631 (N_19631,N_12777,N_12608);
nand U19632 (N_19632,N_13267,N_13447);
and U19633 (N_19633,N_12584,N_13249);
or U19634 (N_19634,N_12756,N_14540);
and U19635 (N_19635,N_12147,N_12663);
nand U19636 (N_19636,N_13930,N_15002);
xnor U19637 (N_19637,N_13558,N_14925);
and U19638 (N_19638,N_15634,N_13285);
nand U19639 (N_19639,N_14415,N_13745);
nor U19640 (N_19640,N_13481,N_15829);
or U19641 (N_19641,N_13944,N_12896);
xnor U19642 (N_19642,N_14603,N_14086);
or U19643 (N_19643,N_13502,N_14556);
or U19644 (N_19644,N_12847,N_12559);
nand U19645 (N_19645,N_15461,N_14886);
and U19646 (N_19646,N_14812,N_12186);
xor U19647 (N_19647,N_15500,N_15905);
xnor U19648 (N_19648,N_13575,N_15506);
and U19649 (N_19649,N_13211,N_15082);
nand U19650 (N_19650,N_13402,N_14802);
or U19651 (N_19651,N_14603,N_14813);
nor U19652 (N_19652,N_14524,N_15207);
or U19653 (N_19653,N_13583,N_13092);
nor U19654 (N_19654,N_13285,N_14774);
xnor U19655 (N_19655,N_13516,N_13814);
nor U19656 (N_19656,N_15606,N_14383);
and U19657 (N_19657,N_14696,N_13694);
or U19658 (N_19658,N_14785,N_14492);
and U19659 (N_19659,N_12791,N_14368);
or U19660 (N_19660,N_12757,N_14298);
nand U19661 (N_19661,N_12553,N_15779);
or U19662 (N_19662,N_13469,N_12914);
or U19663 (N_19663,N_12361,N_13561);
xor U19664 (N_19664,N_14200,N_13253);
or U19665 (N_19665,N_13119,N_12659);
xnor U19666 (N_19666,N_15838,N_15748);
nor U19667 (N_19667,N_12814,N_13870);
nor U19668 (N_19668,N_12392,N_14133);
nor U19669 (N_19669,N_13250,N_12520);
nand U19670 (N_19670,N_12861,N_13616);
nor U19671 (N_19671,N_12522,N_15127);
and U19672 (N_19672,N_13728,N_12644);
or U19673 (N_19673,N_13905,N_15206);
and U19674 (N_19674,N_12122,N_14282);
and U19675 (N_19675,N_13426,N_12791);
or U19676 (N_19676,N_13571,N_15424);
nor U19677 (N_19677,N_14626,N_15779);
xnor U19678 (N_19678,N_12067,N_14444);
or U19679 (N_19679,N_14070,N_14442);
nand U19680 (N_19680,N_15154,N_13240);
and U19681 (N_19681,N_15473,N_14899);
nand U19682 (N_19682,N_14658,N_15053);
xor U19683 (N_19683,N_15049,N_12764);
and U19684 (N_19684,N_13838,N_14447);
nor U19685 (N_19685,N_13873,N_14802);
or U19686 (N_19686,N_14888,N_15756);
xor U19687 (N_19687,N_15930,N_13586);
or U19688 (N_19688,N_14839,N_15121);
and U19689 (N_19689,N_12677,N_14026);
or U19690 (N_19690,N_12520,N_13630);
xor U19691 (N_19691,N_12241,N_14232);
or U19692 (N_19692,N_14692,N_15106);
or U19693 (N_19693,N_15094,N_14187);
nor U19694 (N_19694,N_13089,N_13663);
nor U19695 (N_19695,N_13624,N_15108);
nor U19696 (N_19696,N_14135,N_13610);
and U19697 (N_19697,N_15946,N_14943);
xor U19698 (N_19698,N_13154,N_13995);
or U19699 (N_19699,N_14847,N_13617);
xnor U19700 (N_19700,N_15190,N_15960);
nand U19701 (N_19701,N_13917,N_13074);
nor U19702 (N_19702,N_13498,N_15559);
and U19703 (N_19703,N_14648,N_12583);
or U19704 (N_19704,N_14101,N_13274);
and U19705 (N_19705,N_15539,N_12560);
nand U19706 (N_19706,N_14323,N_12428);
or U19707 (N_19707,N_15582,N_13361);
or U19708 (N_19708,N_14311,N_12438);
or U19709 (N_19709,N_12143,N_15413);
nand U19710 (N_19710,N_13950,N_12443);
xnor U19711 (N_19711,N_15984,N_15555);
and U19712 (N_19712,N_12043,N_13301);
nand U19713 (N_19713,N_15048,N_12990);
nand U19714 (N_19714,N_12777,N_12579);
or U19715 (N_19715,N_13019,N_15517);
xnor U19716 (N_19716,N_13331,N_12957);
xnor U19717 (N_19717,N_13366,N_15465);
and U19718 (N_19718,N_14313,N_14039);
xor U19719 (N_19719,N_12890,N_15537);
nor U19720 (N_19720,N_14097,N_13624);
and U19721 (N_19721,N_15977,N_15566);
xor U19722 (N_19722,N_12931,N_12184);
nand U19723 (N_19723,N_15535,N_14064);
nand U19724 (N_19724,N_13507,N_13362);
nand U19725 (N_19725,N_12939,N_12725);
nand U19726 (N_19726,N_13266,N_12778);
or U19727 (N_19727,N_15345,N_15143);
xnor U19728 (N_19728,N_15273,N_13659);
xor U19729 (N_19729,N_15398,N_14633);
or U19730 (N_19730,N_12339,N_15497);
and U19731 (N_19731,N_14203,N_13329);
nand U19732 (N_19732,N_13289,N_13820);
nand U19733 (N_19733,N_12733,N_15020);
and U19734 (N_19734,N_14692,N_15822);
or U19735 (N_19735,N_12378,N_15644);
or U19736 (N_19736,N_12981,N_12653);
nand U19737 (N_19737,N_15228,N_14746);
nand U19738 (N_19738,N_14979,N_13147);
or U19739 (N_19739,N_15289,N_14106);
or U19740 (N_19740,N_15459,N_15940);
and U19741 (N_19741,N_14088,N_13993);
xnor U19742 (N_19742,N_15854,N_14291);
or U19743 (N_19743,N_13156,N_14441);
or U19744 (N_19744,N_13175,N_14166);
or U19745 (N_19745,N_12214,N_14520);
or U19746 (N_19746,N_13700,N_14581);
xnor U19747 (N_19747,N_12994,N_12367);
xnor U19748 (N_19748,N_15571,N_14715);
nor U19749 (N_19749,N_15108,N_12768);
or U19750 (N_19750,N_15105,N_15094);
nand U19751 (N_19751,N_15285,N_15821);
nor U19752 (N_19752,N_14325,N_14585);
xnor U19753 (N_19753,N_15210,N_13442);
or U19754 (N_19754,N_12043,N_13956);
nand U19755 (N_19755,N_15736,N_15527);
and U19756 (N_19756,N_13065,N_15615);
and U19757 (N_19757,N_12772,N_15106);
nand U19758 (N_19758,N_12400,N_12004);
nand U19759 (N_19759,N_12011,N_14649);
and U19760 (N_19760,N_12667,N_14129);
and U19761 (N_19761,N_15238,N_15154);
or U19762 (N_19762,N_15193,N_15840);
and U19763 (N_19763,N_13981,N_12665);
nand U19764 (N_19764,N_13660,N_12813);
or U19765 (N_19765,N_12538,N_12729);
nor U19766 (N_19766,N_15097,N_12600);
xor U19767 (N_19767,N_13433,N_15318);
nor U19768 (N_19768,N_12113,N_14843);
xnor U19769 (N_19769,N_12621,N_15699);
xnor U19770 (N_19770,N_13777,N_13542);
nand U19771 (N_19771,N_13297,N_15168);
xnor U19772 (N_19772,N_15864,N_15831);
nand U19773 (N_19773,N_14589,N_14895);
nand U19774 (N_19774,N_13594,N_13858);
nor U19775 (N_19775,N_12962,N_14002);
nor U19776 (N_19776,N_14640,N_15242);
or U19777 (N_19777,N_14072,N_12657);
nand U19778 (N_19778,N_14179,N_13647);
nor U19779 (N_19779,N_15340,N_15597);
or U19780 (N_19780,N_15252,N_13686);
xor U19781 (N_19781,N_15289,N_15869);
xor U19782 (N_19782,N_14526,N_12730);
nand U19783 (N_19783,N_13088,N_12147);
or U19784 (N_19784,N_12740,N_15090);
or U19785 (N_19785,N_13056,N_13743);
nand U19786 (N_19786,N_12602,N_15457);
and U19787 (N_19787,N_13960,N_12547);
or U19788 (N_19788,N_13142,N_12537);
and U19789 (N_19789,N_15558,N_14997);
nor U19790 (N_19790,N_13106,N_13264);
and U19791 (N_19791,N_14341,N_13714);
and U19792 (N_19792,N_12019,N_12580);
nand U19793 (N_19793,N_14005,N_12351);
nand U19794 (N_19794,N_12192,N_15652);
or U19795 (N_19795,N_15178,N_13393);
xnor U19796 (N_19796,N_13615,N_14378);
nor U19797 (N_19797,N_15535,N_15943);
xnor U19798 (N_19798,N_12869,N_12043);
nor U19799 (N_19799,N_13450,N_15237);
xnor U19800 (N_19800,N_12005,N_13827);
nand U19801 (N_19801,N_14753,N_12218);
and U19802 (N_19802,N_15423,N_13001);
or U19803 (N_19803,N_14158,N_15882);
nor U19804 (N_19804,N_15130,N_15079);
nand U19805 (N_19805,N_12798,N_13947);
xnor U19806 (N_19806,N_12962,N_14517);
xor U19807 (N_19807,N_12409,N_14319);
xnor U19808 (N_19808,N_12383,N_14118);
nand U19809 (N_19809,N_14704,N_14178);
nand U19810 (N_19810,N_15211,N_15651);
nand U19811 (N_19811,N_13999,N_13402);
or U19812 (N_19812,N_13641,N_12810);
nor U19813 (N_19813,N_15146,N_14516);
nand U19814 (N_19814,N_14372,N_14034);
and U19815 (N_19815,N_15661,N_15250);
or U19816 (N_19816,N_14263,N_13294);
or U19817 (N_19817,N_13029,N_15783);
or U19818 (N_19818,N_14022,N_14058);
and U19819 (N_19819,N_12074,N_15058);
or U19820 (N_19820,N_14719,N_13161);
nor U19821 (N_19821,N_14767,N_15108);
nand U19822 (N_19822,N_13883,N_12346);
or U19823 (N_19823,N_15052,N_13006);
nand U19824 (N_19824,N_14428,N_13577);
or U19825 (N_19825,N_13039,N_14902);
nand U19826 (N_19826,N_15671,N_14027);
nand U19827 (N_19827,N_12536,N_13022);
or U19828 (N_19828,N_14290,N_13794);
nor U19829 (N_19829,N_15503,N_13923);
xnor U19830 (N_19830,N_15254,N_14807);
and U19831 (N_19831,N_14218,N_13793);
nor U19832 (N_19832,N_13621,N_15594);
nand U19833 (N_19833,N_15073,N_15071);
xor U19834 (N_19834,N_12793,N_13948);
or U19835 (N_19835,N_14997,N_15948);
and U19836 (N_19836,N_12801,N_12954);
or U19837 (N_19837,N_15275,N_15283);
or U19838 (N_19838,N_13990,N_14159);
and U19839 (N_19839,N_12285,N_14733);
xor U19840 (N_19840,N_13156,N_14531);
nand U19841 (N_19841,N_15489,N_14432);
nor U19842 (N_19842,N_13819,N_14264);
and U19843 (N_19843,N_12726,N_15075);
nor U19844 (N_19844,N_15531,N_13003);
xnor U19845 (N_19845,N_12644,N_13384);
xnor U19846 (N_19846,N_13020,N_15401);
and U19847 (N_19847,N_15932,N_12183);
nand U19848 (N_19848,N_13868,N_15684);
xnor U19849 (N_19849,N_13262,N_15342);
or U19850 (N_19850,N_13157,N_12770);
xor U19851 (N_19851,N_15288,N_14355);
xnor U19852 (N_19852,N_14537,N_13346);
and U19853 (N_19853,N_15091,N_14111);
or U19854 (N_19854,N_12854,N_14426);
or U19855 (N_19855,N_13040,N_12880);
nand U19856 (N_19856,N_13376,N_14125);
xnor U19857 (N_19857,N_15937,N_13385);
and U19858 (N_19858,N_14289,N_14138);
and U19859 (N_19859,N_12639,N_12783);
or U19860 (N_19860,N_14358,N_13275);
or U19861 (N_19861,N_12629,N_14780);
nor U19862 (N_19862,N_13918,N_14204);
nor U19863 (N_19863,N_13041,N_12085);
xnor U19864 (N_19864,N_12188,N_13174);
and U19865 (N_19865,N_13421,N_12833);
xor U19866 (N_19866,N_14793,N_15548);
xnor U19867 (N_19867,N_14042,N_15923);
nand U19868 (N_19868,N_12547,N_14431);
and U19869 (N_19869,N_15880,N_12622);
nand U19870 (N_19870,N_14204,N_15144);
or U19871 (N_19871,N_12649,N_12132);
nand U19872 (N_19872,N_15327,N_15818);
and U19873 (N_19873,N_14721,N_12238);
nand U19874 (N_19874,N_15808,N_14845);
xor U19875 (N_19875,N_13986,N_15995);
xor U19876 (N_19876,N_13839,N_13015);
nand U19877 (N_19877,N_14930,N_12905);
nor U19878 (N_19878,N_14327,N_13089);
or U19879 (N_19879,N_15624,N_15745);
nor U19880 (N_19880,N_12185,N_13593);
and U19881 (N_19881,N_15753,N_12923);
or U19882 (N_19882,N_14497,N_14663);
and U19883 (N_19883,N_14607,N_12435);
nand U19884 (N_19884,N_12558,N_13830);
or U19885 (N_19885,N_12068,N_13630);
or U19886 (N_19886,N_15823,N_14484);
and U19887 (N_19887,N_14265,N_13236);
xor U19888 (N_19888,N_12755,N_14127);
and U19889 (N_19889,N_12309,N_13040);
and U19890 (N_19890,N_13646,N_14076);
or U19891 (N_19891,N_15949,N_15799);
xor U19892 (N_19892,N_13946,N_12950);
and U19893 (N_19893,N_13436,N_12533);
xnor U19894 (N_19894,N_14988,N_13892);
nor U19895 (N_19895,N_12967,N_14367);
nand U19896 (N_19896,N_15344,N_13189);
or U19897 (N_19897,N_15283,N_14804);
nor U19898 (N_19898,N_13822,N_13334);
nor U19899 (N_19899,N_14352,N_15657);
xor U19900 (N_19900,N_14904,N_13444);
nor U19901 (N_19901,N_12731,N_12118);
nand U19902 (N_19902,N_13135,N_14436);
nand U19903 (N_19903,N_15339,N_12095);
and U19904 (N_19904,N_14985,N_12741);
nand U19905 (N_19905,N_13312,N_14400);
and U19906 (N_19906,N_15945,N_12447);
nand U19907 (N_19907,N_12776,N_14075);
nand U19908 (N_19908,N_12365,N_12848);
and U19909 (N_19909,N_13539,N_13150);
nand U19910 (N_19910,N_12170,N_15660);
or U19911 (N_19911,N_14083,N_14887);
nand U19912 (N_19912,N_14771,N_12023);
xor U19913 (N_19913,N_12380,N_12506);
or U19914 (N_19914,N_13240,N_12268);
nand U19915 (N_19915,N_13558,N_13684);
nor U19916 (N_19916,N_14870,N_14606);
and U19917 (N_19917,N_12404,N_12745);
and U19918 (N_19918,N_12839,N_12771);
or U19919 (N_19919,N_13928,N_12284);
or U19920 (N_19920,N_14169,N_15777);
nand U19921 (N_19921,N_12830,N_12199);
and U19922 (N_19922,N_15429,N_15548);
or U19923 (N_19923,N_12851,N_12356);
and U19924 (N_19924,N_14807,N_12229);
nand U19925 (N_19925,N_12399,N_15409);
and U19926 (N_19926,N_12120,N_15454);
and U19927 (N_19927,N_13270,N_12357);
nor U19928 (N_19928,N_12395,N_15886);
or U19929 (N_19929,N_13416,N_13177);
nand U19930 (N_19930,N_13247,N_13511);
or U19931 (N_19931,N_14647,N_12916);
or U19932 (N_19932,N_12509,N_15246);
or U19933 (N_19933,N_14450,N_15810);
xnor U19934 (N_19934,N_14216,N_15393);
nand U19935 (N_19935,N_14487,N_14243);
nor U19936 (N_19936,N_15939,N_12902);
xnor U19937 (N_19937,N_12757,N_15199);
xor U19938 (N_19938,N_13205,N_15741);
and U19939 (N_19939,N_15757,N_13455);
xnor U19940 (N_19940,N_14843,N_12141);
nand U19941 (N_19941,N_15777,N_14564);
nor U19942 (N_19942,N_14855,N_13145);
and U19943 (N_19943,N_12648,N_14733);
xnor U19944 (N_19944,N_13454,N_13487);
or U19945 (N_19945,N_12268,N_13632);
and U19946 (N_19946,N_14819,N_13093);
or U19947 (N_19947,N_12094,N_12616);
and U19948 (N_19948,N_14310,N_12856);
nand U19949 (N_19949,N_12079,N_13050);
or U19950 (N_19950,N_14844,N_14655);
nand U19951 (N_19951,N_14087,N_15877);
and U19952 (N_19952,N_13817,N_12420);
nand U19953 (N_19953,N_15332,N_12008);
xor U19954 (N_19954,N_12057,N_12330);
and U19955 (N_19955,N_15177,N_14002);
nor U19956 (N_19956,N_14257,N_12519);
nor U19957 (N_19957,N_13440,N_12526);
and U19958 (N_19958,N_15620,N_14975);
and U19959 (N_19959,N_12076,N_13366);
nor U19960 (N_19960,N_13466,N_14295);
xnor U19961 (N_19961,N_14401,N_13261);
or U19962 (N_19962,N_12919,N_15353);
xor U19963 (N_19963,N_14096,N_12608);
nand U19964 (N_19964,N_13473,N_12016);
or U19965 (N_19965,N_13677,N_13134);
or U19966 (N_19966,N_12058,N_15510);
and U19967 (N_19967,N_13155,N_12674);
nor U19968 (N_19968,N_13189,N_12190);
or U19969 (N_19969,N_13448,N_12060);
nand U19970 (N_19970,N_13949,N_14865);
xor U19971 (N_19971,N_14638,N_12357);
xnor U19972 (N_19972,N_13415,N_15056);
nor U19973 (N_19973,N_13281,N_12624);
xnor U19974 (N_19974,N_13755,N_15721);
and U19975 (N_19975,N_13304,N_15230);
xnor U19976 (N_19976,N_14287,N_15173);
or U19977 (N_19977,N_13250,N_13775);
and U19978 (N_19978,N_12104,N_14492);
nand U19979 (N_19979,N_13053,N_14088);
and U19980 (N_19980,N_12580,N_13814);
xnor U19981 (N_19981,N_13148,N_14859);
or U19982 (N_19982,N_15972,N_12085);
xnor U19983 (N_19983,N_12757,N_12685);
or U19984 (N_19984,N_14593,N_14535);
nand U19985 (N_19985,N_13390,N_12634);
or U19986 (N_19986,N_14637,N_13229);
xor U19987 (N_19987,N_13031,N_15400);
and U19988 (N_19988,N_12874,N_15392);
and U19989 (N_19989,N_13692,N_12907);
and U19990 (N_19990,N_14399,N_13623);
or U19991 (N_19991,N_12432,N_15790);
xnor U19992 (N_19992,N_13815,N_15069);
and U19993 (N_19993,N_14957,N_15417);
or U19994 (N_19994,N_15336,N_15456);
nand U19995 (N_19995,N_15521,N_15471);
nor U19996 (N_19996,N_13421,N_13130);
and U19997 (N_19997,N_12469,N_15557);
and U19998 (N_19998,N_12464,N_15075);
xnor U19999 (N_19999,N_13069,N_14596);
and UO_0 (O_0,N_16298,N_17402);
nor UO_1 (O_1,N_17333,N_16514);
nand UO_2 (O_2,N_19232,N_18132);
nand UO_3 (O_3,N_19903,N_18442);
xnor UO_4 (O_4,N_17991,N_16247);
or UO_5 (O_5,N_18651,N_18818);
nand UO_6 (O_6,N_18860,N_18647);
nor UO_7 (O_7,N_19510,N_16627);
nor UO_8 (O_8,N_18584,N_19220);
and UO_9 (O_9,N_16273,N_16338);
or UO_10 (O_10,N_19503,N_18317);
nor UO_11 (O_11,N_16733,N_19476);
or UO_12 (O_12,N_17646,N_18744);
or UO_13 (O_13,N_19245,N_19109);
xnor UO_14 (O_14,N_18617,N_16941);
or UO_15 (O_15,N_16234,N_16766);
nor UO_16 (O_16,N_16208,N_17808);
or UO_17 (O_17,N_18940,N_19635);
and UO_18 (O_18,N_16928,N_17972);
nor UO_19 (O_19,N_18875,N_17967);
and UO_20 (O_20,N_16626,N_17424);
or UO_21 (O_21,N_16493,N_19872);
nor UO_22 (O_22,N_16566,N_18152);
nor UO_23 (O_23,N_18861,N_19848);
or UO_24 (O_24,N_16997,N_18887);
or UO_25 (O_25,N_16448,N_16686);
nor UO_26 (O_26,N_19382,N_18610);
and UO_27 (O_27,N_19904,N_18440);
or UO_28 (O_28,N_17412,N_17536);
nand UO_29 (O_29,N_16707,N_18947);
nand UO_30 (O_30,N_16994,N_18948);
xnor UO_31 (O_31,N_17057,N_19969);
xor UO_32 (O_32,N_17896,N_18742);
nor UO_33 (O_33,N_19357,N_19972);
xnor UO_34 (O_34,N_19808,N_17533);
or UO_35 (O_35,N_19280,N_18984);
or UO_36 (O_36,N_19582,N_16782);
nand UO_37 (O_37,N_19707,N_18364);
or UO_38 (O_38,N_17210,N_17769);
nand UO_39 (O_39,N_18561,N_17734);
nand UO_40 (O_40,N_19802,N_17188);
nand UO_41 (O_41,N_16584,N_16717);
nand UO_42 (O_42,N_17226,N_18746);
nand UO_43 (O_43,N_16126,N_18320);
or UO_44 (O_44,N_18527,N_18218);
or UO_45 (O_45,N_18923,N_16718);
xor UO_46 (O_46,N_19636,N_18715);
or UO_47 (O_47,N_17785,N_19266);
nor UO_48 (O_48,N_16492,N_17451);
and UO_49 (O_49,N_18542,N_17575);
or UO_50 (O_50,N_16039,N_16947);
or UO_51 (O_51,N_19423,N_19682);
xor UO_52 (O_52,N_16855,N_18662);
xnor UO_53 (O_53,N_16524,N_16094);
nand UO_54 (O_54,N_16155,N_16025);
xor UO_55 (O_55,N_16968,N_16682);
xor UO_56 (O_56,N_18119,N_16802);
and UO_57 (O_57,N_18820,N_16370);
nand UO_58 (O_58,N_19076,N_18750);
xor UO_59 (O_59,N_16114,N_16328);
or UO_60 (O_60,N_16647,N_19666);
nand UO_61 (O_61,N_19161,N_17583);
and UO_62 (O_62,N_17483,N_16895);
and UO_63 (O_63,N_17731,N_17974);
and UO_64 (O_64,N_19826,N_18104);
nor UO_65 (O_65,N_18234,N_19955);
and UO_66 (O_66,N_17288,N_16249);
xnor UO_67 (O_67,N_18379,N_19966);
and UO_68 (O_68,N_18450,N_19933);
and UO_69 (O_69,N_18386,N_17134);
xor UO_70 (O_70,N_19971,N_17678);
nand UO_71 (O_71,N_19104,N_18654);
xnor UO_72 (O_72,N_16981,N_19814);
xor UO_73 (O_73,N_18675,N_18613);
xor UO_74 (O_74,N_19304,N_17624);
xor UO_75 (O_75,N_17085,N_17743);
nor UO_76 (O_76,N_18811,N_16023);
nand UO_77 (O_77,N_17309,N_17863);
and UO_78 (O_78,N_19347,N_18928);
nand UO_79 (O_79,N_17066,N_16455);
and UO_80 (O_80,N_16656,N_19276);
nor UO_81 (O_81,N_17529,N_17736);
nand UO_82 (O_82,N_18391,N_17756);
and UO_83 (O_83,N_18376,N_16055);
nand UO_84 (O_84,N_19586,N_16013);
nand UO_85 (O_85,N_19996,N_17659);
and UO_86 (O_86,N_18255,N_17366);
or UO_87 (O_87,N_18232,N_16471);
nor UO_88 (O_88,N_16194,N_19163);
nand UO_89 (O_89,N_17651,N_17006);
or UO_90 (O_90,N_17029,N_17056);
or UO_91 (O_91,N_19370,N_16794);
or UO_92 (O_92,N_17881,N_16784);
and UO_93 (O_93,N_16589,N_18288);
nor UO_94 (O_94,N_19087,N_17822);
and UO_95 (O_95,N_17071,N_16893);
and UO_96 (O_96,N_17194,N_19239);
nand UO_97 (O_97,N_19345,N_16887);
nor UO_98 (O_98,N_18127,N_16595);
xnor UO_99 (O_99,N_19138,N_17013);
and UO_100 (O_100,N_19354,N_19557);
nand UO_101 (O_101,N_16363,N_17541);
and UO_102 (O_102,N_16268,N_18186);
nand UO_103 (O_103,N_18692,N_19467);
nor UO_104 (O_104,N_18471,N_18991);
nand UO_105 (O_105,N_18595,N_18738);
nand UO_106 (O_106,N_17389,N_18642);
nor UO_107 (O_107,N_16381,N_18992);
nor UO_108 (O_108,N_17707,N_19925);
nand UO_109 (O_109,N_17298,N_17216);
nand UO_110 (O_110,N_17561,N_18373);
and UO_111 (O_111,N_16619,N_17538);
nand UO_112 (O_112,N_19386,N_19287);
or UO_113 (O_113,N_18029,N_19600);
xor UO_114 (O_114,N_17098,N_16164);
xnor UO_115 (O_115,N_19783,N_17574);
nand UO_116 (O_116,N_17203,N_17213);
or UO_117 (O_117,N_16266,N_16553);
or UO_118 (O_118,N_17305,N_19900);
or UO_119 (O_119,N_17694,N_18352);
nand UO_120 (O_120,N_19615,N_17016);
nor UO_121 (O_121,N_18405,N_17160);
or UO_122 (O_122,N_17643,N_18925);
nor UO_123 (O_123,N_17344,N_18888);
xor UO_124 (O_124,N_18694,N_17207);
nand UO_125 (O_125,N_16853,N_16953);
or UO_126 (O_126,N_17695,N_16144);
nor UO_127 (O_127,N_19927,N_18351);
xnor UO_128 (O_128,N_19218,N_18519);
nand UO_129 (O_129,N_17633,N_19241);
and UO_130 (O_130,N_16478,N_18849);
nor UO_131 (O_131,N_19203,N_19738);
nor UO_132 (O_132,N_17944,N_18125);
nor UO_133 (O_133,N_19319,N_17360);
or UO_134 (O_134,N_16759,N_18688);
nor UO_135 (O_135,N_18775,N_16675);
nand UO_136 (O_136,N_19843,N_16007);
nand UO_137 (O_137,N_17973,N_19639);
xnor UO_138 (O_138,N_19272,N_16916);
nor UO_139 (O_139,N_17457,N_18553);
nand UO_140 (O_140,N_18250,N_17843);
nor UO_141 (O_141,N_16068,N_19834);
or UO_142 (O_142,N_17848,N_18074);
xor UO_143 (O_143,N_16623,N_19924);
nand UO_144 (O_144,N_16557,N_16588);
or UO_145 (O_145,N_17742,N_18087);
nor UO_146 (O_146,N_19856,N_16952);
or UO_147 (O_147,N_19111,N_18392);
nor UO_148 (O_148,N_17327,N_18309);
nor UO_149 (O_149,N_19518,N_16245);
nor UO_150 (O_150,N_19871,N_19351);
or UO_151 (O_151,N_19727,N_16629);
nand UO_152 (O_152,N_19146,N_17631);
or UO_153 (O_153,N_19982,N_18235);
xor UO_154 (O_154,N_16187,N_17928);
nor UO_155 (O_155,N_19458,N_17115);
or UO_156 (O_156,N_16520,N_17338);
or UO_157 (O_157,N_17431,N_17872);
or UO_158 (O_158,N_16350,N_19751);
xnor UO_159 (O_159,N_16667,N_17139);
xor UO_160 (O_160,N_18963,N_16475);
xor UO_161 (O_161,N_16958,N_16533);
and UO_162 (O_162,N_16185,N_18375);
nand UO_163 (O_163,N_19095,N_18518);
nor UO_164 (O_164,N_17004,N_19836);
or UO_165 (O_165,N_19916,N_17386);
and UO_166 (O_166,N_19571,N_17480);
and UO_167 (O_167,N_18431,N_17603);
or UO_168 (O_168,N_19005,N_18753);
xor UO_169 (O_169,N_18945,N_19689);
or UO_170 (O_170,N_16665,N_19711);
or UO_171 (O_171,N_18059,N_19951);
nor UO_172 (O_172,N_16391,N_19516);
and UO_173 (O_173,N_19793,N_16490);
or UO_174 (O_174,N_19238,N_17452);
and UO_175 (O_175,N_16909,N_17051);
nor UO_176 (O_176,N_16112,N_18611);
and UO_177 (O_177,N_18318,N_18190);
and UO_178 (O_178,N_17238,N_18578);
nor UO_179 (O_179,N_17901,N_19494);
or UO_180 (O_180,N_18293,N_17249);
or UO_181 (O_181,N_16380,N_19395);
xnor UO_182 (O_182,N_16318,N_19781);
nand UO_183 (O_183,N_19658,N_16424);
xnor UO_184 (O_184,N_19380,N_18955);
xor UO_185 (O_185,N_18745,N_16955);
xor UO_186 (O_186,N_17163,N_18917);
and UO_187 (O_187,N_19375,N_19741);
or UO_188 (O_188,N_16767,N_19497);
and UO_189 (O_189,N_19544,N_18126);
and UO_190 (O_190,N_17754,N_17543);
nor UO_191 (O_191,N_17450,N_19874);
nand UO_192 (O_192,N_18428,N_16084);
nor UO_193 (O_193,N_16119,N_17995);
nor UO_194 (O_194,N_16302,N_17670);
or UO_195 (O_195,N_16749,N_17415);
and UO_196 (O_196,N_18426,N_17351);
nor UO_197 (O_197,N_19909,N_19660);
nand UO_198 (O_198,N_18652,N_19122);
nand UO_199 (O_199,N_18129,N_16697);
nand UO_200 (O_200,N_17579,N_19767);
and UO_201 (O_201,N_17816,N_18106);
or UO_202 (O_202,N_17177,N_19963);
nor UO_203 (O_203,N_18280,N_19393);
xnor UO_204 (O_204,N_16961,N_19500);
and UO_205 (O_205,N_17234,N_18377);
nand UO_206 (O_206,N_19022,N_19726);
and UO_207 (O_207,N_17825,N_16790);
or UO_208 (O_208,N_17141,N_19399);
xnor UO_209 (O_209,N_18490,N_17231);
nand UO_210 (O_210,N_18000,N_18404);
and UO_211 (O_211,N_19278,N_18821);
nor UO_212 (O_212,N_16724,N_17322);
xnor UO_213 (O_213,N_19961,N_16314);
nor UO_214 (O_214,N_17729,N_16622);
and UO_215 (O_215,N_17151,N_18165);
xnor UO_216 (O_216,N_18761,N_18025);
nor UO_217 (O_217,N_16414,N_17965);
nor UO_218 (O_218,N_19021,N_19550);
nor UO_219 (O_219,N_17927,N_18054);
nand UO_220 (O_220,N_16573,N_18649);
nor UO_221 (O_221,N_19542,N_19250);
nor UO_222 (O_222,N_16931,N_19353);
nand UO_223 (O_223,N_17737,N_16356);
nand UO_224 (O_224,N_19329,N_19774);
xnor UO_225 (O_225,N_17688,N_17024);
and UO_226 (O_226,N_19739,N_17073);
or UO_227 (O_227,N_19130,N_18965);
nor UO_228 (O_228,N_18813,N_16906);
xor UO_229 (O_229,N_19643,N_16601);
and UO_230 (O_230,N_17684,N_16347);
xor UO_231 (O_231,N_16293,N_19166);
xor UO_232 (O_232,N_18409,N_19405);
xnor UO_233 (O_233,N_19030,N_17011);
or UO_234 (O_234,N_19192,N_16924);
or UO_235 (O_235,N_18683,N_16648);
xnor UO_236 (O_236,N_16546,N_19686);
or UO_237 (O_237,N_19536,N_16699);
xnor UO_238 (O_238,N_16215,N_17943);
xnor UO_239 (O_239,N_19528,N_19387);
and UO_240 (O_240,N_18046,N_18912);
and UO_241 (O_241,N_18339,N_19140);
xnor UO_242 (O_242,N_16828,N_18277);
nor UO_243 (O_243,N_17094,N_18449);
nand UO_244 (O_244,N_16516,N_19057);
xor UO_245 (O_245,N_19162,N_17542);
nor UO_246 (O_246,N_16419,N_16105);
nand UO_247 (O_247,N_17985,N_16526);
and UO_248 (O_248,N_18764,N_16681);
or UO_249 (O_249,N_19367,N_17661);
nand UO_250 (O_250,N_16317,N_19705);
or UO_251 (O_251,N_18146,N_19374);
and UO_252 (O_252,N_16894,N_18222);
and UO_253 (O_253,N_18329,N_19850);
nand UO_254 (O_254,N_19746,N_18008);
nor UO_255 (O_255,N_19828,N_19522);
or UO_256 (O_256,N_17381,N_17993);
nand UO_257 (O_257,N_18982,N_19930);
or UO_258 (O_258,N_17597,N_18458);
or UO_259 (O_259,N_16040,N_17107);
nor UO_260 (O_260,N_16725,N_19053);
or UO_261 (O_261,N_17500,N_17470);
nor UO_262 (O_262,N_16115,N_17776);
nand UO_263 (O_263,N_16796,N_16509);
nand UO_264 (O_264,N_16214,N_19548);
xnor UO_265 (O_265,N_18278,N_19837);
nand UO_266 (O_266,N_16436,N_16210);
xnor UO_267 (O_267,N_17393,N_17607);
nand UO_268 (O_268,N_16570,N_19919);
or UO_269 (O_269,N_19532,N_18242);
nor UO_270 (O_270,N_18804,N_16218);
and UO_271 (O_271,N_18942,N_19419);
or UO_272 (O_272,N_19784,N_19125);
and UO_273 (O_273,N_16616,N_16104);
and UO_274 (O_274,N_19194,N_19785);
and UO_275 (O_275,N_17961,N_19009);
or UO_276 (O_276,N_17002,N_17026);
nand UO_277 (O_277,N_17311,N_17491);
nand UO_278 (O_278,N_17889,N_16653);
or UO_279 (O_279,N_17175,N_16045);
xnor UO_280 (O_280,N_19569,N_16081);
xnor UO_281 (O_281,N_17990,N_19806);
nand UO_282 (O_282,N_16163,N_17458);
and UO_283 (O_283,N_16299,N_18871);
and UO_284 (O_284,N_18850,N_19803);
or UO_285 (O_285,N_18932,N_19294);
or UO_286 (O_286,N_18814,N_19431);
nand UO_287 (O_287,N_17998,N_19152);
xnor UO_288 (O_288,N_16713,N_16945);
nand UO_289 (O_289,N_17448,N_19385);
nand UO_290 (O_290,N_16392,N_16954);
and UO_291 (O_291,N_19948,N_17949);
or UO_292 (O_292,N_18084,N_18673);
and UO_293 (O_293,N_18239,N_19846);
nor UO_294 (O_294,N_18279,N_17193);
or UO_295 (O_295,N_16563,N_17113);
xnor UO_296 (O_296,N_19936,N_16960);
or UO_297 (O_297,N_17099,N_19149);
and UO_298 (O_298,N_19409,N_18953);
nand UO_299 (O_299,N_16582,N_18201);
or UO_300 (O_300,N_18549,N_18975);
nand UO_301 (O_301,N_19195,N_17042);
or UO_302 (O_302,N_17317,N_17110);
nand UO_303 (O_303,N_17104,N_18225);
xnor UO_304 (O_304,N_17941,N_16495);
xor UO_305 (O_305,N_19570,N_17955);
nor UO_306 (O_306,N_17429,N_19379);
nand UO_307 (O_307,N_19762,N_16680);
or UO_308 (O_308,N_18107,N_18809);
nor UO_309 (O_309,N_17422,N_18196);
xnor UO_310 (O_310,N_17053,N_19403);
nand UO_311 (O_311,N_17558,N_16452);
or UO_312 (O_312,N_19868,N_17609);
nand UO_313 (O_313,N_17198,N_18946);
xor UO_314 (O_314,N_18093,N_16548);
and UO_315 (O_315,N_17208,N_16592);
xor UO_316 (O_316,N_17531,N_19350);
nand UO_317 (O_317,N_18643,N_16650);
nand UO_318 (O_318,N_16948,N_17138);
xnor UO_319 (O_319,N_19451,N_16216);
or UO_320 (O_320,N_18677,N_16240);
nor UO_321 (O_321,N_16572,N_16715);
or UO_322 (O_322,N_16578,N_16684);
nor UO_323 (O_323,N_18302,N_16474);
or UO_324 (O_324,N_18915,N_18934);
or UO_325 (O_325,N_17159,N_19970);
nor UO_326 (O_326,N_17873,N_19112);
and UO_327 (O_327,N_17930,N_18602);
or UO_328 (O_328,N_18728,N_16118);
nand UO_329 (O_329,N_19134,N_16064);
or UO_330 (O_330,N_18039,N_18052);
or UO_331 (O_331,N_17576,N_18212);
nand UO_332 (O_332,N_19251,N_18112);
nor UO_333 (O_333,N_18395,N_19240);
and UO_334 (O_334,N_19067,N_19401);
xnor UO_335 (O_335,N_16951,N_16556);
nand UO_336 (O_336,N_16366,N_18701);
nor UO_337 (O_337,N_19277,N_17751);
or UO_338 (O_338,N_18921,N_18719);
nor UO_339 (O_339,N_19252,N_17068);
or UO_340 (O_340,N_19747,N_18272);
nand UO_341 (O_341,N_16295,N_17384);
or UO_342 (O_342,N_17503,N_16037);
and UO_343 (O_343,N_16833,N_17489);
and UO_344 (O_344,N_19444,N_19014);
and UO_345 (O_345,N_18240,N_18733);
and UO_346 (O_346,N_19941,N_18920);
nand UO_347 (O_347,N_17619,N_19857);
and UO_348 (O_348,N_19681,N_16923);
xnor UO_349 (O_349,N_17766,N_16538);
nor UO_350 (O_350,N_19072,N_17587);
and UO_351 (O_351,N_16649,N_16705);
or UO_352 (O_352,N_16652,N_18937);
xor UO_353 (O_353,N_16165,N_19421);
nor UO_354 (O_354,N_19299,N_17981);
nor UO_355 (O_355,N_17664,N_18485);
and UO_356 (O_356,N_19480,N_17919);
nor UO_357 (O_357,N_16036,N_16985);
or UO_358 (O_358,N_18755,N_19263);
or UO_359 (O_359,N_19511,N_19884);
or UO_360 (O_360,N_17586,N_19359);
nand UO_361 (O_361,N_16322,N_17813);
nor UO_362 (O_362,N_17246,N_17388);
xnor UO_363 (O_363,N_16464,N_17701);
xor UO_364 (O_364,N_17720,N_17711);
and UO_365 (O_365,N_17436,N_18935);
nand UO_366 (O_366,N_19291,N_17329);
nor UO_367 (O_367,N_18273,N_19206);
and UO_368 (O_368,N_17553,N_16330);
or UO_369 (O_369,N_17969,N_18384);
or UO_370 (O_370,N_16227,N_16691);
or UO_371 (O_371,N_18962,N_18062);
nand UO_372 (O_372,N_16515,N_17650);
xnor UO_373 (O_373,N_18640,N_18723);
or UO_374 (O_374,N_18762,N_19674);
or UO_375 (O_375,N_16237,N_17685);
and UO_376 (O_376,N_16624,N_16761);
nand UO_377 (O_377,N_19113,N_16964);
and UO_378 (O_378,N_17035,N_19179);
nor UO_379 (O_379,N_18015,N_17025);
nand UO_380 (O_380,N_17798,N_19876);
and UO_381 (O_381,N_17601,N_18170);
or UO_382 (O_382,N_16312,N_18178);
xor UO_383 (O_383,N_17263,N_17183);
nand UO_384 (O_384,N_16445,N_19025);
and UO_385 (O_385,N_17088,N_19913);
and UO_386 (O_386,N_16438,N_16096);
and UO_387 (O_387,N_16612,N_19957);
nand UO_388 (O_388,N_18536,N_16884);
nor UO_389 (O_389,N_17636,N_19816);
or UO_390 (O_390,N_16000,N_16217);
nand UO_391 (O_391,N_18388,N_19036);
and UO_392 (O_392,N_16087,N_19144);
xor UO_393 (O_393,N_17276,N_18687);
nand UO_394 (O_394,N_19530,N_18055);
xnor UO_395 (O_395,N_19224,N_18492);
xor UO_396 (O_396,N_18362,N_16325);
and UO_397 (O_397,N_17572,N_19468);
xnor UO_398 (O_398,N_19879,N_18774);
nand UO_399 (O_399,N_17773,N_16260);
nor UO_400 (O_400,N_16944,N_17325);
nand UO_401 (O_401,N_16617,N_19160);
xor UO_402 (O_402,N_19665,N_18626);
xor UO_403 (O_403,N_18835,N_18822);
and UO_404 (O_404,N_17888,N_18704);
nand UO_405 (O_405,N_18416,N_16848);
or UO_406 (O_406,N_19519,N_16869);
and UO_407 (O_407,N_17794,N_18073);
nor UO_408 (O_408,N_17672,N_18780);
nor UO_409 (O_409,N_17842,N_16992);
nor UO_410 (O_410,N_16810,N_18324);
or UO_411 (O_411,N_17080,N_19221);
or UO_412 (O_412,N_17780,N_19268);
nor UO_413 (O_413,N_19855,N_18569);
or UO_414 (O_414,N_17931,N_19034);
and UO_415 (O_415,N_16145,N_17815);
xnor UO_416 (O_416,N_16028,N_18686);
and UO_417 (O_417,N_18631,N_16743);
and UO_418 (O_418,N_16372,N_18070);
and UO_419 (O_419,N_16897,N_19987);
or UO_420 (O_420,N_17462,N_19302);
or UO_421 (O_421,N_16321,N_17341);
nor UO_422 (O_422,N_18368,N_17730);
nand UO_423 (O_423,N_17850,N_17865);
nand UO_424 (O_424,N_16676,N_17790);
nand UO_425 (O_425,N_18144,N_16800);
xor UO_426 (O_426,N_19653,N_17937);
or UO_427 (O_427,N_18724,N_19605);
and UO_428 (O_428,N_18973,N_19820);
nor UO_429 (O_429,N_19490,N_17963);
nor UO_430 (O_430,N_16387,N_19186);
or UO_431 (O_431,N_17120,N_19853);
or UO_432 (O_432,N_17566,N_17912);
xor UO_433 (O_433,N_18333,N_19776);
nor UO_434 (O_434,N_16877,N_18354);
nor UO_435 (O_435,N_19967,N_17656);
or UO_436 (O_436,N_18434,N_16426);
nand UO_437 (O_437,N_18505,N_17005);
nor UO_438 (O_438,N_17019,N_18323);
xnor UO_439 (O_439,N_16002,N_19466);
or UO_440 (O_440,N_19981,N_18035);
nor UO_441 (O_441,N_19844,N_17675);
and UO_442 (O_442,N_17611,N_16341);
and UO_443 (O_443,N_17408,N_16521);
and UO_444 (O_444,N_16517,N_19701);
nor UO_445 (O_445,N_18024,N_18653);
nor UO_446 (O_446,N_16175,N_18343);
nor UO_447 (O_447,N_18616,N_19552);
or UO_448 (O_448,N_19181,N_17867);
and UO_449 (O_449,N_16903,N_18964);
nor UO_450 (O_450,N_16890,N_19825);
nor UO_451 (O_451,N_18769,N_18619);
nor UO_452 (O_452,N_16362,N_17443);
or UO_453 (O_453,N_17326,N_16080);
nor UO_454 (O_454,N_16267,N_19811);
and UO_455 (O_455,N_17710,N_18766);
or UO_456 (O_456,N_16501,N_18398);
or UO_457 (O_457,N_17047,N_19603);
xor UO_458 (O_458,N_19566,N_16460);
and UO_459 (O_459,N_19920,N_17271);
and UO_460 (O_460,N_19995,N_19633);
nand UO_461 (O_461,N_16644,N_17811);
xor UO_462 (O_462,N_19190,N_17287);
nand UO_463 (O_463,N_19756,N_19398);
nor UO_464 (O_464,N_16729,N_16611);
xnor UO_465 (O_465,N_19817,N_17250);
nor UO_466 (O_466,N_19343,N_17778);
nor UO_467 (O_467,N_17713,N_19108);
or UO_468 (O_468,N_16930,N_16326);
and UO_469 (O_469,N_17223,N_19895);
xor UO_470 (O_470,N_16631,N_17939);
and UO_471 (O_471,N_16360,N_18028);
xnor UO_472 (O_472,N_19943,N_18105);
xnor UO_473 (O_473,N_17083,N_16798);
nor UO_474 (O_474,N_19614,N_16870);
or UO_475 (O_475,N_19634,N_17373);
nand UO_476 (O_476,N_17078,N_17994);
nor UO_477 (O_477,N_19048,N_17602);
nor UO_478 (O_478,N_18496,N_18633);
nand UO_479 (O_479,N_16821,N_18552);
nand UO_480 (O_480,N_16815,N_19117);
or UO_481 (O_481,N_18003,N_19769);
and UO_482 (O_482,N_19944,N_16220);
nand UO_483 (O_483,N_16026,N_18756);
nor UO_484 (O_484,N_19568,N_16562);
and UO_485 (O_485,N_16433,N_18990);
xnor UO_486 (O_486,N_17511,N_18729);
nand UO_487 (O_487,N_18331,N_17127);
nand UO_488 (O_488,N_19988,N_16465);
xor UO_489 (O_489,N_19651,N_19680);
or UO_490 (O_490,N_16505,N_19471);
and UO_491 (O_491,N_17178,N_16001);
and UO_492 (O_492,N_16694,N_18475);
xnor UO_493 (O_493,N_17340,N_16343);
and UO_494 (O_494,N_16176,N_18638);
or UO_495 (O_495,N_18164,N_19644);
or UO_496 (O_496,N_19952,N_18883);
or UO_497 (O_497,N_18316,N_19199);
xor UO_498 (O_498,N_18983,N_19139);
xor UO_499 (O_499,N_18441,N_19407);
nor UO_500 (O_500,N_17274,N_18791);
or UO_501 (O_501,N_16528,N_17644);
nand UO_502 (O_502,N_19050,N_18038);
nor UO_503 (O_503,N_19647,N_18538);
nand UO_504 (O_504,N_19587,N_18710);
and UO_505 (O_505,N_19243,N_16450);
nor UO_506 (O_506,N_18205,N_18369);
nand UO_507 (O_507,N_16447,N_16728);
xor UO_508 (O_508,N_18177,N_17032);
nor UO_509 (O_509,N_17758,N_18844);
or UO_510 (O_510,N_19003,N_16639);
nor UO_511 (O_511,N_16281,N_19325);
or UO_512 (O_512,N_16287,N_16744);
xnor UO_513 (O_513,N_18124,N_19410);
nand UO_514 (O_514,N_16136,N_18670);
xor UO_515 (O_515,N_16597,N_17864);
nand UO_516 (O_516,N_16052,N_16807);
nor UO_517 (O_517,N_18418,N_16873);
xnor UO_518 (O_518,N_16050,N_16915);
xnor UO_519 (O_519,N_16383,N_17236);
or UO_520 (O_520,N_16120,N_18944);
nor UO_521 (O_521,N_17819,N_18266);
xor UO_522 (O_522,N_19931,N_17281);
or UO_523 (O_523,N_17495,N_18005);
and UO_524 (O_524,N_17996,N_17279);
nand UO_525 (O_525,N_19863,N_19284);
nand UO_526 (O_526,N_19051,N_18466);
xor UO_527 (O_527,N_17866,N_17709);
nor UO_528 (O_528,N_17782,N_17404);
and UO_529 (O_529,N_18787,N_16486);
nand UO_530 (O_530,N_19156,N_18090);
xnor UO_531 (O_531,N_16522,N_16880);
or UO_532 (O_532,N_18862,N_19649);
and UO_533 (O_533,N_18727,N_19324);
nand UO_534 (O_534,N_16043,N_19870);
xnor UO_535 (O_535,N_18634,N_17296);
xnor UO_536 (O_536,N_17655,N_16861);
or UO_537 (O_537,N_19188,N_17008);
or UO_538 (O_538,N_17674,N_18906);
nand UO_539 (O_539,N_17526,N_18913);
and UO_540 (O_540,N_18497,N_16334);
and UO_541 (O_541,N_17206,N_19608);
xor UO_542 (O_542,N_17932,N_16283);
or UO_543 (O_543,N_18641,N_17613);
nor UO_544 (O_544,N_19435,N_16090);
xnor UO_545 (O_545,N_16142,N_17810);
nor UO_546 (O_546,N_18001,N_17145);
xnor UO_547 (O_547,N_19133,N_17109);
and UO_548 (O_548,N_16342,N_18604);
nor UO_549 (O_549,N_16730,N_19829);
nor UO_550 (O_550,N_16071,N_16732);
nor UO_551 (O_551,N_17804,N_18315);
and UO_552 (O_552,N_18183,N_18889);
nand UO_553 (O_553,N_16757,N_19154);
nand UO_554 (O_554,N_18572,N_16201);
nor UO_555 (O_555,N_18993,N_19699);
or UO_556 (O_556,N_19724,N_18770);
or UO_557 (O_557,N_17394,N_19233);
or UO_558 (O_558,N_18420,N_17934);
and UO_559 (O_559,N_16021,N_19599);
nand UO_560 (O_560,N_19178,N_16238);
nor UO_561 (O_561,N_19907,N_19706);
xnor UO_562 (O_562,N_17922,N_17312);
nor UO_563 (O_563,N_17308,N_19013);
xor UO_564 (O_564,N_16444,N_18749);
nand UO_565 (O_565,N_16172,N_19672);
xnor UO_566 (O_566,N_18174,N_16024);
or UO_567 (O_567,N_17258,N_17831);
or UO_568 (O_568,N_16329,N_17473);
and UO_569 (O_569,N_17925,N_18080);
xor UO_570 (O_570,N_17984,N_19368);
and UO_571 (O_571,N_17131,N_18978);
xor UO_572 (O_572,N_19237,N_18743);
xor UO_573 (O_573,N_19775,N_19765);
or UO_574 (O_574,N_17708,N_17809);
and UO_575 (O_575,N_19159,N_16769);
nand UO_576 (O_576,N_19400,N_17744);
nor UO_577 (O_577,N_19486,N_17803);
and UO_578 (O_578,N_18195,N_19612);
or UO_579 (O_579,N_16716,N_19759);
xor UO_580 (O_580,N_17852,N_19906);
nand UO_581 (O_581,N_17723,N_18043);
or UO_582 (O_582,N_16324,N_18892);
xnor UO_583 (O_583,N_17041,N_19383);
and UO_584 (O_584,N_17343,N_19959);
nand UO_585 (O_585,N_17580,N_17801);
and UO_586 (O_586,N_17764,N_18436);
or UO_587 (O_587,N_18589,N_16259);
nand UO_588 (O_588,N_16224,N_16345);
and UO_589 (O_589,N_17001,N_16147);
nor UO_590 (O_590,N_19833,N_19645);
nor UO_591 (O_591,N_18899,N_19667);
or UO_592 (O_592,N_18128,N_19892);
or UO_593 (O_593,N_17383,N_16735);
xor UO_594 (O_594,N_17826,N_18380);
xor UO_595 (O_595,N_19521,N_16411);
nand UO_596 (O_596,N_19505,N_16469);
nor UO_597 (O_597,N_18263,N_19623);
nand UO_598 (O_598,N_19800,N_17833);
xnor UO_599 (O_599,N_17445,N_19443);
and UO_600 (O_600,N_18712,N_16154);
or UO_601 (O_601,N_18460,N_18045);
and UO_602 (O_602,N_18854,N_18976);
nand UO_603 (O_603,N_19052,N_19056);
nor UO_604 (O_604,N_18481,N_17721);
and UO_605 (O_605,N_17046,N_18163);
nor UO_606 (O_606,N_18310,N_19734);
or UO_607 (O_607,N_17680,N_16559);
and UO_608 (O_608,N_19523,N_17446);
and UO_609 (O_609,N_17725,N_19234);
nand UO_610 (O_610,N_19061,N_16835);
xnor UO_611 (O_611,N_19580,N_17502);
xor UO_612 (O_612,N_17007,N_16376);
nor UO_613 (O_613,N_16384,N_17036);
nand UO_614 (O_614,N_19714,N_19809);
and UO_615 (O_615,N_18511,N_16943);
or UO_616 (O_616,N_19551,N_16858);
nand UO_617 (O_617,N_19049,N_16975);
xor UO_618 (O_618,N_17087,N_18435);
xor UO_619 (O_619,N_18668,N_18394);
and UO_620 (O_620,N_19448,N_19483);
xor UO_621 (O_621,N_16161,N_16671);
nor UO_622 (O_622,N_16091,N_17823);
or UO_623 (O_623,N_18632,N_18545);
nand UO_624 (O_624,N_18531,N_18717);
nor UO_625 (O_625,N_18758,N_19097);
xor UO_626 (O_626,N_19805,N_16907);
and UO_627 (O_627,N_18064,N_18198);
nor UO_628 (O_628,N_18340,N_18599);
xor UO_629 (O_629,N_18211,N_18684);
nand UO_630 (O_630,N_16579,N_19591);
nand UO_631 (O_631,N_17257,N_16708);
xnor UO_632 (O_632,N_16290,N_19716);
xor UO_633 (O_633,N_16365,N_17796);
or UO_634 (O_634,N_16423,N_16035);
or UO_635 (O_635,N_16241,N_18289);
xnor UO_636 (O_636,N_17358,N_17439);
xor UO_637 (O_637,N_16405,N_19222);
xnor UO_638 (O_638,N_19770,N_17269);
nor UO_639 (O_639,N_19341,N_17063);
nor UO_640 (O_640,N_19029,N_18254);
and UO_641 (O_641,N_19616,N_17942);
xor UO_642 (O_642,N_18197,N_19896);
or UO_643 (O_643,N_18081,N_16248);
nand UO_644 (O_644,N_19498,N_18168);
nor UO_645 (O_645,N_17550,N_16046);
nor UO_646 (O_646,N_19479,N_17054);
xnor UO_647 (O_647,N_16927,N_17968);
nand UO_648 (O_648,N_18357,N_17505);
xor UO_649 (O_649,N_17398,N_16519);
or UO_650 (O_650,N_16417,N_19356);
or UO_651 (O_651,N_19202,N_16171);
nand UO_652 (O_652,N_17420,N_18834);
and UO_653 (O_653,N_19196,N_18894);
and UO_654 (O_654,N_16881,N_16108);
xnor UO_655 (O_655,N_19554,N_16636);
and UO_656 (O_656,N_16698,N_16965);
or UO_657 (O_657,N_18390,N_19177);
or UO_658 (O_658,N_19093,N_18609);
nand UO_659 (O_659,N_16377,N_17565);
xor UO_660 (O_660,N_16292,N_18740);
and UO_661 (O_661,N_17775,N_18644);
xnor UO_662 (O_662,N_17509,N_16212);
xnor UO_663 (O_663,N_17009,N_17557);
and UO_664 (O_664,N_18200,N_18004);
and UO_665 (O_665,N_17982,N_19491);
xnor UO_666 (O_666,N_16552,N_18016);
nor UO_667 (O_667,N_18274,N_18031);
or UO_668 (O_668,N_16966,N_18257);
nor UO_669 (O_669,N_16353,N_17570);
nand UO_670 (O_670,N_16306,N_17610);
and UO_671 (O_671,N_18941,N_19804);
nand UO_672 (O_672,N_17567,N_17233);
xnor UO_673 (O_673,N_17746,N_18017);
or UO_674 (O_674,N_16130,N_16738);
and UO_675 (O_675,N_19363,N_19997);
or UO_676 (O_676,N_17285,N_18338);
or UO_677 (O_677,N_18540,N_16067);
nand UO_678 (O_678,N_17130,N_19625);
and UO_679 (O_679,N_16849,N_16993);
xnor UO_680 (O_680,N_16932,N_19905);
or UO_681 (O_681,N_17853,N_17827);
or UO_682 (O_682,N_18453,N_18452);
nor UO_683 (O_683,N_18548,N_18265);
nand UO_684 (O_684,N_18703,N_18896);
and UO_685 (O_685,N_18448,N_17714);
nor UO_686 (O_686,N_16008,N_18096);
and UO_687 (O_687,N_19627,N_17126);
xor UO_688 (O_688,N_19054,N_19567);
or UO_689 (O_689,N_17487,N_17239);
or UO_690 (O_690,N_17952,N_18614);
or UO_691 (O_691,N_16101,N_17875);
nor UO_692 (O_692,N_17465,N_18173);
and UO_693 (O_693,N_18706,N_18476);
and UO_694 (O_694,N_18571,N_18714);
xnor UO_695 (O_695,N_19964,N_18401);
nand UO_696 (O_696,N_17592,N_16284);
nor UO_697 (O_697,N_18459,N_17467);
nand UO_698 (O_698,N_16585,N_17092);
xor UO_699 (O_699,N_18494,N_16088);
nor UO_700 (O_700,N_17741,N_18474);
xor UO_701 (O_701,N_17828,N_17844);
and UO_702 (O_702,N_17548,N_17978);
nor UO_703 (O_703,N_18044,N_18773);
and UO_704 (O_704,N_18981,N_16209);
or UO_705 (O_705,N_18456,N_19183);
and UO_706 (O_706,N_17372,N_16785);
or UO_707 (O_707,N_19378,N_19211);
nor UO_708 (O_708,N_16874,N_17962);
and UO_709 (O_709,N_16957,N_18792);
nor UO_710 (O_710,N_19891,N_19556);
nand UO_711 (O_711,N_19439,N_18526);
nor UO_712 (O_712,N_19339,N_19121);
nand UO_713 (O_713,N_18524,N_16280);
xnor UO_714 (O_714,N_16852,N_18491);
nor UO_715 (O_715,N_18328,N_19038);
nor UO_716 (O_716,N_17508,N_19915);
nor UO_717 (O_717,N_16760,N_16213);
or UO_718 (O_718,N_16956,N_17129);
or UO_719 (O_719,N_16371,N_16432);
xor UO_720 (O_720,N_16561,N_17292);
xnor UO_721 (O_721,N_18698,N_16139);
nand UO_722 (O_722,N_19371,N_18816);
nand UO_723 (O_723,N_19084,N_17365);
xnor UO_724 (O_724,N_17350,N_19235);
and UO_725 (O_725,N_17370,N_19404);
xnor UO_726 (O_726,N_17604,N_19590);
nand UO_727 (O_727,N_18381,N_19274);
xor UO_728 (O_728,N_17902,N_18248);
nor UO_729 (O_729,N_19901,N_16819);
nand UO_730 (O_730,N_16607,N_17879);
and UO_731 (O_731,N_17442,N_16089);
nor UO_732 (O_732,N_16427,N_16487);
nor UO_733 (O_733,N_17173,N_18305);
and UO_734 (O_734,N_19348,N_16463);
or UO_735 (O_735,N_17235,N_16456);
nand UO_736 (O_736,N_17052,N_19640);
xnor UO_737 (O_737,N_16315,N_17517);
or UO_738 (O_738,N_17481,N_18135);
nor UO_739 (O_739,N_17379,N_18027);
or UO_740 (O_740,N_19265,N_17118);
nand UO_741 (O_741,N_16996,N_16279);
and UO_742 (O_742,N_17368,N_17217);
nand UO_743 (O_743,N_19772,N_18089);
nand UO_744 (O_744,N_19089,N_16540);
nand UO_745 (O_745,N_16827,N_19529);
or UO_746 (O_746,N_19594,N_17152);
and UO_747 (O_747,N_17428,N_18502);
nor UO_748 (O_748,N_16576,N_19719);
nand UO_749 (O_749,N_17256,N_19172);
and UO_750 (O_750,N_18461,N_18483);
nor UO_751 (O_751,N_19470,N_17102);
or UO_752 (O_752,N_18863,N_17691);
nor UO_753 (O_753,N_16777,N_19755);
nor UO_754 (O_754,N_16673,N_17037);
xor UO_755 (O_755,N_19002,N_16851);
or UO_756 (O_756,N_17212,N_18831);
or UO_757 (O_757,N_16093,N_16973);
and UO_758 (O_758,N_18806,N_19259);
and UO_759 (O_759,N_18182,N_16571);
and UO_760 (O_760,N_19381,N_17880);
or UO_761 (O_761,N_17180,N_18767);
xor UO_762 (O_762,N_18630,N_19983);
or UO_763 (O_763,N_16277,N_19798);
xor UO_764 (O_764,N_18546,N_16976);
xor UO_765 (O_765,N_16831,N_19187);
or UO_766 (O_766,N_19327,N_19606);
and UO_767 (O_767,N_17146,N_16320);
xnor UO_768 (O_768,N_17933,N_18330);
nand UO_769 (O_769,N_19396,N_18645);
xor UO_770 (O_770,N_19637,N_18216);
and UO_771 (O_771,N_16613,N_18711);
nor UO_772 (O_772,N_18891,N_16141);
or UO_773 (O_773,N_17679,N_16041);
nor UO_774 (O_774,N_16554,N_19305);
nand UO_775 (O_775,N_17407,N_16116);
or UO_776 (O_776,N_18952,N_16049);
and UO_777 (O_777,N_16892,N_18370);
or UO_778 (O_778,N_18908,N_19007);
or UO_779 (O_779,N_17176,N_16230);
xnor UO_780 (O_780,N_19742,N_17241);
xor UO_781 (O_781,N_16135,N_18901);
or UO_782 (O_782,N_19962,N_18154);
or UO_783 (O_783,N_17706,N_16022);
nand UO_784 (O_784,N_18931,N_18271);
nor UO_785 (O_785,N_17855,N_19425);
xnor UO_786 (O_786,N_18056,N_18741);
nor UO_787 (O_787,N_19619,N_16271);
nor UO_788 (O_788,N_16567,N_16539);
xnor UO_789 (O_789,N_19465,N_18812);
nor UO_790 (O_790,N_18999,N_17914);
xnor UO_791 (O_791,N_18424,N_17497);
or UO_792 (O_792,N_19256,N_17642);
nand UO_793 (O_793,N_17286,N_18040);
or UO_794 (O_794,N_16421,N_17409);
or UO_795 (O_795,N_17728,N_19940);
nor UO_796 (O_796,N_19558,N_19757);
and UO_797 (O_797,N_17248,N_17090);
nand UO_798 (O_798,N_17314,N_18180);
xor UO_799 (O_799,N_19129,N_16786);
nand UO_800 (O_800,N_19020,N_16660);
xnor UO_801 (O_801,N_17562,N_16899);
nor UO_802 (O_802,N_18032,N_16183);
nor UO_803 (O_803,N_17648,N_18554);
xnor UO_804 (O_804,N_16709,N_19389);
nor UO_805 (O_805,N_17444,N_19749);
nor UO_806 (O_806,N_17380,N_19426);
nand UO_807 (O_807,N_18203,N_17514);
nor UO_808 (O_808,N_19153,N_18406);
nor UO_809 (O_809,N_16657,N_18447);
and UO_810 (O_810,N_19397,N_18725);
and UO_811 (O_811,N_16754,N_18366);
and UO_812 (O_812,N_16276,N_18117);
nand UO_813 (O_813,N_18872,N_16581);
or UO_814 (O_814,N_16536,N_16434);
nor UO_815 (O_815,N_17168,N_17211);
and UO_816 (O_816,N_16574,N_17310);
and UO_817 (O_817,N_16125,N_16408);
or UO_818 (O_818,N_17647,N_19338);
nand UO_819 (O_819,N_16866,N_19068);
xor UO_820 (O_820,N_16304,N_16753);
nor UO_821 (O_821,N_19703,N_18130);
xor UO_822 (O_822,N_16117,N_16479);
xor UO_823 (O_823,N_16645,N_18313);
nand UO_824 (O_824,N_19881,N_16674);
and UO_825 (O_825,N_19894,N_18971);
xnor UO_826 (O_826,N_18680,N_16386);
nand UO_827 (O_827,N_17187,N_18805);
xnor UO_828 (O_828,N_17564,N_19932);
nor UO_829 (O_829,N_19512,N_18083);
nor UO_830 (O_830,N_17048,N_16813);
xor UO_831 (O_831,N_19698,N_18314);
and UO_832 (O_832,N_16587,N_19143);
or UO_833 (O_833,N_16132,N_18281);
nand UO_834 (O_834,N_19033,N_17017);
or UO_835 (O_835,N_16710,N_18219);
xnor UO_836 (O_836,N_17584,N_19286);
nor UO_837 (O_837,N_18870,N_16919);
nand UO_838 (O_838,N_19326,N_19255);
nor UO_839 (O_839,N_17980,N_16349);
and UO_840 (O_840,N_16661,N_18301);
xor UO_841 (O_841,N_17549,N_17021);
nor UO_842 (O_842,N_16772,N_18397);
nor UO_843 (O_843,N_19581,N_18592);
or UO_844 (O_844,N_16555,N_19300);
and UO_845 (O_845,N_17957,N_19917);
xnor UO_846 (O_846,N_18194,N_19533);
xnor UO_847 (O_847,N_18836,N_19675);
nand UO_848 (O_848,N_18097,N_16061);
nor UO_849 (O_849,N_17752,N_17155);
and UO_850 (O_850,N_19115,N_16140);
nor UO_851 (O_851,N_17121,N_19191);
nor UO_852 (O_852,N_19429,N_16307);
xor UO_853 (O_853,N_17845,N_16991);
or UO_854 (O_854,N_16246,N_18079);
and UO_855 (O_855,N_17304,N_18312);
nor UO_856 (O_856,N_19956,N_19416);
or UO_857 (O_857,N_18162,N_16838);
or UO_858 (O_858,N_19150,N_16319);
nand UO_859 (O_859,N_19432,N_18776);
and UO_860 (O_860,N_17858,N_19737);
nand UO_861 (O_861,N_18202,N_16097);
and UO_862 (O_862,N_18138,N_16805);
nand UO_863 (O_863,N_17638,N_16275);
nor UO_864 (O_864,N_16461,N_18866);
and UO_865 (O_865,N_17201,N_19492);
or UO_866 (O_866,N_18547,N_19118);
nand UO_867 (O_867,N_19229,N_18586);
nor UO_868 (O_868,N_19460,N_17354);
nand UO_869 (O_869,N_19440,N_17618);
xnor UO_870 (O_870,N_19671,N_19847);
nand UO_871 (O_871,N_19754,N_17621);
nand UO_872 (O_872,N_19670,N_18346);
or UO_873 (O_873,N_19037,N_18768);
and UO_874 (O_874,N_17954,N_18156);
nor UO_875 (O_875,N_18360,N_16060);
xor UO_876 (O_876,N_19219,N_18784);
nor UO_877 (O_877,N_16685,N_18480);
nor UO_878 (O_878,N_19602,N_16003);
xor UO_879 (O_879,N_19822,N_17988);
nor UO_880 (O_880,N_19346,N_17022);
or UO_881 (O_881,N_18311,N_17218);
nor UO_882 (O_882,N_19697,N_16978);
and UO_883 (O_883,N_19978,N_17654);
and UO_884 (O_884,N_16393,N_17038);
xor UO_885 (O_885,N_18399,N_18628);
xor UO_886 (O_886,N_19715,N_17806);
nand UO_887 (O_887,N_18879,N_16285);
nand UO_888 (O_888,N_16543,N_17289);
nand UO_889 (O_889,N_19949,N_16669);
nor UO_890 (O_890,N_17167,N_18856);
or UO_891 (O_891,N_16449,N_19331);
nand UO_892 (O_892,N_16795,N_18606);
nand UO_893 (O_893,N_19099,N_19208);
xnor UO_894 (O_894,N_19540,N_19561);
xor UO_895 (O_895,N_17971,N_18210);
nand UO_896 (O_896,N_18495,N_16936);
or UO_897 (O_897,N_18810,N_18076);
xnor UO_898 (O_898,N_19226,N_18002);
nor UO_899 (O_899,N_18826,N_17485);
xnor UO_900 (O_900,N_16435,N_17687);
nand UO_901 (O_901,N_18136,N_16359);
and UO_902 (O_902,N_17552,N_16620);
and UO_903 (O_903,N_19729,N_17240);
or UO_904 (O_904,N_17911,N_19562);
nor UO_905 (O_905,N_19790,N_18109);
and UO_906 (O_906,N_16453,N_18646);
xor UO_907 (O_907,N_17738,N_18666);
xor UO_908 (O_908,N_16316,N_18430);
nor UO_909 (O_909,N_16527,N_18100);
and UO_910 (O_910,N_16446,N_16797);
or UO_911 (O_911,N_17588,N_16221);
nand UO_912 (O_912,N_17172,N_17768);
nand UO_913 (O_913,N_16162,N_19630);
xnor UO_914 (O_914,N_16764,N_16911);
xor UO_915 (O_915,N_19733,N_19780);
xor UO_916 (O_916,N_17568,N_18468);
nand UO_917 (O_917,N_18367,N_16073);
nor UO_918 (O_918,N_17471,N_17390);
nand UO_919 (O_919,N_18179,N_18996);
nand UO_920 (O_920,N_19712,N_16482);
nand UO_921 (O_921,N_18221,N_16984);
nand UO_922 (O_922,N_16967,N_17573);
nor UO_923 (O_923,N_16019,N_19488);
or UO_924 (O_924,N_17031,N_19722);
nand UO_925 (O_925,N_16178,N_19463);
and UO_926 (O_926,N_16929,N_17913);
or UO_927 (O_927,N_17077,N_16666);
or UO_928 (O_928,N_17660,N_16845);
nand UO_929 (O_929,N_17058,N_16205);
xnor UO_930 (O_930,N_19593,N_18258);
xnor UO_931 (O_931,N_17425,N_19027);
xor UO_932 (O_932,N_16470,N_19047);
xnor UO_933 (O_933,N_18185,N_19889);
and UO_934 (O_934,N_17200,N_17641);
nand UO_935 (O_935,N_17349,N_16020);
nand UO_936 (O_936,N_17426,N_17323);
and UO_937 (O_937,N_19090,N_17762);
nor UO_938 (O_938,N_16742,N_16337);
xnor UO_939 (O_939,N_19306,N_16904);
xnor UO_940 (O_940,N_18103,N_19501);
nor UO_941 (O_941,N_16908,N_17455);
and UO_942 (O_942,N_16127,N_16910);
nand UO_943 (O_943,N_18778,N_18660);
and UO_944 (O_944,N_19958,N_16768);
nor UO_945 (O_945,N_19391,N_17629);
and UO_946 (O_946,N_18669,N_16651);
or UO_947 (O_947,N_17895,N_18374);
xnor UO_948 (O_948,N_17356,N_16791);
and UO_949 (O_949,N_17569,N_19763);
xnor UO_950 (O_950,N_18708,N_19126);
nor UO_951 (O_951,N_18620,N_18462);
nor UO_952 (O_952,N_19572,N_19823);
nand UO_953 (O_953,N_17966,N_17940);
nor UO_954 (O_954,N_17499,N_18269);
nor UO_955 (O_955,N_16783,N_17532);
nor UO_956 (O_956,N_17142,N_19127);
or UO_957 (O_957,N_19546,N_16106);
and UO_958 (O_958,N_17521,N_17181);
nor UO_959 (O_959,N_17581,N_19012);
and UO_960 (O_960,N_17716,N_18520);
or UO_961 (O_961,N_19992,N_19531);
or UO_962 (O_962,N_19424,N_16355);
nor UO_963 (O_963,N_17759,N_16532);
nor UO_964 (O_964,N_19831,N_19632);
xnor UO_965 (O_965,N_16498,N_17103);
xnor UO_966 (O_966,N_16621,N_16740);
nor UO_967 (O_967,N_17441,N_18237);
nor UO_968 (O_968,N_18217,N_17835);
nor UO_969 (O_969,N_17012,N_19060);
or UO_970 (O_970,N_18911,N_19815);
nor UO_971 (O_971,N_16457,N_17834);
and UO_972 (O_972,N_16425,N_19254);
nand UO_973 (O_973,N_19702,N_19976);
and UO_974 (O_974,N_17625,N_16066);
xor UO_975 (O_975,N_18148,N_18500);
nor UO_976 (O_976,N_18624,N_19624);
nand UO_977 (O_977,N_19771,N_18661);
xor UO_978 (O_978,N_18122,N_16841);
xnor UO_979 (O_979,N_18588,N_17150);
and UO_980 (O_980,N_19642,N_18754);
and UO_981 (O_981,N_18927,N_17190);
nor UO_982 (O_982,N_18011,N_19585);
and UO_983 (O_983,N_18718,N_17626);
and UO_984 (O_984,N_18842,N_18389);
xnor UO_985 (O_985,N_16397,N_17628);
nand UO_986 (O_986,N_19298,N_18007);
and UO_987 (O_987,N_17371,N_16282);
nand UO_988 (O_988,N_19142,N_16233);
nor UO_989 (O_989,N_18022,N_17101);
xnor UO_990 (O_990,N_19116,N_19044);
xnor UO_991 (O_991,N_16095,N_17627);
and UO_992 (O_992,N_16369,N_18140);
nor UO_993 (O_993,N_16918,N_18851);
and UO_994 (O_994,N_17696,N_16692);
nor UO_995 (O_995,N_18479,N_16197);
and UO_996 (O_996,N_18533,N_19136);
nor UO_997 (O_997,N_19912,N_18116);
nand UO_998 (O_998,N_16252,N_18099);
and UO_999 (O_999,N_18843,N_17634);
or UO_1000 (O_1000,N_19520,N_17414);
nand UO_1001 (O_1001,N_17049,N_18510);
nand UO_1002 (O_1002,N_19878,N_19275);
nand UO_1003 (O_1003,N_16885,N_19358);
or UO_1004 (O_1004,N_18118,N_17484);
or UO_1005 (O_1005,N_17221,N_16779);
and UO_1006 (O_1006,N_17945,N_19392);
nor UO_1007 (O_1007,N_18878,N_19764);
or UO_1008 (O_1008,N_19412,N_18199);
or UO_1009 (O_1009,N_16507,N_19360);
xor UO_1010 (O_1010,N_16270,N_17923);
nand UO_1011 (O_1011,N_17331,N_19750);
nor UO_1012 (O_1012,N_18726,N_17266);
xor UO_1013 (O_1013,N_18034,N_18256);
or UO_1014 (O_1014,N_17106,N_18014);
and UO_1015 (O_1015,N_16473,N_19650);
xnor UO_1016 (O_1016,N_19975,N_16378);
xor UO_1017 (O_1017,N_17143,N_19549);
xnor UO_1018 (O_1018,N_19882,N_19310);
nor UO_1019 (O_1019,N_18782,N_17293);
nor UO_1020 (O_1020,N_17270,N_16723);
nor UO_1021 (O_1021,N_17018,N_16072);
nand UO_1022 (O_1022,N_17571,N_16603);
or UO_1023 (O_1023,N_19628,N_17692);
or UO_1024 (O_1024,N_16770,N_17657);
nor UO_1025 (O_1025,N_19509,N_18721);
or UO_1026 (O_1026,N_18874,N_18663);
nor UO_1027 (O_1027,N_17537,N_17307);
nor UO_1028 (O_1028,N_18648,N_19946);
nor UO_1029 (O_1029,N_18969,N_17887);
or UO_1030 (O_1030,N_18469,N_18432);
nor UO_1031 (O_1031,N_17352,N_16672);
or UO_1032 (O_1032,N_19565,N_19810);
and UO_1033 (O_1033,N_18396,N_17936);
nor UO_1034 (O_1034,N_18033,N_18383);
nand UO_1035 (O_1035,N_16181,N_18656);
nor UO_1036 (O_1036,N_19058,N_17133);
xnor UO_1037 (O_1037,N_17324,N_16364);
nor UO_1038 (O_1038,N_17987,N_16015);
nand UO_1039 (O_1039,N_16822,N_17461);
xnor UO_1040 (O_1040,N_19877,N_17637);
and UO_1041 (O_1041,N_17144,N_18151);
xor UO_1042 (O_1042,N_18534,N_18241);
or UO_1043 (O_1043,N_16272,N_18344);
and UO_1044 (O_1044,N_17171,N_18759);
xnor UO_1045 (O_1045,N_17898,N_19867);
nor UO_1046 (O_1046,N_16012,N_18916);
and UO_1047 (O_1047,N_17948,N_19228);
nand UO_1048 (O_1048,N_16374,N_17926);
xnor UO_1049 (O_1049,N_19758,N_18472);
and UO_1050 (O_1050,N_17518,N_18425);
and UO_1051 (O_1051,N_19659,N_16477);
xor UO_1052 (O_1052,N_19308,N_16150);
xnor UO_1053 (O_1053,N_16166,N_19661);
or UO_1054 (O_1054,N_17437,N_19459);
xnor UO_1055 (O_1055,N_16054,N_18939);
and UO_1056 (O_1056,N_19954,N_19262);
and UO_1057 (O_1057,N_17761,N_19766);
and UO_1058 (O_1058,N_19017,N_16078);
nor UO_1059 (O_1059,N_19875,N_18228);
nand UO_1060 (O_1060,N_19062,N_16188);
xor UO_1061 (O_1061,N_19019,N_17477);
or UO_1062 (O_1062,N_18707,N_16988);
nor UO_1063 (O_1063,N_16198,N_19103);
and UO_1064 (O_1064,N_19897,N_16289);
and UO_1065 (O_1065,N_18757,N_17045);
nand UO_1066 (O_1066,N_18506,N_19514);
nor UO_1067 (O_1067,N_19427,N_17774);
nor UO_1068 (O_1068,N_19434,N_18342);
or UO_1069 (O_1069,N_18243,N_17745);
nand UO_1070 (O_1070,N_16480,N_19687);
xor UO_1071 (O_1071,N_18414,N_18233);
or UO_1072 (O_1072,N_18565,N_17591);
and UO_1073 (O_1073,N_16168,N_16938);
nor UO_1074 (O_1074,N_18041,N_16018);
and UO_1075 (O_1075,N_16286,N_17284);
nand UO_1076 (O_1076,N_18412,N_16484);
xnor UO_1077 (O_1077,N_18113,N_18612);
or UO_1078 (O_1078,N_19641,N_18061);
or UO_1079 (O_1079,N_16399,N_18347);
nor UO_1080 (O_1080,N_18422,N_17900);
or UO_1081 (O_1081,N_19110,N_18341);
xor UO_1082 (O_1082,N_16720,N_18230);
xnor UO_1083 (O_1083,N_18443,N_17447);
and UO_1084 (O_1084,N_16763,N_16946);
xnor UO_1085 (O_1085,N_16615,N_18427);
nand UO_1086 (O_1086,N_16602,N_17787);
xnor UO_1087 (O_1087,N_17137,N_18171);
nor UO_1088 (O_1088,N_16857,N_17294);
xnor UO_1089 (O_1089,N_19464,N_18830);
xor UO_1090 (O_1090,N_18798,N_19885);
nand UO_1091 (O_1091,N_19886,N_18672);
nor UO_1092 (O_1092,N_17182,N_19085);
and UO_1093 (O_1093,N_19838,N_16922);
and UO_1094 (O_1094,N_18215,N_18147);
nand UO_1095 (O_1095,N_17319,N_19646);
nand UO_1096 (O_1096,N_17757,N_19942);
xnor UO_1097 (O_1097,N_17632,N_19873);
xnor UO_1098 (O_1098,N_18294,N_16825);
nand UO_1099 (O_1099,N_18149,N_16395);
xor UO_1100 (O_1100,N_16590,N_17179);
and UO_1101 (O_1101,N_18114,N_19537);
nand UO_1102 (O_1102,N_19253,N_16983);
nor UO_1103 (O_1103,N_19617,N_18363);
nand UO_1104 (O_1104,N_18659,N_18886);
nand UO_1105 (O_1105,N_16722,N_16499);
nor UO_1106 (O_1106,N_18731,N_19455);
xnor UO_1107 (O_1107,N_17337,N_18345);
xor UO_1108 (O_1108,N_17608,N_19433);
or UO_1109 (O_1109,N_18493,N_19288);
xnor UO_1110 (O_1110,N_17237,N_16635);
nor UO_1111 (O_1111,N_17157,N_19713);
xnor UO_1112 (O_1112,N_17228,N_16939);
or UO_1113 (O_1113,N_16038,N_16375);
nand UO_1114 (O_1114,N_18781,N_18876);
nor UO_1115 (O_1115,N_19517,N_19736);
nor UO_1116 (O_1116,N_18650,N_17799);
nor UO_1117 (O_1117,N_16357,N_18356);
nor UO_1118 (O_1118,N_19887,N_19760);
and UO_1119 (O_1119,N_18115,N_16630);
nor UO_1120 (O_1120,N_16591,N_17535);
nand UO_1121 (O_1121,N_17884,N_19926);
and UO_1122 (O_1122,N_16496,N_19898);
nand UO_1123 (O_1123,N_18803,N_16872);
xor UO_1124 (O_1124,N_16190,N_18023);
and UO_1125 (O_1125,N_19631,N_17739);
or UO_1126 (O_1126,N_17427,N_17123);
nor UO_1127 (O_1127,N_17254,N_19289);
nor UO_1128 (O_1128,N_16755,N_19574);
nand UO_1129 (O_1129,N_17956,N_18512);
xnor UO_1130 (O_1130,N_18608,N_16491);
xnor UO_1131 (O_1131,N_18832,N_17367);
nor UO_1132 (O_1132,N_19493,N_16604);
nand UO_1133 (O_1133,N_17718,N_19461);
nand UO_1134 (O_1134,N_17528,N_16860);
nor UO_1135 (O_1135,N_17667,N_16817);
nand UO_1136 (O_1136,N_16896,N_18783);
xnor UO_1137 (O_1137,N_17469,N_18133);
and UO_1138 (O_1138,N_16346,N_16752);
nor UO_1139 (O_1139,N_17681,N_17306);
xor UO_1140 (O_1140,N_17905,N_19676);
and UO_1141 (O_1141,N_16816,N_17671);
and UO_1142 (O_1142,N_18411,N_19720);
nor UO_1143 (O_1143,N_17846,N_18825);
and UO_1144 (O_1144,N_16806,N_19320);
and UO_1145 (O_1145,N_19890,N_17958);
nor UO_1146 (O_1146,N_18929,N_17086);
or UO_1147 (O_1147,N_19010,N_16062);
nor UO_1148 (O_1148,N_17252,N_16206);
nand UO_1149 (O_1149,N_16258,N_19173);
and UO_1150 (O_1150,N_19694,N_18300);
or UO_1151 (O_1151,N_17189,N_16780);
or UO_1152 (O_1152,N_17406,N_18249);
nor UO_1153 (O_1153,N_19842,N_19066);
or UO_1154 (O_1154,N_19787,N_16006);
xor UO_1155 (O_1155,N_16500,N_19579);
xor UO_1156 (O_1156,N_19303,N_17174);
nand UO_1157 (O_1157,N_19174,N_19070);
nand UO_1158 (O_1158,N_17540,N_16412);
nand UO_1159 (O_1159,N_18139,N_18445);
nor UO_1160 (O_1160,N_17060,N_19621);
nand UO_1161 (O_1161,N_17876,N_17050);
nand UO_1162 (O_1162,N_18482,N_18150);
xor UO_1163 (O_1163,N_18702,N_17612);
nor UO_1164 (O_1164,N_16494,N_19883);
xor UO_1165 (O_1165,N_17870,N_18522);
nand UO_1166 (O_1166,N_18760,N_19080);
or UO_1167 (O_1167,N_17559,N_19679);
xnor UO_1168 (O_1168,N_17219,N_19355);
or UO_1169 (O_1169,N_18796,N_17299);
nand UO_1170 (O_1170,N_17732,N_18385);
nand UO_1171 (O_1171,N_16308,N_19789);
nor UO_1172 (O_1172,N_16173,N_16809);
nand UO_1173 (O_1173,N_18455,N_18622);
and UO_1174 (O_1174,N_18454,N_18623);
or UO_1175 (O_1175,N_16253,N_17516);
xnor UO_1176 (O_1176,N_19730,N_16236);
nor UO_1177 (O_1177,N_17345,N_17432);
xor UO_1178 (O_1178,N_18541,N_18037);
or UO_1179 (O_1179,N_17666,N_18042);
or UO_1180 (O_1180,N_16823,N_19799);
and UO_1181 (O_1181,N_17105,N_17878);
nand UO_1182 (O_1182,N_19124,N_18869);
xor UO_1183 (O_1183,N_18191,N_19945);
and UO_1184 (O_1184,N_19950,N_19474);
or UO_1185 (O_1185,N_18596,N_19290);
and UO_1186 (O_1186,N_18337,N_17015);
nor UO_1187 (O_1187,N_18997,N_16803);
or UO_1188 (O_1188,N_19322,N_17336);
or UO_1189 (O_1189,N_16231,N_16508);
nand UO_1190 (O_1190,N_18021,N_16431);
xnor UO_1191 (O_1191,N_18930,N_18799);
and UO_1192 (O_1192,N_19485,N_19695);
and UO_1193 (O_1193,N_18348,N_16203);
nand UO_1194 (O_1194,N_16410,N_19333);
and UO_1195 (O_1195,N_18600,N_19246);
and UO_1196 (O_1196,N_16195,N_16867);
nand UO_1197 (O_1197,N_19691,N_18979);
or UO_1198 (O_1198,N_17125,N_19989);
or UO_1199 (O_1199,N_18213,N_18537);
and UO_1200 (O_1200,N_17946,N_16401);
nor UO_1201 (O_1201,N_17836,N_18513);
nor UO_1202 (O_1202,N_18857,N_19994);
xor UO_1203 (O_1203,N_19794,N_19869);
nor UO_1204 (O_1204,N_16726,N_18665);
nor UO_1205 (O_1205,N_19311,N_16051);
and UO_1206 (O_1206,N_18110,N_18259);
nor UO_1207 (O_1207,N_16265,N_19777);
nand UO_1208 (O_1208,N_18735,N_19105);
nor UO_1209 (O_1209,N_16033,N_19812);
xnor UO_1210 (O_1210,N_17947,N_18470);
nor UO_1211 (O_1211,N_17959,N_18204);
xnor UO_1212 (O_1212,N_17251,N_16053);
and UO_1213 (O_1213,N_16092,N_17530);
and UO_1214 (O_1214,N_16987,N_18036);
nand UO_1215 (O_1215,N_18507,N_16982);
and UO_1216 (O_1216,N_19064,N_17302);
xor UO_1217 (O_1217,N_17195,N_17976);
nor UO_1218 (O_1218,N_19321,N_18551);
nand UO_1219 (O_1219,N_17149,N_16949);
nand UO_1220 (O_1220,N_19575,N_18484);
xor UO_1221 (O_1221,N_18153,N_17525);
nor UO_1222 (O_1222,N_18802,N_19656);
and UO_1223 (O_1223,N_19184,N_16102);
and UO_1224 (O_1224,N_18786,N_18841);
xnor UO_1225 (O_1225,N_19073,N_17417);
and UO_1226 (O_1226,N_17396,N_18539);
xnor UO_1227 (O_1227,N_17064,N_19157);
or UO_1228 (O_1228,N_16830,N_16643);
and UO_1229 (O_1229,N_18282,N_19663);
and UO_1230 (O_1230,N_19001,N_18297);
and UO_1231 (O_1231,N_18403,N_16196);
and UO_1232 (O_1232,N_16787,N_17615);
nor UO_1233 (O_1233,N_18693,N_16871);
or UO_1234 (O_1234,N_17617,N_19797);
or UO_1235 (O_1235,N_17154,N_19301);
nand UO_1236 (O_1236,N_19538,N_19830);
nand UO_1237 (O_1237,N_17658,N_16303);
xor UO_1238 (O_1238,N_16074,N_18270);
and UO_1239 (O_1239,N_18986,N_16110);
nor UO_1240 (O_1240,N_17712,N_16688);
nand UO_1241 (O_1241,N_18625,N_19472);
xnor UO_1242 (O_1242,N_19131,N_17039);
xor UO_1243 (O_1243,N_16719,N_17539);
and UO_1244 (O_1244,N_17856,N_19081);
nand UO_1245 (O_1245,N_19369,N_19502);
and UO_1246 (O_1246,N_19418,N_16100);
xor UO_1247 (O_1247,N_17463,N_18882);
or UO_1248 (O_1248,N_18587,N_16523);
nor UO_1249 (O_1249,N_16358,N_18838);
xor UO_1250 (O_1250,N_17456,N_17273);
nor UO_1251 (O_1251,N_19618,N_16633);
nand UO_1252 (O_1252,N_18563,N_19335);
nand UO_1253 (O_1253,N_17277,N_16625);
nor UO_1254 (O_1254,N_19862,N_17740);
and UO_1255 (O_1255,N_16242,N_18904);
nor UO_1256 (O_1256,N_16331,N_19469);
xor UO_1257 (O_1257,N_17112,N_16679);
nor UO_1258 (O_1258,N_19768,N_16032);
or UO_1259 (O_1259,N_19200,N_16382);
or UO_1260 (O_1260,N_18868,N_18048);
xor UO_1261 (O_1261,N_18131,N_17639);
nand UO_1262 (O_1262,N_16792,N_16148);
nand UO_1263 (O_1263,N_17378,N_18085);
nor UO_1264 (O_1264,N_17916,N_19937);
or UO_1265 (O_1265,N_17377,N_17395);
or UO_1266 (O_1266,N_17851,N_18734);
and UO_1267 (O_1267,N_19732,N_19524);
or UO_1268 (O_1268,N_18517,N_18881);
and UO_1269 (O_1269,N_18172,N_18509);
and UO_1270 (O_1270,N_19230,N_18193);
and UO_1271 (O_1271,N_17779,N_17028);
xnor UO_1272 (O_1272,N_17382,N_19071);
xnor UO_1273 (O_1273,N_16568,N_17283);
xnor UO_1274 (O_1274,N_18890,N_17117);
xor UO_1275 (O_1275,N_18576,N_19336);
nor UO_1276 (O_1276,N_18467,N_19171);
nand UO_1277 (O_1277,N_17702,N_19708);
nand UO_1278 (O_1278,N_17578,N_19000);
nand UO_1279 (O_1279,N_17596,N_18478);
nand UO_1280 (O_1280,N_16832,N_17820);
or UO_1281 (O_1281,N_16998,N_19102);
nand UO_1282 (O_1282,N_18557,N_16113);
nand UO_1283 (O_1283,N_16059,N_18532);
and UO_1284 (O_1284,N_17332,N_18716);
nor UO_1285 (O_1285,N_19041,N_18286);
xnor UO_1286 (O_1286,N_17147,N_19953);
and UO_1287 (O_1287,N_16914,N_19584);
xor UO_1288 (O_1288,N_18655,N_17791);
or UO_1289 (O_1289,N_19677,N_18918);
nor UO_1290 (O_1290,N_16774,N_17454);
nor UO_1291 (O_1291,N_16917,N_18486);
xnor UO_1292 (O_1292,N_16596,N_19040);
xor UO_1293 (O_1293,N_18295,N_18690);
or UO_1294 (O_1294,N_18327,N_18088);
xor UO_1295 (O_1295,N_18499,N_19979);
nor UO_1296 (O_1296,N_18515,N_16441);
nor UO_1297 (O_1297,N_17829,N_16191);
nor UO_1298 (O_1298,N_18094,N_18575);
xnor UO_1299 (O_1299,N_16940,N_17169);
nor UO_1300 (O_1300,N_18417,N_16980);
xor UO_1301 (O_1301,N_19841,N_18914);
xor UO_1302 (O_1302,N_17084,N_18949);
xnor UO_1303 (O_1303,N_17645,N_19445);
or UO_1304 (O_1304,N_16179,N_19296);
and UO_1305 (O_1305,N_17339,N_19074);
or UO_1306 (O_1306,N_16879,N_18577);
or UO_1307 (O_1307,N_19752,N_18730);
xnor UO_1308 (O_1308,N_18291,N_19069);
xor UO_1309 (O_1309,N_17209,N_19236);
xor UO_1310 (O_1310,N_16972,N_16990);
or UO_1311 (O_1311,N_18938,N_18795);
xor UO_1312 (O_1312,N_17244,N_19031);
or UO_1313 (O_1313,N_19261,N_16547);
or UO_1314 (O_1314,N_17259,N_19543);
or UO_1315 (O_1315,N_19668,N_16481);
or UO_1316 (O_1316,N_16193,N_18898);
or UO_1317 (O_1317,N_19525,N_19786);
xor UO_1318 (O_1318,N_16274,N_17097);
nand UO_1319 (O_1319,N_17689,N_17067);
nor UO_1320 (O_1320,N_16856,N_17316);
xnor UO_1321 (O_1321,N_19620,N_16430);
or UO_1322 (O_1322,N_17582,N_16264);
and UO_1323 (O_1323,N_17493,N_18252);
xnor UO_1324 (O_1324,N_18072,N_16138);
nand UO_1325 (O_1325,N_16693,N_17347);
or UO_1326 (O_1326,N_19059,N_16122);
and UO_1327 (O_1327,N_17423,N_17727);
or UO_1328 (O_1328,N_16107,N_18181);
or UO_1329 (O_1329,N_16646,N_18905);
nand UO_1330 (O_1330,N_18415,N_19438);
or UO_1331 (O_1331,N_17225,N_19317);
nand UO_1332 (O_1332,N_18285,N_17605);
nand UO_1333 (O_1333,N_17070,N_18852);
xnor UO_1334 (O_1334,N_17315,N_17812);
xnor UO_1335 (O_1335,N_17614,N_18157);
or UO_1336 (O_1336,N_16687,N_19453);
xor UO_1337 (O_1337,N_17034,N_19323);
or UO_1338 (O_1338,N_19700,N_19454);
nand UO_1339 (O_1339,N_16301,N_19939);
or UO_1340 (O_1340,N_16255,N_16842);
and UO_1341 (O_1341,N_16005,N_19377);
nand UO_1342 (O_1342,N_19638,N_17119);
xor UO_1343 (O_1343,N_18053,N_18574);
xnor UO_1344 (O_1344,N_19696,N_19583);
and UO_1345 (O_1345,N_19725,N_17267);
nand UO_1346 (O_1346,N_17095,N_19026);
and UO_1347 (O_1347,N_17165,N_19180);
and UO_1348 (O_1348,N_19215,N_16016);
nand UO_1349 (O_1349,N_17577,N_19819);
xor UO_1350 (O_1350,N_16057,N_17265);
nand UO_1351 (O_1351,N_18713,N_17772);
or UO_1352 (O_1352,N_16811,N_18184);
or UO_1353 (O_1353,N_16506,N_18676);
nor UO_1354 (O_1354,N_19388,N_17554);
or UO_1355 (O_1355,N_19077,N_16677);
or UO_1356 (O_1356,N_16745,N_19854);
or UO_1357 (O_1357,N_17970,N_17303);
and UO_1358 (O_1358,N_18583,N_19922);
or UO_1359 (O_1359,N_19496,N_19205);
xor UO_1360 (O_1360,N_19024,N_16912);
or UO_1361 (O_1361,N_16420,N_17227);
or UO_1362 (O_1362,N_16225,N_16641);
and UO_1363 (O_1363,N_19168,N_18010);
or UO_1364 (O_1364,N_19297,N_17199);
nand UO_1365 (O_1365,N_16177,N_19176);
xor UO_1366 (O_1366,N_17677,N_19840);
and UO_1367 (O_1367,N_17435,N_19918);
and UO_1368 (O_1368,N_19655,N_19313);
xor UO_1369 (O_1369,N_16098,N_17749);
and UO_1370 (O_1370,N_18800,N_19683);
nand UO_1371 (O_1371,N_17733,N_18437);
xor UO_1372 (O_1372,N_18166,N_16634);
or UO_1373 (O_1373,N_18739,N_18943);
xnor UO_1374 (O_1374,N_17374,N_19318);
xnor UO_1375 (O_1375,N_16900,N_18839);
xnor UO_1376 (O_1376,N_18419,N_16801);
xnor UO_1377 (O_1377,N_17297,N_17387);
nand UO_1378 (O_1378,N_16756,N_17832);
nand UO_1379 (O_1379,N_17156,N_18958);
and UO_1380 (O_1380,N_19446,N_18322);
xor UO_1381 (O_1381,N_19213,N_19709);
or UO_1382 (O_1382,N_16403,N_16462);
or UO_1383 (O_1383,N_16878,N_17760);
xnor UO_1384 (O_1384,N_19065,N_19910);
nor UO_1385 (O_1385,N_18298,N_17546);
and UO_1386 (O_1386,N_19947,N_16789);
nor UO_1387 (O_1387,N_17862,N_19710);
or UO_1388 (O_1388,N_16714,N_17964);
nor UO_1389 (O_1389,N_17838,N_16750);
or UO_1390 (O_1390,N_17295,N_17560);
xor UO_1391 (O_1391,N_19373,N_18102);
nand UO_1392 (O_1392,N_19267,N_16935);
or UO_1393 (O_1393,N_19860,N_16336);
or UO_1394 (O_1394,N_19504,N_18355);
or UO_1395 (O_1395,N_17693,N_16388);
or UO_1396 (O_1396,N_17789,N_19366);
and UO_1397 (O_1397,N_19923,N_16580);
nand UO_1398 (O_1398,N_17929,N_19559);
or UO_1399 (O_1399,N_19980,N_17556);
or UO_1400 (O_1400,N_19123,N_16721);
xor UO_1401 (O_1401,N_17430,N_18451);
nor UO_1402 (O_1402,N_17492,N_16269);
and UO_1403 (O_1403,N_16969,N_17903);
xnor UO_1404 (O_1404,N_18657,N_16340);
nand UO_1405 (O_1405,N_16913,N_17000);
xnor UO_1406 (O_1406,N_16659,N_17401);
and UO_1407 (O_1407,N_16637,N_16565);
or UO_1408 (O_1408,N_17877,N_17891);
nor UO_1409 (O_1409,N_19807,N_18777);
or UO_1410 (O_1410,N_16428,N_16564);
xnor UO_1411 (O_1411,N_17494,N_16075);
nor UO_1412 (O_1412,N_19693,N_18926);
nand UO_1413 (O_1413,N_16009,N_16663);
xor UO_1414 (O_1414,N_17504,N_17594);
nand UO_1415 (O_1415,N_17918,N_16047);
xnor UO_1416 (O_1416,N_17781,N_16352);
nor UO_1417 (O_1417,N_19657,N_19185);
xor UO_1418 (O_1418,N_17705,N_17205);
xor UO_1419 (O_1419,N_17111,N_18220);
and UO_1420 (O_1420,N_18562,N_17268);
and UO_1421 (O_1421,N_16541,N_19578);
nor UO_1422 (O_1422,N_18287,N_18837);
and UO_1423 (O_1423,N_19145,N_18120);
nor UO_1424 (O_1424,N_17100,N_19376);
or UO_1425 (O_1425,N_18597,N_16926);
xnor UO_1426 (O_1426,N_18283,N_18429);
nor UO_1427 (O_1427,N_18877,N_17805);
or UO_1428 (O_1428,N_17860,N_16525);
nand UO_1429 (O_1429,N_18464,N_17453);
or UO_1430 (O_1430,N_18709,N_18995);
xnor UO_1431 (O_1431,N_16404,N_16875);
or UO_1432 (O_1432,N_17590,N_17069);
xnor UO_1433 (O_1433,N_17255,N_16065);
and UO_1434 (O_1434,N_17357,N_18564);
nor UO_1435 (O_1435,N_16605,N_19555);
xnor UO_1436 (O_1436,N_19016,N_19456);
or UO_1437 (O_1437,N_16642,N_18977);
nor UO_1438 (O_1438,N_19004,N_18421);
or UO_1439 (O_1439,N_16313,N_19270);
nor UO_1440 (O_1440,N_19613,N_19604);
nor UO_1441 (O_1441,N_18590,N_16153);
nand UO_1442 (O_1442,N_16199,N_17348);
nand UO_1443 (O_1443,N_17055,N_19141);
and UO_1444 (O_1444,N_16077,N_18060);
or UO_1445 (O_1445,N_16257,N_17953);
nor UO_1446 (O_1446,N_17640,N_16778);
or UO_1447 (O_1447,N_16776,N_18407);
nand UO_1448 (O_1448,N_17158,N_17748);
nor UO_1449 (O_1449,N_19678,N_18188);
nor UO_1450 (O_1450,N_19120,N_19731);
xnor UO_1451 (O_1451,N_16440,N_19851);
or UO_1452 (O_1452,N_16701,N_17222);
and UO_1453 (O_1453,N_18566,N_17132);
or UO_1454 (O_1454,N_17622,N_17802);
or UO_1455 (O_1455,N_19292,N_18223);
nand UO_1456 (O_1456,N_19547,N_16747);
or UO_1457 (O_1457,N_16223,N_16158);
and UO_1458 (O_1458,N_18077,N_18123);
nand UO_1459 (O_1459,N_18444,N_16186);
nand UO_1460 (O_1460,N_16159,N_18303);
xor UO_1461 (O_1461,N_19217,N_17229);
xnor UO_1462 (O_1462,N_19450,N_18897);
or UO_1463 (O_1463,N_17897,N_17589);
nand UO_1464 (O_1464,N_18959,N_18408);
or UO_1465 (O_1465,N_16379,N_18961);
nand UO_1466 (O_1466,N_16296,N_19165);
xor UO_1467 (O_1467,N_16736,N_18267);
nand UO_1468 (O_1468,N_16662,N_18678);
nand UO_1469 (O_1469,N_16229,N_19328);
nor UO_1470 (O_1470,N_19495,N_16294);
and UO_1471 (O_1471,N_17392,N_16748);
and UO_1472 (O_1472,N_19449,N_17040);
xnor UO_1473 (O_1473,N_16250,N_17313);
or UO_1474 (O_1474,N_16468,N_18629);
or UO_1475 (O_1475,N_19394,N_17376);
xnor UO_1476 (O_1476,N_16921,N_17418);
xnor UO_1477 (O_1477,N_17821,N_17771);
xnor UO_1478 (O_1478,N_16121,N_16655);
nor UO_1479 (O_1479,N_18155,N_16004);
and UO_1480 (O_1480,N_19482,N_16545);
nand UO_1481 (O_1481,N_19977,N_16560);
or UO_1482 (O_1482,N_19622,N_16550);
nor UO_1483 (O_1483,N_18960,N_19607);
nor UO_1484 (O_1484,N_18111,N_18098);
or UO_1485 (O_1485,N_17513,N_17837);
xnor UO_1486 (O_1486,N_17061,N_17854);
or UO_1487 (O_1487,N_19534,N_16808);
xnor UO_1488 (O_1488,N_17245,N_17524);
nor UO_1489 (O_1489,N_18521,N_18736);
nand UO_1490 (O_1490,N_16608,N_18779);
or UO_1491 (O_1491,N_18637,N_19484);
xnor UO_1492 (O_1492,N_17291,N_18530);
and UO_1493 (O_1493,N_19094,N_16737);
nand UO_1494 (O_1494,N_16544,N_18167);
and UO_1495 (O_1495,N_16704,N_18350);
xor UO_1496 (O_1496,N_19342,N_19101);
or UO_1497 (O_1497,N_16076,N_18679);
or UO_1498 (O_1498,N_17747,N_19990);
and UO_1499 (O_1499,N_18550,N_16846);
or UO_1500 (O_1500,N_16416,N_18498);
and UO_1501 (O_1501,N_19283,N_16703);
or UO_1502 (O_1502,N_17397,N_18065);
nand UO_1503 (O_1503,N_16836,N_17673);
or UO_1504 (O_1504,N_17797,N_16751);
xnor UO_1505 (O_1505,N_16535,N_18700);
nand UO_1506 (O_1506,N_16031,N_19609);
and UO_1507 (O_1507,N_16606,N_16180);
and UO_1508 (O_1508,N_19723,N_18853);
nor UO_1509 (O_1509,N_17662,N_19417);
and UO_1510 (O_1510,N_16854,N_17215);
and UO_1511 (O_1511,N_16614,N_18581);
and UO_1512 (O_1512,N_18121,N_19032);
nand UO_1513 (O_1513,N_17989,N_19197);
nand UO_1514 (O_1514,N_18815,N_16598);
nand UO_1515 (O_1515,N_18737,N_19452);
or UO_1516 (O_1516,N_16583,N_19148);
and UO_1517 (O_1517,N_18667,N_16850);
nor UO_1518 (O_1518,N_16202,N_16504);
and UO_1519 (O_1519,N_18828,N_18410);
nor UO_1520 (O_1520,N_19865,N_16586);
nand UO_1521 (O_1521,N_19242,N_18292);
nor UO_1522 (O_1522,N_18438,N_16251);
nand UO_1523 (O_1523,N_17519,N_19349);
and UO_1524 (O_1524,N_17767,N_17717);
nand UO_1525 (O_1525,N_19258,N_16530);
or UO_1526 (O_1526,N_17334,N_18819);
nand UO_1527 (O_1527,N_18353,N_18603);
and UO_1528 (O_1528,N_19893,N_17683);
xor UO_1529 (O_1529,N_17698,N_18145);
and UO_1530 (O_1530,N_17081,N_16454);
nor UO_1531 (O_1531,N_16327,N_18247);
and UO_1532 (O_1532,N_17148,N_17894);
or UO_1533 (O_1533,N_17362,N_17986);
or UO_1534 (O_1534,N_16683,N_16888);
or UO_1535 (O_1535,N_19717,N_18771);
xnor UO_1536 (O_1536,N_18827,N_17924);
and UO_1537 (O_1537,N_19309,N_18101);
or UO_1538 (O_1538,N_16937,N_19384);
and UO_1539 (O_1539,N_19721,N_18846);
nand UO_1540 (O_1540,N_19973,N_18159);
or UO_1541 (O_1541,N_17753,N_16056);
and UO_1542 (O_1542,N_19796,N_16131);
or UO_1543 (O_1543,N_17938,N_18785);
xnor UO_1544 (O_1544,N_19487,N_19128);
xnor UO_1545 (O_1545,N_18956,N_18051);
xnor UO_1546 (O_1546,N_16762,N_16128);
nor UO_1547 (O_1547,N_17635,N_16632);
and UO_1548 (O_1548,N_17161,N_16351);
xor UO_1549 (O_1549,N_17868,N_16654);
or UO_1550 (O_1550,N_19372,N_16518);
and UO_1551 (O_1551,N_18664,N_17857);
xnor UO_1552 (O_1552,N_18019,N_17330);
nor UO_1553 (O_1553,N_17479,N_16344);
or UO_1554 (O_1554,N_19092,N_17468);
nor UO_1555 (O_1555,N_17686,N_17507);
nand UO_1556 (O_1556,N_17795,N_17075);
nor UO_1557 (O_1557,N_17027,N_17136);
and UO_1558 (O_1558,N_17355,N_17871);
xor UO_1559 (O_1559,N_16027,N_16891);
or UO_1560 (O_1560,N_16775,N_16394);
nor UO_1561 (O_1561,N_16226,N_18236);
or UO_1562 (O_1562,N_18307,N_18158);
or UO_1563 (O_1563,N_18161,N_19273);
or UO_1564 (O_1564,N_18372,N_19588);
nand UO_1565 (O_1565,N_19998,N_19428);
nor UO_1566 (O_1566,N_16300,N_17153);
and UO_1567 (O_1567,N_19539,N_17220);
xor UO_1568 (O_1568,N_17765,N_18903);
nor UO_1569 (O_1569,N_17419,N_16549);
nand UO_1570 (O_1570,N_17700,N_19086);
nor UO_1571 (O_1571,N_16123,N_19986);
xnor UO_1572 (O_1572,N_16610,N_16695);
nor UO_1573 (O_1573,N_16422,N_19315);
or UO_1574 (O_1574,N_17703,N_19654);
and UO_1575 (O_1575,N_18290,N_17230);
and UO_1576 (O_1576,N_18321,N_19415);
and UO_1577 (O_1577,N_19824,N_18752);
xor UO_1578 (O_1578,N_17478,N_19114);
or UO_1579 (O_1579,N_16844,N_16156);
nand UO_1580 (O_1580,N_16111,N_17915);
and UO_1581 (O_1581,N_19652,N_18400);
nand UO_1582 (O_1582,N_19859,N_17369);
or UO_1583 (O_1583,N_19155,N_16824);
nor UO_1584 (O_1584,N_18968,N_17886);
nor UO_1585 (O_1585,N_17999,N_17282);
xor UO_1586 (O_1586,N_16143,N_19499);
xor UO_1587 (O_1587,N_18336,N_16335);
nor UO_1588 (O_1588,N_18066,N_17082);
nor UO_1589 (O_1589,N_18361,N_18763);
and UO_1590 (O_1590,N_19170,N_17869);
xnor UO_1591 (O_1591,N_18050,N_16418);
and UO_1592 (O_1592,N_19743,N_16843);
nor UO_1593 (O_1593,N_19748,N_18801);
or UO_1594 (O_1594,N_17262,N_19960);
and UO_1595 (O_1595,N_17074,N_18319);
xor UO_1596 (O_1596,N_17606,N_16406);
nor UO_1597 (O_1597,N_18808,N_17003);
or UO_1598 (O_1598,N_16373,N_18067);
or UO_1599 (O_1599,N_17792,N_19035);
or UO_1600 (O_1600,N_19560,N_16905);
and UO_1601 (O_1601,N_17043,N_19413);
nand UO_1602 (O_1602,N_17783,N_18378);
nor UO_1603 (O_1603,N_19189,N_19249);
or UO_1604 (O_1604,N_16485,N_17204);
nor UO_1605 (O_1605,N_19597,N_17044);
and UO_1606 (O_1606,N_18817,N_18514);
nor UO_1607 (O_1607,N_16664,N_18922);
nor UO_1608 (O_1608,N_16109,N_18697);
and UO_1609 (O_1609,N_17510,N_18615);
or UO_1610 (O_1610,N_18078,N_17399);
xor UO_1611 (O_1611,N_18671,N_17261);
or UO_1612 (O_1612,N_16069,N_19098);
xor UO_1613 (O_1613,N_17840,N_18880);
xnor UO_1614 (O_1614,N_19365,N_16310);
or UO_1615 (O_1615,N_19704,N_18012);
nor UO_1616 (O_1616,N_19791,N_16184);
xor UO_1617 (O_1617,N_16537,N_16309);
xnor UO_1618 (O_1618,N_18580,N_19626);
nor UO_1619 (O_1619,N_19411,N_17830);
or UO_1620 (O_1620,N_19008,N_19447);
or UO_1621 (O_1621,N_16864,N_19515);
nor UO_1622 (O_1622,N_19595,N_18910);
nor UO_1623 (O_1623,N_18751,N_17506);
and UO_1624 (O_1624,N_17328,N_19227);
nor UO_1625 (O_1625,N_18873,N_17490);
nand UO_1626 (O_1626,N_16254,N_16288);
and UO_1627 (O_1627,N_18966,N_19462);
nand UO_1628 (O_1628,N_19137,N_16174);
nand UO_1629 (O_1629,N_19545,N_17921);
and UO_1630 (O_1630,N_19745,N_19082);
or UO_1631 (O_1631,N_17400,N_16531);
and UO_1632 (O_1632,N_16099,N_16010);
nor UO_1633 (O_1633,N_18143,N_18299);
or UO_1634 (O_1634,N_16962,N_17975);
nor UO_1635 (O_1635,N_17534,N_16812);
nand UO_1636 (O_1636,N_18207,N_18465);
and UO_1637 (O_1637,N_19792,N_16354);
or UO_1638 (O_1638,N_17977,N_17997);
or UO_1639 (O_1639,N_16758,N_18192);
and UO_1640 (O_1640,N_18334,N_17917);
xnor UO_1641 (O_1641,N_17770,N_18463);
and UO_1642 (O_1642,N_17162,N_16886);
xnor UO_1643 (O_1643,N_18682,N_16593);
nand UO_1644 (O_1644,N_17839,N_18618);
nor UO_1645 (O_1645,N_17224,N_19147);
and UO_1646 (O_1646,N_16711,N_16297);
and UO_1647 (O_1647,N_17676,N_16628);
xor UO_1648 (O_1648,N_17522,N_18705);
nor UO_1649 (O_1649,N_16690,N_18244);
xnor UO_1650 (O_1650,N_17630,N_19107);
and UO_1651 (O_1651,N_17649,N_18276);
nor UO_1652 (O_1652,N_16847,N_17403);
xnor UO_1653 (O_1653,N_17690,N_16829);
xor UO_1654 (O_1654,N_16476,N_17616);
and UO_1655 (O_1655,N_16995,N_19011);
xnor UO_1656 (O_1656,N_18895,N_19437);
xor UO_1657 (O_1657,N_18924,N_16451);
nor UO_1658 (O_1658,N_17882,N_17385);
or UO_1659 (O_1659,N_17030,N_19985);
nor UO_1660 (O_1660,N_18591,N_16609);
nor UO_1661 (O_1661,N_18909,N_16262);
xor UO_1662 (O_1662,N_17960,N_19167);
or UO_1663 (O_1663,N_19735,N_18446);
nand UO_1664 (O_1664,N_16311,N_16746);
and UO_1665 (O_1665,N_18797,N_17520);
nor UO_1666 (O_1666,N_19314,N_18972);
nor UO_1667 (O_1667,N_17527,N_16085);
nand UO_1668 (O_1668,N_17335,N_17108);
or UO_1669 (O_1669,N_16534,N_18504);
xnor UO_1670 (O_1670,N_17482,N_19045);
and UO_1671 (O_1671,N_17859,N_19921);
or UO_1672 (O_1672,N_19592,N_19541);
nand UO_1673 (O_1673,N_17474,N_17476);
nor UO_1674 (O_1674,N_18246,N_18864);
nor UO_1675 (O_1675,N_19018,N_16999);
nor UO_1676 (O_1676,N_17093,N_19965);
xnor UO_1677 (O_1677,N_19214,N_17653);
nand UO_1678 (O_1678,N_19899,N_18069);
nor UO_1679 (O_1679,N_19207,N_19293);
nor UO_1680 (O_1680,N_17232,N_19669);
nor UO_1681 (O_1681,N_17814,N_19075);
nand UO_1682 (O_1682,N_19204,N_19526);
and UO_1683 (O_1683,N_19934,N_19577);
xor UO_1684 (O_1684,N_18579,N_17904);
and UO_1685 (O_1685,N_17185,N_19055);
and UO_1686 (O_1686,N_18229,N_16569);
nor UO_1687 (O_1687,N_18987,N_17272);
or UO_1688 (O_1688,N_18224,N_18020);
or UO_1689 (O_1689,N_18789,N_19023);
nor UO_1690 (O_1690,N_18160,N_18823);
nor UO_1691 (O_1691,N_18503,N_19914);
nor UO_1692 (O_1692,N_17320,N_16151);
or UO_1693 (O_1693,N_18691,N_18169);
xor UO_1694 (O_1694,N_19845,N_16182);
nand UO_1695 (O_1695,N_18075,N_17515);
nand UO_1696 (O_1696,N_18994,N_19928);
or UO_1697 (O_1697,N_18238,N_18989);
nor UO_1698 (O_1698,N_19564,N_16799);
or UO_1699 (O_1699,N_19248,N_19420);
and UO_1700 (O_1700,N_18794,N_18681);
xor UO_1701 (O_1701,N_19028,N_16137);
xnor UO_1702 (O_1702,N_19100,N_16859);
nand UO_1703 (O_1703,N_17264,N_17214);
xor UO_1704 (O_1704,N_17438,N_18957);
or UO_1705 (O_1705,N_18790,N_17124);
nand UO_1706 (O_1706,N_18275,N_16235);
xor UO_1707 (O_1707,N_18260,N_16385);
nand UO_1708 (O_1708,N_18528,N_16558);
xor UO_1709 (O_1709,N_18720,N_17072);
nor UO_1710 (O_1710,N_18598,N_16488);
and UO_1711 (O_1711,N_19993,N_16638);
nand UO_1712 (O_1712,N_16739,N_19402);
xor UO_1713 (O_1713,N_18047,N_18251);
nor UO_1714 (O_1714,N_16170,N_19175);
or UO_1715 (O_1715,N_19601,N_17979);
nand UO_1716 (O_1716,N_18058,N_18593);
nand UO_1717 (O_1717,N_18433,N_18457);
xnor UO_1718 (O_1718,N_19390,N_19692);
xnor UO_1719 (O_1719,N_17906,N_17321);
nor UO_1720 (O_1720,N_17433,N_18559);
and UO_1721 (O_1721,N_17464,N_16781);
nand UO_1722 (O_1722,N_18214,N_17020);
and UO_1723 (O_1723,N_19231,N_19866);
nand UO_1724 (O_1724,N_16413,N_19999);
nor UO_1725 (O_1725,N_19664,N_17364);
or UO_1726 (O_1726,N_18855,N_18793);
nand UO_1727 (O_1727,N_18558,N_16149);
or UO_1728 (O_1728,N_18840,N_19527);
nor UO_1729 (O_1729,N_16788,N_16542);
nand UO_1730 (O_1730,N_17301,N_16889);
nor UO_1731 (O_1731,N_16070,N_17669);
or UO_1732 (O_1732,N_19442,N_17786);
nor UO_1733 (O_1733,N_16409,N_19281);
or UO_1734 (O_1734,N_16134,N_17699);
and UO_1735 (O_1735,N_17793,N_16200);
and UO_1736 (O_1736,N_19406,N_16407);
nand UO_1737 (O_1737,N_19106,N_17715);
or UO_1738 (O_1738,N_18560,N_18998);
and UO_1739 (O_1739,N_18142,N_19135);
or UO_1740 (O_1740,N_17413,N_16402);
xnor UO_1741 (O_1741,N_16442,N_19312);
and UO_1742 (O_1742,N_16668,N_17849);
nor UO_1743 (O_1743,N_19212,N_16863);
and UO_1744 (O_1744,N_16167,N_17719);
xor UO_1745 (O_1745,N_17817,N_16934);
nor UO_1746 (O_1746,N_18951,N_18980);
xor UO_1747 (O_1747,N_18489,N_19198);
xnor UO_1748 (O_1748,N_18954,N_17405);
and UO_1749 (O_1749,N_17253,N_18296);
nand UO_1750 (O_1750,N_18208,N_18082);
or UO_1751 (O_1751,N_19282,N_17563);
xor UO_1752 (O_1752,N_18325,N_19648);
and UO_1753 (O_1753,N_17555,N_17486);
nand UO_1754 (O_1754,N_16868,N_19788);
or UO_1755 (O_1755,N_19507,N_19573);
nor UO_1756 (O_1756,N_16771,N_18833);
and UO_1757 (O_1757,N_17346,N_19888);
nor UO_1758 (O_1758,N_18477,N_18635);
or UO_1759 (O_1759,N_17361,N_16204);
nor UO_1760 (O_1760,N_19481,N_17170);
nor UO_1761 (O_1761,N_18865,N_19795);
and UO_1762 (O_1762,N_17192,N_16959);
xnor UO_1763 (O_1763,N_18845,N_17197);
nor UO_1764 (O_1764,N_18245,N_16734);
xnor UO_1765 (O_1765,N_16971,N_16974);
nor UO_1766 (O_1766,N_16058,N_16034);
and UO_1767 (O_1767,N_17363,N_19441);
nand UO_1768 (O_1768,N_19718,N_16979);
nor UO_1769 (O_1769,N_18382,N_19473);
nand UO_1770 (O_1770,N_19295,N_19818);
and UO_1771 (O_1771,N_17908,N_18824);
xnor UO_1772 (O_1772,N_16511,N_17665);
or UO_1773 (O_1773,N_18829,N_16079);
and UO_1774 (O_1774,N_17883,N_16368);
xor UO_1775 (O_1775,N_16773,N_17096);
nand UO_1776 (O_1776,N_19260,N_19576);
xnor UO_1777 (O_1777,N_16706,N_19408);
xor UO_1778 (O_1778,N_16793,N_16011);
nand UO_1779 (O_1779,N_16443,N_18529);
or UO_1780 (O_1780,N_16512,N_18627);
or UO_1781 (O_1781,N_18268,N_16865);
or UO_1782 (O_1782,N_17375,N_19773);
nand UO_1783 (O_1783,N_16529,N_18226);
or UO_1784 (O_1784,N_19662,N_19991);
or UO_1785 (O_1785,N_16970,N_16348);
xnor UO_1786 (O_1786,N_18985,N_17724);
nand UO_1787 (O_1787,N_18018,N_16670);
xor UO_1788 (O_1788,N_17682,N_18371);
xor UO_1789 (O_1789,N_17598,N_17697);
nor UO_1790 (O_1790,N_17824,N_16902);
or UO_1791 (O_1791,N_18189,N_17726);
nand UO_1792 (O_1792,N_19091,N_17909);
nor UO_1793 (O_1793,N_17512,N_18227);
and UO_1794 (O_1794,N_17704,N_19015);
nor UO_1795 (O_1795,N_19849,N_19436);
or UO_1796 (O_1796,N_16497,N_19968);
xor UO_1797 (O_1797,N_18807,N_19629);
nand UO_1798 (O_1798,N_16291,N_17114);
xor UO_1799 (O_1799,N_16228,N_16731);
nor UO_1800 (O_1800,N_18092,N_19761);
nand UO_1801 (O_1801,N_17599,N_19740);
nand UO_1802 (O_1802,N_18091,N_17593);
xor UO_1803 (O_1803,N_16700,N_16029);
or UO_1804 (O_1804,N_18332,N_17300);
xnor UO_1805 (O_1805,N_16876,N_16243);
and UO_1806 (O_1806,N_16146,N_17722);
or UO_1807 (O_1807,N_18141,N_18206);
xor UO_1808 (O_1808,N_16030,N_16658);
nand UO_1809 (O_1809,N_18473,N_17278);
and UO_1810 (O_1810,N_18068,N_19225);
nor UO_1811 (O_1811,N_19835,N_16600);
nor UO_1812 (O_1812,N_19414,N_16942);
xor UO_1813 (O_1813,N_16222,N_18988);
nor UO_1814 (O_1814,N_18639,N_17065);
or UO_1815 (O_1815,N_17116,N_19475);
or UO_1816 (O_1816,N_18359,N_17243);
nand UO_1817 (O_1817,N_19330,N_17907);
and UO_1818 (O_1818,N_18108,N_16367);
or UO_1819 (O_1819,N_19477,N_19728);
and UO_1820 (O_1820,N_17847,N_18009);
xor UO_1821 (O_1821,N_17079,N_18902);
nand UO_1822 (O_1822,N_19779,N_18393);
xor UO_1823 (O_1823,N_17449,N_17275);
nand UO_1824 (O_1824,N_18543,N_16323);
nor UO_1825 (O_1825,N_18525,N_16765);
nand UO_1826 (O_1826,N_16804,N_16986);
or UO_1827 (O_1827,N_19457,N_17735);
or UO_1828 (O_1828,N_17184,N_19193);
and UO_1829 (O_1829,N_17014,N_19852);
nor UO_1830 (O_1830,N_18423,N_16640);
xnor UO_1831 (O_1831,N_18696,N_16219);
and UO_1832 (O_1832,N_17874,N_18933);
nand UO_1833 (O_1833,N_19307,N_17410);
and UO_1834 (O_1834,N_17585,N_18488);
nor UO_1835 (O_1835,N_16361,N_16263);
xnor UO_1836 (O_1836,N_18535,N_18175);
or UO_1837 (O_1837,N_18501,N_19753);
nand UO_1838 (O_1838,N_18264,N_19216);
nor UO_1839 (O_1839,N_16458,N_17488);
nand UO_1840 (O_1840,N_16472,N_17600);
and UO_1841 (O_1841,N_17890,N_17523);
and UO_1842 (O_1842,N_16862,N_19334);
nor UO_1843 (O_1843,N_16818,N_16192);
or UO_1844 (O_1844,N_19088,N_16920);
or UO_1845 (O_1845,N_19201,N_18335);
and UO_1846 (O_1846,N_18134,N_18568);
xor UO_1847 (O_1847,N_17059,N_16063);
nor UO_1848 (O_1848,N_19778,N_18919);
nand UO_1849 (O_1849,N_19247,N_16989);
or UO_1850 (O_1850,N_17459,N_19610);
and UO_1851 (O_1851,N_17807,N_17496);
xnor UO_1852 (O_1852,N_16014,N_16502);
or UO_1853 (O_1853,N_17544,N_18284);
and UO_1854 (O_1854,N_17777,N_16489);
nor UO_1855 (O_1855,N_18848,N_18950);
nand UO_1856 (O_1856,N_18071,N_18636);
nor UO_1857 (O_1857,N_16396,N_18607);
xor UO_1858 (O_1858,N_18523,N_18137);
or UO_1859 (O_1859,N_19611,N_16333);
nor UO_1860 (O_1860,N_17951,N_19782);
nor UO_1861 (O_1861,N_17841,N_18570);
nand UO_1862 (O_1862,N_16261,N_17342);
and UO_1863 (O_1863,N_19151,N_16901);
xnor UO_1864 (O_1864,N_18095,N_19223);
xor UO_1865 (O_1865,N_17421,N_16678);
nand UO_1866 (O_1866,N_17818,N_19257);
or UO_1867 (O_1867,N_16278,N_16211);
nor UO_1868 (O_1868,N_19908,N_19096);
and UO_1869 (O_1869,N_16950,N_17595);
or UO_1870 (O_1870,N_18057,N_16042);
nor UO_1871 (O_1871,N_19513,N_17010);
or UO_1872 (O_1872,N_19827,N_18732);
nor UO_1873 (O_1873,N_18858,N_17755);
and UO_1874 (O_1874,N_16696,N_18006);
xor UO_1875 (O_1875,N_16256,N_18231);
or UO_1876 (O_1876,N_17466,N_16575);
and UO_1877 (O_1877,N_16467,N_17140);
or UO_1878 (O_1878,N_19984,N_18605);
nand UO_1879 (O_1879,N_17475,N_18555);
nand UO_1880 (O_1880,N_19673,N_16840);
nor UO_1881 (O_1881,N_18262,N_18747);
nor UO_1882 (O_1882,N_16727,N_16189);
and UO_1883 (O_1883,N_18349,N_19535);
nand UO_1884 (O_1884,N_19158,N_17091);
nand UO_1885 (O_1885,N_19688,N_19911);
xnor UO_1886 (O_1886,N_18176,N_18884);
and UO_1887 (O_1887,N_17135,N_19039);
nand UO_1888 (O_1888,N_18439,N_16577);
and UO_1889 (O_1889,N_17498,N_16837);
nand UO_1890 (O_1890,N_17784,N_17910);
xor UO_1891 (O_1891,N_16834,N_16925);
and UO_1892 (O_1892,N_19563,N_17668);
or UO_1893 (O_1893,N_19938,N_17416);
xor UO_1894 (O_1894,N_17547,N_18487);
nand UO_1895 (O_1895,N_18365,N_17411);
or UO_1896 (O_1896,N_19209,N_16551);
or UO_1897 (O_1897,N_18358,N_18788);
nor UO_1898 (O_1898,N_16898,N_17460);
and UO_1899 (O_1899,N_19164,N_16510);
or UO_1900 (O_1900,N_16086,N_18695);
nor UO_1901 (O_1901,N_16466,N_19043);
and UO_1902 (O_1902,N_18187,N_19506);
nor UO_1903 (O_1903,N_19690,N_18304);
and UO_1904 (O_1904,N_16503,N_18722);
and UO_1905 (O_1905,N_17260,N_19422);
nand UO_1906 (O_1906,N_18885,N_19269);
nand UO_1907 (O_1907,N_16437,N_17885);
nand UO_1908 (O_1908,N_18685,N_16429);
nor UO_1909 (O_1909,N_16459,N_19361);
nand UO_1910 (O_1910,N_17128,N_16839);
or UO_1911 (O_1911,N_16483,N_18699);
or UO_1912 (O_1912,N_17935,N_17920);
or UO_1913 (O_1913,N_18567,N_18621);
xor UO_1914 (O_1914,N_16439,N_16618);
xnor UO_1915 (O_1915,N_16048,N_19478);
or UO_1916 (O_1916,N_19344,N_18544);
nand UO_1917 (O_1917,N_17892,N_19430);
nand UO_1918 (O_1918,N_17950,N_16124);
nand UO_1919 (O_1919,N_16305,N_18970);
xnor UO_1920 (O_1920,N_17620,N_16712);
nor UO_1921 (O_1921,N_18326,N_19006);
xor UO_1922 (O_1922,N_18573,N_18508);
or UO_1923 (O_1923,N_19685,N_19935);
nand UO_1924 (O_1924,N_16082,N_17280);
and UO_1925 (O_1925,N_19744,N_16160);
and UO_1926 (O_1926,N_17663,N_19553);
or UO_1927 (O_1927,N_17202,N_19244);
xnor UO_1928 (O_1928,N_18893,N_18867);
and UO_1929 (O_1929,N_18748,N_16977);
xnor UO_1930 (O_1930,N_17652,N_18306);
nand UO_1931 (O_1931,N_19119,N_17186);
nor UO_1932 (O_1932,N_17023,N_18308);
xnor UO_1933 (O_1933,N_19858,N_18030);
nor UO_1934 (O_1934,N_16933,N_16826);
or UO_1935 (O_1935,N_19684,N_18063);
xor UO_1936 (O_1936,N_19801,N_16882);
nand UO_1937 (O_1937,N_17247,N_17788);
nand UO_1938 (O_1938,N_19598,N_16883);
or UO_1939 (O_1939,N_16814,N_19589);
xnor UO_1940 (O_1940,N_18900,N_18847);
nor UO_1941 (O_1941,N_19279,N_16390);
nand UO_1942 (O_1942,N_17623,N_17899);
or UO_1943 (O_1943,N_16415,N_17983);
nand UO_1944 (O_1944,N_19079,N_16599);
nand UO_1945 (O_1945,N_17501,N_18674);
xnor UO_1946 (O_1946,N_19974,N_18387);
and UO_1947 (O_1947,N_19364,N_19340);
or UO_1948 (O_1948,N_17992,N_16169);
or UO_1949 (O_1949,N_19132,N_19864);
xor UO_1950 (O_1950,N_18402,N_19813);
nand UO_1951 (O_1951,N_19210,N_17750);
nand UO_1952 (O_1952,N_18086,N_17763);
xor UO_1953 (O_1953,N_17191,N_16339);
nor UO_1954 (O_1954,N_16239,N_17440);
and UO_1955 (O_1955,N_16398,N_18601);
nor UO_1956 (O_1956,N_19083,N_19046);
nor UO_1957 (O_1957,N_18967,N_19902);
nand UO_1958 (O_1958,N_18765,N_18658);
and UO_1959 (O_1959,N_17122,N_16133);
nand UO_1960 (O_1960,N_16741,N_19337);
nand UO_1961 (O_1961,N_19182,N_16513);
and UO_1962 (O_1962,N_17062,N_16963);
or UO_1963 (O_1963,N_17290,N_17861);
and UO_1964 (O_1964,N_16152,N_19169);
nor UO_1965 (O_1965,N_16044,N_18689);
xor UO_1966 (O_1966,N_18585,N_17391);
or UO_1967 (O_1967,N_18582,N_18907);
or UO_1968 (O_1968,N_16389,N_18556);
or UO_1969 (O_1969,N_18859,N_17551);
or UO_1970 (O_1970,N_18936,N_17242);
nor UO_1971 (O_1971,N_16232,N_19832);
and UO_1972 (O_1972,N_19929,N_17318);
or UO_1973 (O_1973,N_19264,N_17434);
nor UO_1974 (O_1974,N_16129,N_19042);
nand UO_1975 (O_1975,N_16103,N_19596);
and UO_1976 (O_1976,N_19821,N_18253);
or UO_1977 (O_1977,N_18261,N_19861);
xnor UO_1978 (O_1978,N_19362,N_17353);
and UO_1979 (O_1979,N_19078,N_18026);
and UO_1980 (O_1980,N_17545,N_17033);
xnor UO_1981 (O_1981,N_19332,N_19285);
or UO_1982 (O_1982,N_18594,N_16820);
or UO_1983 (O_1983,N_17800,N_16332);
nand UO_1984 (O_1984,N_16594,N_16207);
and UO_1985 (O_1985,N_19063,N_18974);
and UO_1986 (O_1986,N_17166,N_19316);
and UO_1987 (O_1987,N_17164,N_16400);
nor UO_1988 (O_1988,N_16689,N_19839);
or UO_1989 (O_1989,N_18013,N_19508);
nor UO_1990 (O_1990,N_19489,N_19880);
or UO_1991 (O_1991,N_17359,N_18772);
xnor UO_1992 (O_1992,N_18516,N_16244);
xor UO_1993 (O_1993,N_18413,N_17076);
xnor UO_1994 (O_1994,N_17196,N_17089);
or UO_1995 (O_1995,N_16157,N_18049);
nand UO_1996 (O_1996,N_17472,N_16702);
nand UO_1997 (O_1997,N_19352,N_19271);
or UO_1998 (O_1998,N_16017,N_18209);
and UO_1999 (O_1999,N_17893,N_16083);
and UO_2000 (O_2000,N_17271,N_16795);
nor UO_2001 (O_2001,N_17143,N_16990);
and UO_2002 (O_2002,N_18099,N_17388);
nor UO_2003 (O_2003,N_16864,N_17515);
or UO_2004 (O_2004,N_19145,N_18975);
and UO_2005 (O_2005,N_18910,N_16256);
xor UO_2006 (O_2006,N_17224,N_19988);
nor UO_2007 (O_2007,N_18396,N_16061);
nor UO_2008 (O_2008,N_18980,N_18029);
nor UO_2009 (O_2009,N_17676,N_18519);
xor UO_2010 (O_2010,N_18915,N_16807);
nor UO_2011 (O_2011,N_16764,N_16721);
nor UO_2012 (O_2012,N_19960,N_19455);
nor UO_2013 (O_2013,N_19942,N_16545);
and UO_2014 (O_2014,N_17778,N_16875);
xor UO_2015 (O_2015,N_18789,N_19045);
or UO_2016 (O_2016,N_19948,N_16643);
or UO_2017 (O_2017,N_16088,N_19931);
and UO_2018 (O_2018,N_19037,N_16326);
xnor UO_2019 (O_2019,N_16676,N_17384);
or UO_2020 (O_2020,N_18316,N_18187);
xnor UO_2021 (O_2021,N_16103,N_18574);
nor UO_2022 (O_2022,N_17193,N_17839);
nand UO_2023 (O_2023,N_18646,N_18846);
and UO_2024 (O_2024,N_16379,N_16786);
or UO_2025 (O_2025,N_19444,N_18604);
xor UO_2026 (O_2026,N_18403,N_17063);
nand UO_2027 (O_2027,N_19863,N_19699);
nand UO_2028 (O_2028,N_17929,N_17614);
or UO_2029 (O_2029,N_19843,N_18993);
xnor UO_2030 (O_2030,N_18986,N_18188);
xnor UO_2031 (O_2031,N_19573,N_18101);
or UO_2032 (O_2032,N_18477,N_17148);
nor UO_2033 (O_2033,N_17554,N_19597);
nor UO_2034 (O_2034,N_19671,N_17893);
and UO_2035 (O_2035,N_16673,N_18507);
xor UO_2036 (O_2036,N_18835,N_19725);
or UO_2037 (O_2037,N_16833,N_17593);
and UO_2038 (O_2038,N_19665,N_19622);
or UO_2039 (O_2039,N_19517,N_17709);
or UO_2040 (O_2040,N_16356,N_19762);
xor UO_2041 (O_2041,N_16604,N_17638);
nor UO_2042 (O_2042,N_18733,N_18086);
and UO_2043 (O_2043,N_19737,N_18711);
or UO_2044 (O_2044,N_16593,N_18404);
nor UO_2045 (O_2045,N_19111,N_19426);
nor UO_2046 (O_2046,N_17180,N_16426);
nand UO_2047 (O_2047,N_16613,N_16077);
xnor UO_2048 (O_2048,N_19551,N_19097);
nand UO_2049 (O_2049,N_16832,N_18853);
or UO_2050 (O_2050,N_19665,N_19750);
xnor UO_2051 (O_2051,N_19861,N_17681);
xnor UO_2052 (O_2052,N_16305,N_16067);
nor UO_2053 (O_2053,N_19709,N_17431);
or UO_2054 (O_2054,N_17754,N_19899);
or UO_2055 (O_2055,N_17493,N_18762);
nand UO_2056 (O_2056,N_19804,N_18028);
or UO_2057 (O_2057,N_16391,N_17915);
nor UO_2058 (O_2058,N_18969,N_19302);
xor UO_2059 (O_2059,N_18441,N_18296);
or UO_2060 (O_2060,N_18740,N_16382);
or UO_2061 (O_2061,N_18750,N_18110);
and UO_2062 (O_2062,N_16860,N_18449);
nor UO_2063 (O_2063,N_19837,N_16955);
xnor UO_2064 (O_2064,N_18536,N_19935);
nor UO_2065 (O_2065,N_19341,N_18442);
and UO_2066 (O_2066,N_17822,N_18682);
or UO_2067 (O_2067,N_18186,N_18242);
and UO_2068 (O_2068,N_18198,N_19472);
and UO_2069 (O_2069,N_18474,N_18301);
and UO_2070 (O_2070,N_17331,N_16275);
and UO_2071 (O_2071,N_16779,N_16374);
or UO_2072 (O_2072,N_16436,N_16155);
nand UO_2073 (O_2073,N_19482,N_18455);
and UO_2074 (O_2074,N_16323,N_17843);
xnor UO_2075 (O_2075,N_19381,N_17884);
or UO_2076 (O_2076,N_17071,N_18023);
nor UO_2077 (O_2077,N_17740,N_17106);
xor UO_2078 (O_2078,N_17094,N_18564);
xnor UO_2079 (O_2079,N_17927,N_17899);
and UO_2080 (O_2080,N_16564,N_19765);
xnor UO_2081 (O_2081,N_19871,N_19994);
nand UO_2082 (O_2082,N_16119,N_16410);
xnor UO_2083 (O_2083,N_16968,N_17972);
nand UO_2084 (O_2084,N_16472,N_18426);
xor UO_2085 (O_2085,N_17640,N_16455);
nand UO_2086 (O_2086,N_16112,N_17286);
or UO_2087 (O_2087,N_18712,N_17136);
or UO_2088 (O_2088,N_19159,N_19632);
xor UO_2089 (O_2089,N_16226,N_18061);
nor UO_2090 (O_2090,N_19239,N_19690);
and UO_2091 (O_2091,N_18158,N_16306);
nor UO_2092 (O_2092,N_19609,N_18445);
nor UO_2093 (O_2093,N_19555,N_16445);
nand UO_2094 (O_2094,N_16880,N_17828);
xor UO_2095 (O_2095,N_17744,N_18629);
or UO_2096 (O_2096,N_19069,N_16378);
xor UO_2097 (O_2097,N_17178,N_16439);
nand UO_2098 (O_2098,N_18660,N_17933);
and UO_2099 (O_2099,N_19662,N_17171);
and UO_2100 (O_2100,N_16909,N_19115);
and UO_2101 (O_2101,N_16660,N_16539);
nor UO_2102 (O_2102,N_16910,N_17337);
or UO_2103 (O_2103,N_16515,N_18405);
nand UO_2104 (O_2104,N_17972,N_18578);
nand UO_2105 (O_2105,N_16961,N_17219);
nor UO_2106 (O_2106,N_16819,N_16817);
and UO_2107 (O_2107,N_18381,N_16829);
xor UO_2108 (O_2108,N_18841,N_16341);
or UO_2109 (O_2109,N_19742,N_16969);
or UO_2110 (O_2110,N_19769,N_19036);
nor UO_2111 (O_2111,N_19606,N_17630);
and UO_2112 (O_2112,N_18139,N_16034);
nand UO_2113 (O_2113,N_17369,N_18057);
and UO_2114 (O_2114,N_16594,N_19088);
and UO_2115 (O_2115,N_18203,N_19158);
and UO_2116 (O_2116,N_19409,N_19169);
nor UO_2117 (O_2117,N_16651,N_18531);
or UO_2118 (O_2118,N_17491,N_19962);
nor UO_2119 (O_2119,N_16036,N_19708);
or UO_2120 (O_2120,N_18817,N_19368);
nand UO_2121 (O_2121,N_17300,N_19378);
nor UO_2122 (O_2122,N_18582,N_17449);
or UO_2123 (O_2123,N_17988,N_16248);
and UO_2124 (O_2124,N_19468,N_19972);
nor UO_2125 (O_2125,N_17417,N_18455);
xor UO_2126 (O_2126,N_18298,N_18982);
or UO_2127 (O_2127,N_16237,N_16020);
nor UO_2128 (O_2128,N_16313,N_16316);
nor UO_2129 (O_2129,N_19854,N_16910);
nand UO_2130 (O_2130,N_18095,N_18196);
xnor UO_2131 (O_2131,N_19572,N_17479);
or UO_2132 (O_2132,N_17814,N_16122);
and UO_2133 (O_2133,N_19098,N_16680);
nor UO_2134 (O_2134,N_16804,N_19411);
or UO_2135 (O_2135,N_18427,N_18578);
nor UO_2136 (O_2136,N_19558,N_17535);
xnor UO_2137 (O_2137,N_17521,N_18431);
xnor UO_2138 (O_2138,N_18382,N_18881);
or UO_2139 (O_2139,N_17470,N_19202);
xnor UO_2140 (O_2140,N_16589,N_17181);
or UO_2141 (O_2141,N_18488,N_18657);
xnor UO_2142 (O_2142,N_17756,N_16106);
nand UO_2143 (O_2143,N_18993,N_19633);
nand UO_2144 (O_2144,N_17483,N_19736);
nor UO_2145 (O_2145,N_18072,N_17969);
and UO_2146 (O_2146,N_17352,N_18580);
xnor UO_2147 (O_2147,N_19449,N_16314);
nor UO_2148 (O_2148,N_18359,N_18904);
and UO_2149 (O_2149,N_18680,N_16268);
and UO_2150 (O_2150,N_16837,N_16121);
nor UO_2151 (O_2151,N_17038,N_17440);
nand UO_2152 (O_2152,N_17409,N_19462);
xor UO_2153 (O_2153,N_16129,N_17532);
nand UO_2154 (O_2154,N_19954,N_16089);
nand UO_2155 (O_2155,N_16947,N_18978);
and UO_2156 (O_2156,N_16960,N_18278);
nor UO_2157 (O_2157,N_18736,N_16731);
or UO_2158 (O_2158,N_17061,N_16257);
and UO_2159 (O_2159,N_18574,N_18700);
and UO_2160 (O_2160,N_16764,N_18284);
nand UO_2161 (O_2161,N_17637,N_16496);
nand UO_2162 (O_2162,N_18104,N_17801);
nand UO_2163 (O_2163,N_18563,N_16370);
and UO_2164 (O_2164,N_17312,N_17653);
xnor UO_2165 (O_2165,N_18932,N_19745);
nor UO_2166 (O_2166,N_18239,N_18833);
nor UO_2167 (O_2167,N_16734,N_16209);
nand UO_2168 (O_2168,N_19872,N_19373);
xor UO_2169 (O_2169,N_17872,N_19745);
nor UO_2170 (O_2170,N_19558,N_17272);
xor UO_2171 (O_2171,N_16712,N_18142);
xor UO_2172 (O_2172,N_16648,N_16934);
xor UO_2173 (O_2173,N_17628,N_18654);
nand UO_2174 (O_2174,N_18011,N_19614);
nor UO_2175 (O_2175,N_18522,N_18791);
nand UO_2176 (O_2176,N_18771,N_17172);
or UO_2177 (O_2177,N_19853,N_19820);
nand UO_2178 (O_2178,N_18637,N_18047);
or UO_2179 (O_2179,N_18923,N_17135);
nand UO_2180 (O_2180,N_16871,N_17336);
nor UO_2181 (O_2181,N_16777,N_16487);
or UO_2182 (O_2182,N_16895,N_18786);
xnor UO_2183 (O_2183,N_19243,N_17450);
xor UO_2184 (O_2184,N_18143,N_16525);
and UO_2185 (O_2185,N_18046,N_17091);
or UO_2186 (O_2186,N_19605,N_16307);
or UO_2187 (O_2187,N_19505,N_18217);
or UO_2188 (O_2188,N_18725,N_16815);
xnor UO_2189 (O_2189,N_18473,N_17775);
nand UO_2190 (O_2190,N_18601,N_18684);
nand UO_2191 (O_2191,N_16724,N_16802);
or UO_2192 (O_2192,N_18824,N_18831);
or UO_2193 (O_2193,N_18540,N_19534);
nand UO_2194 (O_2194,N_19714,N_17373);
xnor UO_2195 (O_2195,N_16509,N_19023);
and UO_2196 (O_2196,N_17466,N_16692);
or UO_2197 (O_2197,N_18281,N_16715);
xor UO_2198 (O_2198,N_18301,N_19197);
or UO_2199 (O_2199,N_19955,N_18747);
nand UO_2200 (O_2200,N_18582,N_17780);
or UO_2201 (O_2201,N_16033,N_16575);
xnor UO_2202 (O_2202,N_16345,N_19463);
nor UO_2203 (O_2203,N_18030,N_19271);
nand UO_2204 (O_2204,N_16685,N_16663);
and UO_2205 (O_2205,N_16234,N_19585);
or UO_2206 (O_2206,N_16678,N_17242);
nand UO_2207 (O_2207,N_19947,N_18532);
nor UO_2208 (O_2208,N_17007,N_18346);
xnor UO_2209 (O_2209,N_17200,N_16169);
and UO_2210 (O_2210,N_19823,N_19170);
xnor UO_2211 (O_2211,N_16462,N_19328);
or UO_2212 (O_2212,N_16369,N_19300);
and UO_2213 (O_2213,N_18236,N_19864);
nand UO_2214 (O_2214,N_16580,N_17194);
nand UO_2215 (O_2215,N_16988,N_19408);
and UO_2216 (O_2216,N_18495,N_16960);
nor UO_2217 (O_2217,N_16221,N_18689);
nand UO_2218 (O_2218,N_17683,N_18475);
and UO_2219 (O_2219,N_19692,N_16190);
nand UO_2220 (O_2220,N_18025,N_17748);
xnor UO_2221 (O_2221,N_17297,N_17816);
xnor UO_2222 (O_2222,N_18060,N_16668);
nor UO_2223 (O_2223,N_18847,N_17901);
nand UO_2224 (O_2224,N_18914,N_19798);
nor UO_2225 (O_2225,N_19781,N_18851);
nand UO_2226 (O_2226,N_19843,N_18167);
and UO_2227 (O_2227,N_19062,N_17074);
or UO_2228 (O_2228,N_17738,N_17101);
xnor UO_2229 (O_2229,N_17731,N_19292);
or UO_2230 (O_2230,N_16102,N_16359);
nor UO_2231 (O_2231,N_19403,N_16640);
or UO_2232 (O_2232,N_19735,N_18802);
nor UO_2233 (O_2233,N_18281,N_18661);
or UO_2234 (O_2234,N_16886,N_19329);
and UO_2235 (O_2235,N_17372,N_18089);
xnor UO_2236 (O_2236,N_16972,N_19451);
nand UO_2237 (O_2237,N_16450,N_17839);
nand UO_2238 (O_2238,N_18032,N_17371);
nand UO_2239 (O_2239,N_18369,N_18584);
and UO_2240 (O_2240,N_18053,N_16903);
nor UO_2241 (O_2241,N_18348,N_19146);
and UO_2242 (O_2242,N_17129,N_18606);
and UO_2243 (O_2243,N_18211,N_18862);
xnor UO_2244 (O_2244,N_19475,N_19993);
xnor UO_2245 (O_2245,N_17352,N_16157);
or UO_2246 (O_2246,N_18211,N_16541);
xnor UO_2247 (O_2247,N_16552,N_18553);
and UO_2248 (O_2248,N_19424,N_18866);
nand UO_2249 (O_2249,N_19092,N_16301);
xor UO_2250 (O_2250,N_18270,N_19541);
nor UO_2251 (O_2251,N_18567,N_18949);
nand UO_2252 (O_2252,N_18991,N_19662);
or UO_2253 (O_2253,N_17344,N_16118);
xnor UO_2254 (O_2254,N_17327,N_18503);
and UO_2255 (O_2255,N_17037,N_17288);
xor UO_2256 (O_2256,N_17410,N_18269);
nor UO_2257 (O_2257,N_19720,N_19465);
nand UO_2258 (O_2258,N_18071,N_16163);
and UO_2259 (O_2259,N_17404,N_16854);
nand UO_2260 (O_2260,N_19134,N_19448);
and UO_2261 (O_2261,N_19414,N_19221);
or UO_2262 (O_2262,N_19895,N_18412);
xnor UO_2263 (O_2263,N_19080,N_19185);
nand UO_2264 (O_2264,N_17435,N_19181);
and UO_2265 (O_2265,N_19422,N_16265);
nor UO_2266 (O_2266,N_18787,N_17425);
or UO_2267 (O_2267,N_19919,N_19610);
or UO_2268 (O_2268,N_16195,N_16797);
and UO_2269 (O_2269,N_17359,N_19121);
nand UO_2270 (O_2270,N_19278,N_19114);
or UO_2271 (O_2271,N_19452,N_19532);
xor UO_2272 (O_2272,N_16618,N_17032);
nor UO_2273 (O_2273,N_19827,N_17777);
xor UO_2274 (O_2274,N_18635,N_17400);
nand UO_2275 (O_2275,N_17503,N_18135);
and UO_2276 (O_2276,N_18756,N_19516);
and UO_2277 (O_2277,N_19987,N_19594);
nand UO_2278 (O_2278,N_17112,N_16952);
or UO_2279 (O_2279,N_18286,N_18719);
nor UO_2280 (O_2280,N_18607,N_16780);
or UO_2281 (O_2281,N_19130,N_16903);
nand UO_2282 (O_2282,N_19473,N_19844);
nand UO_2283 (O_2283,N_17558,N_16541);
nand UO_2284 (O_2284,N_19610,N_17309);
or UO_2285 (O_2285,N_17968,N_18794);
xnor UO_2286 (O_2286,N_18944,N_16663);
nand UO_2287 (O_2287,N_16102,N_19085);
xnor UO_2288 (O_2288,N_19702,N_19520);
nand UO_2289 (O_2289,N_18353,N_19009);
nor UO_2290 (O_2290,N_18169,N_19949);
nand UO_2291 (O_2291,N_19439,N_18722);
xor UO_2292 (O_2292,N_19199,N_16940);
nand UO_2293 (O_2293,N_16843,N_18157);
nand UO_2294 (O_2294,N_18871,N_18343);
xor UO_2295 (O_2295,N_16823,N_18889);
xor UO_2296 (O_2296,N_16665,N_17467);
nor UO_2297 (O_2297,N_19754,N_16000);
nor UO_2298 (O_2298,N_16737,N_17498);
or UO_2299 (O_2299,N_16310,N_16610);
and UO_2300 (O_2300,N_18737,N_18734);
nand UO_2301 (O_2301,N_19691,N_19829);
nor UO_2302 (O_2302,N_19651,N_18954);
nor UO_2303 (O_2303,N_18974,N_19598);
or UO_2304 (O_2304,N_18936,N_16663);
xnor UO_2305 (O_2305,N_18126,N_19179);
nand UO_2306 (O_2306,N_19021,N_18975);
or UO_2307 (O_2307,N_19167,N_17935);
nor UO_2308 (O_2308,N_17849,N_16735);
nor UO_2309 (O_2309,N_16864,N_16013);
nand UO_2310 (O_2310,N_17174,N_18284);
or UO_2311 (O_2311,N_17500,N_16147);
and UO_2312 (O_2312,N_17311,N_16137);
or UO_2313 (O_2313,N_16469,N_18057);
nor UO_2314 (O_2314,N_19064,N_17408);
nand UO_2315 (O_2315,N_19287,N_16554);
and UO_2316 (O_2316,N_17340,N_16102);
nor UO_2317 (O_2317,N_19334,N_16516);
xor UO_2318 (O_2318,N_19406,N_16305);
and UO_2319 (O_2319,N_19205,N_18607);
and UO_2320 (O_2320,N_19003,N_17635);
and UO_2321 (O_2321,N_17369,N_18456);
or UO_2322 (O_2322,N_17035,N_16625);
nor UO_2323 (O_2323,N_18962,N_19174);
and UO_2324 (O_2324,N_16726,N_19556);
and UO_2325 (O_2325,N_16663,N_18424);
or UO_2326 (O_2326,N_18297,N_17635);
and UO_2327 (O_2327,N_18426,N_16889);
or UO_2328 (O_2328,N_17936,N_18420);
and UO_2329 (O_2329,N_18873,N_17203);
nand UO_2330 (O_2330,N_17576,N_19590);
and UO_2331 (O_2331,N_17819,N_19471);
and UO_2332 (O_2332,N_17061,N_18002);
and UO_2333 (O_2333,N_16145,N_19779);
xnor UO_2334 (O_2334,N_16946,N_17772);
xnor UO_2335 (O_2335,N_17628,N_16303);
or UO_2336 (O_2336,N_18090,N_17143);
nor UO_2337 (O_2337,N_18504,N_19530);
or UO_2338 (O_2338,N_17035,N_17544);
xnor UO_2339 (O_2339,N_19672,N_17817);
xor UO_2340 (O_2340,N_19811,N_18614);
or UO_2341 (O_2341,N_17640,N_17880);
xnor UO_2342 (O_2342,N_16517,N_17278);
xor UO_2343 (O_2343,N_17738,N_18216);
nand UO_2344 (O_2344,N_17952,N_16228);
xnor UO_2345 (O_2345,N_18396,N_19513);
nor UO_2346 (O_2346,N_19182,N_17996);
nand UO_2347 (O_2347,N_18967,N_19717);
xor UO_2348 (O_2348,N_19742,N_16574);
xor UO_2349 (O_2349,N_16862,N_19564);
and UO_2350 (O_2350,N_16824,N_19469);
nor UO_2351 (O_2351,N_19580,N_17300);
nor UO_2352 (O_2352,N_19116,N_19414);
nor UO_2353 (O_2353,N_18379,N_18016);
or UO_2354 (O_2354,N_18375,N_19211);
xor UO_2355 (O_2355,N_16006,N_17291);
nor UO_2356 (O_2356,N_18310,N_18992);
or UO_2357 (O_2357,N_16257,N_19945);
or UO_2358 (O_2358,N_18118,N_16061);
and UO_2359 (O_2359,N_19971,N_17481);
and UO_2360 (O_2360,N_17462,N_16034);
nor UO_2361 (O_2361,N_16034,N_16903);
nand UO_2362 (O_2362,N_19025,N_18721);
nand UO_2363 (O_2363,N_16992,N_16204);
or UO_2364 (O_2364,N_17426,N_16981);
xnor UO_2365 (O_2365,N_17261,N_16164);
or UO_2366 (O_2366,N_16004,N_18775);
nand UO_2367 (O_2367,N_17895,N_17940);
nand UO_2368 (O_2368,N_16327,N_16964);
or UO_2369 (O_2369,N_16983,N_17238);
xor UO_2370 (O_2370,N_18531,N_19601);
nor UO_2371 (O_2371,N_19497,N_17588);
nand UO_2372 (O_2372,N_16419,N_16739);
xor UO_2373 (O_2373,N_16283,N_17048);
and UO_2374 (O_2374,N_16405,N_16134);
xor UO_2375 (O_2375,N_19676,N_19208);
xor UO_2376 (O_2376,N_19949,N_18920);
or UO_2377 (O_2377,N_19403,N_19274);
nand UO_2378 (O_2378,N_19402,N_17679);
nand UO_2379 (O_2379,N_16455,N_17260);
xnor UO_2380 (O_2380,N_16346,N_17516);
xor UO_2381 (O_2381,N_16135,N_17678);
nor UO_2382 (O_2382,N_19729,N_19234);
xnor UO_2383 (O_2383,N_17674,N_19930);
nor UO_2384 (O_2384,N_17355,N_17188);
nand UO_2385 (O_2385,N_18129,N_18446);
nor UO_2386 (O_2386,N_17669,N_16317);
and UO_2387 (O_2387,N_17929,N_16944);
nand UO_2388 (O_2388,N_17695,N_19071);
or UO_2389 (O_2389,N_16147,N_18923);
nand UO_2390 (O_2390,N_16038,N_16712);
nand UO_2391 (O_2391,N_19008,N_19619);
xor UO_2392 (O_2392,N_19252,N_19690);
nor UO_2393 (O_2393,N_17474,N_16703);
nor UO_2394 (O_2394,N_18604,N_17655);
nor UO_2395 (O_2395,N_18047,N_16854);
nand UO_2396 (O_2396,N_18455,N_18877);
xor UO_2397 (O_2397,N_18901,N_16896);
nor UO_2398 (O_2398,N_19376,N_19968);
nor UO_2399 (O_2399,N_18424,N_18694);
or UO_2400 (O_2400,N_19207,N_16178);
and UO_2401 (O_2401,N_17614,N_18591);
or UO_2402 (O_2402,N_18524,N_19434);
xnor UO_2403 (O_2403,N_19021,N_16072);
nand UO_2404 (O_2404,N_19114,N_19221);
xnor UO_2405 (O_2405,N_19592,N_19080);
nor UO_2406 (O_2406,N_17657,N_17570);
nand UO_2407 (O_2407,N_18083,N_19107);
nor UO_2408 (O_2408,N_18207,N_17870);
and UO_2409 (O_2409,N_19547,N_18721);
xor UO_2410 (O_2410,N_19310,N_18644);
or UO_2411 (O_2411,N_17971,N_19246);
or UO_2412 (O_2412,N_16320,N_16986);
xnor UO_2413 (O_2413,N_16093,N_19420);
nand UO_2414 (O_2414,N_17344,N_16117);
or UO_2415 (O_2415,N_17261,N_16730);
xnor UO_2416 (O_2416,N_17496,N_18822);
nand UO_2417 (O_2417,N_19647,N_19521);
nor UO_2418 (O_2418,N_19689,N_19543);
nor UO_2419 (O_2419,N_16935,N_18039);
or UO_2420 (O_2420,N_18506,N_18877);
or UO_2421 (O_2421,N_18852,N_17262);
and UO_2422 (O_2422,N_17137,N_17406);
xnor UO_2423 (O_2423,N_19539,N_18788);
nor UO_2424 (O_2424,N_18269,N_16941);
and UO_2425 (O_2425,N_17525,N_16789);
and UO_2426 (O_2426,N_18445,N_16765);
xor UO_2427 (O_2427,N_18495,N_17778);
or UO_2428 (O_2428,N_17943,N_16982);
nand UO_2429 (O_2429,N_18106,N_19574);
xnor UO_2430 (O_2430,N_18049,N_17382);
or UO_2431 (O_2431,N_17410,N_16593);
nor UO_2432 (O_2432,N_17860,N_16038);
and UO_2433 (O_2433,N_17801,N_18655);
nor UO_2434 (O_2434,N_16362,N_19155);
xor UO_2435 (O_2435,N_17279,N_18853);
xor UO_2436 (O_2436,N_18681,N_19743);
nand UO_2437 (O_2437,N_19108,N_17933);
and UO_2438 (O_2438,N_19500,N_18139);
nor UO_2439 (O_2439,N_18862,N_17452);
xor UO_2440 (O_2440,N_17819,N_16283);
nor UO_2441 (O_2441,N_17612,N_19170);
nor UO_2442 (O_2442,N_17899,N_19984);
and UO_2443 (O_2443,N_16481,N_19738);
and UO_2444 (O_2444,N_19419,N_18205);
xor UO_2445 (O_2445,N_17615,N_17697);
xnor UO_2446 (O_2446,N_16456,N_17660);
xnor UO_2447 (O_2447,N_18428,N_18501);
nor UO_2448 (O_2448,N_16797,N_18453);
nand UO_2449 (O_2449,N_18962,N_19972);
nand UO_2450 (O_2450,N_19329,N_19467);
or UO_2451 (O_2451,N_19145,N_16961);
nand UO_2452 (O_2452,N_18471,N_19612);
nand UO_2453 (O_2453,N_16857,N_17245);
or UO_2454 (O_2454,N_18614,N_19205);
nand UO_2455 (O_2455,N_18487,N_19130);
or UO_2456 (O_2456,N_16130,N_16177);
and UO_2457 (O_2457,N_17581,N_17594);
xor UO_2458 (O_2458,N_17994,N_19517);
xnor UO_2459 (O_2459,N_17102,N_19346);
nor UO_2460 (O_2460,N_18806,N_16403);
nor UO_2461 (O_2461,N_19058,N_17016);
nor UO_2462 (O_2462,N_17484,N_19525);
xnor UO_2463 (O_2463,N_19571,N_17630);
and UO_2464 (O_2464,N_16217,N_19407);
nand UO_2465 (O_2465,N_16421,N_16565);
xor UO_2466 (O_2466,N_19916,N_18308);
xnor UO_2467 (O_2467,N_16177,N_19037);
and UO_2468 (O_2468,N_18179,N_16215);
nand UO_2469 (O_2469,N_18625,N_17417);
nand UO_2470 (O_2470,N_17788,N_18427);
or UO_2471 (O_2471,N_19288,N_18094);
and UO_2472 (O_2472,N_17393,N_18434);
xnor UO_2473 (O_2473,N_18367,N_17415);
xor UO_2474 (O_2474,N_18081,N_16826);
or UO_2475 (O_2475,N_19600,N_18304);
nor UO_2476 (O_2476,N_19354,N_17024);
nor UO_2477 (O_2477,N_17916,N_16004);
nand UO_2478 (O_2478,N_17764,N_18174);
and UO_2479 (O_2479,N_19348,N_19392);
nand UO_2480 (O_2480,N_18530,N_16744);
xnor UO_2481 (O_2481,N_16537,N_17826);
and UO_2482 (O_2482,N_16774,N_17819);
or UO_2483 (O_2483,N_18939,N_17648);
nor UO_2484 (O_2484,N_17135,N_18009);
nand UO_2485 (O_2485,N_17128,N_19640);
and UO_2486 (O_2486,N_18572,N_19011);
nor UO_2487 (O_2487,N_19445,N_19634);
and UO_2488 (O_2488,N_19148,N_16378);
xnor UO_2489 (O_2489,N_18140,N_17100);
or UO_2490 (O_2490,N_17534,N_17521);
and UO_2491 (O_2491,N_18643,N_16575);
or UO_2492 (O_2492,N_19443,N_18315);
and UO_2493 (O_2493,N_17724,N_16739);
nor UO_2494 (O_2494,N_16572,N_17860);
xnor UO_2495 (O_2495,N_16839,N_18235);
nor UO_2496 (O_2496,N_19880,N_18364);
and UO_2497 (O_2497,N_19961,N_16681);
nand UO_2498 (O_2498,N_18789,N_19210);
nand UO_2499 (O_2499,N_16395,N_19691);
endmodule