module basic_3000_30000_3500_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_2800,In_2418);
or U1 (N_1,In_1704,In_2818);
xor U2 (N_2,In_2788,In_1771);
nand U3 (N_3,In_2178,In_703);
and U4 (N_4,In_1807,In_1229);
nor U5 (N_5,In_310,In_1431);
xnor U6 (N_6,In_210,In_2291);
or U7 (N_7,In_284,In_1866);
nand U8 (N_8,In_1044,In_1976);
nor U9 (N_9,In_1712,In_2652);
or U10 (N_10,In_1565,In_2315);
xnor U11 (N_11,In_713,In_2486);
nand U12 (N_12,In_1908,In_2298);
or U13 (N_13,In_653,In_2766);
or U14 (N_14,In_1511,In_2245);
nor U15 (N_15,In_574,In_1102);
nand U16 (N_16,In_1223,In_171);
xnor U17 (N_17,In_61,In_763);
nor U18 (N_18,In_2757,In_2600);
or U19 (N_19,In_329,In_618);
xor U20 (N_20,In_971,In_247);
and U21 (N_21,In_1330,In_532);
and U22 (N_22,In_2306,In_997);
and U23 (N_23,In_2344,In_590);
xor U24 (N_24,In_1854,In_2759);
and U25 (N_25,In_1774,In_119);
and U26 (N_26,In_641,In_2790);
or U27 (N_27,In_2347,In_2176);
and U28 (N_28,In_133,In_2712);
nand U29 (N_29,In_1245,In_593);
or U30 (N_30,In_1574,In_963);
and U31 (N_31,In_1715,In_475);
nor U32 (N_32,In_2342,In_792);
and U33 (N_33,In_968,In_2743);
or U34 (N_34,In_67,In_880);
nor U35 (N_35,In_2936,In_1372);
nor U36 (N_36,In_366,In_2067);
nand U37 (N_37,In_12,In_1040);
nor U38 (N_38,In_2762,In_1210);
xor U39 (N_39,In_510,In_2475);
or U40 (N_40,In_665,In_414);
nor U41 (N_41,In_1277,In_2419);
nand U42 (N_42,In_2211,In_422);
nand U43 (N_43,In_1031,In_160);
or U44 (N_44,In_634,In_1775);
xnor U45 (N_45,In_1512,In_1247);
nand U46 (N_46,In_1527,In_798);
xnor U47 (N_47,In_2625,In_1256);
or U48 (N_48,In_251,In_1241);
or U49 (N_49,In_636,In_996);
nor U50 (N_50,In_2927,In_1325);
and U51 (N_51,In_2324,In_545);
nand U52 (N_52,In_1896,In_1417);
nor U53 (N_53,In_2695,In_323);
nand U54 (N_54,In_2983,In_2720);
nand U55 (N_55,In_1575,In_728);
nor U56 (N_56,In_1536,In_660);
xnor U57 (N_57,In_1239,In_2497);
nor U58 (N_58,In_2514,In_2887);
and U59 (N_59,In_2133,In_2705);
nand U60 (N_60,In_1713,In_169);
or U61 (N_61,In_2167,In_933);
xnor U62 (N_62,In_443,In_132);
nand U63 (N_63,In_1455,In_1062);
xnor U64 (N_64,In_2183,In_2040);
nor U65 (N_65,In_554,In_1990);
nor U66 (N_66,In_43,In_1488);
nor U67 (N_67,In_1861,In_836);
nand U68 (N_68,In_1649,In_1781);
and U69 (N_69,In_1370,In_70);
xor U70 (N_70,In_2478,In_2048);
nor U71 (N_71,In_1625,In_733);
nor U72 (N_72,In_1928,In_1419);
or U73 (N_73,In_2860,In_2437);
or U74 (N_74,In_2467,In_1394);
nand U75 (N_75,In_2161,In_1738);
xor U76 (N_76,In_570,In_2714);
nor U77 (N_77,In_1793,In_2699);
or U78 (N_78,In_751,In_2856);
nor U79 (N_79,In_395,In_1197);
xor U80 (N_80,In_1810,In_1399);
nand U81 (N_81,In_1754,In_1028);
or U82 (N_82,In_1349,In_1489);
nor U83 (N_83,In_1054,In_2726);
xor U84 (N_84,In_2237,In_2281);
or U85 (N_85,In_32,In_1189);
nor U86 (N_86,In_2287,In_2939);
and U87 (N_87,In_2279,In_527);
or U88 (N_88,In_635,In_1334);
nand U89 (N_89,In_2541,In_692);
or U90 (N_90,In_1406,In_2100);
or U91 (N_91,In_373,In_312);
nor U92 (N_92,In_1145,In_2422);
xnor U93 (N_93,In_998,In_2620);
or U94 (N_94,In_2058,In_2103);
or U95 (N_95,In_2775,In_226);
and U96 (N_96,In_1675,In_2485);
nor U97 (N_97,In_1018,In_1113);
nand U98 (N_98,In_1042,In_2973);
and U99 (N_99,In_2544,In_427);
nand U100 (N_100,In_435,In_288);
nand U101 (N_101,In_2734,In_122);
and U102 (N_102,In_1448,In_120);
xor U103 (N_103,In_222,In_45);
and U104 (N_104,In_1260,In_212);
and U105 (N_105,In_1280,In_899);
or U106 (N_106,In_51,In_748);
and U107 (N_107,In_1800,In_598);
or U108 (N_108,In_377,In_2593);
nand U109 (N_109,In_791,In_215);
and U110 (N_110,In_890,In_594);
nand U111 (N_111,In_1446,In_1127);
and U112 (N_112,In_1445,In_2149);
xor U113 (N_113,In_1064,In_477);
xor U114 (N_114,In_764,In_1550);
xor U115 (N_115,In_901,In_1526);
nor U116 (N_116,In_237,In_1502);
and U117 (N_117,In_604,In_2651);
nand U118 (N_118,In_388,In_805);
xor U119 (N_119,In_2522,In_196);
xor U120 (N_120,In_906,In_2851);
nand U121 (N_121,In_1170,In_2380);
and U122 (N_122,In_1882,In_2524);
nand U123 (N_123,In_1120,In_1172);
and U124 (N_124,In_2633,In_1601);
nand U125 (N_125,In_1281,In_1524);
and U126 (N_126,In_2138,In_603);
or U127 (N_127,In_1732,In_769);
nand U128 (N_128,In_1842,In_375);
and U129 (N_129,In_694,In_995);
nor U130 (N_130,In_567,In_1594);
nor U131 (N_131,In_1870,In_2559);
and U132 (N_132,In_528,In_2533);
xor U133 (N_133,In_1272,In_1549);
or U134 (N_134,In_143,In_1750);
nor U135 (N_135,In_650,In_961);
nand U136 (N_136,In_956,In_178);
xor U137 (N_137,In_1714,In_81);
xor U138 (N_138,In_1193,In_2221);
nor U139 (N_139,In_1737,In_107);
and U140 (N_140,In_26,In_1288);
and U141 (N_141,In_1533,In_253);
nand U142 (N_142,In_304,In_106);
and U143 (N_143,In_8,In_1961);
nor U144 (N_144,In_2504,In_981);
and U145 (N_145,In_589,In_951);
xnor U146 (N_146,In_2045,In_260);
or U147 (N_147,In_519,In_924);
nand U148 (N_148,In_2729,In_2961);
nor U149 (N_149,In_2822,In_1099);
nand U150 (N_150,In_2038,In_658);
xor U151 (N_151,In_10,In_52);
xnor U152 (N_152,In_1420,In_1418);
nor U153 (N_153,In_2715,In_1400);
nand U154 (N_154,In_2055,In_195);
xnor U155 (N_155,In_423,In_159);
xnor U156 (N_156,In_1667,In_967);
nand U157 (N_157,In_2389,In_217);
nor U158 (N_158,In_599,In_1289);
nor U159 (N_159,In_1530,In_2144);
and U160 (N_160,In_279,In_2438);
or U161 (N_161,In_903,In_1639);
xnor U162 (N_162,In_202,In_1112);
nand U163 (N_163,In_1571,In_441);
and U164 (N_164,In_2654,In_674);
nand U165 (N_165,In_333,In_1593);
nand U166 (N_166,In_1760,In_2442);
nand U167 (N_167,In_2261,In_1080);
or U168 (N_168,In_2453,In_2171);
nand U169 (N_169,In_706,In_1303);
nor U170 (N_170,In_1382,In_898);
nand U171 (N_171,In_2374,In_1162);
or U172 (N_172,In_675,In_1006);
and U173 (N_173,In_36,In_2891);
nand U174 (N_174,In_1825,In_2343);
and U175 (N_175,In_1230,In_60);
and U176 (N_176,In_2918,In_2028);
and U177 (N_177,In_2693,In_1336);
nand U178 (N_178,In_2831,In_1930);
nor U179 (N_179,In_1381,In_2606);
nor U180 (N_180,In_2558,In_117);
or U181 (N_181,In_1066,In_186);
nor U182 (N_182,In_2203,In_2041);
nand U183 (N_183,In_408,In_2976);
nor U184 (N_184,In_308,In_2139);
or U185 (N_185,In_977,In_2719);
or U186 (N_186,In_2907,In_1378);
or U187 (N_187,In_2368,In_608);
or U188 (N_188,In_1873,In_1857);
and U189 (N_189,In_2676,In_768);
or U190 (N_190,In_2596,In_1504);
nand U191 (N_191,In_2321,In_2154);
or U192 (N_192,In_297,In_2543);
or U193 (N_193,In_1353,In_2553);
nor U194 (N_194,In_2166,In_1173);
or U195 (N_195,In_2925,In_18);
or U196 (N_196,In_2303,In_2220);
or U197 (N_197,In_1368,In_1492);
or U198 (N_198,In_1019,In_2771);
and U199 (N_199,In_1942,In_2156);
xor U200 (N_200,In_1208,In_166);
nand U201 (N_201,In_2375,In_824);
and U202 (N_202,In_620,In_1206);
xor U203 (N_203,In_1853,In_2034);
and U204 (N_204,In_2039,In_1318);
xnor U205 (N_205,In_701,In_664);
or U206 (N_206,In_121,In_1890);
xnor U207 (N_207,In_524,In_2022);
or U208 (N_208,In_887,In_190);
nand U209 (N_209,In_1126,In_2458);
or U210 (N_210,In_978,In_685);
nor U211 (N_211,In_2824,In_1618);
and U212 (N_212,In_1947,In_817);
or U213 (N_213,In_1885,In_638);
nand U214 (N_214,In_1183,In_294);
xor U215 (N_215,In_2899,In_1159);
xor U216 (N_216,In_1143,In_1723);
and U217 (N_217,In_1731,In_2531);
xnor U218 (N_218,In_490,In_2960);
nor U219 (N_219,In_563,In_93);
and U220 (N_220,In_2090,In_1643);
or U221 (N_221,In_2382,In_2284);
or U222 (N_222,In_275,In_964);
and U223 (N_223,In_103,In_337);
xnor U224 (N_224,In_396,In_1875);
or U225 (N_225,In_405,In_2568);
xnor U226 (N_226,In_55,In_155);
nor U227 (N_227,In_2312,In_790);
and U228 (N_228,In_320,In_897);
and U229 (N_229,In_1827,In_2980);
or U230 (N_230,In_75,In_2909);
or U231 (N_231,In_272,In_2802);
xor U232 (N_232,In_95,In_2366);
and U233 (N_233,In_1185,In_208);
xnor U234 (N_234,In_2104,In_1175);
and U235 (N_235,In_2940,In_610);
and U236 (N_236,In_867,In_846);
and U237 (N_237,In_381,In_2113);
nor U238 (N_238,In_1435,In_1878);
xor U239 (N_239,In_2666,In_1196);
or U240 (N_240,In_2194,In_1812);
nand U241 (N_241,In_2701,In_1652);
xnor U242 (N_242,In_838,In_2560);
or U243 (N_243,In_1912,In_2622);
xnor U244 (N_244,In_1478,In_2425);
nand U245 (N_245,In_1889,In_2737);
nand U246 (N_246,In_515,In_2008);
and U247 (N_247,In_2175,In_2096);
and U248 (N_248,In_2069,In_934);
nand U249 (N_249,In_718,In_1000);
and U250 (N_250,In_1236,In_2185);
xnor U251 (N_251,In_1943,In_1579);
xor U252 (N_252,In_2172,In_2739);
nand U253 (N_253,In_2981,In_2057);
nor U254 (N_254,In_2920,In_1474);
nor U255 (N_255,In_109,In_1266);
or U256 (N_256,In_1033,In_2957);
or U257 (N_257,In_1538,In_572);
nand U258 (N_258,In_989,In_1225);
nor U259 (N_259,In_1790,In_484);
nor U260 (N_260,In_2763,In_514);
xnor U261 (N_261,In_236,In_986);
nand U262 (N_262,In_2598,In_2123);
nor U263 (N_263,In_560,In_1415);
nor U264 (N_264,In_2356,In_2711);
nor U265 (N_265,In_1003,In_1220);
nor U266 (N_266,In_2327,In_172);
and U267 (N_267,In_1458,In_227);
or U268 (N_268,In_2772,In_2603);
or U269 (N_269,In_2607,In_2669);
xor U270 (N_270,In_2345,In_46);
and U271 (N_271,In_1058,In_271);
or U272 (N_272,In_2256,In_311);
nor U273 (N_273,In_1572,In_1114);
nor U274 (N_274,In_613,In_2253);
nor U275 (N_275,In_2482,In_386);
nand U276 (N_276,In_2371,In_1546);
or U277 (N_277,In_1547,In_2736);
or U278 (N_278,In_2446,In_1111);
and U279 (N_279,In_873,In_170);
nand U280 (N_280,In_1043,In_1024);
or U281 (N_281,In_605,In_966);
xor U282 (N_282,In_2833,In_1139);
nor U283 (N_283,In_2906,In_2958);
or U284 (N_284,In_1994,In_1498);
nand U285 (N_285,In_2503,In_256);
xor U286 (N_286,In_1864,In_2963);
nand U287 (N_287,In_2546,In_1321);
nor U288 (N_288,In_2443,In_1200);
nand U289 (N_289,In_2902,In_2148);
and U290 (N_290,In_1250,In_682);
nand U291 (N_291,In_2884,In_2357);
or U292 (N_292,In_40,In_2997);
xnor U293 (N_293,In_1887,In_1469);
xor U294 (N_294,In_2026,In_878);
or U295 (N_295,In_761,In_182);
nand U296 (N_296,In_2410,In_565);
nor U297 (N_297,In_128,In_73);
nor U298 (N_298,In_185,In_1217);
nor U299 (N_299,In_1609,In_156);
or U300 (N_300,In_595,In_164);
and U301 (N_301,In_1104,In_1385);
xnor U302 (N_302,In_1863,In_1525);
nand U303 (N_303,In_1228,In_723);
and U304 (N_304,In_785,In_2785);
nor U305 (N_305,In_447,In_1467);
and U306 (N_306,In_2498,In_2180);
and U307 (N_307,In_990,In_319);
or U308 (N_308,In_1906,In_911);
xor U309 (N_309,In_406,In_601);
nor U310 (N_310,In_2885,In_1679);
and U311 (N_311,In_278,In_1059);
and U312 (N_312,In_436,In_1508);
or U313 (N_313,In_1296,In_2992);
and U314 (N_314,In_361,In_2621);
nor U315 (N_315,In_2730,In_2082);
xnor U316 (N_316,In_513,In_98);
xor U317 (N_317,In_1782,In_2416);
nor U318 (N_318,In_953,In_2826);
nand U319 (N_319,In_1171,In_1464);
and U320 (N_320,In_2573,In_2257);
xnor U321 (N_321,In_561,In_207);
nand U322 (N_322,In_1721,In_1891);
xnor U323 (N_323,In_181,In_434);
nand U324 (N_324,In_238,In_1117);
nand U325 (N_325,In_2434,In_1946);
nand U326 (N_326,In_1057,In_1360);
nand U327 (N_327,In_632,In_2488);
nor U328 (N_328,In_619,In_1954);
nor U329 (N_329,In_2076,In_473);
nand U330 (N_330,In_1268,In_896);
xnor U331 (N_331,In_710,In_1327);
nor U332 (N_332,In_2555,In_662);
nand U333 (N_333,In_828,In_1563);
and U334 (N_334,In_57,In_1687);
xnor U335 (N_335,In_2217,In_1299);
nor U336 (N_336,In_2332,In_240);
and U337 (N_337,In_1991,In_2519);
xor U338 (N_338,In_1515,In_2011);
nor U339 (N_339,In_411,In_2445);
xor U340 (N_340,In_535,In_2223);
nand U341 (N_341,In_779,In_152);
xor U342 (N_342,In_2777,In_2879);
or U343 (N_343,In_2612,In_283);
nand U344 (N_344,In_439,In_2629);
xor U345 (N_345,In_2878,In_1328);
nand U346 (N_346,In_1603,In_876);
and U347 (N_347,In_1025,In_600);
and U348 (N_348,In_1851,In_365);
nand U349 (N_349,In_2271,In_1374);
or U350 (N_350,In_2116,In_1633);
or U351 (N_351,In_1030,In_258);
or U352 (N_352,In_340,In_2530);
or U353 (N_353,In_47,In_1985);
xor U354 (N_354,In_2584,In_2289);
nor U355 (N_355,In_2862,In_2043);
xnor U356 (N_356,In_1796,In_2349);
or U357 (N_357,In_2866,In_1460);
nand U358 (N_358,In_2904,In_2009);
or U359 (N_359,In_2074,In_2896);
or U360 (N_360,In_1672,In_2428);
nand U361 (N_361,In_1880,In_657);
xnor U362 (N_362,In_2440,In_1957);
xnor U363 (N_363,In_220,In_2461);
nor U364 (N_364,In_1638,In_1022);
xnor U365 (N_365,In_877,In_2258);
nand U366 (N_366,In_1926,In_485);
nor U367 (N_367,In_1442,In_352);
xor U368 (N_368,In_1707,In_2362);
xor U369 (N_369,In_2994,In_735);
and U370 (N_370,In_1518,In_2858);
nor U371 (N_371,In_1219,In_1555);
nor U372 (N_372,In_654,In_673);
or U373 (N_373,In_1537,In_1751);
or U374 (N_374,In_2218,In_1739);
or U375 (N_375,In_1283,In_1823);
or U376 (N_376,In_1514,In_640);
or U377 (N_377,In_2575,In_2665);
and U378 (N_378,In_232,In_1822);
nand U379 (N_379,In_520,In_2044);
or U380 (N_380,In_2337,In_0);
xor U381 (N_381,In_1364,In_1065);
xor U382 (N_382,In_962,In_2863);
nor U383 (N_383,In_2017,In_920);
or U384 (N_384,In_2982,In_1981);
nand U385 (N_385,In_287,In_2092);
or U386 (N_386,In_1309,In_2995);
nor U387 (N_387,In_1699,In_1867);
and U388 (N_388,In_745,In_400);
or U389 (N_389,In_869,In_1007);
and U390 (N_390,In_94,In_2713);
xor U391 (N_391,In_1710,In_1129);
nor U392 (N_392,In_711,In_131);
nand U393 (N_393,In_752,In_1501);
nor U394 (N_394,In_1520,In_1740);
xnor U395 (N_395,In_2641,In_1094);
nand U396 (N_396,In_1214,In_1304);
xor U397 (N_397,In_1623,In_2153);
nand U398 (N_398,In_1995,In_2682);
and U399 (N_399,In_1921,In_233);
or U400 (N_400,In_2226,In_1244);
and U401 (N_401,In_1125,In_360);
nor U402 (N_402,In_15,In_894);
xor U403 (N_403,In_2035,In_2984);
and U404 (N_404,In_900,In_1499);
or U405 (N_405,In_913,In_1137);
nor U406 (N_406,In_30,In_1074);
or U407 (N_407,In_1375,In_7);
nand U408 (N_408,In_689,In_843);
xor U409 (N_409,In_2319,In_1859);
nand U410 (N_410,In_2807,In_2264);
nand U411 (N_411,In_1118,In_41);
nand U412 (N_412,In_1519,In_633);
xnor U413 (N_413,In_2805,In_1454);
nand U414 (N_414,In_1082,In_725);
nand U415 (N_415,In_458,In_2242);
nor U416 (N_416,In_2774,In_193);
xor U417 (N_417,In_2535,In_1227);
nor U418 (N_418,In_2151,In_1128);
nand U419 (N_419,In_1544,In_1668);
nand U420 (N_420,In_2949,In_2212);
nand U421 (N_421,In_1224,In_812);
nor U422 (N_422,In_1300,In_778);
and U423 (N_423,In_1993,In_292);
nor U424 (N_424,In_489,In_722);
and U425 (N_425,In_628,In_1337);
or U426 (N_426,In_539,In_2455);
nor U427 (N_427,In_879,In_1310);
nor U428 (N_428,In_48,In_2260);
nand U429 (N_429,In_1980,In_1267);
and U430 (N_430,In_77,In_1688);
xor U431 (N_431,In_25,In_1323);
and U432 (N_432,In_2406,In_2731);
nor U433 (N_433,In_1910,In_402);
xor U434 (N_434,In_2480,In_562);
or U435 (N_435,In_1932,In_2868);
and U436 (N_436,In_2454,In_2943);
nand U437 (N_437,In_2283,In_690);
nand U438 (N_438,In_2019,In_465);
nor U439 (N_439,In_114,In_2081);
or U440 (N_440,In_87,In_2106);
nor U441 (N_441,In_2733,In_2302);
nand U442 (N_442,In_2814,In_917);
or U443 (N_443,In_2971,In_2191);
xor U444 (N_444,In_2664,In_448);
nand U445 (N_445,In_1487,In_1509);
nand U446 (N_446,In_776,In_2201);
nor U447 (N_447,In_645,In_1925);
nand U448 (N_448,In_1,In_642);
xor U449 (N_449,In_2411,In_2532);
nand U450 (N_450,In_707,In_2931);
or U451 (N_451,In_2948,In_2249);
or U452 (N_452,In_125,In_1295);
or U453 (N_453,In_1726,In_980);
and U454 (N_454,In_2660,In_1763);
xnor U455 (N_455,In_1453,In_2238);
nand U456 (N_456,In_765,In_1002);
xor U457 (N_457,In_1806,In_2721);
nand U458 (N_458,In_854,In_2024);
nor U459 (N_459,In_575,In_1226);
nor U460 (N_460,In_2572,In_428);
and U461 (N_461,In_2134,In_1392);
and U462 (N_462,In_437,In_63);
nor U463 (N_463,In_1068,In_1262);
nand U464 (N_464,In_2601,In_766);
and U465 (N_465,In_147,In_927);
nor U466 (N_466,In_586,In_1429);
nand U467 (N_467,In_2259,In_580);
nor U468 (N_468,In_127,In_54);
or U469 (N_469,In_1722,In_597);
or U470 (N_470,In_1384,In_2003);
nand U471 (N_471,In_2547,In_2400);
nand U472 (N_472,In_24,In_712);
and U473 (N_473,In_1081,In_397);
nor U474 (N_474,In_2657,In_252);
or U475 (N_475,In_1179,In_883);
nor U476 (N_476,In_2334,In_409);
xor U477 (N_477,In_2079,In_2658);
nor U478 (N_478,In_584,In_2838);
and U479 (N_479,In_2846,In_2589);
nand U480 (N_480,In_1640,In_866);
or U481 (N_481,In_1157,In_2397);
nor U482 (N_482,In_2689,In_2213);
xor U483 (N_483,In_872,In_833);
or U484 (N_484,In_941,In_2921);
nor U485 (N_485,In_1147,In_1450);
or U486 (N_486,In_2781,In_1341);
nand U487 (N_487,In_2108,In_68);
nor U488 (N_488,In_616,In_426);
xor U489 (N_489,In_248,In_2588);
and U490 (N_490,In_702,In_2487);
nor U491 (N_491,In_362,In_2893);
and U492 (N_492,In_2409,In_1794);
and U493 (N_493,In_2192,In_1831);
and U494 (N_494,In_2764,In_550);
and U495 (N_495,In_332,In_2094);
and U496 (N_496,In_1849,In_909);
nand U497 (N_497,In_626,In_2797);
nand U498 (N_498,In_681,In_1899);
and U499 (N_499,In_136,In_1577);
xnor U500 (N_500,In_721,In_255);
and U501 (N_501,In_1339,In_2470);
nor U502 (N_502,In_2912,In_2989);
or U503 (N_503,In_2084,In_2209);
nor U504 (N_504,In_1573,In_1115);
nand U505 (N_505,In_2977,In_2095);
and U506 (N_506,In_2872,In_2549);
nor U507 (N_507,In_959,In_392);
and U508 (N_508,In_786,In_2494);
and U509 (N_509,In_2534,In_1342);
or U510 (N_510,In_749,In_985);
xor U511 (N_511,In_2029,In_2361);
or U512 (N_512,In_173,In_2523);
nor U513 (N_513,In_530,In_1862);
and U514 (N_514,In_265,In_2427);
and U515 (N_515,In_1461,In_922);
xor U516 (N_516,In_2965,In_62);
or U517 (N_517,In_223,In_2052);
nor U518 (N_518,In_501,In_1037);
nand U519 (N_519,In_2962,In_425);
or U520 (N_520,In_2071,In_1746);
xnor U521 (N_521,In_1592,In_556);
or U522 (N_522,In_551,In_1380);
nand U523 (N_523,In_2832,In_2304);
or U524 (N_524,In_2617,In_1351);
and U525 (N_525,In_2305,In_1922);
nor U526 (N_526,In_2012,In_2146);
xor U527 (N_527,In_915,In_1651);
nor U528 (N_528,In_1069,In_1124);
or U529 (N_529,In_1876,In_289);
and U530 (N_530,In_531,In_2252);
nor U531 (N_531,In_2817,In_1316);
and U532 (N_532,In_803,In_2507);
nor U533 (N_533,In_2173,In_343);
and U534 (N_534,In_826,In_80);
or U535 (N_535,In_2137,In_4);
xnor U536 (N_536,In_2966,In_2854);
xnor U537 (N_537,In_468,In_1077);
nor U538 (N_538,In_431,In_2004);
or U539 (N_539,In_2758,In_2270);
nor U540 (N_540,In_1616,In_891);
xor U541 (N_541,In_1620,In_1619);
and U542 (N_542,In_359,In_1051);
nor U543 (N_543,In_1913,In_1730);
or U544 (N_544,In_1729,In_2248);
xor U545 (N_545,In_440,In_2619);
and U546 (N_546,In_498,In_1088);
nand U547 (N_547,In_335,In_949);
nor U548 (N_548,In_2649,In_89);
and U549 (N_549,In_2360,In_2561);
and U550 (N_550,In_242,In_285);
xnor U551 (N_551,In_17,In_2552);
or U552 (N_552,In_568,In_796);
xor U553 (N_553,In_379,In_676);
xor U554 (N_554,In_1658,In_417);
nor U555 (N_555,In_179,In_2867);
xnor U556 (N_556,In_157,In_2563);
xnor U557 (N_557,In_2413,In_2608);
xor U558 (N_558,In_246,In_1929);
nand U559 (N_559,In_1881,In_1727);
or U560 (N_560,In_1329,In_1109);
or U561 (N_561,In_184,In_1108);
nor U562 (N_562,In_2126,In_130);
nor U563 (N_563,In_1084,In_2938);
nor U564 (N_564,In_2582,In_502);
nand U565 (N_565,In_2680,In_2892);
or U566 (N_566,In_1142,In_1931);
or U567 (N_567,In_1083,In_204);
xnor U568 (N_568,In_2569,In_918);
or U569 (N_569,In_715,In_1982);
or U570 (N_570,In_705,In_1004);
xnor U571 (N_571,In_943,In_1868);
or U572 (N_572,In_760,In_952);
xor U573 (N_573,In_2604,In_2010);
xor U574 (N_574,In_2755,In_588);
nor U575 (N_575,In_669,In_1012);
xnor U576 (N_576,In_2791,In_1567);
or U577 (N_577,In_1797,In_2186);
xnor U578 (N_578,In_1358,In_2087);
nor U579 (N_579,In_2325,In_2450);
or U580 (N_580,In_1144,In_2770);
and U581 (N_581,In_244,In_538);
and U582 (N_582,In_1343,In_1359);
nand U583 (N_583,In_1089,In_2614);
and U584 (N_584,In_577,In_1933);
nor U585 (N_585,In_1869,In_1416);
nor U586 (N_586,In_787,In_585);
nand U587 (N_587,In_1554,In_1067);
and U588 (N_588,In_1009,In_2060);
xnor U589 (N_589,In_935,In_21);
and U590 (N_590,In_1365,In_1252);
and U591 (N_591,In_2778,In_2656);
nand U592 (N_592,In_413,In_2511);
nor U593 (N_593,In_401,In_2244);
and U594 (N_594,In_2554,In_1169);
nor U595 (N_595,In_2871,In_2586);
nand U596 (N_596,In_2567,In_2810);
nand U597 (N_597,In_2447,In_2521);
xor U598 (N_598,In_2968,In_2230);
nor U599 (N_599,In_948,In_885);
and U600 (N_600,In_1920,In_2353);
or U601 (N_601,In_2355,In_2101);
or U602 (N_602,In_1379,In_2005);
and U603 (N_603,In_2492,In_811);
nor U604 (N_604,In_737,In_1456);
or U605 (N_605,In_1940,In_286);
xnor U606 (N_606,In_857,In_1485);
or U607 (N_607,In_523,In_1122);
or U608 (N_608,In_1749,In_6);
nand U609 (N_609,In_2578,In_2636);
nor U610 (N_610,In_2182,In_1466);
nand U611 (N_611,In_2147,In_1258);
or U612 (N_612,In_1596,In_2114);
xnor U613 (N_613,In_1778,In_1808);
nand U614 (N_614,In_1050,In_1235);
xor U615 (N_615,In_677,In_1205);
and U616 (N_616,In_2585,In_680);
nand U617 (N_617,In_988,In_347);
xor U618 (N_618,In_2895,In_2783);
and U619 (N_619,In_2272,In_1291);
and U620 (N_620,In_1011,In_438);
nand U621 (N_621,In_2922,In_2670);
nand U622 (N_622,In_738,In_1457);
xnor U623 (N_623,In_2728,In_321);
nand U624 (N_624,In_369,In_2974);
nand U625 (N_625,In_1070,In_840);
nor U626 (N_626,In_932,In_1839);
xor U627 (N_627,In_1100,In_793);
nand U628 (N_628,In_651,In_2187);
xnor U629 (N_629,In_1564,In_802);
nor U630 (N_630,In_1053,In_1350);
and U631 (N_631,In_1422,In_462);
nand U632 (N_632,In_553,In_807);
xnor U633 (N_633,In_1645,In_731);
xor U634 (N_634,In_2216,In_1837);
xor U635 (N_635,In_2373,In_487);
or U636 (N_636,In_2128,In_1388);
nor U637 (N_637,In_2241,In_110);
xnor U638 (N_638,In_2269,In_2704);
nand U639 (N_639,In_2827,In_541);
or U640 (N_640,In_2557,In_2990);
or U641 (N_641,In_1874,In_1010);
nand U642 (N_642,In_1393,In_85);
nand U643 (N_643,In_954,In_2352);
nor U644 (N_644,In_262,In_1424);
nor U645 (N_645,In_2634,In_263);
nor U646 (N_646,In_2150,In_259);
or U647 (N_647,In_2295,In_1276);
and U648 (N_648,In_2502,In_1934);
nor U649 (N_649,In_2449,In_982);
nor U650 (N_650,In_559,In_1871);
nand U651 (N_651,In_145,In_1698);
nand U652 (N_652,In_1079,In_974);
xor U653 (N_653,In_2288,In_234);
nor U654 (N_654,In_1786,In_1302);
nor U655 (N_655,In_2602,In_719);
nand U656 (N_656,In_2299,In_419);
xor U657 (N_657,In_1606,In_1809);
xnor U658 (N_658,In_2402,In_1785);
xnor U659 (N_659,In_1804,In_699);
or U660 (N_660,In_1317,In_2335);
nor U661 (N_661,In_886,In_23);
xnor U662 (N_662,In_1752,In_1614);
and U663 (N_663,In_1354,In_2369);
xor U664 (N_664,In_578,In_809);
nand U665 (N_665,In_1204,In_2426);
and U666 (N_666,In_1634,In_1192);
and U667 (N_667,In_2111,In_2077);
nand U668 (N_668,In_2801,In_307);
and U669 (N_669,In_730,In_1149);
nand U670 (N_670,In_1376,In_2367);
or U671 (N_671,In_2840,In_606);
nor U672 (N_672,In_2049,In_2667);
or U673 (N_673,In_432,In_810);
or U674 (N_674,In_370,In_2756);
nor U675 (N_675,In_1017,In_33);
or U676 (N_676,In_1834,In_1548);
nand U677 (N_677,In_534,In_257);
and U678 (N_678,In_2107,In_2414);
nand U679 (N_679,In_1348,In_2451);
xnor U680 (N_680,In_969,In_2391);
and U681 (N_681,In_637,In_134);
nor U682 (N_682,In_1473,In_1313);
xor U683 (N_683,In_460,In_1026);
and U684 (N_684,In_1897,In_587);
nor U685 (N_685,In_1938,In_322);
nand U686 (N_686,In_1286,In_546);
xnor U687 (N_687,In_2477,In_1986);
nor U688 (N_688,In_2509,In_2037);
nor U689 (N_689,In_2659,In_2508);
and U690 (N_690,In_1056,In_525);
and U691 (N_691,In_695,In_2932);
nand U692 (N_692,In_2661,In_1152);
and U693 (N_693,In_1755,In_91);
and U694 (N_694,In_346,In_946);
xor U695 (N_695,In_1158,In_591);
and U696 (N_696,In_2160,In_1340);
nand U697 (N_697,In_1331,In_1765);
nand U698 (N_698,In_2472,In_1369);
or U699 (N_699,In_1582,In_2707);
or U700 (N_700,In_1034,In_1581);
nand U701 (N_701,In_717,In_2155);
nand U702 (N_702,In_1167,In_2933);
or U703 (N_703,In_2341,In_1734);
nand U704 (N_704,In_1543,In_2754);
or U705 (N_705,In_318,In_1848);
nor U706 (N_706,In_2310,In_2329);
nor U707 (N_707,In_108,In_2512);
nand U708 (N_708,In_276,In_2204);
and U709 (N_709,In_1768,In_2696);
and U710 (N_710,In_2722,In_2174);
or U711 (N_711,In_2460,In_1491);
or U712 (N_712,In_552,In_2528);
and U713 (N_713,In_720,In_2481);
xor U714 (N_714,In_2812,In_1506);
and U715 (N_715,In_1148,In_2782);
and U716 (N_716,In_2363,In_2339);
or U717 (N_717,In_2372,In_2955);
or U718 (N_718,In_2803,In_1676);
or U719 (N_719,In_1654,In_1720);
xor U720 (N_720,In_940,In_2972);
nor U721 (N_721,In_1098,In_2916);
nand U722 (N_722,In_1029,In_2313);
nand U723 (N_723,In_1072,In_910);
and U724 (N_724,In_2206,In_2590);
nor U725 (N_725,In_936,In_1194);
nor U726 (N_726,In_2692,In_2493);
or U727 (N_727,In_2277,In_2317);
xnor U728 (N_728,In_1559,In_1659);
and U729 (N_729,In_868,In_199);
and U730 (N_730,In_2469,In_1036);
or U731 (N_731,In_2200,In_2875);
nand U732 (N_732,In_495,In_162);
or U733 (N_733,In_1636,In_916);
nor U734 (N_734,In_72,In_1153);
or U735 (N_735,In_1269,In_153);
nand U736 (N_736,In_1311,In_2266);
xnor U737 (N_737,In_2565,In_1607);
xor U738 (N_738,In_2110,In_2250);
or U739 (N_739,In_1275,In_2457);
nor U740 (N_740,In_2850,In_1937);
xor U741 (N_741,In_2744,In_78);
and U742 (N_742,In_203,In_2207);
nand U743 (N_743,In_2830,In_2592);
nor U744 (N_744,In_2742,In_2393);
and U745 (N_745,In_76,In_771);
and U746 (N_746,In_2,In_2326);
and U747 (N_747,In_1123,In_1249);
xnor U748 (N_748,In_1716,In_1745);
or U749 (N_749,In_2491,In_313);
xnor U750 (N_750,In_1207,In_105);
xnor U751 (N_751,In_960,In_1974);
and U752 (N_752,In_2181,In_296);
or U753 (N_753,In_1819,In_2290);
or U754 (N_754,In_2385,In_1216);
and U755 (N_755,In_557,In_615);
or U756 (N_756,In_1718,In_773);
and U757 (N_757,In_1591,In_542);
xor U758 (N_758,In_2836,In_1798);
nand U759 (N_759,In_2117,In_1306);
or U760 (N_760,In_2903,In_1703);
and U761 (N_761,In_1784,In_2351);
xor U762 (N_762,In_2746,In_338);
nand U763 (N_763,In_767,In_1107);
and U764 (N_764,In_13,In_2613);
or U765 (N_765,In_1815,In_351);
nand U766 (N_766,In_889,In_2929);
xor U767 (N_767,In_49,In_1558);
xnor U768 (N_768,In_2923,In_543);
and U769 (N_769,In_1187,In_929);
xor U770 (N_770,In_2479,In_1692);
xnor U771 (N_771,In_2789,In_2033);
xnor U772 (N_772,In_66,In_454);
or U773 (N_773,In_1894,In_2417);
xor U774 (N_774,In_500,In_2441);
nor U775 (N_775,In_2650,In_1315);
or U776 (N_776,In_1138,In_2224);
and U777 (N_777,In_912,In_1174);
xnor U778 (N_778,In_2579,In_2359);
nand U779 (N_779,In_137,In_757);
xnor U780 (N_780,In_2748,In_958);
nor U781 (N_781,In_403,In_1407);
nor U782 (N_782,In_747,In_1078);
nand U783 (N_783,In_1503,In_382);
and U784 (N_784,In_830,In_1725);
nand U785 (N_785,In_2273,In_1562);
or U786 (N_786,In_1789,In_1398);
nor U787 (N_787,In_1232,In_1140);
nand U788 (N_788,In_1190,In_2420);
nand U789 (N_789,In_421,In_697);
xor U790 (N_790,In_2328,In_1841);
nor U791 (N_791,In_479,In_2179);
xnor U792 (N_792,In_858,In_1835);
nor U793 (N_793,In_753,In_1404);
xnor U794 (N_794,In_2276,In_2580);
and U795 (N_795,In_1346,In_1046);
nand U796 (N_796,In_442,In_2468);
or U797 (N_797,In_991,In_1637);
nand U798 (N_798,In_1248,In_1673);
nor U799 (N_799,In_2143,In_1850);
nand U800 (N_800,In_688,In_2403);
or U801 (N_801,In_2959,In_201);
xor U802 (N_802,In_1569,In_1624);
xor U803 (N_803,In_2145,In_2761);
or U804 (N_804,In_740,In_1150);
nand U805 (N_805,In_2718,In_1599);
nand U806 (N_806,In_1091,In_1852);
nor U807 (N_807,In_65,In_2489);
nand U808 (N_808,In_533,In_494);
nor U809 (N_809,In_2433,In_2828);
and U810 (N_810,In_661,In_921);
nor U811 (N_811,In_493,In_2080);
or U812 (N_812,In_2675,In_1132);
and U813 (N_813,In_463,In_2566);
xor U814 (N_814,In_1027,In_947);
xor U815 (N_815,In_1020,In_630);
and U816 (N_816,In_1237,In_2490);
nand U817 (N_817,In_1955,In_2421);
xnor U818 (N_818,In_1677,In_1635);
or U819 (N_819,In_1983,In_2820);
nand U820 (N_820,In_950,In_1924);
nor U821 (N_821,In_1630,In_1626);
and U822 (N_822,In_254,In_174);
xnor U823 (N_823,In_1254,In_804);
and U824 (N_824,In_571,In_2864);
and U825 (N_825,In_2140,In_853);
or U826 (N_826,In_862,In_762);
xnor U827 (N_827,In_2016,In_345);
xor U828 (N_828,In_2112,In_2645);
and U829 (N_829,In_609,In_2999);
nor U830 (N_830,In_2571,In_871);
and U831 (N_831,In_1163,In_2027);
nor U832 (N_832,In_1361,In_1709);
nand U833 (N_833,In_1307,In_488);
or U834 (N_834,In_1708,In_1483);
nand U835 (N_835,In_191,In_1008);
nor U836 (N_836,In_931,In_2804);
xnor U837 (N_837,In_2063,In_218);
nand U838 (N_838,In_69,In_420);
nor U839 (N_839,In_249,In_2611);
nand U840 (N_840,In_2889,In_2520);
or U841 (N_841,In_1949,In_746);
and U842 (N_842,In_341,In_1680);
nor U843 (N_843,In_1918,In_1186);
or U844 (N_844,In_1693,In_874);
and U845 (N_845,In_1770,In_1160);
nor U846 (N_846,In_1772,In_1218);
or U847 (N_847,In_326,In_1556);
xnor U848 (N_848,In_847,In_2545);
nand U849 (N_849,In_1711,In_1093);
nor U850 (N_850,In_1253,In_2835);
or U851 (N_851,In_112,In_2322);
nor U852 (N_852,In_1998,In_2798);
and U853 (N_853,In_2865,In_2251);
nor U854 (N_854,In_1462,In_1801);
nor U855 (N_855,In_2632,In_2773);
nor U856 (N_856,In_2431,In_2066);
and U857 (N_857,In_2577,In_2510);
and U858 (N_858,In_2053,In_2626);
or U859 (N_859,In_1979,In_20);
nand U860 (N_860,In_464,In_281);
and U861 (N_861,In_2668,In_2765);
and U862 (N_862,In_1877,In_844);
xor U863 (N_863,In_2255,In_1297);
xor U864 (N_864,In_1314,In_334);
nor U865 (N_865,In_50,In_2120);
nand U866 (N_866,In_2880,In_74);
or U867 (N_867,In_1741,In_353);
and U868 (N_868,In_1188,In_2919);
xnor U869 (N_869,In_993,In_2861);
xnor U870 (N_870,In_2115,In_623);
or U871 (N_871,In_1557,In_1956);
nand U872 (N_872,In_328,In_1917);
and U873 (N_873,In_1182,In_2888);
or U874 (N_874,In_2690,In_1589);
and U875 (N_875,In_1747,In_1724);
nand U876 (N_876,In_2845,In_566);
and U877 (N_877,In_1178,In_451);
or U878 (N_878,In_1076,In_211);
nand U879 (N_879,In_1165,In_1830);
nand U880 (N_880,In_1689,In_229);
and U881 (N_881,In_1950,In_1685);
xnor U882 (N_882,In_1893,In_902);
and U883 (N_883,In_1855,In_2097);
or U884 (N_884,In_2189,In_2673);
nand U885 (N_885,In_926,In_2127);
nor U886 (N_886,In_2125,In_1240);
and U887 (N_887,In_1613,In_228);
and U888 (N_888,In_693,In_2691);
xor U889 (N_889,In_656,In_188);
nor U890 (N_890,In_2702,In_839);
or U891 (N_891,In_348,In_1602);
or U892 (N_892,In_2643,In_1423);
nor U893 (N_893,In_2537,In_2869);
nand U894 (N_894,In_1847,In_486);
xnor U895 (N_895,In_445,In_1611);
or U896 (N_896,In_424,In_1795);
or U897 (N_897,In_2275,In_1901);
nor U898 (N_898,In_2542,In_1274);
and U899 (N_899,In_1598,In_1553);
nand U900 (N_900,In_2934,In_576);
nor U901 (N_901,In_2911,In_1953);
nand U902 (N_902,In_999,In_2709);
xor U903 (N_903,In_455,In_1484);
nand U904 (N_904,In_780,In_2749);
and U905 (N_905,In_1761,In_1345);
or U906 (N_906,In_2583,In_2118);
xor U907 (N_907,In_1439,In_2540);
and U908 (N_908,In_544,In_327);
or U909 (N_909,In_1627,In_1164);
nand U910 (N_910,In_2527,In_2119);
or U911 (N_911,In_729,In_391);
and U912 (N_912,In_101,In_2001);
and U913 (N_913,In_2639,In_2164);
xnor U914 (N_914,In_739,In_845);
and U915 (N_915,In_2376,In_1363);
and U916 (N_916,In_716,In_1628);
nand U917 (N_917,In_2466,In_1792);
nand U918 (N_918,In_339,In_1540);
xor U919 (N_919,In_206,In_1437);
nand U920 (N_920,In_2296,In_2130);
xor U921 (N_921,In_1285,In_2930);
xnor U922 (N_922,In_683,In_274);
xor U923 (N_923,In_163,In_2474);
nand U924 (N_924,In_2821,In_1531);
and U925 (N_925,In_1641,In_393);
nand U926 (N_926,In_2623,In_2476);
nor U927 (N_927,In_1261,In_1060);
nand U928 (N_928,In_3,In_2050);
and U929 (N_929,In_945,In_1648);
or U930 (N_930,In_1776,In_97);
nand U931 (N_931,In_1409,In_2637);
and U932 (N_932,In_822,In_2951);
nor U933 (N_933,In_516,In_2853);
or U934 (N_934,In_1838,In_1308);
nor U935 (N_935,In_295,In_1650);
and U936 (N_936,In_2177,In_2631);
xnor U937 (N_937,In_2574,In_727);
or U938 (N_938,In_355,In_126);
or U939 (N_939,In_1071,In_659);
or U940 (N_940,In_1472,In_1888);
xor U941 (N_941,In_2883,In_1691);
nand U942 (N_942,In_1935,In_325);
or U943 (N_943,In_698,In_418);
xnor U944 (N_944,In_2942,In_104);
xnor U945 (N_945,In_529,In_1696);
and U946 (N_946,In_742,In_2517);
xor U947 (N_947,In_1597,In_1231);
and U948 (N_948,In_2404,In_2196);
nor U949 (N_949,In_2597,In_135);
nand U950 (N_950,In_1803,In_2062);
nand U951 (N_951,In_1390,In_1073);
nand U952 (N_952,In_848,In_1757);
and U953 (N_953,In_2199,In_1201);
nand U954 (N_954,In_2910,In_2390);
and U955 (N_955,In_888,In_2513);
nand U956 (N_956,In_2065,In_2975);
nand U957 (N_957,In_1802,In_1005);
xor U958 (N_958,In_2168,In_1326);
nand U959 (N_959,In_1493,In_1039);
xor U960 (N_960,In_42,In_2698);
or U961 (N_961,In_2842,In_349);
xor U962 (N_962,In_471,In_564);
nor U963 (N_963,In_1683,In_453);
nand U964 (N_964,In_383,In_282);
and U965 (N_965,In_2687,In_938);
nand U966 (N_966,In_1821,In_2377);
nor U967 (N_967,In_2587,In_1779);
or U968 (N_968,In_2935,In_2484);
and U969 (N_969,In_1141,In_1939);
xor U970 (N_970,In_503,In_759);
nand U971 (N_971,In_611,In_1941);
xor U972 (N_972,In_2784,In_1021);
xnor U973 (N_973,In_2292,In_2913);
and U974 (N_974,In_1660,In_2439);
and U975 (N_975,In_183,In_239);
and U976 (N_976,In_1669,In_2210);
nand U977 (N_977,In_1434,In_138);
or U978 (N_978,In_2727,In_496);
and U979 (N_979,In_882,In_356);
nor U980 (N_980,In_1049,In_1278);
xor U981 (N_981,In_1600,In_1570);
or U982 (N_982,In_280,In_92);
and U983 (N_983,In_2031,In_1764);
xnor U984 (N_984,In_2121,In_129);
and U985 (N_985,In_1480,In_2677);
nand U986 (N_986,In_2886,In_243);
nand U987 (N_987,In_2301,In_2640);
and U988 (N_988,In_221,In_2760);
and U989 (N_989,In_1213,In_1013);
nor U990 (N_990,In_1914,In_389);
xor U991 (N_991,In_666,In_649);
or U992 (N_992,In_1413,In_2064);
and U993 (N_993,In_1063,In_970);
nor U994 (N_994,In_2870,In_818);
nand U995 (N_995,In_293,In_1700);
nand U996 (N_996,In_2638,In_2809);
xor U997 (N_997,In_1287,In_1690);
and U998 (N_998,In_1284,In_1966);
and U999 (N_999,In_1706,In_923);
nor U1000 (N_1000,In_1055,In_2671);
nand U1001 (N_1001,In_2229,In_925);
xor U1002 (N_1002,In_39,In_2423);
and U1003 (N_1003,In_1886,In_2091);
nand U1004 (N_1004,In_1662,In_506);
and U1005 (N_1005,In_1119,In_511);
and U1006 (N_1006,In_1697,In_892);
or U1007 (N_1007,In_1106,In_1742);
nand U1008 (N_1008,In_1970,In_1161);
and U1009 (N_1009,In_2348,In_1221);
nor U1010 (N_1010,In_2717,In_1136);
nand U1011 (N_1011,In_1090,In_2330);
nand U1012 (N_1012,In_2914,In_1265);
or U1013 (N_1013,In_1246,In_2239);
or U1014 (N_1014,In_1061,In_2340);
and U1015 (N_1015,In_1883,In_1631);
xor U1016 (N_1016,In_2370,In_1818);
and U1017 (N_1017,In_1666,In_1975);
nor U1018 (N_1018,In_2394,In_621);
and U1019 (N_1019,In_1684,In_452);
or U1020 (N_1020,In_842,In_512);
nor U1021 (N_1021,In_569,In_306);
or U1022 (N_1022,In_1780,In_536);
nand U1023 (N_1023,In_756,In_115);
nand U1024 (N_1024,In_2162,In_816);
xnor U1025 (N_1025,In_2630,In_1824);
and U1026 (N_1026,In_113,In_1443);
nand U1027 (N_1027,In_410,In_1086);
or U1028 (N_1028,In_1048,In_1753);
xor U1029 (N_1029,In_357,In_467);
nor U1030 (N_1030,In_1915,In_189);
nor U1031 (N_1031,In_517,In_1121);
nand U1032 (N_1032,In_2834,In_904);
and U1033 (N_1033,In_350,In_2267);
or U1034 (N_1034,In_2882,In_893);
xnor U1035 (N_1035,In_622,In_2848);
xor U1036 (N_1036,In_1701,In_521);
nor U1037 (N_1037,In_2020,In_1561);
or U1038 (N_1038,In_2816,In_1181);
xor U1039 (N_1039,In_225,In_2815);
nand U1040 (N_1040,In_71,In_1438);
nand U1041 (N_1041,In_2085,In_2723);
nand U1042 (N_1042,In_1255,In_2599);
nor U1043 (N_1043,In_1972,In_581);
or U1044 (N_1044,In_1496,In_775);
or U1045 (N_1045,In_140,In_736);
nand U1046 (N_1046,In_540,In_1096);
and U1047 (N_1047,In_2859,In_1184);
or U1048 (N_1048,In_875,In_1656);
and U1049 (N_1049,In_124,In_744);
nand U1050 (N_1050,In_1402,In_547);
and U1051 (N_1051,In_1756,In_1948);
or U1052 (N_1052,In_2021,In_1414);
and U1053 (N_1053,In_2526,In_1911);
or U1054 (N_1054,In_1748,In_1198);
xnor U1055 (N_1055,In_231,In_2991);
or U1056 (N_1056,In_895,In_2852);
and U1057 (N_1057,In_504,In_755);
xnor U1058 (N_1058,In_2937,In_2235);
or U1059 (N_1059,In_2581,In_2628);
xnor U1060 (N_1060,In_629,In_2901);
or U1061 (N_1061,In_450,In_34);
and U1062 (N_1062,In_200,In_2681);
nor U1063 (N_1063,In_1967,In_631);
nand U1064 (N_1064,In_1105,In_2036);
xor U1065 (N_1065,In_2663,In_149);
and U1066 (N_1066,In_1305,In_2365);
xnor U1067 (N_1067,In_154,In_2928);
nand U1068 (N_1068,In_870,In_2684);
and U1069 (N_1069,In_2648,In_789);
nor U1070 (N_1070,In_679,In_2336);
nor U1071 (N_1071,In_407,In_2358);
nand U1072 (N_1072,In_219,In_829);
nand U1073 (N_1073,In_1777,In_1811);
nor U1074 (N_1074,In_2131,In_2293);
xor U1075 (N_1075,In_2897,In_1215);
and U1076 (N_1076,In_2779,In_1590);
xnor U1077 (N_1077,In_2398,In_2685);
nand U1078 (N_1078,In_2768,In_2072);
nor U1079 (N_1079,In_2662,In_1829);
and U1080 (N_1080,In_31,In_1909);
xnor U1081 (N_1081,In_1500,In_1279);
nand U1082 (N_1082,In_367,In_979);
nand U1083 (N_1083,In_2309,In_1356);
nor U1084 (N_1084,In_2890,In_16);
or U1085 (N_1085,In_1452,In_2740);
nand U1086 (N_1086,In_884,In_823);
nor U1087 (N_1087,In_2941,In_2350);
and U1088 (N_1088,In_881,In_277);
nand U1089 (N_1089,In_1156,In_146);
and U1090 (N_1090,In_834,In_548);
xnor U1091 (N_1091,In_314,In_639);
or U1092 (N_1092,In_2105,In_2499);
or U1093 (N_1093,In_1783,In_2738);
or U1094 (N_1094,In_1357,In_1016);
xnor U1095 (N_1095,In_1960,In_783);
and U1096 (N_1096,In_1522,In_849);
nand U1097 (N_1097,In_1664,In_2529);
or U1098 (N_1098,In_342,In_1817);
nand U1099 (N_1099,In_2947,In_1832);
or U1100 (N_1100,In_56,In_27);
or U1101 (N_1101,In_205,In_627);
or U1102 (N_1102,In_795,In_2448);
or U1103 (N_1103,In_142,In_794);
nand U1104 (N_1104,In_1642,In_2338);
nor U1105 (N_1105,In_1545,In_2908);
nor U1106 (N_1106,In_1644,In_2208);
and U1107 (N_1107,In_2605,In_1202);
nor U1108 (N_1108,In_1840,In_1858);
nor U1109 (N_1109,In_1373,In_1270);
nor U1110 (N_1110,In_2471,In_774);
and U1111 (N_1111,In_2462,In_2386);
nor U1112 (N_1112,In_404,In_841);
nor U1113 (N_1113,In_148,In_305);
and U1114 (N_1114,In_2165,In_2135);
nor U1115 (N_1115,In_976,In_1945);
nor U1116 (N_1116,In_2388,In_1521);
nor U1117 (N_1117,In_1257,In_2741);
xnor U1118 (N_1118,In_2998,In_100);
nand U1119 (N_1119,In_1999,In_1134);
and U1120 (N_1120,In_647,In_1203);
or U1121 (N_1121,In_781,In_743);
nand U1122 (N_1122,In_37,In_398);
and U1123 (N_1123,In_2769,In_2706);
and U1124 (N_1124,In_1095,In_1432);
nand U1125 (N_1125,In_2642,In_2282);
xnor U1126 (N_1126,In_2412,In_2548);
or U1127 (N_1127,In_2384,In_2653);
xor U1128 (N_1128,In_815,In_1377);
xnor U1129 (N_1129,In_2068,In_1397);
and U1130 (N_1130,In_667,In_1647);
and U1131 (N_1131,In_1510,In_2227);
or U1132 (N_1132,In_2059,In_1542);
and U1133 (N_1133,In_1552,In_1743);
xnor U1134 (N_1134,In_2032,In_175);
or U1135 (N_1135,In_141,In_2190);
nand U1136 (N_1136,In_2401,In_2263);
and U1137 (N_1137,In_602,In_1312);
nor U1138 (N_1138,In_364,In_1655);
nor U1139 (N_1139,In_470,In_1529);
xnor U1140 (N_1140,In_2354,In_1259);
and U1141 (N_1141,In_2978,In_2436);
xnor U1142 (N_1142,In_2222,In_714);
or U1143 (N_1143,In_526,In_390);
and U1144 (N_1144,In_2395,In_2307);
or U1145 (N_1145,In_1411,In_192);
nand U1146 (N_1146,In_930,In_1465);
xor U1147 (N_1147,In_2225,In_2679);
or U1148 (N_1148,In_315,In_53);
xnor U1149 (N_1149,In_2316,In_1900);
or U1150 (N_1150,In_2061,In_750);
or U1151 (N_1151,In_2188,In_1996);
nand U1152 (N_1152,In_1290,In_1436);
xor U1153 (N_1153,In_1805,In_480);
and U1154 (N_1154,In_537,In_919);
and U1155 (N_1155,In_2042,In_2170);
nor U1156 (N_1156,In_2109,In_372);
nand U1157 (N_1157,In_852,In_2697);
nand U1158 (N_1158,In_777,In_2946);
or U1159 (N_1159,In_508,In_2320);
nand U1160 (N_1160,In_1646,In_1539);
or U1161 (N_1161,In_1180,In_2102);
xor U1162 (N_1162,In_1430,In_1944);
nand U1163 (N_1163,In_1632,In_2124);
and U1164 (N_1164,In_2198,In_549);
or U1165 (N_1165,In_2926,In_2799);
nand U1166 (N_1166,In_1773,In_1023);
or U1167 (N_1167,In_939,In_724);
or U1168 (N_1168,In_2268,In_2950);
xnor U1169 (N_1169,In_797,In_1168);
or U1170 (N_1170,In_2158,In_2839);
xnor U1171 (N_1171,In_1087,In_1844);
nor U1172 (N_1172,In_1904,In_309);
xor U1173 (N_1173,In_808,In_1610);
xor U1174 (N_1174,In_2967,In_394);
xnor U1175 (N_1175,In_429,In_2184);
nor U1176 (N_1176,In_123,In_1528);
nand U1177 (N_1177,In_1962,In_1155);
nor U1178 (N_1178,In_344,In_2609);
xor U1179 (N_1179,In_928,In_2088);
and U1180 (N_1180,In_865,In_1001);
nor U1181 (N_1181,In_1451,In_1663);
or U1182 (N_1182,In_1146,In_1787);
nor U1183 (N_1183,In_2463,In_1992);
xor U1184 (N_1184,In_2505,In_2506);
or U1185 (N_1185,In_2323,In_2776);
xor U1186 (N_1186,In_1041,In_2576);
or U1187 (N_1187,In_2083,In_2294);
xor U1188 (N_1188,In_2688,In_399);
or U1189 (N_1189,In_607,In_1767);
nor U1190 (N_1190,In_1389,In_331);
nand U1191 (N_1191,In_1333,In_583);
nor U1192 (N_1192,In_819,In_2993);
xor U1193 (N_1193,In_2525,In_457);
nor U1194 (N_1194,In_1661,In_1860);
or U1195 (N_1195,In_2813,In_267);
nand U1196 (N_1196,In_83,In_522);
xnor U1197 (N_1197,In_1273,In_2751);
or U1198 (N_1198,In_1583,In_643);
xor U1199 (N_1199,In_187,In_2030);
xor U1200 (N_1200,In_1293,In_1735);
and U1201 (N_1201,In_1856,In_832);
or U1202 (N_1202,In_1014,In_1759);
or U1203 (N_1203,In_624,In_1578);
nand U1204 (N_1204,In_772,In_1344);
nor U1205 (N_1205,In_88,In_2159);
and U1206 (N_1206,In_1560,In_216);
nor U1207 (N_1207,In_2099,In_1212);
or U1208 (N_1208,In_1371,In_2285);
nand U1209 (N_1209,In_2556,In_11);
or U1210 (N_1210,In_1362,In_5);
or U1211 (N_1211,In_316,In_1820);
xor U1212 (N_1212,In_984,In_2945);
nor U1213 (N_1213,In_2047,In_481);
nor U1214 (N_1214,In_1324,In_1605);
and U1215 (N_1215,In_2829,In_433);
nor U1216 (N_1216,In_2025,In_1903);
xnor U1217 (N_1217,In_82,In_482);
or U1218 (N_1218,In_2825,In_2710);
or U1219 (N_1219,In_518,In_1052);
or U1220 (N_1220,In_2129,In_1766);
nand U1221 (N_1221,In_579,In_330);
or U1222 (N_1222,In_96,In_387);
or U1223 (N_1223,In_2392,In_573);
nor U1224 (N_1224,In_1387,In_973);
nand U1225 (N_1225,In_1532,In_2318);
xnor U1226 (N_1226,In_1681,In_2564);
nand U1227 (N_1227,In_1513,In_754);
and U1228 (N_1228,In_1110,In_2986);
nand U1229 (N_1229,In_139,In_907);
nand U1230 (N_1230,In_2725,In_198);
xnor U1231 (N_1231,In_1355,In_2236);
nand U1232 (N_1232,In_855,In_2855);
and U1233 (N_1233,In_1233,In_1584);
xor U1234 (N_1234,In_1497,In_2881);
or U1235 (N_1235,In_1872,In_1977);
or U1236 (N_1236,In_415,In_1898);
or U1237 (N_1237,In_2424,In_2311);
xnor U1238 (N_1238,In_2954,In_58);
or U1239 (N_1239,In_1032,In_2595);
nor U1240 (N_1240,In_831,In_1209);
nor U1241 (N_1241,In_1705,In_1843);
xnor U1242 (N_1242,In_499,In_814);
and U1243 (N_1243,In_1923,In_700);
nand U1244 (N_1244,In_2787,In_102);
and U1245 (N_1245,In_732,In_1470);
or U1246 (N_1246,In_472,In_2231);
and U1247 (N_1247,In_358,In_741);
nor U1248 (N_1248,In_2618,In_354);
nand U1249 (N_1249,In_2459,In_1116);
nand U1250 (N_1250,In_99,In_35);
or U1251 (N_1251,In_2013,In_2429);
or U1252 (N_1252,In_2023,In_2841);
nand U1253 (N_1253,In_19,In_860);
and U1254 (N_1254,In_1320,In_235);
nor U1255 (N_1255,In_2157,In_1665);
and U1256 (N_1256,In_1332,In_1845);
nand U1257 (N_1257,In_1133,In_2240);
nor U1258 (N_1258,In_1987,In_1166);
nor U1259 (N_1259,In_270,In_1969);
xnor U1260 (N_1260,In_261,In_2387);
or U1261 (N_1261,In_1686,In_1828);
xor U1262 (N_1262,In_2278,In_1482);
or U1263 (N_1263,In_1895,In_1386);
or U1264 (N_1264,In_1495,In_158);
xor U1265 (N_1265,In_614,In_2415);
xor U1266 (N_1266,In_1617,In_2616);
nand U1267 (N_1267,In_2247,In_1440);
or U1268 (N_1268,In_2246,In_612);
xor U1269 (N_1269,In_1047,In_2735);
xnor U1270 (N_1270,In_1045,In_555);
and U1271 (N_1271,In_2808,In_1251);
xor U1272 (N_1272,In_1426,In_2624);
nand U1273 (N_1273,In_2364,In_194);
or U1274 (N_1274,In_2627,In_446);
nor U1275 (N_1275,In_965,In_1177);
or U1276 (N_1276,In_456,In_1865);
nand U1277 (N_1277,In_1927,In_2193);
nor U1278 (N_1278,In_444,In_1585);
or U1279 (N_1279,In_2086,In_1092);
and U1280 (N_1280,In_1958,In_1744);
nor U1281 (N_1281,In_1264,In_2956);
and U1282 (N_1282,In_2002,In_1580);
xnor U1283 (N_1283,In_2915,In_644);
xnor U1284 (N_1284,In_1383,In_1622);
or U1285 (N_1285,In_704,In_1621);
nor U1286 (N_1286,In_2214,In_2905);
nand U1287 (N_1287,In_14,In_1997);
or U1288 (N_1288,In_1615,In_2849);
nor U1289 (N_1289,In_625,In_1421);
xnor U1290 (N_1290,In_835,In_478);
or U1291 (N_1291,In_176,In_59);
nand U1292 (N_1292,In_1135,In_2964);
nor U1293 (N_1293,In_469,In_2399);
or U1294 (N_1294,In_2857,In_800);
nand U1295 (N_1295,In_2538,In_1405);
nand U1296 (N_1296,In_2006,In_2132);
nor U1297 (N_1297,In_86,In_1595);
nor U1298 (N_1298,In_1907,In_264);
and U1299 (N_1299,In_2136,In_79);
and U1300 (N_1300,In_1507,In_937);
nand U1301 (N_1301,In_994,In_2142);
nand U1302 (N_1302,In_2873,In_1959);
nand U1303 (N_1303,In_2501,In_165);
xor U1304 (N_1304,In_1717,In_1447);
xnor U1305 (N_1305,In_1814,In_2073);
or U1306 (N_1306,In_1101,In_825);
or U1307 (N_1307,In_461,In_2408);
or U1308 (N_1308,In_144,In_336);
nand U1309 (N_1309,In_1678,In_301);
nand U1310 (N_1310,In_2098,In_2786);
xor U1311 (N_1311,In_1352,In_2780);
nor U1312 (N_1312,In_412,In_474);
nand U1313 (N_1313,In_1576,In_1211);
nor U1314 (N_1314,In_459,In_1401);
nor U1315 (N_1315,In_2683,In_2141);
xnor U1316 (N_1316,In_1736,In_2686);
and U1317 (N_1317,In_1477,In_2732);
xor U1318 (N_1318,In_2518,In_1984);
nor U1319 (N_1319,In_1568,In_2396);
xor U1320 (N_1320,In_2900,In_1131);
nor U1321 (N_1321,In_2647,In_1682);
nand U1322 (N_1322,In_596,In_1587);
xnor U1323 (N_1323,In_363,In_1154);
or U1324 (N_1324,In_2430,In_1670);
nand U1325 (N_1325,In_908,In_2197);
nand U1326 (N_1326,In_376,In_161);
and U1327 (N_1327,In_806,In_726);
nor U1328 (N_1328,In_670,In_449);
nor U1329 (N_1329,In_1769,In_1505);
xnor U1330 (N_1330,In_687,In_2495);
or U1331 (N_1331,In_2262,In_1097);
nand U1332 (N_1332,In_861,In_2444);
xnor U1333 (N_1333,In_1816,In_1604);
nand U1334 (N_1334,In_957,In_1879);
or U1335 (N_1335,In_2843,In_1222);
nand U1336 (N_1336,In_2635,In_2122);
and U1337 (N_1337,In_2202,In_1151);
and U1338 (N_1338,In_1486,In_2894);
or U1339 (N_1339,In_1884,In_799);
or U1340 (N_1340,In_1403,In_1475);
or U1341 (N_1341,In_696,In_1292);
nand U1342 (N_1342,In_273,In_209);
and U1343 (N_1343,In_483,In_770);
and U1344 (N_1344,In_558,In_684);
nor U1345 (N_1345,In_507,In_2562);
nand U1346 (N_1346,In_1902,In_2550);
nand U1347 (N_1347,In_416,In_2234);
nand U1348 (N_1348,In_2747,In_1695);
nand U1349 (N_1349,In_1015,In_992);
nand U1350 (N_1350,In_368,In_38);
nand U1351 (N_1351,In_1234,In_2452);
and U1352 (N_1352,In_671,In_2308);
or U1353 (N_1353,In_1702,In_1608);
or U1354 (N_1354,In_2753,In_2465);
or U1355 (N_1355,In_1366,In_2570);
nand U1356 (N_1356,In_709,In_652);
and U1357 (N_1357,In_2473,In_2806);
nor U1358 (N_1358,In_1671,In_491);
and U1359 (N_1359,In_655,In_1833);
and U1360 (N_1360,In_2297,In_2254);
or U1361 (N_1361,In_1523,In_1425);
nor U1362 (N_1362,In_1199,In_1535);
xnor U1363 (N_1363,In_2979,In_1988);
or U1364 (N_1364,In_1653,In_22);
nor U1365 (N_1365,In_1588,In_1813);
nor U1366 (N_1366,In_374,In_1338);
nor U1367 (N_1367,In_1238,In_2515);
nand U1368 (N_1368,In_1657,In_801);
xor U1369 (N_1369,In_2847,In_2381);
nand U1370 (N_1370,In_384,In_2169);
xor U1371 (N_1371,In_151,In_1762);
nor U1372 (N_1372,In_430,In_827);
nor U1373 (N_1373,In_1951,In_914);
nand U1374 (N_1374,In_2000,In_2678);
xor U1375 (N_1375,In_837,In_1490);
and U1376 (N_1376,In_1799,In_1195);
and U1377 (N_1377,In_1586,In_1395);
nand U1378 (N_1378,In_975,In_582);
nor U1379 (N_1379,In_2944,In_788);
or U1380 (N_1380,In_1719,In_2070);
and U1381 (N_1381,In_2018,In_2346);
nor U1382 (N_1382,In_268,In_298);
and U1383 (N_1383,In_1263,In_1396);
and U1384 (N_1384,In_944,In_1301);
xnor U1385 (N_1385,In_466,In_1551);
nand U1386 (N_1386,In_2610,In_2054);
or U1387 (N_1387,In_2152,In_2700);
xnor U1388 (N_1388,In_2876,In_303);
nor U1389 (N_1389,In_1035,In_1836);
or U1390 (N_1390,In_2015,In_734);
nand U1391 (N_1391,In_1294,In_2988);
nor U1392 (N_1392,In_668,In_850);
xnor U1393 (N_1393,In_245,In_300);
or U1394 (N_1394,In_1971,In_2970);
nand U1395 (N_1395,In_2379,In_197);
or U1396 (N_1396,In_2716,In_2985);
or U1397 (N_1397,In_851,In_592);
or U1398 (N_1398,In_2228,In_1964);
nand U1399 (N_1399,In_2215,In_1916);
xnor U1400 (N_1400,In_84,In_324);
and U1401 (N_1401,In_820,In_1892);
xor U1402 (N_1402,In_1936,In_821);
nor U1403 (N_1403,In_1517,In_1978);
and U1404 (N_1404,In_2752,In_2724);
nor U1405 (N_1405,In_2500,In_782);
nor U1406 (N_1406,In_371,In_1674);
xnor U1407 (N_1407,In_2837,In_2898);
and U1408 (N_1408,In_1085,In_2093);
nand U1409 (N_1409,In_2551,In_1463);
nor U1410 (N_1410,In_2243,In_2280);
nand U1411 (N_1411,In_2496,In_2819);
and U1412 (N_1412,In_2265,In_1968);
and U1413 (N_1413,In_2464,In_1758);
xnor U1414 (N_1414,In_2969,In_177);
nand U1415 (N_1415,In_2219,In_1298);
nand U1416 (N_1416,In_1989,In_672);
nor U1417 (N_1417,In_2331,In_44);
xor U1418 (N_1418,In_2516,In_90);
and U1419 (N_1419,In_2874,In_1612);
nor U1420 (N_1420,In_856,In_2163);
and U1421 (N_1421,In_2435,In_942);
xnor U1422 (N_1422,In_2195,In_224);
and U1423 (N_1423,In_708,In_269);
nand U1424 (N_1424,In_1243,In_250);
xnor U1425 (N_1425,In_2456,In_9);
nor U1426 (N_1426,In_2591,In_2536);
nor U1427 (N_1427,In_2646,In_1534);
and U1428 (N_1428,In_1629,In_1905);
nor U1429 (N_1429,In_646,In_2407);
and U1430 (N_1430,In_1479,In_2811);
nand U1431 (N_1431,In_1973,In_1412);
and U1432 (N_1432,In_2014,In_905);
xor U1433 (N_1433,In_1471,In_213);
or U1434 (N_1434,In_2796,In_1541);
or U1435 (N_1435,In_663,In_2539);
nand U1436 (N_1436,In_2795,In_2996);
xor U1437 (N_1437,In_1242,In_1038);
and U1438 (N_1438,In_686,In_2952);
or U1439 (N_1439,In_1075,In_1952);
and U1440 (N_1440,In_29,In_1449);
or U1441 (N_1441,In_180,In_167);
and U1442 (N_1442,In_955,In_214);
and U1443 (N_1443,In_1468,In_299);
or U1444 (N_1444,In_317,In_385);
nand U1445 (N_1445,In_302,In_1191);
nor U1446 (N_1446,In_2046,In_2056);
or U1447 (N_1447,In_509,In_1319);
and U1448 (N_1448,In_1433,In_1441);
nor U1449 (N_1449,In_1408,In_1826);
nand U1450 (N_1450,In_1476,In_1733);
or U1451 (N_1451,In_1410,In_1322);
nand U1452 (N_1452,In_2750,In_1459);
nor U1453 (N_1453,In_758,In_1282);
nand U1454 (N_1454,In_2767,In_2924);
nand U1455 (N_1455,In_2007,In_492);
and U1456 (N_1456,In_983,In_2794);
nor U1457 (N_1457,In_859,In_1428);
and U1458 (N_1458,In_1963,In_2286);
nand U1459 (N_1459,In_1391,In_1516);
or U1460 (N_1460,In_1367,In_2300);
nor U1461 (N_1461,In_1335,In_2205);
nor U1462 (N_1462,In_1919,In_691);
xnor U1463 (N_1463,In_2674,In_2333);
nand U1464 (N_1464,In_1728,In_2075);
xnor U1465 (N_1465,In_2078,In_230);
nor U1466 (N_1466,In_64,In_2655);
nand U1467 (N_1467,In_1103,In_2615);
xnor U1468 (N_1468,In_2378,In_1481);
nor U1469 (N_1469,In_1965,In_2708);
nand U1470 (N_1470,In_2314,In_2823);
nand U1471 (N_1471,In_505,In_648);
xor U1472 (N_1472,In_972,In_2274);
and U1473 (N_1473,In_1176,In_863);
nand U1474 (N_1474,In_2644,In_1791);
nand U1475 (N_1475,In_987,In_150);
nand U1476 (N_1476,In_2987,In_2953);
nand U1477 (N_1477,In_864,In_241);
or U1478 (N_1478,In_2745,In_2594);
or U1479 (N_1479,In_813,In_2383);
and U1480 (N_1480,In_2233,In_291);
xor U1481 (N_1481,In_378,In_1788);
and U1482 (N_1482,In_476,In_784);
nand U1483 (N_1483,In_1566,In_2232);
nand U1484 (N_1484,In_2792,In_2703);
nand U1485 (N_1485,In_1271,In_1427);
xor U1486 (N_1486,In_2405,In_2089);
and U1487 (N_1487,In_2694,In_1347);
and U1488 (N_1488,In_1846,In_290);
xor U1489 (N_1489,In_2917,In_2844);
nor U1490 (N_1490,In_1494,In_2672);
xor U1491 (N_1491,In_1130,In_28);
nand U1492 (N_1492,In_118,In_380);
and U1493 (N_1493,In_168,In_111);
nand U1494 (N_1494,In_1694,In_617);
xor U1495 (N_1495,In_116,In_2432);
and U1496 (N_1496,In_266,In_2483);
nor U1497 (N_1497,In_2051,In_678);
nand U1498 (N_1498,In_1444,In_2877);
nand U1499 (N_1499,In_497,In_2793);
or U1500 (N_1500,In_577,In_1982);
xor U1501 (N_1501,In_1377,In_1271);
nand U1502 (N_1502,In_2481,In_91);
xnor U1503 (N_1503,In_2201,In_71);
and U1504 (N_1504,In_663,In_2401);
or U1505 (N_1505,In_601,In_1536);
xnor U1506 (N_1506,In_1217,In_551);
nor U1507 (N_1507,In_1443,In_1924);
nor U1508 (N_1508,In_257,In_2581);
nand U1509 (N_1509,In_76,In_1492);
nor U1510 (N_1510,In_864,In_1704);
nor U1511 (N_1511,In_1516,In_126);
or U1512 (N_1512,In_2153,In_2206);
and U1513 (N_1513,In_358,In_81);
nor U1514 (N_1514,In_2199,In_503);
nand U1515 (N_1515,In_26,In_1894);
or U1516 (N_1516,In_2422,In_1373);
or U1517 (N_1517,In_2624,In_745);
or U1518 (N_1518,In_1426,In_2514);
or U1519 (N_1519,In_1629,In_208);
nor U1520 (N_1520,In_1520,In_2016);
and U1521 (N_1521,In_968,In_543);
and U1522 (N_1522,In_1577,In_21);
nand U1523 (N_1523,In_2100,In_2984);
and U1524 (N_1524,In_131,In_1750);
nand U1525 (N_1525,In_2602,In_2699);
xnor U1526 (N_1526,In_455,In_2299);
and U1527 (N_1527,In_1192,In_780);
and U1528 (N_1528,In_270,In_2104);
nor U1529 (N_1529,In_1043,In_2917);
nand U1530 (N_1530,In_567,In_290);
nor U1531 (N_1531,In_683,In_2451);
nand U1532 (N_1532,In_803,In_2469);
xnor U1533 (N_1533,In_1445,In_1404);
and U1534 (N_1534,In_16,In_421);
xor U1535 (N_1535,In_1665,In_2382);
nor U1536 (N_1536,In_772,In_280);
and U1537 (N_1537,In_2438,In_1479);
xnor U1538 (N_1538,In_745,In_749);
nand U1539 (N_1539,In_2494,In_1424);
nand U1540 (N_1540,In_302,In_1225);
xnor U1541 (N_1541,In_213,In_2500);
and U1542 (N_1542,In_1169,In_2941);
or U1543 (N_1543,In_40,In_2858);
xnor U1544 (N_1544,In_748,In_293);
nand U1545 (N_1545,In_1670,In_2339);
nor U1546 (N_1546,In_2881,In_1435);
nand U1547 (N_1547,In_1857,In_2318);
and U1548 (N_1548,In_895,In_989);
and U1549 (N_1549,In_41,In_890);
and U1550 (N_1550,In_1826,In_1222);
or U1551 (N_1551,In_1911,In_129);
xnor U1552 (N_1552,In_2274,In_2548);
xor U1553 (N_1553,In_603,In_1265);
nand U1554 (N_1554,In_344,In_2651);
nand U1555 (N_1555,In_657,In_1915);
nand U1556 (N_1556,In_1616,In_2697);
xor U1557 (N_1557,In_405,In_2268);
or U1558 (N_1558,In_2283,In_2532);
nor U1559 (N_1559,In_1548,In_939);
nor U1560 (N_1560,In_2718,In_821);
xnor U1561 (N_1561,In_1578,In_1427);
nand U1562 (N_1562,In_2064,In_1931);
or U1563 (N_1563,In_1836,In_510);
nor U1564 (N_1564,In_2644,In_2471);
and U1565 (N_1565,In_1609,In_1177);
nand U1566 (N_1566,In_1025,In_217);
and U1567 (N_1567,In_1281,In_921);
nor U1568 (N_1568,In_2425,In_1615);
or U1569 (N_1569,In_851,In_1109);
and U1570 (N_1570,In_312,In_1415);
or U1571 (N_1571,In_146,In_2753);
nor U1572 (N_1572,In_256,In_1349);
xnor U1573 (N_1573,In_1345,In_658);
nor U1574 (N_1574,In_1511,In_1650);
nand U1575 (N_1575,In_2945,In_1619);
or U1576 (N_1576,In_2329,In_599);
nand U1577 (N_1577,In_606,In_564);
nor U1578 (N_1578,In_2089,In_1328);
xnor U1579 (N_1579,In_370,In_373);
nor U1580 (N_1580,In_127,In_1511);
or U1581 (N_1581,In_688,In_1837);
and U1582 (N_1582,In_2426,In_2850);
xnor U1583 (N_1583,In_550,In_1349);
and U1584 (N_1584,In_825,In_1397);
nor U1585 (N_1585,In_2040,In_841);
nor U1586 (N_1586,In_1125,In_1920);
or U1587 (N_1587,In_1771,In_1322);
nand U1588 (N_1588,In_2771,In_2333);
xnor U1589 (N_1589,In_776,In_1657);
and U1590 (N_1590,In_350,In_1074);
nand U1591 (N_1591,In_2419,In_1599);
or U1592 (N_1592,In_644,In_650);
or U1593 (N_1593,In_1573,In_10);
xnor U1594 (N_1594,In_1937,In_1942);
nor U1595 (N_1595,In_1202,In_968);
nand U1596 (N_1596,In_845,In_1910);
xor U1597 (N_1597,In_1949,In_1514);
or U1598 (N_1598,In_2709,In_1367);
or U1599 (N_1599,In_1135,In_516);
or U1600 (N_1600,In_1007,In_1051);
nand U1601 (N_1601,In_784,In_2320);
nand U1602 (N_1602,In_2381,In_2409);
or U1603 (N_1603,In_1274,In_1176);
and U1604 (N_1604,In_1504,In_2422);
nand U1605 (N_1605,In_1960,In_773);
nand U1606 (N_1606,In_2928,In_1907);
or U1607 (N_1607,In_2022,In_1575);
or U1608 (N_1608,In_652,In_2580);
and U1609 (N_1609,In_1886,In_777);
or U1610 (N_1610,In_481,In_2252);
and U1611 (N_1611,In_1625,In_524);
and U1612 (N_1612,In_2855,In_1188);
xor U1613 (N_1613,In_1983,In_2130);
or U1614 (N_1614,In_2617,In_79);
or U1615 (N_1615,In_2060,In_52);
nand U1616 (N_1616,In_2898,In_2222);
or U1617 (N_1617,In_801,In_1081);
xnor U1618 (N_1618,In_1031,In_2918);
nand U1619 (N_1619,In_2379,In_2102);
xor U1620 (N_1620,In_903,In_2185);
or U1621 (N_1621,In_477,In_2706);
nor U1622 (N_1622,In_2315,In_2949);
nor U1623 (N_1623,In_2903,In_439);
and U1624 (N_1624,In_659,In_1980);
and U1625 (N_1625,In_217,In_1561);
xnor U1626 (N_1626,In_2651,In_2744);
or U1627 (N_1627,In_1194,In_1281);
nand U1628 (N_1628,In_1352,In_133);
and U1629 (N_1629,In_126,In_1751);
xor U1630 (N_1630,In_863,In_1555);
nor U1631 (N_1631,In_879,In_2877);
nand U1632 (N_1632,In_359,In_2756);
nor U1633 (N_1633,In_1806,In_825);
xnor U1634 (N_1634,In_1409,In_2765);
or U1635 (N_1635,In_2477,In_2701);
nor U1636 (N_1636,In_2929,In_1153);
or U1637 (N_1637,In_1498,In_2715);
xnor U1638 (N_1638,In_1449,In_670);
nand U1639 (N_1639,In_1449,In_1150);
and U1640 (N_1640,In_0,In_666);
xor U1641 (N_1641,In_2591,In_514);
nand U1642 (N_1642,In_983,In_2402);
nand U1643 (N_1643,In_915,In_681);
nand U1644 (N_1644,In_158,In_248);
nor U1645 (N_1645,In_1906,In_1978);
or U1646 (N_1646,In_580,In_2735);
or U1647 (N_1647,In_128,In_1379);
and U1648 (N_1648,In_2530,In_1362);
and U1649 (N_1649,In_2467,In_826);
nand U1650 (N_1650,In_1868,In_1795);
or U1651 (N_1651,In_2512,In_332);
xnor U1652 (N_1652,In_436,In_2369);
nor U1653 (N_1653,In_1273,In_1953);
nand U1654 (N_1654,In_2877,In_191);
nor U1655 (N_1655,In_2597,In_1386);
nor U1656 (N_1656,In_1278,In_25);
nor U1657 (N_1657,In_2485,In_2705);
nand U1658 (N_1658,In_1704,In_1453);
and U1659 (N_1659,In_1036,In_2711);
nor U1660 (N_1660,In_921,In_1386);
nor U1661 (N_1661,In_1214,In_2585);
xnor U1662 (N_1662,In_507,In_2468);
or U1663 (N_1663,In_103,In_1404);
nand U1664 (N_1664,In_2305,In_424);
nand U1665 (N_1665,In_1142,In_1246);
or U1666 (N_1666,In_181,In_1574);
and U1667 (N_1667,In_2815,In_143);
xnor U1668 (N_1668,In_1409,In_2622);
xnor U1669 (N_1669,In_433,In_713);
xor U1670 (N_1670,In_1108,In_2439);
xnor U1671 (N_1671,In_2719,In_1930);
and U1672 (N_1672,In_1127,In_2533);
nand U1673 (N_1673,In_558,In_1385);
xnor U1674 (N_1674,In_2268,In_189);
nor U1675 (N_1675,In_1245,In_1498);
or U1676 (N_1676,In_2167,In_1465);
nand U1677 (N_1677,In_1831,In_35);
and U1678 (N_1678,In_2631,In_1160);
nand U1679 (N_1679,In_946,In_319);
nor U1680 (N_1680,In_319,In_1757);
nand U1681 (N_1681,In_1992,In_358);
and U1682 (N_1682,In_1127,In_4);
xnor U1683 (N_1683,In_734,In_1732);
xor U1684 (N_1684,In_7,In_1336);
nor U1685 (N_1685,In_601,In_760);
nand U1686 (N_1686,In_83,In_551);
xor U1687 (N_1687,In_2856,In_77);
and U1688 (N_1688,In_67,In_45);
and U1689 (N_1689,In_63,In_2371);
or U1690 (N_1690,In_2267,In_322);
xnor U1691 (N_1691,In_1551,In_933);
xnor U1692 (N_1692,In_2176,In_2203);
nor U1693 (N_1693,In_2908,In_1215);
nor U1694 (N_1694,In_53,In_2086);
nor U1695 (N_1695,In_669,In_878);
and U1696 (N_1696,In_2567,In_1051);
nor U1697 (N_1697,In_2727,In_390);
nor U1698 (N_1698,In_2266,In_2479);
nand U1699 (N_1699,In_1810,In_470);
or U1700 (N_1700,In_339,In_500);
or U1701 (N_1701,In_168,In_1191);
nor U1702 (N_1702,In_2583,In_1015);
nand U1703 (N_1703,In_2715,In_1580);
nor U1704 (N_1704,In_1155,In_1119);
and U1705 (N_1705,In_2818,In_1911);
nand U1706 (N_1706,In_2279,In_1959);
or U1707 (N_1707,In_2837,In_2369);
nand U1708 (N_1708,In_1751,In_2762);
nor U1709 (N_1709,In_744,In_1931);
and U1710 (N_1710,In_25,In_189);
nand U1711 (N_1711,In_1197,In_2419);
xnor U1712 (N_1712,In_1069,In_1848);
nor U1713 (N_1713,In_482,In_1772);
and U1714 (N_1714,In_173,In_606);
nor U1715 (N_1715,In_1293,In_2429);
nand U1716 (N_1716,In_2077,In_1072);
or U1717 (N_1717,In_1283,In_263);
nor U1718 (N_1718,In_380,In_2899);
nor U1719 (N_1719,In_404,In_615);
and U1720 (N_1720,In_39,In_1167);
or U1721 (N_1721,In_198,In_2900);
xnor U1722 (N_1722,In_1849,In_2462);
nand U1723 (N_1723,In_1068,In_510);
and U1724 (N_1724,In_2259,In_142);
and U1725 (N_1725,In_2564,In_391);
xor U1726 (N_1726,In_193,In_1984);
nand U1727 (N_1727,In_1050,In_2961);
and U1728 (N_1728,In_2930,In_1680);
or U1729 (N_1729,In_2837,In_1593);
nand U1730 (N_1730,In_378,In_613);
or U1731 (N_1731,In_2043,In_1596);
xor U1732 (N_1732,In_879,In_603);
or U1733 (N_1733,In_2393,In_2114);
nor U1734 (N_1734,In_304,In_2058);
nand U1735 (N_1735,In_2379,In_1641);
or U1736 (N_1736,In_2498,In_258);
xnor U1737 (N_1737,In_2496,In_1344);
and U1738 (N_1738,In_182,In_1227);
or U1739 (N_1739,In_2007,In_2811);
xor U1740 (N_1740,In_1888,In_60);
nor U1741 (N_1741,In_1459,In_2886);
xnor U1742 (N_1742,In_2804,In_2651);
xor U1743 (N_1743,In_1776,In_376);
xnor U1744 (N_1744,In_1802,In_172);
nor U1745 (N_1745,In_138,In_1918);
or U1746 (N_1746,In_1239,In_2796);
nor U1747 (N_1747,In_2277,In_1136);
and U1748 (N_1748,In_669,In_2147);
or U1749 (N_1749,In_1794,In_1142);
xor U1750 (N_1750,In_702,In_1046);
nand U1751 (N_1751,In_1267,In_1695);
nand U1752 (N_1752,In_616,In_311);
nor U1753 (N_1753,In_2037,In_417);
xnor U1754 (N_1754,In_2957,In_1973);
nand U1755 (N_1755,In_1500,In_1501);
nor U1756 (N_1756,In_541,In_964);
xor U1757 (N_1757,In_1212,In_1889);
and U1758 (N_1758,In_2409,In_393);
or U1759 (N_1759,In_944,In_2032);
xnor U1760 (N_1760,In_1161,In_1679);
or U1761 (N_1761,In_568,In_2809);
xor U1762 (N_1762,In_224,In_1635);
xnor U1763 (N_1763,In_1333,In_2035);
nand U1764 (N_1764,In_2938,In_1471);
nand U1765 (N_1765,In_104,In_2230);
nor U1766 (N_1766,In_1321,In_2004);
nand U1767 (N_1767,In_2727,In_418);
and U1768 (N_1768,In_1126,In_2974);
nor U1769 (N_1769,In_258,In_1245);
nor U1770 (N_1770,In_2344,In_2332);
nor U1771 (N_1771,In_1323,In_2356);
and U1772 (N_1772,In_2445,In_2136);
nand U1773 (N_1773,In_2393,In_1227);
xnor U1774 (N_1774,In_2068,In_144);
xor U1775 (N_1775,In_19,In_2749);
nand U1776 (N_1776,In_723,In_846);
or U1777 (N_1777,In_913,In_331);
nor U1778 (N_1778,In_1245,In_213);
or U1779 (N_1779,In_1893,In_2425);
nor U1780 (N_1780,In_1261,In_375);
nand U1781 (N_1781,In_1262,In_1801);
and U1782 (N_1782,In_1120,In_59);
nand U1783 (N_1783,In_338,In_2123);
xor U1784 (N_1784,In_2060,In_2408);
nor U1785 (N_1785,In_2524,In_2253);
nor U1786 (N_1786,In_328,In_651);
nor U1787 (N_1787,In_2085,In_1163);
or U1788 (N_1788,In_1178,In_2425);
or U1789 (N_1789,In_2696,In_2768);
xnor U1790 (N_1790,In_2774,In_2187);
nor U1791 (N_1791,In_962,In_2484);
xor U1792 (N_1792,In_331,In_1168);
nor U1793 (N_1793,In_642,In_779);
or U1794 (N_1794,In_2321,In_695);
or U1795 (N_1795,In_722,In_1743);
nor U1796 (N_1796,In_2048,In_859);
xnor U1797 (N_1797,In_417,In_2536);
nand U1798 (N_1798,In_2196,In_2657);
nand U1799 (N_1799,In_1869,In_1139);
xnor U1800 (N_1800,In_2341,In_460);
or U1801 (N_1801,In_368,In_1304);
nor U1802 (N_1802,In_741,In_384);
and U1803 (N_1803,In_1717,In_2904);
or U1804 (N_1804,In_1338,In_2104);
nor U1805 (N_1805,In_103,In_610);
nor U1806 (N_1806,In_2135,In_721);
nor U1807 (N_1807,In_2613,In_1725);
or U1808 (N_1808,In_908,In_1710);
nor U1809 (N_1809,In_796,In_94);
nand U1810 (N_1810,In_2771,In_391);
and U1811 (N_1811,In_2253,In_459);
nor U1812 (N_1812,In_358,In_296);
xnor U1813 (N_1813,In_1560,In_1228);
nor U1814 (N_1814,In_2973,In_807);
nor U1815 (N_1815,In_990,In_2144);
or U1816 (N_1816,In_290,In_2086);
or U1817 (N_1817,In_2623,In_2518);
or U1818 (N_1818,In_525,In_1503);
and U1819 (N_1819,In_690,In_1880);
or U1820 (N_1820,In_579,In_1959);
or U1821 (N_1821,In_1830,In_1123);
nor U1822 (N_1822,In_2414,In_1215);
and U1823 (N_1823,In_2842,In_1274);
and U1824 (N_1824,In_2894,In_1717);
nor U1825 (N_1825,In_1438,In_1156);
or U1826 (N_1826,In_2174,In_690);
and U1827 (N_1827,In_2420,In_1893);
nor U1828 (N_1828,In_156,In_1144);
xor U1829 (N_1829,In_1252,In_2403);
or U1830 (N_1830,In_1780,In_1226);
xor U1831 (N_1831,In_734,In_1023);
nand U1832 (N_1832,In_215,In_38);
nand U1833 (N_1833,In_2022,In_2079);
xor U1834 (N_1834,In_2426,In_289);
nand U1835 (N_1835,In_1064,In_2922);
and U1836 (N_1836,In_2606,In_24);
xor U1837 (N_1837,In_824,In_2558);
or U1838 (N_1838,In_2602,In_1245);
or U1839 (N_1839,In_1948,In_1274);
xor U1840 (N_1840,In_1895,In_1229);
or U1841 (N_1841,In_1429,In_1972);
nor U1842 (N_1842,In_2734,In_2193);
nor U1843 (N_1843,In_2267,In_1083);
nor U1844 (N_1844,In_374,In_1448);
nor U1845 (N_1845,In_996,In_2064);
or U1846 (N_1846,In_2532,In_168);
or U1847 (N_1847,In_1379,In_1507);
xor U1848 (N_1848,In_2059,In_2825);
nor U1849 (N_1849,In_2021,In_2198);
xor U1850 (N_1850,In_2701,In_1653);
nand U1851 (N_1851,In_844,In_1675);
nor U1852 (N_1852,In_2588,In_1);
or U1853 (N_1853,In_546,In_1466);
and U1854 (N_1854,In_1681,In_2975);
and U1855 (N_1855,In_2708,In_97);
nor U1856 (N_1856,In_629,In_1000);
nand U1857 (N_1857,In_2631,In_1186);
and U1858 (N_1858,In_1638,In_2741);
or U1859 (N_1859,In_2205,In_2291);
or U1860 (N_1860,In_1854,In_1085);
nand U1861 (N_1861,In_320,In_1502);
nand U1862 (N_1862,In_1879,In_268);
xor U1863 (N_1863,In_1929,In_1727);
nor U1864 (N_1864,In_909,In_2935);
nor U1865 (N_1865,In_2035,In_1512);
nand U1866 (N_1866,In_614,In_267);
and U1867 (N_1867,In_962,In_2815);
and U1868 (N_1868,In_1042,In_2062);
and U1869 (N_1869,In_2782,In_724);
xor U1870 (N_1870,In_1875,In_704);
nand U1871 (N_1871,In_501,In_2276);
nor U1872 (N_1872,In_2758,In_890);
xnor U1873 (N_1873,In_374,In_294);
and U1874 (N_1874,In_909,In_1043);
xor U1875 (N_1875,In_989,In_1143);
nor U1876 (N_1876,In_1593,In_2134);
nor U1877 (N_1877,In_729,In_2942);
xnor U1878 (N_1878,In_1980,In_1548);
and U1879 (N_1879,In_1881,In_701);
or U1880 (N_1880,In_2704,In_2993);
and U1881 (N_1881,In_899,In_2991);
and U1882 (N_1882,In_2116,In_554);
nor U1883 (N_1883,In_334,In_1059);
nor U1884 (N_1884,In_704,In_1343);
xor U1885 (N_1885,In_383,In_1383);
or U1886 (N_1886,In_965,In_2535);
nor U1887 (N_1887,In_600,In_915);
xnor U1888 (N_1888,In_1361,In_1736);
nand U1889 (N_1889,In_1904,In_652);
xnor U1890 (N_1890,In_697,In_193);
and U1891 (N_1891,In_2844,In_480);
nor U1892 (N_1892,In_163,In_1458);
or U1893 (N_1893,In_1905,In_1889);
nand U1894 (N_1894,In_1614,In_501);
or U1895 (N_1895,In_1552,In_1768);
or U1896 (N_1896,In_2575,In_438);
and U1897 (N_1897,In_1056,In_1253);
nor U1898 (N_1898,In_757,In_2335);
or U1899 (N_1899,In_1366,In_685);
and U1900 (N_1900,In_2366,In_1347);
nand U1901 (N_1901,In_1848,In_1989);
nand U1902 (N_1902,In_2994,In_10);
or U1903 (N_1903,In_2200,In_2032);
or U1904 (N_1904,In_2316,In_2687);
or U1905 (N_1905,In_1968,In_1977);
nor U1906 (N_1906,In_2863,In_2813);
or U1907 (N_1907,In_2214,In_157);
xor U1908 (N_1908,In_764,In_1453);
xnor U1909 (N_1909,In_780,In_282);
xnor U1910 (N_1910,In_2727,In_2789);
xor U1911 (N_1911,In_2437,In_2404);
xnor U1912 (N_1912,In_1329,In_203);
xnor U1913 (N_1913,In_2009,In_258);
and U1914 (N_1914,In_599,In_1692);
xnor U1915 (N_1915,In_91,In_610);
and U1916 (N_1916,In_2851,In_545);
nand U1917 (N_1917,In_1825,In_1987);
nand U1918 (N_1918,In_1906,In_1112);
xor U1919 (N_1919,In_269,In_815);
or U1920 (N_1920,In_600,In_632);
xor U1921 (N_1921,In_2677,In_1308);
nand U1922 (N_1922,In_2128,In_291);
nor U1923 (N_1923,In_497,In_820);
nand U1924 (N_1924,In_1912,In_1281);
nand U1925 (N_1925,In_1102,In_537);
or U1926 (N_1926,In_2971,In_1916);
nor U1927 (N_1927,In_2750,In_2755);
nor U1928 (N_1928,In_1255,In_1325);
nor U1929 (N_1929,In_229,In_2587);
nor U1930 (N_1930,In_1036,In_1265);
nor U1931 (N_1931,In_1377,In_495);
nand U1932 (N_1932,In_2112,In_2649);
or U1933 (N_1933,In_279,In_1622);
and U1934 (N_1934,In_806,In_361);
or U1935 (N_1935,In_1681,In_386);
xor U1936 (N_1936,In_2628,In_2144);
nand U1937 (N_1937,In_1730,In_130);
nor U1938 (N_1938,In_835,In_2621);
nor U1939 (N_1939,In_751,In_2942);
xor U1940 (N_1940,In_1895,In_1164);
nor U1941 (N_1941,In_2267,In_1755);
or U1942 (N_1942,In_2897,In_807);
nor U1943 (N_1943,In_1863,In_2390);
nand U1944 (N_1944,In_2368,In_1447);
and U1945 (N_1945,In_412,In_1562);
or U1946 (N_1946,In_2916,In_2693);
nand U1947 (N_1947,In_2819,In_311);
and U1948 (N_1948,In_1336,In_2989);
xor U1949 (N_1949,In_1233,In_333);
or U1950 (N_1950,In_2524,In_1463);
xor U1951 (N_1951,In_1373,In_489);
nand U1952 (N_1952,In_315,In_2309);
or U1953 (N_1953,In_2145,In_578);
nand U1954 (N_1954,In_2457,In_363);
or U1955 (N_1955,In_1999,In_1216);
or U1956 (N_1956,In_424,In_464);
or U1957 (N_1957,In_2860,In_406);
or U1958 (N_1958,In_656,In_828);
or U1959 (N_1959,In_911,In_1128);
and U1960 (N_1960,In_1001,In_427);
xnor U1961 (N_1961,In_2154,In_2159);
nor U1962 (N_1962,In_22,In_2294);
and U1963 (N_1963,In_232,In_2985);
nor U1964 (N_1964,In_2719,In_579);
nor U1965 (N_1965,In_2095,In_757);
nor U1966 (N_1966,In_2292,In_1075);
and U1967 (N_1967,In_2563,In_182);
and U1968 (N_1968,In_1485,In_2704);
nand U1969 (N_1969,In_1690,In_1338);
and U1970 (N_1970,In_1842,In_18);
or U1971 (N_1971,In_990,In_2733);
nand U1972 (N_1972,In_1846,In_2452);
or U1973 (N_1973,In_1242,In_1013);
nand U1974 (N_1974,In_1960,In_148);
nor U1975 (N_1975,In_1214,In_322);
nand U1976 (N_1976,In_2104,In_2383);
or U1977 (N_1977,In_129,In_1142);
nor U1978 (N_1978,In_897,In_904);
and U1979 (N_1979,In_2353,In_83);
nand U1980 (N_1980,In_2901,In_2467);
and U1981 (N_1981,In_206,In_1130);
nand U1982 (N_1982,In_761,In_2333);
and U1983 (N_1983,In_159,In_617);
nand U1984 (N_1984,In_1286,In_1676);
xor U1985 (N_1985,In_1664,In_2441);
and U1986 (N_1986,In_609,In_1511);
nor U1987 (N_1987,In_690,In_235);
nand U1988 (N_1988,In_1675,In_1883);
or U1989 (N_1989,In_952,In_124);
xnor U1990 (N_1990,In_2555,In_1458);
xor U1991 (N_1991,In_2263,In_2719);
nor U1992 (N_1992,In_1225,In_967);
and U1993 (N_1993,In_2573,In_2043);
or U1994 (N_1994,In_2587,In_805);
or U1995 (N_1995,In_325,In_2448);
nand U1996 (N_1996,In_2070,In_846);
and U1997 (N_1997,In_470,In_2661);
or U1998 (N_1998,In_18,In_1509);
nand U1999 (N_1999,In_1878,In_1876);
nand U2000 (N_2000,In_2006,In_2639);
nor U2001 (N_2001,In_1932,In_2111);
xnor U2002 (N_2002,In_2733,In_1222);
nor U2003 (N_2003,In_931,In_254);
nand U2004 (N_2004,In_481,In_1994);
and U2005 (N_2005,In_1032,In_2748);
nor U2006 (N_2006,In_766,In_2219);
nand U2007 (N_2007,In_1973,In_1364);
nor U2008 (N_2008,In_225,In_673);
and U2009 (N_2009,In_203,In_262);
nand U2010 (N_2010,In_411,In_380);
and U2011 (N_2011,In_2504,In_32);
or U2012 (N_2012,In_78,In_1263);
or U2013 (N_2013,In_590,In_717);
nor U2014 (N_2014,In_1581,In_2920);
nand U2015 (N_2015,In_2122,In_2264);
nor U2016 (N_2016,In_257,In_2781);
nor U2017 (N_2017,In_2771,In_326);
xnor U2018 (N_2018,In_1010,In_1018);
nand U2019 (N_2019,In_262,In_2178);
nor U2020 (N_2020,In_916,In_607);
nor U2021 (N_2021,In_1060,In_1243);
nor U2022 (N_2022,In_697,In_1352);
nor U2023 (N_2023,In_107,In_1402);
xnor U2024 (N_2024,In_1866,In_1447);
nand U2025 (N_2025,In_2671,In_281);
nor U2026 (N_2026,In_1248,In_520);
or U2027 (N_2027,In_2861,In_2740);
nand U2028 (N_2028,In_2881,In_2188);
and U2029 (N_2029,In_969,In_1074);
or U2030 (N_2030,In_1937,In_1196);
nor U2031 (N_2031,In_951,In_248);
nand U2032 (N_2032,In_1910,In_2828);
or U2033 (N_2033,In_341,In_1742);
nand U2034 (N_2034,In_2338,In_2614);
or U2035 (N_2035,In_444,In_2920);
and U2036 (N_2036,In_2162,In_2791);
or U2037 (N_2037,In_585,In_1519);
nand U2038 (N_2038,In_2776,In_684);
nor U2039 (N_2039,In_2934,In_1397);
xor U2040 (N_2040,In_2262,In_1611);
and U2041 (N_2041,In_632,In_1639);
nand U2042 (N_2042,In_2331,In_944);
xor U2043 (N_2043,In_1720,In_1938);
nor U2044 (N_2044,In_20,In_1607);
and U2045 (N_2045,In_2853,In_1990);
nor U2046 (N_2046,In_1437,In_1021);
or U2047 (N_2047,In_1142,In_2300);
nand U2048 (N_2048,In_657,In_1714);
nand U2049 (N_2049,In_930,In_2773);
xnor U2050 (N_2050,In_2787,In_2728);
and U2051 (N_2051,In_2128,In_926);
nor U2052 (N_2052,In_2579,In_1338);
or U2053 (N_2053,In_2093,In_1899);
or U2054 (N_2054,In_1337,In_2667);
nor U2055 (N_2055,In_2556,In_1700);
nand U2056 (N_2056,In_1462,In_253);
xor U2057 (N_2057,In_870,In_1582);
and U2058 (N_2058,In_1467,In_1988);
xor U2059 (N_2059,In_2578,In_1035);
nand U2060 (N_2060,In_1916,In_240);
xor U2061 (N_2061,In_971,In_941);
xor U2062 (N_2062,In_1217,In_2342);
nand U2063 (N_2063,In_1993,In_1303);
or U2064 (N_2064,In_2192,In_1418);
and U2065 (N_2065,In_2495,In_2461);
xnor U2066 (N_2066,In_1591,In_2526);
and U2067 (N_2067,In_2096,In_404);
or U2068 (N_2068,In_1512,In_2118);
xnor U2069 (N_2069,In_2362,In_1511);
nand U2070 (N_2070,In_1558,In_1459);
or U2071 (N_2071,In_2925,In_217);
and U2072 (N_2072,In_2134,In_866);
xnor U2073 (N_2073,In_133,In_2506);
or U2074 (N_2074,In_324,In_2147);
xnor U2075 (N_2075,In_1318,In_2521);
nor U2076 (N_2076,In_415,In_92);
nand U2077 (N_2077,In_1436,In_2865);
nand U2078 (N_2078,In_2636,In_2371);
nor U2079 (N_2079,In_1327,In_2039);
or U2080 (N_2080,In_663,In_252);
or U2081 (N_2081,In_1444,In_2849);
xnor U2082 (N_2082,In_2380,In_2107);
and U2083 (N_2083,In_2619,In_2902);
xor U2084 (N_2084,In_1416,In_1529);
xor U2085 (N_2085,In_2675,In_25);
xor U2086 (N_2086,In_2199,In_1574);
nand U2087 (N_2087,In_1095,In_443);
xnor U2088 (N_2088,In_2744,In_1557);
nand U2089 (N_2089,In_2809,In_60);
nand U2090 (N_2090,In_2850,In_2407);
nand U2091 (N_2091,In_617,In_926);
xnor U2092 (N_2092,In_2432,In_2703);
nor U2093 (N_2093,In_671,In_151);
and U2094 (N_2094,In_1928,In_2820);
nor U2095 (N_2095,In_2506,In_947);
nand U2096 (N_2096,In_231,In_1682);
xnor U2097 (N_2097,In_1328,In_1783);
nand U2098 (N_2098,In_741,In_1310);
xnor U2099 (N_2099,In_218,In_260);
and U2100 (N_2100,In_555,In_884);
and U2101 (N_2101,In_639,In_1855);
or U2102 (N_2102,In_2589,In_1363);
xnor U2103 (N_2103,In_1690,In_2389);
xnor U2104 (N_2104,In_848,In_480);
or U2105 (N_2105,In_1356,In_1528);
nand U2106 (N_2106,In_1789,In_1169);
nor U2107 (N_2107,In_2103,In_613);
nor U2108 (N_2108,In_765,In_1489);
nand U2109 (N_2109,In_1911,In_1826);
nand U2110 (N_2110,In_2302,In_1063);
nand U2111 (N_2111,In_2663,In_1517);
or U2112 (N_2112,In_401,In_902);
and U2113 (N_2113,In_0,In_200);
xor U2114 (N_2114,In_394,In_2284);
or U2115 (N_2115,In_666,In_2756);
nand U2116 (N_2116,In_2305,In_1284);
nor U2117 (N_2117,In_938,In_2203);
and U2118 (N_2118,In_392,In_2080);
nor U2119 (N_2119,In_545,In_1348);
or U2120 (N_2120,In_709,In_1873);
nand U2121 (N_2121,In_1614,In_2381);
nor U2122 (N_2122,In_2967,In_1023);
nor U2123 (N_2123,In_630,In_2576);
nand U2124 (N_2124,In_1187,In_1046);
and U2125 (N_2125,In_666,In_2604);
and U2126 (N_2126,In_2750,In_2530);
nand U2127 (N_2127,In_2392,In_1316);
nand U2128 (N_2128,In_428,In_2603);
or U2129 (N_2129,In_1002,In_2907);
xor U2130 (N_2130,In_1155,In_847);
and U2131 (N_2131,In_1459,In_1152);
nor U2132 (N_2132,In_1912,In_198);
xor U2133 (N_2133,In_929,In_1689);
or U2134 (N_2134,In_758,In_446);
or U2135 (N_2135,In_1966,In_314);
nand U2136 (N_2136,In_1561,In_1816);
xnor U2137 (N_2137,In_1496,In_28);
nand U2138 (N_2138,In_239,In_14);
nor U2139 (N_2139,In_346,In_1831);
nor U2140 (N_2140,In_2266,In_1418);
nor U2141 (N_2141,In_2107,In_2331);
or U2142 (N_2142,In_1549,In_1350);
xor U2143 (N_2143,In_2323,In_1026);
nand U2144 (N_2144,In_1727,In_2919);
or U2145 (N_2145,In_2636,In_1166);
xor U2146 (N_2146,In_2500,In_2097);
or U2147 (N_2147,In_2805,In_1441);
or U2148 (N_2148,In_2160,In_1284);
and U2149 (N_2149,In_2389,In_2975);
nand U2150 (N_2150,In_1967,In_447);
nor U2151 (N_2151,In_1702,In_2759);
nand U2152 (N_2152,In_678,In_1187);
and U2153 (N_2153,In_1045,In_567);
nor U2154 (N_2154,In_606,In_1644);
xnor U2155 (N_2155,In_2397,In_2389);
nand U2156 (N_2156,In_830,In_2108);
xnor U2157 (N_2157,In_672,In_1568);
and U2158 (N_2158,In_489,In_1146);
or U2159 (N_2159,In_1748,In_879);
and U2160 (N_2160,In_2857,In_798);
nand U2161 (N_2161,In_1439,In_648);
nor U2162 (N_2162,In_10,In_356);
nor U2163 (N_2163,In_599,In_621);
xnor U2164 (N_2164,In_54,In_1697);
nor U2165 (N_2165,In_2004,In_1343);
and U2166 (N_2166,In_119,In_2519);
xnor U2167 (N_2167,In_88,In_239);
or U2168 (N_2168,In_1635,In_1203);
or U2169 (N_2169,In_1357,In_827);
and U2170 (N_2170,In_2411,In_1024);
or U2171 (N_2171,In_2188,In_759);
nor U2172 (N_2172,In_446,In_1679);
or U2173 (N_2173,In_1967,In_2746);
nand U2174 (N_2174,In_717,In_1292);
nand U2175 (N_2175,In_688,In_2454);
or U2176 (N_2176,In_2703,In_1508);
or U2177 (N_2177,In_525,In_196);
nor U2178 (N_2178,In_1109,In_2774);
xnor U2179 (N_2179,In_1844,In_284);
and U2180 (N_2180,In_1100,In_2074);
or U2181 (N_2181,In_134,In_727);
or U2182 (N_2182,In_364,In_859);
and U2183 (N_2183,In_2832,In_2652);
nand U2184 (N_2184,In_2391,In_1391);
or U2185 (N_2185,In_2620,In_2299);
nor U2186 (N_2186,In_1737,In_1459);
nand U2187 (N_2187,In_1146,In_164);
nand U2188 (N_2188,In_628,In_2572);
nand U2189 (N_2189,In_2566,In_828);
nand U2190 (N_2190,In_2554,In_771);
nand U2191 (N_2191,In_1461,In_2619);
and U2192 (N_2192,In_631,In_2417);
nor U2193 (N_2193,In_1921,In_1419);
nand U2194 (N_2194,In_2898,In_2450);
nor U2195 (N_2195,In_540,In_1861);
nor U2196 (N_2196,In_1219,In_1235);
and U2197 (N_2197,In_2658,In_2310);
nand U2198 (N_2198,In_2064,In_2934);
xor U2199 (N_2199,In_2914,In_1220);
and U2200 (N_2200,In_2212,In_1828);
xnor U2201 (N_2201,In_382,In_1346);
and U2202 (N_2202,In_2503,In_683);
xnor U2203 (N_2203,In_160,In_609);
nor U2204 (N_2204,In_2,In_1948);
nor U2205 (N_2205,In_1229,In_2636);
nand U2206 (N_2206,In_1994,In_2436);
nor U2207 (N_2207,In_2858,In_2600);
xor U2208 (N_2208,In_1624,In_1258);
nor U2209 (N_2209,In_7,In_2641);
nand U2210 (N_2210,In_1484,In_2053);
or U2211 (N_2211,In_1341,In_535);
nor U2212 (N_2212,In_1019,In_2895);
nand U2213 (N_2213,In_926,In_2522);
and U2214 (N_2214,In_2022,In_17);
nand U2215 (N_2215,In_96,In_2378);
nand U2216 (N_2216,In_702,In_848);
nor U2217 (N_2217,In_2437,In_2598);
nand U2218 (N_2218,In_1189,In_1246);
nand U2219 (N_2219,In_2815,In_2791);
or U2220 (N_2220,In_2713,In_2206);
nand U2221 (N_2221,In_642,In_2577);
and U2222 (N_2222,In_2981,In_948);
and U2223 (N_2223,In_2489,In_1863);
and U2224 (N_2224,In_427,In_404);
or U2225 (N_2225,In_710,In_679);
xor U2226 (N_2226,In_1222,In_1673);
nor U2227 (N_2227,In_274,In_334);
xor U2228 (N_2228,In_845,In_2235);
and U2229 (N_2229,In_2536,In_2635);
nor U2230 (N_2230,In_2856,In_1928);
nand U2231 (N_2231,In_989,In_1898);
nand U2232 (N_2232,In_2282,In_2170);
xor U2233 (N_2233,In_1478,In_235);
and U2234 (N_2234,In_1217,In_1622);
or U2235 (N_2235,In_419,In_2410);
xor U2236 (N_2236,In_1111,In_83);
nor U2237 (N_2237,In_2220,In_443);
xor U2238 (N_2238,In_771,In_1279);
xnor U2239 (N_2239,In_28,In_2316);
nand U2240 (N_2240,In_1572,In_2712);
or U2241 (N_2241,In_2106,In_2834);
or U2242 (N_2242,In_2690,In_2990);
nand U2243 (N_2243,In_2345,In_2116);
or U2244 (N_2244,In_2315,In_2598);
nand U2245 (N_2245,In_2590,In_2473);
and U2246 (N_2246,In_82,In_2518);
xor U2247 (N_2247,In_68,In_1969);
and U2248 (N_2248,In_1532,In_1950);
nor U2249 (N_2249,In_34,In_1183);
nand U2250 (N_2250,In_1689,In_1658);
or U2251 (N_2251,In_2937,In_2822);
and U2252 (N_2252,In_1559,In_1737);
nand U2253 (N_2253,In_2080,In_1230);
and U2254 (N_2254,In_2236,In_516);
or U2255 (N_2255,In_200,In_2151);
and U2256 (N_2256,In_1163,In_192);
and U2257 (N_2257,In_1377,In_808);
nor U2258 (N_2258,In_1033,In_2588);
xor U2259 (N_2259,In_686,In_1688);
or U2260 (N_2260,In_1559,In_1579);
or U2261 (N_2261,In_389,In_2038);
xnor U2262 (N_2262,In_2672,In_2027);
nand U2263 (N_2263,In_414,In_2379);
or U2264 (N_2264,In_204,In_1477);
nor U2265 (N_2265,In_988,In_1041);
xor U2266 (N_2266,In_2629,In_1203);
nand U2267 (N_2267,In_1392,In_2439);
nand U2268 (N_2268,In_819,In_2505);
nor U2269 (N_2269,In_2065,In_1506);
nor U2270 (N_2270,In_1009,In_18);
nor U2271 (N_2271,In_1327,In_803);
xor U2272 (N_2272,In_185,In_2967);
nand U2273 (N_2273,In_2838,In_1883);
nand U2274 (N_2274,In_2298,In_1562);
and U2275 (N_2275,In_463,In_213);
xnor U2276 (N_2276,In_2042,In_2818);
nor U2277 (N_2277,In_1976,In_1559);
or U2278 (N_2278,In_609,In_2085);
and U2279 (N_2279,In_515,In_2248);
or U2280 (N_2280,In_667,In_316);
or U2281 (N_2281,In_2236,In_273);
nor U2282 (N_2282,In_1002,In_1989);
xor U2283 (N_2283,In_2836,In_79);
and U2284 (N_2284,In_590,In_1948);
xor U2285 (N_2285,In_2932,In_583);
or U2286 (N_2286,In_2421,In_954);
nand U2287 (N_2287,In_2784,In_1816);
and U2288 (N_2288,In_50,In_791);
or U2289 (N_2289,In_1049,In_2469);
or U2290 (N_2290,In_2585,In_895);
xnor U2291 (N_2291,In_410,In_588);
nor U2292 (N_2292,In_1034,In_1037);
nor U2293 (N_2293,In_710,In_80);
nand U2294 (N_2294,In_799,In_1754);
and U2295 (N_2295,In_1367,In_869);
xnor U2296 (N_2296,In_2053,In_2530);
and U2297 (N_2297,In_1281,In_2115);
or U2298 (N_2298,In_150,In_2392);
nand U2299 (N_2299,In_1165,In_2976);
and U2300 (N_2300,In_165,In_1248);
xor U2301 (N_2301,In_2658,In_2076);
and U2302 (N_2302,In_1488,In_922);
or U2303 (N_2303,In_2188,In_1923);
xor U2304 (N_2304,In_474,In_724);
or U2305 (N_2305,In_1962,In_1275);
nor U2306 (N_2306,In_492,In_179);
or U2307 (N_2307,In_680,In_780);
or U2308 (N_2308,In_1889,In_2153);
xnor U2309 (N_2309,In_2670,In_863);
nor U2310 (N_2310,In_350,In_562);
or U2311 (N_2311,In_1307,In_2029);
xnor U2312 (N_2312,In_131,In_1179);
nand U2313 (N_2313,In_2563,In_1886);
or U2314 (N_2314,In_442,In_929);
or U2315 (N_2315,In_2497,In_487);
or U2316 (N_2316,In_379,In_2136);
or U2317 (N_2317,In_603,In_536);
and U2318 (N_2318,In_371,In_519);
nor U2319 (N_2319,In_2614,In_1545);
and U2320 (N_2320,In_2127,In_744);
xor U2321 (N_2321,In_2864,In_1833);
xnor U2322 (N_2322,In_1264,In_182);
nand U2323 (N_2323,In_1528,In_2877);
and U2324 (N_2324,In_2216,In_2373);
nand U2325 (N_2325,In_1606,In_2600);
nand U2326 (N_2326,In_1340,In_1987);
xnor U2327 (N_2327,In_252,In_2722);
xor U2328 (N_2328,In_196,In_708);
nor U2329 (N_2329,In_302,In_1211);
nor U2330 (N_2330,In_2305,In_1361);
nand U2331 (N_2331,In_1143,In_916);
xor U2332 (N_2332,In_898,In_752);
nor U2333 (N_2333,In_2058,In_1795);
and U2334 (N_2334,In_1509,In_949);
nand U2335 (N_2335,In_1740,In_907);
xor U2336 (N_2336,In_169,In_2451);
nand U2337 (N_2337,In_2013,In_2193);
xnor U2338 (N_2338,In_1170,In_184);
xnor U2339 (N_2339,In_1037,In_1979);
or U2340 (N_2340,In_2179,In_1873);
xor U2341 (N_2341,In_998,In_190);
or U2342 (N_2342,In_2228,In_1086);
or U2343 (N_2343,In_1687,In_1943);
nor U2344 (N_2344,In_2937,In_2640);
xnor U2345 (N_2345,In_1367,In_135);
or U2346 (N_2346,In_2705,In_1655);
nand U2347 (N_2347,In_2182,In_617);
or U2348 (N_2348,In_2821,In_2648);
and U2349 (N_2349,In_823,In_267);
xnor U2350 (N_2350,In_341,In_2100);
nand U2351 (N_2351,In_1582,In_1407);
or U2352 (N_2352,In_212,In_904);
nand U2353 (N_2353,In_473,In_61);
nor U2354 (N_2354,In_716,In_961);
and U2355 (N_2355,In_1020,In_290);
and U2356 (N_2356,In_200,In_2905);
xor U2357 (N_2357,In_2336,In_425);
xnor U2358 (N_2358,In_1250,In_2094);
nor U2359 (N_2359,In_2617,In_2540);
nor U2360 (N_2360,In_73,In_1620);
nand U2361 (N_2361,In_2926,In_2942);
or U2362 (N_2362,In_1640,In_982);
nand U2363 (N_2363,In_2379,In_2224);
or U2364 (N_2364,In_1530,In_2137);
nor U2365 (N_2365,In_2923,In_1442);
nor U2366 (N_2366,In_2187,In_1297);
nand U2367 (N_2367,In_705,In_604);
xor U2368 (N_2368,In_703,In_1194);
or U2369 (N_2369,In_1637,In_594);
and U2370 (N_2370,In_1034,In_53);
and U2371 (N_2371,In_484,In_706);
xor U2372 (N_2372,In_665,In_2634);
nor U2373 (N_2373,In_1317,In_1982);
nor U2374 (N_2374,In_287,In_2237);
nor U2375 (N_2375,In_376,In_1015);
xnor U2376 (N_2376,In_1790,In_1504);
and U2377 (N_2377,In_50,In_2541);
or U2378 (N_2378,In_711,In_1514);
xnor U2379 (N_2379,In_2105,In_1012);
and U2380 (N_2380,In_859,In_2962);
or U2381 (N_2381,In_2194,In_990);
and U2382 (N_2382,In_557,In_2992);
nand U2383 (N_2383,In_430,In_1616);
nor U2384 (N_2384,In_1850,In_124);
nand U2385 (N_2385,In_2752,In_817);
xor U2386 (N_2386,In_197,In_2994);
and U2387 (N_2387,In_1974,In_1781);
and U2388 (N_2388,In_242,In_1834);
and U2389 (N_2389,In_1678,In_2413);
and U2390 (N_2390,In_1358,In_2081);
and U2391 (N_2391,In_1599,In_2705);
nor U2392 (N_2392,In_1146,In_720);
or U2393 (N_2393,In_399,In_1490);
nor U2394 (N_2394,In_669,In_1820);
nor U2395 (N_2395,In_798,In_889);
nand U2396 (N_2396,In_272,In_1630);
and U2397 (N_2397,In_2589,In_2383);
nand U2398 (N_2398,In_628,In_2104);
and U2399 (N_2399,In_1661,In_2953);
nand U2400 (N_2400,In_559,In_1173);
nand U2401 (N_2401,In_1103,In_1224);
or U2402 (N_2402,In_1192,In_1003);
and U2403 (N_2403,In_2082,In_847);
or U2404 (N_2404,In_2003,In_1509);
nand U2405 (N_2405,In_2544,In_453);
or U2406 (N_2406,In_2852,In_2483);
or U2407 (N_2407,In_2996,In_2108);
nor U2408 (N_2408,In_1278,In_33);
or U2409 (N_2409,In_145,In_2406);
or U2410 (N_2410,In_1878,In_2030);
and U2411 (N_2411,In_2008,In_912);
xnor U2412 (N_2412,In_1729,In_1714);
and U2413 (N_2413,In_4,In_1602);
nand U2414 (N_2414,In_2405,In_604);
nand U2415 (N_2415,In_246,In_832);
nor U2416 (N_2416,In_97,In_2230);
nand U2417 (N_2417,In_181,In_1354);
xor U2418 (N_2418,In_2523,In_316);
nand U2419 (N_2419,In_310,In_2194);
nor U2420 (N_2420,In_1276,In_509);
nor U2421 (N_2421,In_1816,In_238);
nand U2422 (N_2422,In_2750,In_1165);
xor U2423 (N_2423,In_1086,In_4);
nor U2424 (N_2424,In_2661,In_1176);
and U2425 (N_2425,In_1196,In_1622);
nor U2426 (N_2426,In_235,In_1485);
nand U2427 (N_2427,In_2238,In_1393);
and U2428 (N_2428,In_1528,In_1522);
xor U2429 (N_2429,In_2651,In_1402);
xnor U2430 (N_2430,In_1703,In_372);
nor U2431 (N_2431,In_1001,In_652);
or U2432 (N_2432,In_940,In_547);
and U2433 (N_2433,In_2224,In_1265);
and U2434 (N_2434,In_2371,In_1507);
nand U2435 (N_2435,In_1948,In_497);
or U2436 (N_2436,In_1663,In_225);
or U2437 (N_2437,In_594,In_1063);
nor U2438 (N_2438,In_2005,In_1869);
or U2439 (N_2439,In_370,In_676);
nor U2440 (N_2440,In_2050,In_2663);
xor U2441 (N_2441,In_191,In_2967);
or U2442 (N_2442,In_1277,In_2004);
xnor U2443 (N_2443,In_382,In_1858);
xnor U2444 (N_2444,In_2654,In_1401);
or U2445 (N_2445,In_570,In_229);
nand U2446 (N_2446,In_2892,In_2539);
or U2447 (N_2447,In_1103,In_2560);
and U2448 (N_2448,In_603,In_2830);
or U2449 (N_2449,In_864,In_1811);
xor U2450 (N_2450,In_1000,In_2763);
or U2451 (N_2451,In_1354,In_734);
and U2452 (N_2452,In_2250,In_894);
nor U2453 (N_2453,In_1679,In_129);
nor U2454 (N_2454,In_2940,In_627);
nand U2455 (N_2455,In_1846,In_2360);
nand U2456 (N_2456,In_1384,In_126);
nand U2457 (N_2457,In_928,In_825);
nor U2458 (N_2458,In_2351,In_1100);
and U2459 (N_2459,In_2275,In_2770);
and U2460 (N_2460,In_2518,In_65);
nand U2461 (N_2461,In_2652,In_1563);
nor U2462 (N_2462,In_1488,In_151);
xnor U2463 (N_2463,In_2413,In_653);
or U2464 (N_2464,In_1901,In_2098);
or U2465 (N_2465,In_357,In_1493);
or U2466 (N_2466,In_85,In_756);
xnor U2467 (N_2467,In_125,In_2779);
nor U2468 (N_2468,In_1681,In_2765);
or U2469 (N_2469,In_2837,In_268);
xor U2470 (N_2470,In_2619,In_1429);
nand U2471 (N_2471,In_1028,In_2060);
or U2472 (N_2472,In_1562,In_229);
and U2473 (N_2473,In_467,In_623);
nor U2474 (N_2474,In_312,In_2728);
or U2475 (N_2475,In_2614,In_2229);
nand U2476 (N_2476,In_2917,In_1213);
xnor U2477 (N_2477,In_2983,In_2045);
nand U2478 (N_2478,In_920,In_2890);
nor U2479 (N_2479,In_2078,In_2103);
nor U2480 (N_2480,In_290,In_2827);
nor U2481 (N_2481,In_2345,In_374);
xnor U2482 (N_2482,In_680,In_974);
xnor U2483 (N_2483,In_1018,In_2524);
or U2484 (N_2484,In_177,In_2428);
nand U2485 (N_2485,In_1694,In_845);
nand U2486 (N_2486,In_2847,In_1394);
xor U2487 (N_2487,In_2151,In_859);
nor U2488 (N_2488,In_485,In_1854);
nor U2489 (N_2489,In_100,In_955);
nand U2490 (N_2490,In_613,In_2796);
and U2491 (N_2491,In_2154,In_996);
nor U2492 (N_2492,In_2145,In_2086);
and U2493 (N_2493,In_1803,In_2224);
nand U2494 (N_2494,In_191,In_262);
nand U2495 (N_2495,In_567,In_2973);
xor U2496 (N_2496,In_2676,In_867);
nor U2497 (N_2497,In_341,In_1324);
nand U2498 (N_2498,In_368,In_2317);
nand U2499 (N_2499,In_968,In_379);
or U2500 (N_2500,In_1307,In_1970);
nor U2501 (N_2501,In_1682,In_2290);
and U2502 (N_2502,In_2819,In_860);
nand U2503 (N_2503,In_1733,In_772);
nor U2504 (N_2504,In_1231,In_281);
xnor U2505 (N_2505,In_138,In_517);
xor U2506 (N_2506,In_1808,In_637);
xor U2507 (N_2507,In_2848,In_1276);
nand U2508 (N_2508,In_1065,In_179);
and U2509 (N_2509,In_638,In_2331);
xnor U2510 (N_2510,In_2928,In_811);
nand U2511 (N_2511,In_163,In_1644);
and U2512 (N_2512,In_2957,In_1355);
nand U2513 (N_2513,In_2902,In_681);
nand U2514 (N_2514,In_1318,In_2703);
or U2515 (N_2515,In_525,In_439);
and U2516 (N_2516,In_2894,In_2173);
nor U2517 (N_2517,In_256,In_2488);
nand U2518 (N_2518,In_259,In_2063);
nand U2519 (N_2519,In_1654,In_747);
and U2520 (N_2520,In_488,In_1134);
nand U2521 (N_2521,In_1234,In_2424);
nor U2522 (N_2522,In_2144,In_2666);
and U2523 (N_2523,In_764,In_1657);
nor U2524 (N_2524,In_42,In_1454);
nand U2525 (N_2525,In_2610,In_2638);
or U2526 (N_2526,In_1969,In_1111);
or U2527 (N_2527,In_2936,In_1870);
and U2528 (N_2528,In_2467,In_2319);
xnor U2529 (N_2529,In_1561,In_1142);
and U2530 (N_2530,In_1094,In_761);
nor U2531 (N_2531,In_604,In_571);
nand U2532 (N_2532,In_1291,In_612);
and U2533 (N_2533,In_2712,In_527);
or U2534 (N_2534,In_486,In_689);
nand U2535 (N_2535,In_1051,In_117);
and U2536 (N_2536,In_799,In_1071);
nor U2537 (N_2537,In_170,In_2015);
and U2538 (N_2538,In_372,In_1590);
nand U2539 (N_2539,In_631,In_601);
nand U2540 (N_2540,In_2958,In_1989);
nor U2541 (N_2541,In_1530,In_2586);
nor U2542 (N_2542,In_727,In_1814);
or U2543 (N_2543,In_678,In_1039);
and U2544 (N_2544,In_2628,In_2675);
or U2545 (N_2545,In_2372,In_2423);
nand U2546 (N_2546,In_2071,In_2839);
nand U2547 (N_2547,In_94,In_2602);
nand U2548 (N_2548,In_41,In_2336);
nor U2549 (N_2549,In_2556,In_918);
and U2550 (N_2550,In_751,In_1469);
or U2551 (N_2551,In_2177,In_2539);
nand U2552 (N_2552,In_1577,In_1572);
and U2553 (N_2553,In_135,In_258);
nor U2554 (N_2554,In_2796,In_1492);
or U2555 (N_2555,In_2152,In_2398);
nand U2556 (N_2556,In_404,In_2940);
xnor U2557 (N_2557,In_63,In_2744);
nor U2558 (N_2558,In_1029,In_695);
nor U2559 (N_2559,In_2005,In_2119);
nand U2560 (N_2560,In_2402,In_396);
or U2561 (N_2561,In_2808,In_300);
xor U2562 (N_2562,In_928,In_10);
and U2563 (N_2563,In_2011,In_2770);
xor U2564 (N_2564,In_1939,In_2267);
xor U2565 (N_2565,In_2124,In_2940);
or U2566 (N_2566,In_341,In_257);
or U2567 (N_2567,In_1776,In_2469);
and U2568 (N_2568,In_1945,In_2257);
nor U2569 (N_2569,In_2966,In_734);
xnor U2570 (N_2570,In_2966,In_446);
or U2571 (N_2571,In_2538,In_1563);
xor U2572 (N_2572,In_2879,In_2902);
nand U2573 (N_2573,In_1753,In_1551);
xor U2574 (N_2574,In_2530,In_2498);
or U2575 (N_2575,In_2077,In_2336);
nor U2576 (N_2576,In_552,In_759);
or U2577 (N_2577,In_2863,In_2034);
and U2578 (N_2578,In_2080,In_1522);
and U2579 (N_2579,In_1100,In_2208);
and U2580 (N_2580,In_785,In_1012);
xnor U2581 (N_2581,In_2457,In_682);
xnor U2582 (N_2582,In_1547,In_539);
or U2583 (N_2583,In_1675,In_31);
nor U2584 (N_2584,In_1478,In_706);
and U2585 (N_2585,In_1119,In_2208);
and U2586 (N_2586,In_2599,In_754);
or U2587 (N_2587,In_2446,In_761);
nor U2588 (N_2588,In_642,In_1132);
or U2589 (N_2589,In_1376,In_607);
nor U2590 (N_2590,In_2254,In_1186);
xor U2591 (N_2591,In_2791,In_1003);
nand U2592 (N_2592,In_1868,In_1259);
xor U2593 (N_2593,In_445,In_2692);
and U2594 (N_2594,In_13,In_1666);
nor U2595 (N_2595,In_2578,In_2162);
or U2596 (N_2596,In_67,In_1579);
or U2597 (N_2597,In_2657,In_1427);
nor U2598 (N_2598,In_2317,In_2231);
or U2599 (N_2599,In_404,In_1223);
xnor U2600 (N_2600,In_1100,In_2307);
and U2601 (N_2601,In_1566,In_2261);
nor U2602 (N_2602,In_2905,In_2645);
and U2603 (N_2603,In_2080,In_601);
and U2604 (N_2604,In_2305,In_125);
xnor U2605 (N_2605,In_278,In_1903);
and U2606 (N_2606,In_2606,In_2831);
xor U2607 (N_2607,In_154,In_0);
nand U2608 (N_2608,In_1067,In_1685);
nor U2609 (N_2609,In_2151,In_660);
or U2610 (N_2610,In_542,In_2115);
nand U2611 (N_2611,In_2062,In_849);
nor U2612 (N_2612,In_2213,In_35);
and U2613 (N_2613,In_2941,In_2814);
nor U2614 (N_2614,In_179,In_2843);
and U2615 (N_2615,In_1297,In_1);
nand U2616 (N_2616,In_1654,In_1987);
and U2617 (N_2617,In_136,In_1371);
nor U2618 (N_2618,In_2188,In_705);
nor U2619 (N_2619,In_1519,In_2138);
and U2620 (N_2620,In_198,In_1898);
and U2621 (N_2621,In_2773,In_1645);
xnor U2622 (N_2622,In_404,In_787);
and U2623 (N_2623,In_1721,In_1822);
and U2624 (N_2624,In_1928,In_1470);
nand U2625 (N_2625,In_2557,In_1518);
xor U2626 (N_2626,In_1214,In_137);
nand U2627 (N_2627,In_2185,In_553);
xnor U2628 (N_2628,In_810,In_189);
nor U2629 (N_2629,In_2239,In_526);
nor U2630 (N_2630,In_1113,In_2989);
or U2631 (N_2631,In_1536,In_641);
nand U2632 (N_2632,In_828,In_100);
nor U2633 (N_2633,In_2480,In_1598);
nor U2634 (N_2634,In_1198,In_1289);
or U2635 (N_2635,In_2950,In_1737);
nor U2636 (N_2636,In_1957,In_2957);
nor U2637 (N_2637,In_1348,In_434);
xor U2638 (N_2638,In_1683,In_2166);
or U2639 (N_2639,In_1599,In_1001);
nand U2640 (N_2640,In_2465,In_1939);
nand U2641 (N_2641,In_1755,In_709);
and U2642 (N_2642,In_1247,In_317);
and U2643 (N_2643,In_306,In_2013);
or U2644 (N_2644,In_1464,In_2965);
nand U2645 (N_2645,In_2699,In_549);
and U2646 (N_2646,In_1516,In_418);
nand U2647 (N_2647,In_2732,In_1160);
nand U2648 (N_2648,In_1833,In_2329);
or U2649 (N_2649,In_2289,In_1491);
xor U2650 (N_2650,In_257,In_760);
xnor U2651 (N_2651,In_190,In_703);
xor U2652 (N_2652,In_818,In_2492);
and U2653 (N_2653,In_1685,In_476);
nor U2654 (N_2654,In_2061,In_539);
xnor U2655 (N_2655,In_2071,In_182);
xor U2656 (N_2656,In_569,In_800);
xor U2657 (N_2657,In_1229,In_2293);
nand U2658 (N_2658,In_1202,In_2436);
and U2659 (N_2659,In_105,In_2348);
nor U2660 (N_2660,In_2913,In_1856);
xor U2661 (N_2661,In_1431,In_1561);
nand U2662 (N_2662,In_916,In_639);
nor U2663 (N_2663,In_2299,In_115);
nand U2664 (N_2664,In_597,In_2933);
nand U2665 (N_2665,In_2444,In_829);
nand U2666 (N_2666,In_2464,In_2681);
xnor U2667 (N_2667,In_1509,In_1870);
nor U2668 (N_2668,In_2544,In_318);
xnor U2669 (N_2669,In_1999,In_1567);
nor U2670 (N_2670,In_1473,In_2925);
nand U2671 (N_2671,In_1987,In_796);
or U2672 (N_2672,In_1981,In_1786);
nand U2673 (N_2673,In_2355,In_673);
xnor U2674 (N_2674,In_1497,In_867);
nor U2675 (N_2675,In_484,In_2291);
or U2676 (N_2676,In_1679,In_2945);
nor U2677 (N_2677,In_2897,In_899);
or U2678 (N_2678,In_191,In_593);
xnor U2679 (N_2679,In_737,In_1432);
or U2680 (N_2680,In_525,In_108);
nor U2681 (N_2681,In_2980,In_645);
or U2682 (N_2682,In_2320,In_2099);
nand U2683 (N_2683,In_132,In_2889);
or U2684 (N_2684,In_218,In_1145);
or U2685 (N_2685,In_2809,In_2882);
or U2686 (N_2686,In_568,In_597);
nand U2687 (N_2687,In_374,In_447);
nor U2688 (N_2688,In_2230,In_441);
xnor U2689 (N_2689,In_1638,In_1052);
nor U2690 (N_2690,In_2256,In_278);
nand U2691 (N_2691,In_451,In_2909);
nor U2692 (N_2692,In_611,In_2200);
nor U2693 (N_2693,In_989,In_659);
or U2694 (N_2694,In_2398,In_571);
and U2695 (N_2695,In_2502,In_1301);
or U2696 (N_2696,In_1152,In_2453);
nand U2697 (N_2697,In_371,In_444);
nand U2698 (N_2698,In_178,In_253);
nor U2699 (N_2699,In_1256,In_645);
nor U2700 (N_2700,In_177,In_1300);
or U2701 (N_2701,In_2295,In_2167);
or U2702 (N_2702,In_2023,In_885);
nand U2703 (N_2703,In_1443,In_2308);
and U2704 (N_2704,In_2756,In_2342);
xor U2705 (N_2705,In_2404,In_2139);
or U2706 (N_2706,In_2031,In_2986);
nand U2707 (N_2707,In_713,In_2801);
or U2708 (N_2708,In_1365,In_273);
nor U2709 (N_2709,In_2299,In_131);
or U2710 (N_2710,In_1244,In_272);
or U2711 (N_2711,In_1870,In_1154);
and U2712 (N_2712,In_1899,In_161);
xnor U2713 (N_2713,In_2406,In_998);
or U2714 (N_2714,In_293,In_2527);
xor U2715 (N_2715,In_805,In_1890);
or U2716 (N_2716,In_671,In_2626);
nand U2717 (N_2717,In_2520,In_1839);
xnor U2718 (N_2718,In_1325,In_2585);
xnor U2719 (N_2719,In_1728,In_857);
and U2720 (N_2720,In_547,In_2806);
nor U2721 (N_2721,In_754,In_114);
or U2722 (N_2722,In_1929,In_653);
and U2723 (N_2723,In_2982,In_181);
xnor U2724 (N_2724,In_1893,In_1931);
xnor U2725 (N_2725,In_2360,In_1334);
nand U2726 (N_2726,In_665,In_302);
or U2727 (N_2727,In_1060,In_1945);
or U2728 (N_2728,In_743,In_2572);
nand U2729 (N_2729,In_424,In_574);
nor U2730 (N_2730,In_648,In_460);
or U2731 (N_2731,In_1773,In_139);
and U2732 (N_2732,In_515,In_2571);
xor U2733 (N_2733,In_2571,In_1852);
or U2734 (N_2734,In_2109,In_673);
and U2735 (N_2735,In_1828,In_319);
xnor U2736 (N_2736,In_127,In_1830);
nand U2737 (N_2737,In_707,In_2309);
xor U2738 (N_2738,In_824,In_287);
nand U2739 (N_2739,In_859,In_2203);
nand U2740 (N_2740,In_74,In_2387);
nor U2741 (N_2741,In_89,In_240);
and U2742 (N_2742,In_1425,In_1489);
nor U2743 (N_2743,In_59,In_1156);
or U2744 (N_2744,In_369,In_48);
nand U2745 (N_2745,In_2702,In_603);
and U2746 (N_2746,In_2457,In_2375);
xnor U2747 (N_2747,In_2425,In_1489);
nand U2748 (N_2748,In_2533,In_1427);
or U2749 (N_2749,In_1026,In_2806);
nor U2750 (N_2750,In_97,In_2631);
or U2751 (N_2751,In_2411,In_1099);
nand U2752 (N_2752,In_2852,In_996);
nor U2753 (N_2753,In_2413,In_647);
nand U2754 (N_2754,In_780,In_1978);
and U2755 (N_2755,In_25,In_2116);
and U2756 (N_2756,In_2623,In_1632);
and U2757 (N_2757,In_2550,In_2804);
and U2758 (N_2758,In_1990,In_891);
or U2759 (N_2759,In_909,In_2799);
or U2760 (N_2760,In_2758,In_2008);
nor U2761 (N_2761,In_2755,In_2099);
xor U2762 (N_2762,In_2271,In_2285);
nor U2763 (N_2763,In_20,In_1863);
nor U2764 (N_2764,In_2843,In_1172);
and U2765 (N_2765,In_39,In_1061);
xnor U2766 (N_2766,In_2139,In_2856);
nor U2767 (N_2767,In_1842,In_1088);
or U2768 (N_2768,In_2643,In_327);
xnor U2769 (N_2769,In_1060,In_1082);
and U2770 (N_2770,In_190,In_2512);
xor U2771 (N_2771,In_1531,In_2323);
xor U2772 (N_2772,In_2159,In_424);
and U2773 (N_2773,In_554,In_1619);
and U2774 (N_2774,In_508,In_1334);
nor U2775 (N_2775,In_1902,In_1940);
nor U2776 (N_2776,In_2722,In_1931);
xnor U2777 (N_2777,In_2506,In_2117);
and U2778 (N_2778,In_2117,In_1467);
nand U2779 (N_2779,In_1584,In_1144);
or U2780 (N_2780,In_2348,In_2874);
xnor U2781 (N_2781,In_483,In_2378);
xnor U2782 (N_2782,In_1322,In_2595);
xnor U2783 (N_2783,In_1123,In_2074);
nand U2784 (N_2784,In_2096,In_1293);
or U2785 (N_2785,In_1762,In_1123);
xnor U2786 (N_2786,In_2515,In_1061);
and U2787 (N_2787,In_2920,In_265);
and U2788 (N_2788,In_1346,In_2386);
nand U2789 (N_2789,In_1207,In_2079);
xnor U2790 (N_2790,In_1497,In_5);
nor U2791 (N_2791,In_1758,In_2339);
and U2792 (N_2792,In_638,In_427);
xnor U2793 (N_2793,In_2800,In_1605);
nor U2794 (N_2794,In_426,In_590);
and U2795 (N_2795,In_2082,In_275);
or U2796 (N_2796,In_775,In_1069);
nand U2797 (N_2797,In_250,In_2033);
xor U2798 (N_2798,In_704,In_2719);
nor U2799 (N_2799,In_1459,In_1707);
nand U2800 (N_2800,In_1266,In_2696);
nor U2801 (N_2801,In_338,In_417);
nand U2802 (N_2802,In_2315,In_1768);
nand U2803 (N_2803,In_2336,In_1819);
nand U2804 (N_2804,In_2033,In_1729);
xor U2805 (N_2805,In_2813,In_722);
nor U2806 (N_2806,In_1561,In_1992);
xor U2807 (N_2807,In_1036,In_1360);
nor U2808 (N_2808,In_1067,In_1676);
or U2809 (N_2809,In_313,In_2718);
and U2810 (N_2810,In_764,In_148);
or U2811 (N_2811,In_806,In_792);
xor U2812 (N_2812,In_2100,In_2212);
nor U2813 (N_2813,In_1370,In_590);
xor U2814 (N_2814,In_1795,In_1358);
and U2815 (N_2815,In_2330,In_688);
nand U2816 (N_2816,In_2806,In_1605);
and U2817 (N_2817,In_585,In_574);
and U2818 (N_2818,In_2659,In_1338);
and U2819 (N_2819,In_1325,In_1395);
or U2820 (N_2820,In_2828,In_1651);
and U2821 (N_2821,In_2165,In_1119);
and U2822 (N_2822,In_116,In_859);
nand U2823 (N_2823,In_839,In_1964);
xor U2824 (N_2824,In_413,In_2550);
xnor U2825 (N_2825,In_1501,In_886);
and U2826 (N_2826,In_698,In_1238);
or U2827 (N_2827,In_2202,In_954);
xnor U2828 (N_2828,In_1257,In_1009);
nor U2829 (N_2829,In_2107,In_2704);
nand U2830 (N_2830,In_490,In_878);
nor U2831 (N_2831,In_1360,In_2306);
nand U2832 (N_2832,In_596,In_68);
or U2833 (N_2833,In_1953,In_2087);
or U2834 (N_2834,In_960,In_357);
nand U2835 (N_2835,In_1029,In_1248);
xor U2836 (N_2836,In_68,In_630);
or U2837 (N_2837,In_13,In_1736);
nor U2838 (N_2838,In_2242,In_2560);
nand U2839 (N_2839,In_635,In_579);
and U2840 (N_2840,In_2340,In_605);
nand U2841 (N_2841,In_110,In_2398);
and U2842 (N_2842,In_1239,In_1545);
nor U2843 (N_2843,In_2910,In_2345);
nor U2844 (N_2844,In_25,In_1723);
nor U2845 (N_2845,In_2020,In_98);
nor U2846 (N_2846,In_473,In_146);
nor U2847 (N_2847,In_583,In_997);
nand U2848 (N_2848,In_423,In_1883);
nand U2849 (N_2849,In_1993,In_2918);
or U2850 (N_2850,In_395,In_1330);
or U2851 (N_2851,In_2641,In_2772);
and U2852 (N_2852,In_1395,In_1671);
xor U2853 (N_2853,In_805,In_609);
nor U2854 (N_2854,In_1043,In_757);
nor U2855 (N_2855,In_2124,In_284);
or U2856 (N_2856,In_1925,In_2140);
and U2857 (N_2857,In_566,In_1397);
or U2858 (N_2858,In_1056,In_981);
xor U2859 (N_2859,In_2345,In_2477);
nand U2860 (N_2860,In_49,In_2023);
or U2861 (N_2861,In_487,In_2279);
or U2862 (N_2862,In_920,In_1338);
xnor U2863 (N_2863,In_1503,In_2865);
xnor U2864 (N_2864,In_1484,In_2084);
nor U2865 (N_2865,In_1679,In_131);
nand U2866 (N_2866,In_986,In_1952);
nand U2867 (N_2867,In_2780,In_2446);
nor U2868 (N_2868,In_2091,In_2395);
xor U2869 (N_2869,In_378,In_2826);
nor U2870 (N_2870,In_2699,In_2824);
xnor U2871 (N_2871,In_384,In_2188);
nand U2872 (N_2872,In_2585,In_1409);
and U2873 (N_2873,In_998,In_1327);
or U2874 (N_2874,In_1694,In_2184);
or U2875 (N_2875,In_1567,In_333);
or U2876 (N_2876,In_477,In_1274);
nand U2877 (N_2877,In_2146,In_1733);
xor U2878 (N_2878,In_906,In_274);
xor U2879 (N_2879,In_800,In_2826);
nand U2880 (N_2880,In_2759,In_1171);
nor U2881 (N_2881,In_1943,In_1221);
xnor U2882 (N_2882,In_1897,In_2843);
xnor U2883 (N_2883,In_2027,In_892);
xnor U2884 (N_2884,In_1520,In_367);
nand U2885 (N_2885,In_2370,In_1965);
nor U2886 (N_2886,In_108,In_357);
xor U2887 (N_2887,In_2782,In_1211);
nand U2888 (N_2888,In_2592,In_2143);
nor U2889 (N_2889,In_1544,In_2142);
and U2890 (N_2890,In_983,In_491);
nor U2891 (N_2891,In_19,In_787);
and U2892 (N_2892,In_2221,In_1652);
or U2893 (N_2893,In_2658,In_2888);
nor U2894 (N_2894,In_2037,In_551);
or U2895 (N_2895,In_631,In_1410);
nand U2896 (N_2896,In_403,In_2395);
and U2897 (N_2897,In_528,In_2637);
nand U2898 (N_2898,In_1967,In_1002);
nor U2899 (N_2899,In_2624,In_174);
nor U2900 (N_2900,In_2258,In_2340);
nand U2901 (N_2901,In_1812,In_1291);
or U2902 (N_2902,In_304,In_1605);
and U2903 (N_2903,In_2083,In_2233);
and U2904 (N_2904,In_2500,In_1024);
xor U2905 (N_2905,In_1639,In_1106);
xor U2906 (N_2906,In_1077,In_440);
and U2907 (N_2907,In_2455,In_1525);
nor U2908 (N_2908,In_1702,In_1897);
nand U2909 (N_2909,In_2602,In_717);
and U2910 (N_2910,In_362,In_1438);
nand U2911 (N_2911,In_1136,In_154);
nand U2912 (N_2912,In_32,In_2423);
or U2913 (N_2913,In_2813,In_1025);
nor U2914 (N_2914,In_2131,In_768);
or U2915 (N_2915,In_1393,In_1169);
and U2916 (N_2916,In_2004,In_2478);
nand U2917 (N_2917,In_176,In_4);
or U2918 (N_2918,In_819,In_1474);
xor U2919 (N_2919,In_1115,In_9);
or U2920 (N_2920,In_9,In_1419);
nand U2921 (N_2921,In_298,In_2166);
and U2922 (N_2922,In_416,In_1603);
nand U2923 (N_2923,In_1046,In_2437);
xnor U2924 (N_2924,In_429,In_1902);
nor U2925 (N_2925,In_343,In_434);
and U2926 (N_2926,In_1721,In_1616);
and U2927 (N_2927,In_86,In_1105);
nor U2928 (N_2928,In_1042,In_1337);
nand U2929 (N_2929,In_324,In_226);
or U2930 (N_2930,In_2672,In_270);
nand U2931 (N_2931,In_1350,In_2142);
nor U2932 (N_2932,In_756,In_1661);
or U2933 (N_2933,In_865,In_2907);
xnor U2934 (N_2934,In_1014,In_1128);
nor U2935 (N_2935,In_2287,In_1427);
and U2936 (N_2936,In_10,In_484);
or U2937 (N_2937,In_1778,In_113);
nand U2938 (N_2938,In_2239,In_2678);
nor U2939 (N_2939,In_1305,In_2624);
or U2940 (N_2940,In_707,In_2220);
nor U2941 (N_2941,In_264,In_2659);
nor U2942 (N_2942,In_2854,In_830);
or U2943 (N_2943,In_1469,In_242);
or U2944 (N_2944,In_1394,In_338);
xor U2945 (N_2945,In_1324,In_2267);
xnor U2946 (N_2946,In_958,In_185);
nor U2947 (N_2947,In_324,In_937);
nand U2948 (N_2948,In_1123,In_2865);
nor U2949 (N_2949,In_1018,In_433);
xnor U2950 (N_2950,In_956,In_131);
nor U2951 (N_2951,In_107,In_407);
or U2952 (N_2952,In_2154,In_1236);
xor U2953 (N_2953,In_1679,In_1190);
and U2954 (N_2954,In_2466,In_2321);
nand U2955 (N_2955,In_334,In_2222);
xnor U2956 (N_2956,In_215,In_1037);
xnor U2957 (N_2957,In_2438,In_1888);
xor U2958 (N_2958,In_2931,In_675);
or U2959 (N_2959,In_1563,In_362);
xnor U2960 (N_2960,In_2689,In_2586);
nand U2961 (N_2961,In_1138,In_2052);
xor U2962 (N_2962,In_631,In_2689);
xor U2963 (N_2963,In_1448,In_2509);
and U2964 (N_2964,In_2737,In_154);
xor U2965 (N_2965,In_2912,In_695);
xnor U2966 (N_2966,In_1887,In_2523);
nand U2967 (N_2967,In_1538,In_1324);
xnor U2968 (N_2968,In_2236,In_1055);
xnor U2969 (N_2969,In_2430,In_410);
nand U2970 (N_2970,In_955,In_2029);
xor U2971 (N_2971,In_6,In_1568);
xor U2972 (N_2972,In_850,In_1108);
nand U2973 (N_2973,In_733,In_2716);
and U2974 (N_2974,In_2414,In_226);
nand U2975 (N_2975,In_222,In_1762);
and U2976 (N_2976,In_433,In_2727);
and U2977 (N_2977,In_1967,In_1677);
nor U2978 (N_2978,In_94,In_2756);
and U2979 (N_2979,In_2341,In_1195);
xor U2980 (N_2980,In_1891,In_87);
nand U2981 (N_2981,In_1743,In_2109);
and U2982 (N_2982,In_1531,In_938);
and U2983 (N_2983,In_1364,In_2989);
nor U2984 (N_2984,In_2348,In_948);
nor U2985 (N_2985,In_2423,In_2815);
and U2986 (N_2986,In_965,In_2008);
or U2987 (N_2987,In_747,In_1974);
nand U2988 (N_2988,In_2429,In_1274);
and U2989 (N_2989,In_2873,In_2283);
and U2990 (N_2990,In_605,In_230);
nand U2991 (N_2991,In_2889,In_886);
or U2992 (N_2992,In_1572,In_1031);
nor U2993 (N_2993,In_1186,In_2662);
xor U2994 (N_2994,In_2344,In_2184);
nor U2995 (N_2995,In_1713,In_1467);
or U2996 (N_2996,In_869,In_2679);
nor U2997 (N_2997,In_1922,In_152);
xnor U2998 (N_2998,In_2817,In_1398);
nand U2999 (N_2999,In_1487,In_1821);
or U3000 (N_3000,N_899,N_2983);
and U3001 (N_3001,N_1344,N_1670);
or U3002 (N_3002,N_2768,N_1739);
and U3003 (N_3003,N_2247,N_2510);
and U3004 (N_3004,N_865,N_770);
xor U3005 (N_3005,N_36,N_2897);
and U3006 (N_3006,N_499,N_11);
nor U3007 (N_3007,N_2918,N_1800);
nand U3008 (N_3008,N_771,N_2109);
nand U3009 (N_3009,N_1780,N_278);
xnor U3010 (N_3010,N_1668,N_1267);
nor U3011 (N_3011,N_1880,N_617);
nand U3012 (N_3012,N_1281,N_2513);
or U3013 (N_3013,N_716,N_574);
and U3014 (N_3014,N_1261,N_41);
or U3015 (N_3015,N_1425,N_2865);
nor U3016 (N_3016,N_2051,N_1889);
and U3017 (N_3017,N_1637,N_641);
and U3018 (N_3018,N_501,N_539);
and U3019 (N_3019,N_2959,N_1881);
nand U3020 (N_3020,N_712,N_90);
and U3021 (N_3021,N_2192,N_0);
xnor U3022 (N_3022,N_75,N_2532);
xnor U3023 (N_3023,N_2709,N_2364);
nor U3024 (N_3024,N_2038,N_1480);
nand U3025 (N_3025,N_276,N_2435);
xnor U3026 (N_3026,N_2818,N_2246);
nand U3027 (N_3027,N_2309,N_1536);
nor U3028 (N_3028,N_814,N_2869);
nand U3029 (N_3029,N_165,N_257);
or U3030 (N_3030,N_2490,N_575);
xor U3031 (N_3031,N_599,N_1353);
nand U3032 (N_3032,N_2328,N_1601);
and U3033 (N_3033,N_2224,N_1252);
xnor U3034 (N_3034,N_2162,N_2636);
nand U3035 (N_3035,N_198,N_2941);
nand U3036 (N_3036,N_2703,N_1154);
nand U3037 (N_3037,N_2987,N_1181);
nand U3038 (N_3038,N_1345,N_903);
and U3039 (N_3039,N_1285,N_1634);
nand U3040 (N_3040,N_923,N_654);
nand U3041 (N_3041,N_793,N_2524);
nor U3042 (N_3042,N_1234,N_2862);
or U3043 (N_3043,N_170,N_2137);
or U3044 (N_3044,N_1373,N_1944);
nor U3045 (N_3045,N_996,N_2681);
nor U3046 (N_3046,N_2445,N_767);
xor U3047 (N_3047,N_2846,N_310);
nor U3048 (N_3048,N_16,N_2819);
or U3049 (N_3049,N_91,N_201);
nand U3050 (N_3050,N_1291,N_457);
and U3051 (N_3051,N_2702,N_2405);
xor U3052 (N_3052,N_2997,N_933);
or U3053 (N_3053,N_2775,N_1703);
nand U3054 (N_3054,N_826,N_1374);
nand U3055 (N_3055,N_623,N_727);
and U3056 (N_3056,N_1268,N_1014);
or U3057 (N_3057,N_1764,N_2280);
nand U3058 (N_3058,N_1066,N_629);
nor U3059 (N_3059,N_279,N_281);
nor U3060 (N_3060,N_2883,N_943);
or U3061 (N_3061,N_1886,N_1928);
nor U3062 (N_3062,N_2090,N_34);
xnor U3063 (N_3063,N_1304,N_156);
xnor U3064 (N_3064,N_1969,N_2423);
xor U3065 (N_3065,N_350,N_2848);
and U3066 (N_3066,N_572,N_636);
or U3067 (N_3067,N_2826,N_1189);
or U3068 (N_3068,N_1349,N_2145);
xnor U3069 (N_3069,N_2854,N_2578);
xor U3070 (N_3070,N_1576,N_344);
or U3071 (N_3071,N_2606,N_1130);
and U3072 (N_3072,N_509,N_1009);
xor U3073 (N_3073,N_2528,N_59);
nand U3074 (N_3074,N_2780,N_642);
or U3075 (N_3075,N_2029,N_2529);
nand U3076 (N_3076,N_761,N_2124);
or U3077 (N_3077,N_2482,N_2426);
or U3078 (N_3078,N_2892,N_2620);
nand U3079 (N_3079,N_1057,N_1724);
xor U3080 (N_3080,N_495,N_591);
and U3081 (N_3081,N_567,N_2171);
or U3082 (N_3082,N_2676,N_860);
or U3083 (N_3083,N_1606,N_1947);
and U3084 (N_3084,N_569,N_2824);
and U3085 (N_3085,N_364,N_358);
nand U3086 (N_3086,N_1020,N_2303);
or U3087 (N_3087,N_1572,N_1114);
nor U3088 (N_3088,N_2725,N_604);
and U3089 (N_3089,N_951,N_1006);
xor U3090 (N_3090,N_2632,N_2188);
xnor U3091 (N_3091,N_1805,N_1191);
xor U3092 (N_3092,N_1967,N_2878);
xor U3093 (N_3093,N_1337,N_737);
and U3094 (N_3094,N_573,N_2555);
nand U3095 (N_3095,N_2948,N_404);
and U3096 (N_3096,N_2706,N_1423);
nor U3097 (N_3097,N_1554,N_2164);
and U3098 (N_3098,N_435,N_1610);
xnor U3099 (N_3099,N_587,N_1221);
or U3100 (N_3100,N_498,N_1769);
and U3101 (N_3101,N_63,N_1763);
and U3102 (N_3102,N_1567,N_2004);
nand U3103 (N_3103,N_2996,N_2602);
xor U3104 (N_3104,N_2293,N_1115);
or U3105 (N_3105,N_1549,N_2605);
nor U3106 (N_3106,N_1597,N_297);
nor U3107 (N_3107,N_2789,N_928);
nand U3108 (N_3108,N_1021,N_597);
xor U3109 (N_3109,N_126,N_2402);
nand U3110 (N_3110,N_2122,N_2469);
and U3111 (N_3111,N_1419,N_2412);
nor U3112 (N_3112,N_1022,N_1338);
nand U3113 (N_3113,N_1795,N_2177);
xnor U3114 (N_3114,N_1359,N_52);
nor U3115 (N_3115,N_603,N_242);
and U3116 (N_3116,N_2209,N_18);
xor U3117 (N_3117,N_355,N_1785);
and U3118 (N_3118,N_1163,N_2242);
nor U3119 (N_3119,N_1137,N_902);
or U3120 (N_3120,N_1834,N_2593);
or U3121 (N_3121,N_1542,N_2563);
xor U3122 (N_3122,N_941,N_1086);
nand U3123 (N_3123,N_356,N_2048);
nand U3124 (N_3124,N_2163,N_1919);
or U3125 (N_3125,N_2581,N_1938);
xnor U3126 (N_3126,N_584,N_638);
nand U3127 (N_3127,N_890,N_1034);
or U3128 (N_3128,N_1393,N_2332);
nand U3129 (N_3129,N_78,N_2363);
nor U3130 (N_3130,N_871,N_901);
nand U3131 (N_3131,N_1529,N_129);
or U3132 (N_3132,N_49,N_2075);
nand U3133 (N_3133,N_967,N_1129);
nor U3134 (N_3134,N_1557,N_1629);
nand U3135 (N_3135,N_2037,N_226);
xnor U3136 (N_3136,N_511,N_1272);
nor U3137 (N_3137,N_222,N_1987);
or U3138 (N_3138,N_548,N_1213);
and U3139 (N_3139,N_2118,N_493);
nand U3140 (N_3140,N_740,N_1516);
or U3141 (N_3141,N_2849,N_2320);
nand U3142 (N_3142,N_1408,N_747);
xor U3143 (N_3143,N_1256,N_1485);
or U3144 (N_3144,N_2433,N_492);
xor U3145 (N_3145,N_1429,N_1642);
xor U3146 (N_3146,N_408,N_1173);
nor U3147 (N_3147,N_341,N_1717);
or U3148 (N_3148,N_866,N_606);
nor U3149 (N_3149,N_2723,N_239);
or U3150 (N_3150,N_2175,N_2138);
and U3151 (N_3151,N_1943,N_42);
xor U3152 (N_3152,N_2909,N_2352);
and U3153 (N_3153,N_541,N_2413);
nor U3154 (N_3154,N_2274,N_1794);
nand U3155 (N_3155,N_2530,N_2279);
nand U3156 (N_3156,N_2629,N_1211);
and U3157 (N_3157,N_1327,N_2511);
xor U3158 (N_3158,N_1084,N_1094);
or U3159 (N_3159,N_240,N_1410);
nor U3160 (N_3160,N_1607,N_2060);
and U3161 (N_3161,N_888,N_2131);
or U3162 (N_3162,N_2663,N_2253);
xor U3163 (N_3163,N_458,N_986);
and U3164 (N_3164,N_1831,N_2307);
xnor U3165 (N_3165,N_365,N_2512);
or U3166 (N_3166,N_1604,N_2670);
xor U3167 (N_3167,N_2704,N_1566);
nand U3168 (N_3168,N_1658,N_357);
nor U3169 (N_3169,N_713,N_1915);
or U3170 (N_3170,N_982,N_2659);
nor U3171 (N_3171,N_216,N_2647);
and U3172 (N_3172,N_2944,N_1511);
nand U3173 (N_3173,N_73,N_58);
nor U3174 (N_3174,N_1481,N_1736);
or U3175 (N_3175,N_33,N_1656);
or U3176 (N_3176,N_2764,N_2956);
or U3177 (N_3177,N_2098,N_2820);
nor U3178 (N_3178,N_459,N_328);
or U3179 (N_3179,N_1965,N_625);
or U3180 (N_3180,N_455,N_280);
xnor U3181 (N_3181,N_2639,N_2572);
nand U3182 (N_3182,N_1031,N_152);
or U3183 (N_3183,N_436,N_1602);
or U3184 (N_3184,N_554,N_1766);
xor U3185 (N_3185,N_1517,N_403);
and U3186 (N_3186,N_2757,N_1286);
or U3187 (N_3187,N_2313,N_596);
and U3188 (N_3188,N_2440,N_1294);
nor U3189 (N_3189,N_1519,N_1200);
xor U3190 (N_3190,N_2934,N_926);
and U3191 (N_3191,N_1852,N_1323);
and U3192 (N_3192,N_2615,N_2091);
or U3193 (N_3193,N_1666,N_621);
nor U3194 (N_3194,N_908,N_1814);
and U3195 (N_3195,N_86,N_2054);
xnor U3196 (N_3196,N_815,N_1340);
and U3197 (N_3197,N_1412,N_2014);
and U3198 (N_3198,N_1299,N_749);
or U3199 (N_3199,N_1829,N_2119);
or U3200 (N_3200,N_1004,N_513);
xnor U3201 (N_3201,N_1621,N_2917);
xor U3202 (N_3202,N_2399,N_882);
nor U3203 (N_3203,N_1113,N_934);
nand U3204 (N_3204,N_419,N_652);
nor U3205 (N_3205,N_332,N_2586);
nor U3206 (N_3206,N_1231,N_763);
or U3207 (N_3207,N_735,N_766);
and U3208 (N_3208,N_2385,N_2575);
nor U3209 (N_3209,N_825,N_2990);
or U3210 (N_3210,N_685,N_30);
or U3211 (N_3211,N_679,N_1400);
nand U3212 (N_3212,N_204,N_635);
or U3213 (N_3213,N_443,N_743);
xnor U3214 (N_3214,N_393,N_1433);
or U3215 (N_3215,N_1152,N_568);
or U3216 (N_3216,N_2989,N_1280);
nand U3217 (N_3217,N_1526,N_2305);
nor U3218 (N_3218,N_2002,N_2794);
nor U3219 (N_3219,N_1983,N_1251);
or U3220 (N_3220,N_1882,N_2411);
or U3221 (N_3221,N_904,N_644);
or U3222 (N_3222,N_1184,N_389);
and U3223 (N_3223,N_2227,N_2367);
xor U3224 (N_3224,N_1992,N_2803);
nor U3225 (N_3225,N_2805,N_1594);
nor U3226 (N_3226,N_1099,N_1505);
nor U3227 (N_3227,N_2356,N_1375);
and U3228 (N_3228,N_764,N_1316);
and U3229 (N_3229,N_1239,N_1187);
nand U3230 (N_3230,N_1390,N_31);
xnor U3231 (N_3231,N_1096,N_878);
nand U3232 (N_3232,N_169,N_1755);
xnor U3233 (N_3233,N_2932,N_1539);
and U3234 (N_3234,N_2084,N_2646);
and U3235 (N_3235,N_2617,N_148);
or U3236 (N_3236,N_2302,N_690);
xor U3237 (N_3237,N_699,N_842);
nor U3238 (N_3238,N_2028,N_161);
xor U3239 (N_3239,N_705,N_684);
nand U3240 (N_3240,N_667,N_1756);
xnor U3241 (N_3241,N_831,N_1161);
nor U3242 (N_3242,N_1659,N_2321);
nor U3243 (N_3243,N_1204,N_2106);
and U3244 (N_3244,N_2627,N_2732);
xnor U3245 (N_3245,N_2898,N_1867);
xnor U3246 (N_3246,N_2432,N_1333);
nor U3247 (N_3247,N_2314,N_2452);
nor U3248 (N_3248,N_1553,N_2121);
or U3249 (N_3249,N_2195,N_681);
or U3250 (N_3250,N_744,N_836);
nand U3251 (N_3251,N_2677,N_834);
and U3252 (N_3252,N_1781,N_676);
nor U3253 (N_3253,N_974,N_179);
nor U3254 (N_3254,N_1685,N_1104);
nor U3255 (N_3255,N_1224,N_1145);
xor U3256 (N_3256,N_1907,N_77);
xor U3257 (N_3257,N_2097,N_2782);
nor U3258 (N_3258,N_633,N_118);
nor U3259 (N_3259,N_1738,N_627);
nand U3260 (N_3260,N_489,N_486);
and U3261 (N_3261,N_166,N_1071);
or U3262 (N_3262,N_925,N_670);
nor U3263 (N_3263,N_536,N_2977);
nor U3264 (N_3264,N_2596,N_2889);
nand U3265 (N_3265,N_415,N_1625);
nor U3266 (N_3266,N_2810,N_1247);
nor U3267 (N_3267,N_2476,N_756);
xnor U3268 (N_3268,N_2288,N_1108);
nor U3269 (N_3269,N_2792,N_1876);
nand U3270 (N_3270,N_2635,N_1986);
and U3271 (N_3271,N_391,N_829);
nor U3272 (N_3272,N_277,N_323);
or U3273 (N_3273,N_2222,N_519);
and U3274 (N_3274,N_2760,N_106);
and U3275 (N_3275,N_227,N_1591);
xor U3276 (N_3276,N_2380,N_1850);
and U3277 (N_3277,N_2938,N_1449);
nor U3278 (N_3278,N_480,N_1035);
xor U3279 (N_3279,N_2248,N_1277);
xnor U3280 (N_3280,N_1334,N_2179);
or U3281 (N_3281,N_312,N_2955);
xnor U3282 (N_3282,N_2058,N_2755);
xor U3283 (N_3283,N_311,N_2929);
and U3284 (N_3284,N_558,N_1384);
or U3285 (N_3285,N_725,N_2069);
nor U3286 (N_3286,N_2808,N_2778);
and U3287 (N_3287,N_2527,N_72);
and U3288 (N_3288,N_579,N_1697);
xnor U3289 (N_3289,N_1266,N_1227);
nor U3290 (N_3290,N_1993,N_2430);
and U3291 (N_3291,N_423,N_1863);
nand U3292 (N_3292,N_1711,N_2867);
and U3293 (N_3293,N_640,N_1422);
or U3294 (N_3294,N_2652,N_1883);
nor U3295 (N_3295,N_1787,N_726);
and U3296 (N_3296,N_211,N_2674);
and U3297 (N_3297,N_1705,N_1219);
nand U3298 (N_3298,N_1278,N_1720);
and U3299 (N_3299,N_2348,N_1577);
or U3300 (N_3300,N_230,N_1543);
nand U3301 (N_3301,N_1910,N_2715);
xnor U3302 (N_3302,N_653,N_1649);
or U3303 (N_3303,N_1547,N_2404);
or U3304 (N_3304,N_691,N_2263);
or U3305 (N_3305,N_1328,N_250);
nand U3306 (N_3306,N_1903,N_997);
or U3307 (N_3307,N_409,N_208);
and U3308 (N_3308,N_1148,N_2984);
or U3309 (N_3309,N_1873,N_2945);
xor U3310 (N_3310,N_1744,N_1560);
nand U3311 (N_3311,N_2556,N_159);
nor U3312 (N_3312,N_2836,N_1376);
xor U3313 (N_3313,N_110,N_1141);
xnor U3314 (N_3314,N_2200,N_2216);
nor U3315 (N_3315,N_2160,N_801);
xor U3316 (N_3316,N_267,N_2566);
nand U3317 (N_3317,N_414,N_2238);
and U3318 (N_3318,N_259,N_728);
and U3319 (N_3319,N_2351,N_609);
nor U3320 (N_3320,N_261,N_2410);
nor U3321 (N_3321,N_2916,N_371);
nand U3322 (N_3322,N_2649,N_2338);
xnor U3323 (N_3323,N_2473,N_1460);
xnor U3324 (N_3324,N_2920,N_1798);
nor U3325 (N_3325,N_1467,N_1475);
xnor U3326 (N_3326,N_2599,N_171);
nor U3327 (N_3327,N_1587,N_2454);
and U3328 (N_3328,N_752,N_172);
or U3329 (N_3329,N_1041,N_2126);
xor U3330 (N_3330,N_1469,N_231);
nor U3331 (N_3331,N_1589,N_85);
nand U3332 (N_3332,N_530,N_2459);
or U3333 (N_3333,N_753,N_1156);
and U3334 (N_3334,N_1245,N_1308);
or U3335 (N_3335,N_233,N_282);
nand U3336 (N_3336,N_2043,N_2052);
nand U3337 (N_3337,N_413,N_2498);
xnor U3338 (N_3338,N_1463,N_517);
xnor U3339 (N_3339,N_2077,N_2422);
nor U3340 (N_3340,N_2261,N_1767);
nor U3341 (N_3341,N_1896,N_200);
nor U3342 (N_3342,N_1363,N_1395);
nand U3343 (N_3343,N_714,N_2071);
and U3344 (N_3344,N_556,N_94);
or U3345 (N_3345,N_2841,N_1953);
or U3346 (N_3346,N_37,N_1179);
nor U3347 (N_3347,N_1980,N_2065);
nand U3348 (N_3348,N_2842,N_153);
or U3349 (N_3349,N_1904,N_2449);
or U3350 (N_3350,N_2812,N_334);
nor U3351 (N_3351,N_1578,N_889);
or U3352 (N_3352,N_191,N_1617);
nand U3353 (N_3353,N_619,N_1432);
nand U3354 (N_3354,N_1364,N_1885);
nor U3355 (N_3355,N_700,N_168);
nand U3356 (N_3356,N_2044,N_2531);
or U3357 (N_3357,N_2550,N_922);
and U3358 (N_3358,N_396,N_1731);
nand U3359 (N_3359,N_959,N_613);
xor U3360 (N_3360,N_2939,N_427);
nand U3361 (N_3361,N_2285,N_2493);
xnor U3362 (N_3362,N_2101,N_2229);
nand U3363 (N_3363,N_1974,N_2167);
and U3364 (N_3364,N_2622,N_1263);
and U3365 (N_3365,N_2264,N_1807);
or U3366 (N_3366,N_2902,N_1608);
or U3367 (N_3367,N_2358,N_35);
xnor U3368 (N_3368,N_1030,N_1127);
nor U3369 (N_3369,N_1053,N_481);
or U3370 (N_3370,N_2429,N_616);
or U3371 (N_3371,N_2458,N_2886);
nor U3372 (N_3372,N_2690,N_2169);
and U3373 (N_3373,N_1778,N_2545);
and U3374 (N_3374,N_1136,N_1869);
nand U3375 (N_3375,N_2960,N_1950);
or U3376 (N_3376,N_1097,N_932);
or U3377 (N_3377,N_870,N_1297);
or U3378 (N_3378,N_1428,N_1914);
or U3379 (N_3379,N_2913,N_392);
or U3380 (N_3380,N_1010,N_2788);
and U3381 (N_3381,N_1966,N_167);
nor U3382 (N_3382,N_907,N_1092);
xor U3383 (N_3383,N_1503,N_255);
xor U3384 (N_3384,N_2552,N_2969);
nor U3385 (N_3385,N_2885,N_1196);
nand U3386 (N_3386,N_2018,N_232);
nand U3387 (N_3387,N_1858,N_444);
nand U3388 (N_3388,N_614,N_2991);
nor U3389 (N_3389,N_1217,N_1082);
xor U3390 (N_3390,N_2291,N_2471);
xor U3391 (N_3391,N_1588,N_1321);
nor U3392 (N_3392,N_109,N_893);
or U3393 (N_3393,N_689,N_1595);
xor U3394 (N_3394,N_561,N_433);
nor U3395 (N_3395,N_850,N_2693);
or U3396 (N_3396,N_1678,N_2104);
or U3397 (N_3397,N_1810,N_1216);
nand U3398 (N_3398,N_1747,N_660);
xor U3399 (N_3399,N_1208,N_998);
or U3400 (N_3400,N_432,N_1988);
or U3401 (N_3401,N_809,N_864);
or U3402 (N_3402,N_1128,N_1442);
or U3403 (N_3403,N_43,N_1930);
xor U3404 (N_3404,N_2981,N_2967);
nand U3405 (N_3405,N_438,N_1105);
or U3406 (N_3406,N_2750,N_1754);
and U3407 (N_3407,N_268,N_2793);
nand U3408 (N_3408,N_581,N_1123);
xnor U3409 (N_3409,N_1820,N_1434);
xor U3410 (N_3410,N_1264,N_2249);
xnor U3411 (N_3411,N_586,N_185);
nor U3412 (N_3412,N_1760,N_671);
xnor U3413 (N_3413,N_2543,N_2244);
nand U3414 (N_3414,N_2409,N_315);
and U3415 (N_3415,N_1913,N_1362);
and U3416 (N_3416,N_1713,N_987);
xor U3417 (N_3417,N_299,N_1828);
xnor U3418 (N_3418,N_2685,N_1038);
nor U3419 (N_3419,N_906,N_2203);
nor U3420 (N_3420,N_1813,N_1972);
nand U3421 (N_3421,N_550,N_2392);
and U3422 (N_3422,N_1259,N_2899);
or U3423 (N_3423,N_1922,N_2215);
xnor U3424 (N_3424,N_1631,N_417);
nor U3425 (N_3425,N_610,N_1054);
nand U3426 (N_3426,N_843,N_1859);
nand U3427 (N_3427,N_1962,N_2751);
or U3428 (N_3428,N_802,N_2568);
and U3429 (N_3429,N_2213,N_2083);
xor U3430 (N_3430,N_2191,N_1394);
nand U3431 (N_3431,N_1025,N_2597);
nor U3432 (N_3432,N_2975,N_1825);
xor U3433 (N_3433,N_1894,N_1790);
xnor U3434 (N_3434,N_2278,N_1477);
nand U3435 (N_3435,N_2834,N_2024);
and U3436 (N_3436,N_2508,N_2379);
or U3437 (N_3437,N_1727,N_1933);
nand U3438 (N_3438,N_2073,N_1171);
or U3439 (N_3439,N_2610,N_1050);
nor U3440 (N_3440,N_450,N_2993);
nand U3441 (N_3441,N_844,N_970);
or U3442 (N_3442,N_2110,N_1199);
xnor U3443 (N_3443,N_491,N_225);
nor U3444 (N_3444,N_1201,N_2016);
xnor U3445 (N_3445,N_1538,N_2204);
xnor U3446 (N_3446,N_877,N_1167);
or U3447 (N_3447,N_2500,N_2494);
nand U3448 (N_3448,N_2518,N_1583);
nand U3449 (N_3449,N_1499,N_1326);
and U3450 (N_3450,N_1646,N_983);
or U3451 (N_3451,N_2117,N_2922);
or U3452 (N_3452,N_398,N_1366);
nor U3453 (N_3453,N_2863,N_2265);
nand U3454 (N_3454,N_2446,N_1806);
nand U3455 (N_3455,N_154,N_322);
nor U3456 (N_3456,N_1146,N_1691);
or U3457 (N_3457,N_2728,N_1279);
or U3458 (N_3458,N_23,N_1377);
xnor U3459 (N_3459,N_692,N_2373);
nand U3460 (N_3460,N_2372,N_2587);
xor U3461 (N_3461,N_1635,N_1207);
xnor U3462 (N_3462,N_2190,N_1640);
xnor U3463 (N_3463,N_2270,N_2089);
nand U3464 (N_3464,N_178,N_1169);
xnor U3465 (N_3465,N_1897,N_2995);
nand U3466 (N_3466,N_2377,N_119);
nor U3467 (N_3467,N_721,N_1122);
xor U3468 (N_3468,N_947,N_868);
xnor U3469 (N_3469,N_697,N_2149);
nor U3470 (N_3470,N_2015,N_2840);
nor U3471 (N_3471,N_2856,N_966);
or U3472 (N_3472,N_128,N_38);
and U3473 (N_3473,N_1046,N_1464);
or U3474 (N_3474,N_1212,N_859);
xnor U3475 (N_3475,N_2269,N_862);
nand U3476 (N_3476,N_2957,N_521);
and U3477 (N_3477,N_2507,N_1160);
or U3478 (N_3478,N_991,N_1170);
or U3479 (N_3479,N_2245,N_2174);
nand U3480 (N_3480,N_2623,N_445);
and U3481 (N_3481,N_44,N_979);
nor U3482 (N_3482,N_1409,N_45);
or U3483 (N_3483,N_1679,N_2882);
nand U3484 (N_3484,N_626,N_992);
or U3485 (N_3485,N_2349,N_582);
nand U3486 (N_3486,N_2463,N_2915);
nor U3487 (N_3487,N_3,N_905);
nand U3488 (N_3488,N_1391,N_308);
nor U3489 (N_3489,N_503,N_852);
nor U3490 (N_3490,N_2151,N_807);
nand U3491 (N_3491,N_51,N_2784);
and U3492 (N_3492,N_1223,N_2415);
xnor U3493 (N_3493,N_60,N_2741);
and U3494 (N_3494,N_2478,N_2526);
and U3495 (N_3495,N_2428,N_424);
nand U3496 (N_3496,N_2341,N_762);
or U3497 (N_3497,N_2694,N_769);
and U3498 (N_3498,N_2061,N_123);
nand U3499 (N_3499,N_1112,N_1804);
nor U3500 (N_3500,N_535,N_1476);
nor U3501 (N_3501,N_2154,N_1087);
xnor U3502 (N_3502,N_158,N_533);
or U3503 (N_3503,N_1151,N_577);
or U3504 (N_3504,N_329,N_2731);
nand U3505 (N_3505,N_64,N_1241);
and U3506 (N_3506,N_2665,N_1990);
nor U3507 (N_3507,N_2081,N_2041);
and U3508 (N_3508,N_872,N_39);
nor U3509 (N_3509,N_774,N_687);
nor U3510 (N_3510,N_2608,N_29);
and U3511 (N_3511,N_2085,N_2821);
and U3512 (N_3512,N_2439,N_1995);
and U3513 (N_3513,N_672,N_2339);
and U3514 (N_3514,N_1180,N_2814);
nand U3515 (N_3515,N_2671,N_2055);
nand U3516 (N_3516,N_2408,N_380);
and U3517 (N_3517,N_910,N_2968);
or U3518 (N_3518,N_1765,N_2857);
or U3519 (N_3519,N_1945,N_2912);
or U3520 (N_3520,N_602,N_2218);
or U3521 (N_3521,N_2754,N_2901);
and U3522 (N_3522,N_2100,N_1598);
or U3523 (N_3523,N_918,N_2717);
and U3524 (N_3524,N_1743,N_2485);
xnor U3525 (N_3525,N_1065,N_1770);
or U3526 (N_3526,N_295,N_1808);
xor U3527 (N_3527,N_1905,N_1925);
nor U3528 (N_3528,N_555,N_1195);
and U3529 (N_3529,N_2390,N_1725);
or U3530 (N_3530,N_2514,N_351);
nor U3531 (N_3531,N_189,N_1871);
nand U3532 (N_3532,N_2343,N_741);
xor U3533 (N_3533,N_2963,N_787);
or U3534 (N_3534,N_429,N_1968);
nor U3535 (N_3535,N_2837,N_2749);
nor U3536 (N_3536,N_319,N_520);
and U3537 (N_3537,N_1300,N_2455);
or U3538 (N_3538,N_2734,N_2421);
xor U3539 (N_3539,N_1613,N_1815);
nor U3540 (N_3540,N_2626,N_1638);
nor U3541 (N_3541,N_1982,N_1921);
or U3542 (N_3542,N_2551,N_2953);
and U3543 (N_3543,N_1077,N_1324);
xor U3544 (N_3544,N_1446,N_1948);
nor U3545 (N_3545,N_1138,N_2322);
and U3546 (N_3546,N_1864,N_590);
nor U3547 (N_3547,N_2710,N_2835);
nand U3548 (N_3548,N_260,N_2908);
xnor U3549 (N_3549,N_61,N_1775);
or U3550 (N_3550,N_1109,N_2113);
or U3551 (N_3551,N_1758,N_62);
xnor U3552 (N_3552,N_1149,N_1205);
xor U3553 (N_3553,N_2811,N_452);
nor U3554 (N_3554,N_2226,N_1282);
and U3555 (N_3555,N_1833,N_1370);
nor U3556 (N_3556,N_2416,N_2650);
xnor U3557 (N_3557,N_2006,N_598);
nor U3558 (N_3558,N_1581,N_2894);
nor U3559 (N_3559,N_2070,N_946);
xnor U3560 (N_3560,N_2949,N_1015);
and U3561 (N_3561,N_1655,N_2708);
nor U3562 (N_3562,N_839,N_632);
and U3563 (N_3563,N_2577,N_1562);
nor U3564 (N_3564,N_22,N_1615);
and U3565 (N_3565,N_366,N_2591);
nor U3566 (N_3566,N_1492,N_650);
nand U3567 (N_3567,N_505,N_938);
nor U3568 (N_3568,N_510,N_828);
and U3569 (N_3569,N_2340,N_1325);
or U3570 (N_3570,N_840,N_21);
and U3571 (N_3571,N_327,N_484);
nor U3572 (N_3572,N_1612,N_1142);
nand U3573 (N_3573,N_2225,N_1788);
or U3574 (N_3574,N_1585,N_1541);
nand U3575 (N_3575,N_228,N_2418);
and U3576 (N_3576,N_1389,N_2616);
or U3577 (N_3577,N_659,N_1732);
and U3578 (N_3578,N_117,N_70);
or U3579 (N_3579,N_1088,N_430);
nor U3580 (N_3580,N_1185,N_132);
and U3581 (N_3581,N_2438,N_2711);
nand U3582 (N_3582,N_1317,N_2005);
nor U3583 (N_3583,N_2139,N_1791);
or U3584 (N_3584,N_1246,N_851);
xnor U3585 (N_3585,N_969,N_26);
or U3586 (N_3586,N_348,N_2825);
nor U3587 (N_3587,N_538,N_1520);
nor U3588 (N_3588,N_1571,N_176);
or U3589 (N_3589,N_2951,N_12);
nand U3590 (N_3590,N_2839,N_822);
or U3591 (N_3591,N_751,N_2609);
nor U3592 (N_3592,N_2830,N_1322);
nand U3593 (N_3593,N_116,N_1134);
or U3594 (N_3594,N_263,N_292);
or U3595 (N_3595,N_565,N_1075);
nand U3596 (N_3596,N_2266,N_669);
nor U3597 (N_3597,N_1978,N_53);
or U3598 (N_3598,N_2166,N_531);
xnor U3599 (N_3599,N_2143,N_2895);
nand U3600 (N_3600,N_2795,N_1437);
nand U3601 (N_3601,N_2538,N_2871);
xnor U3602 (N_3602,N_543,N_846);
nand U3603 (N_3603,N_399,N_1348);
nand U3604 (N_3604,N_2420,N_108);
and U3605 (N_3605,N_1551,N_754);
xnor U3606 (N_3606,N_724,N_585);
nor U3607 (N_3607,N_1117,N_2381);
nor U3608 (N_3608,N_2744,N_385);
and U3609 (N_3609,N_2460,N_217);
or U3610 (N_3610,N_576,N_2942);
or U3611 (N_3611,N_69,N_2724);
and U3612 (N_3612,N_1523,N_1570);
xnor U3613 (N_3613,N_658,N_162);
and U3614 (N_3614,N_1402,N_212);
or U3615 (N_3615,N_1932,N_1964);
nand U3616 (N_3616,N_2753,N_1235);
nor U3617 (N_3617,N_2790,N_748);
nand U3618 (N_3618,N_471,N_2653);
xnor U3619 (N_3619,N_395,N_440);
nand U3620 (N_3620,N_1024,N_1120);
or U3621 (N_3621,N_2783,N_808);
or U3622 (N_3622,N_1222,N_2888);
and U3623 (N_3623,N_194,N_522);
xor U3624 (N_3624,N_637,N_2603);
xor U3625 (N_3625,N_731,N_799);
nor U3626 (N_3626,N_83,N_758);
or U3627 (N_3627,N_662,N_1689);
nor U3628 (N_3628,N_303,N_664);
nand U3629 (N_3629,N_847,N_1762);
nand U3630 (N_3630,N_1238,N_1949);
nand U3631 (N_3631,N_1675,N_101);
or U3632 (N_3632,N_916,N_1901);
nor U3633 (N_3633,N_1265,N_65);
xor U3634 (N_3634,N_892,N_197);
or U3635 (N_3635,N_25,N_2360);
nand U3636 (N_3636,N_254,N_607);
or U3637 (N_3637,N_2185,N_1489);
xnor U3638 (N_3638,N_2398,N_2333);
or U3639 (N_3639,N_1522,N_2231);
and U3640 (N_3640,N_841,N_1676);
nor U3641 (N_3641,N_2347,N_2378);
nand U3642 (N_3642,N_2142,N_1479);
xnor U3643 (N_3643,N_1599,N_206);
nand U3644 (N_3644,N_1961,N_2925);
and U3645 (N_3645,N_1600,N_2357);
and U3646 (N_3646,N_594,N_2331);
nor U3647 (N_3647,N_1320,N_1722);
nor U3648 (N_3648,N_2434,N_2644);
nor U3649 (N_3649,N_564,N_2383);
and U3650 (N_3650,N_924,N_155);
xor U3651 (N_3651,N_425,N_141);
nand U3652 (N_3652,N_810,N_378);
and U3653 (N_3653,N_2573,N_1521);
xnor U3654 (N_3654,N_2763,N_2010);
nor U3655 (N_3655,N_2891,N_2877);
and U3656 (N_3656,N_1288,N_107);
or U3657 (N_3657,N_2686,N_1093);
nand U3658 (N_3658,N_1140,N_1575);
nor U3659 (N_3659,N_2008,N_381);
or U3660 (N_3660,N_135,N_1040);
and U3661 (N_3661,N_2743,N_2770);
nor U3662 (N_3662,N_620,N_307);
nand U3663 (N_3663,N_1823,N_1734);
and U3664 (N_3664,N_2000,N_1865);
nand U3665 (N_3665,N_745,N_883);
nor U3666 (N_3666,N_187,N_1509);
nor U3667 (N_3667,N_2050,N_113);
xor U3668 (N_3668,N_1592,N_1927);
xor U3669 (N_3669,N_1777,N_283);
nor U3670 (N_3670,N_940,N_2092);
and U3671 (N_3671,N_559,N_686);
and U3672 (N_3672,N_2624,N_321);
and U3673 (N_3673,N_188,N_1939);
nor U3674 (N_3674,N_1270,N_1111);
and U3675 (N_3675,N_1311,N_2311);
nor U3676 (N_3676,N_2259,N_8);
xnor U3677 (N_3677,N_92,N_1431);
and U3678 (N_3678,N_1741,N_140);
xnor U3679 (N_3679,N_634,N_2643);
xnor U3680 (N_3680,N_1202,N_1019);
or U3681 (N_3681,N_2391,N_2779);
nor U3682 (N_3682,N_1796,N_1435);
and U3683 (N_3683,N_742,N_2914);
nor U3684 (N_3684,N_2712,N_2107);
xnor U3685 (N_3685,N_1531,N_1632);
or U3686 (N_3686,N_1083,N_320);
xnor U3687 (N_3687,N_286,N_1684);
xnor U3688 (N_3688,N_1178,N_1008);
or U3689 (N_3689,N_1845,N_1443);
or U3690 (N_3690,N_2182,N_1002);
or U3691 (N_3691,N_2424,N_1421);
and U3692 (N_3692,N_1455,N_2105);
xor U3693 (N_3693,N_1708,N_1447);
xnor U3694 (N_3694,N_1628,N_1603);
or U3695 (N_3695,N_2306,N_2223);
and U3696 (N_3696,N_474,N_1197);
or U3697 (N_3697,N_2950,N_723);
nor U3698 (N_3698,N_2406,N_1413);
or U3699 (N_3699,N_2148,N_1661);
or U3700 (N_3700,N_2548,N_1540);
or U3701 (N_3701,N_1305,N_1970);
xor U3702 (N_3702,N_302,N_1890);
and U3703 (N_3703,N_1996,N_2);
xor U3704 (N_3704,N_2662,N_2258);
xor U3705 (N_3705,N_2562,N_1855);
xor U3706 (N_3706,N_849,N_2115);
xnor U3707 (N_3707,N_2267,N_2561);
nor U3708 (N_3708,N_2719,N_2417);
and U3709 (N_3709,N_494,N_1593);
nand U3710 (N_3710,N_1683,N_950);
nor U3711 (N_3711,N_696,N_1500);
xnor U3712 (N_3712,N_1426,N_1302);
nand U3713 (N_3713,N_2289,N_2233);
xor U3714 (N_3714,N_353,N_1047);
xor U3715 (N_3715,N_999,N_2806);
nor U3716 (N_3716,N_1751,N_1662);
nand U3717 (N_3717,N_1699,N_2078);
and U3718 (N_3718,N_1651,N_1528);
nor U3719 (N_3719,N_1702,N_125);
xnor U3720 (N_3720,N_2116,N_120);
nor U3721 (N_3721,N_1036,N_2590);
and U3722 (N_3722,N_241,N_900);
nand U3723 (N_3723,N_2099,N_2521);
nor U3724 (N_3724,N_1309,N_2973);
or U3725 (N_3725,N_1942,N_953);
xnor U3726 (N_3726,N_2112,N_2382);
or U3727 (N_3727,N_248,N_1991);
xnor U3728 (N_3728,N_2813,N_2095);
nor U3729 (N_3729,N_806,N_2601);
or U3730 (N_3730,N_412,N_1405);
and U3731 (N_3731,N_1101,N_2132);
and U3732 (N_3732,N_2998,N_2651);
or U3733 (N_3733,N_2325,N_229);
and U3734 (N_3734,N_2506,N_1233);
nand U3735 (N_3735,N_2679,N_1228);
xnor U3736 (N_3736,N_674,N_1644);
nor U3737 (N_3737,N_2181,N_949);
nand U3738 (N_3738,N_963,N_2355);
xor U3739 (N_3739,N_777,N_2850);
nand U3740 (N_3740,N_2815,N_668);
nor U3741 (N_3741,N_1887,N_352);
nand U3742 (N_3742,N_1513,N_258);
xnor U3743 (N_3743,N_2497,N_2619);
nand U3744 (N_3744,N_2658,N_2958);
or U3745 (N_3745,N_848,N_1249);
or U3746 (N_3746,N_431,N_803);
or U3747 (N_3747,N_2640,N_382);
xnor U3748 (N_3748,N_1382,N_1343);
nor U3749 (N_3749,N_2125,N_759);
and U3750 (N_3750,N_256,N_2437);
and U3751 (N_3751,N_2766,N_1074);
nor U3752 (N_3752,N_478,N_1069);
and U3753 (N_3753,N_506,N_622);
or U3754 (N_3754,N_819,N_1611);
nor U3755 (N_3755,N_1301,N_235);
nand U3756 (N_3756,N_249,N_1648);
nor U3757 (N_3757,N_1438,N_955);
nand U3758 (N_3758,N_2198,N_2082);
and U3759 (N_3759,N_1497,N_2873);
xor U3760 (N_3760,N_1878,N_2152);
nor U3761 (N_3761,N_1652,N_562);
and U3762 (N_3762,N_1555,N_2496);
nand U3763 (N_3763,N_2023,N_1534);
or U3764 (N_3764,N_1682,N_1835);
xor U3765 (N_3765,N_1417,N_376);
nand U3766 (N_3766,N_1653,N_2035);
nor U3767 (N_3767,N_2765,N_830);
xnor U3768 (N_3768,N_1623,N_615);
nand U3769 (N_3769,N_605,N_220);
and U3770 (N_3770,N_2491,N_2337);
nor U3771 (N_3771,N_1383,N_964);
nand U3772 (N_3772,N_2465,N_1789);
nand U3773 (N_3773,N_402,N_1918);
nand U3774 (N_3774,N_2489,N_87);
xor U3775 (N_3775,N_2668,N_1470);
nor U3776 (N_3776,N_1843,N_2184);
and U3777 (N_3777,N_2161,N_898);
and U3778 (N_3778,N_2631,N_1070);
nand U3779 (N_3779,N_1368,N_1174);
and U3780 (N_3780,N_1203,N_1546);
and U3781 (N_3781,N_2286,N_122);
nor U3782 (N_3782,N_2298,N_81);
or U3783 (N_3783,N_1103,N_2295);
nand U3784 (N_3784,N_1558,N_1404);
nand U3785 (N_3785,N_2457,N_1811);
nor U3786 (N_3786,N_1225,N_2870);
nand U3787 (N_3787,N_2832,N_2688);
nand U3788 (N_3788,N_739,N_2486);
nand U3789 (N_3789,N_57,N_1660);
xor U3790 (N_3790,N_2739,N_1537);
nor U3791 (N_3791,N_593,N_1565);
or U3792 (N_3792,N_1917,N_2645);
nand U3793 (N_3793,N_2745,N_342);
or U3794 (N_3794,N_1868,N_1461);
nand U3795 (N_3795,N_2595,N_2542);
xnor U3796 (N_3796,N_1295,N_1287);
or U3797 (N_3797,N_407,N_719);
and U3798 (N_3798,N_2936,N_339);
xnor U3799 (N_3799,N_1669,N_1023);
and U3800 (N_3800,N_2064,N_874);
xnor U3801 (N_3801,N_99,N_1742);
xnor U3802 (N_3802,N_2492,N_1639);
and U3803 (N_3803,N_1483,N_1923);
nand U3804 (N_3804,N_224,N_1013);
nor U3805 (N_3805,N_1840,N_1033);
nand U3806 (N_3806,N_1032,N_74);
xnor U3807 (N_3807,N_680,N_2056);
or U3808 (N_3808,N_1144,N_2450);
or U3809 (N_3809,N_1215,N_426);
and U3810 (N_3810,N_1110,N_2150);
xnor U3811 (N_3811,N_2759,N_318);
nor U3812 (N_3812,N_2049,N_2323);
and U3813 (N_3813,N_264,N_706);
nor U3814 (N_3814,N_272,N_1258);
and U3815 (N_3815,N_2228,N_301);
nand U3816 (N_3816,N_975,N_252);
or U3817 (N_3817,N_2933,N_1866);
nor U3818 (N_3818,N_2165,N_146);
nand U3819 (N_3819,N_1872,N_186);
or U3820 (N_3820,N_2461,N_2042);
and U3821 (N_3821,N_2666,N_1812);
xor U3822 (N_3822,N_1959,N_397);
and U3823 (N_3823,N_1462,N_2988);
xnor U3824 (N_3824,N_2656,N_656);
nor U3825 (N_3825,N_2965,N_1975);
nand U3826 (N_3826,N_2786,N_526);
or U3827 (N_3827,N_1677,N_2517);
nor U3828 (N_3828,N_2176,N_1218);
xor U3829 (N_3829,N_1369,N_387);
and U3830 (N_3830,N_234,N_1102);
and U3831 (N_3831,N_1260,N_2588);
or U3832 (N_3832,N_2354,N_2484);
nor U3833 (N_3833,N_1672,N_181);
and U3834 (N_3834,N_1490,N_643);
or U3835 (N_3835,N_2401,N_952);
and U3836 (N_3836,N_390,N_1580);
or U3837 (N_3837,N_980,N_1647);
or U3838 (N_3838,N_1058,N_134);
and U3839 (N_3839,N_1044,N_1076);
nor U3840 (N_3840,N_2251,N_96);
nand U3841 (N_3841,N_734,N_1210);
xnor U3842 (N_3842,N_2370,N_1372);
nand U3843 (N_3843,N_324,N_812);
and U3844 (N_3844,N_2714,N_2844);
xor U3845 (N_3845,N_2281,N_885);
nand U3846 (N_3846,N_2872,N_2893);
and U3847 (N_3847,N_965,N_24);
nand U3848 (N_3848,N_2966,N_1107);
or U3849 (N_3849,N_1028,N_1);
and U3850 (N_3850,N_738,N_142);
or U3851 (N_3851,N_1126,N_2516);
and U3852 (N_3852,N_1803,N_1836);
and U3853 (N_3853,N_1392,N_911);
nor U3854 (N_3854,N_163,N_1119);
nand U3855 (N_3855,N_1875,N_331);
or U3856 (N_3856,N_948,N_1336);
or U3857 (N_3857,N_2612,N_2344);
or U3858 (N_3858,N_1465,N_873);
nor U3859 (N_3859,N_47,N_1339);
nor U3860 (N_3860,N_1645,N_879);
or U3861 (N_3861,N_547,N_1548);
and U3862 (N_3862,N_2986,N_2904);
nor U3863 (N_3863,N_441,N_271);
or U3864 (N_3864,N_875,N_2769);
and U3865 (N_3865,N_2697,N_2747);
or U3866 (N_3866,N_2661,N_288);
and U3867 (N_3867,N_954,N_394);
nor U3868 (N_3868,N_1018,N_1089);
nor U3869 (N_3869,N_379,N_2342);
nor U3870 (N_3870,N_1712,N_2407);
xor U3871 (N_3871,N_2761,N_2505);
nor U3872 (N_3872,N_989,N_2822);
and U3873 (N_3873,N_1862,N_1746);
nand U3874 (N_3874,N_386,N_2495);
and U3875 (N_3875,N_2964,N_2576);
and U3876 (N_3876,N_710,N_1457);
or U3877 (N_3877,N_1049,N_682);
xor U3878 (N_3878,N_1472,N_496);
xnor U3879 (N_3879,N_1730,N_1895);
and U3880 (N_3880,N_2239,N_500);
and U3881 (N_3881,N_1633,N_2232);
xor U3882 (N_3882,N_2114,N_1494);
nand U3883 (N_3883,N_1616,N_1452);
and U3884 (N_3884,N_262,N_1488);
nor U3885 (N_3885,N_1275,N_2057);
xnor U3886 (N_3886,N_2155,N_666);
xnor U3887 (N_3887,N_2194,N_855);
and U3888 (N_3888,N_649,N_1080);
nor U3889 (N_3889,N_2874,N_645);
or U3890 (N_3890,N_972,N_354);
nand U3891 (N_3891,N_549,N_467);
and U3892 (N_3892,N_1837,N_2827);
nand U3893 (N_3893,N_960,N_2781);
xnor U3894 (N_3894,N_2479,N_2499);
and U3895 (N_3895,N_251,N_1341);
nand U3896 (N_3896,N_136,N_174);
and U3897 (N_3897,N_2442,N_2425);
or U3898 (N_3898,N_2301,N_647);
nor U3899 (N_3899,N_2464,N_1929);
xnor U3900 (N_3900,N_446,N_313);
or U3901 (N_3901,N_1379,N_456);
or U3902 (N_3902,N_1761,N_1847);
xor U3903 (N_3903,N_1150,N_832);
or U3904 (N_3904,N_1844,N_2362);
nor U3905 (N_3905,N_9,N_2230);
nand U3906 (N_3906,N_2553,N_363);
nor U3907 (N_3907,N_780,N_1296);
or U3908 (N_3908,N_1192,N_1745);
nor U3909 (N_3909,N_488,N_2158);
and U3910 (N_3910,N_2053,N_2208);
xnor U3911 (N_3911,N_1508,N_374);
nor U3912 (N_3912,N_218,N_2027);
and U3913 (N_3913,N_205,N_1240);
or U3914 (N_3914,N_2729,N_2978);
nand U3915 (N_3915,N_306,N_1686);
or U3916 (N_3916,N_2696,N_957);
xnor U3917 (N_3917,N_2585,N_2034);
or U3918 (N_3918,N_1027,N_2481);
nand U3919 (N_3919,N_2186,N_1784);
xnor U3920 (N_3920,N_2141,N_157);
nand U3921 (N_3921,N_551,N_2436);
xnor U3922 (N_3922,N_95,N_757);
or U3923 (N_3923,N_2799,N_2480);
or U3924 (N_3924,N_1060,N_2648);
nand U3925 (N_3925,N_2752,N_795);
nor U3926 (N_3926,N_2011,N_1237);
xor U3927 (N_3927,N_326,N_2255);
nand U3928 (N_3928,N_2147,N_1106);
and U3929 (N_3929,N_729,N_1723);
and U3930 (N_3930,N_837,N_317);
or U3931 (N_3931,N_1121,N_962);
and U3932 (N_3932,N_2451,N_1176);
nor U3933 (N_3933,N_164,N_2087);
nand U3934 (N_3934,N_542,N_79);
nor U3935 (N_3935,N_1721,N_1830);
or U3936 (N_3936,N_1029,N_410);
and U3937 (N_3937,N_247,N_2804);
nor U3938 (N_3938,N_2019,N_2031);
and U3939 (N_3939,N_127,N_193);
nand U3940 (N_3940,N_304,N_1064);
nor U3941 (N_3941,N_2829,N_497);
nor U3942 (N_3942,N_2026,N_490);
nor U3943 (N_3943,N_121,N_1043);
nand U3944 (N_3944,N_2193,N_1401);
nor U3945 (N_3945,N_2720,N_1414);
or U3946 (N_3946,N_2756,N_2183);
nor U3947 (N_3947,N_540,N_2319);
or U3948 (N_3948,N_1773,N_1118);
or U3949 (N_3949,N_1524,N_2536);
or U3950 (N_3950,N_833,N_779);
and U3951 (N_3951,N_1692,N_1441);
or U3952 (N_3952,N_2943,N_383);
nor U3953 (N_3953,N_333,N_1292);
nand U3954 (N_3954,N_816,N_2103);
and U3955 (N_3955,N_518,N_103);
nand U3956 (N_3956,N_1147,N_2816);
xnor U3957 (N_3957,N_2940,N_2210);
nor U3958 (N_3958,N_2403,N_618);
xnor U3959 (N_3959,N_956,N_1360);
xor U3960 (N_3960,N_1378,N_13);
or U3961 (N_3961,N_2088,N_131);
and U3962 (N_3962,N_2187,N_71);
and U3963 (N_3963,N_732,N_798);
xnor U3964 (N_3964,N_1641,N_1042);
xnor U3965 (N_3965,N_592,N_2722);
nand U3966 (N_3966,N_1584,N_571);
and U3967 (N_3967,N_1346,N_2207);
nor U3968 (N_3968,N_935,N_2072);
xor U3969 (N_3969,N_17,N_1357);
xor U3970 (N_3970,N_104,N_1159);
nor U3971 (N_3971,N_2868,N_600);
xnor U3972 (N_3972,N_346,N_203);
nor U3973 (N_3973,N_2946,N_1451);
nand U3974 (N_3974,N_1448,N_853);
xnor U3975 (N_3975,N_773,N_2673);
and U3976 (N_3976,N_2641,N_1733);
xnor U3977 (N_3977,N_746,N_1512);
nor U3978 (N_3978,N_2937,N_788);
and U3979 (N_3979,N_2268,N_507);
nand U3980 (N_3980,N_1386,N_1257);
nor U3981 (N_3981,N_1486,N_612);
nor U3982 (N_3982,N_2682,N_360);
or U3983 (N_3983,N_56,N_475);
nand U3984 (N_3984,N_27,N_296);
or U3985 (N_3985,N_1935,N_1759);
and U3986 (N_3986,N_1851,N_2855);
xor U3987 (N_3987,N_130,N_2660);
and U3988 (N_3988,N_2079,N_755);
nor U3989 (N_3989,N_984,N_1335);
nand U3990 (N_3990,N_2046,N_2613);
or U3991 (N_3991,N_2594,N_1532);
nor U3992 (N_3992,N_2721,N_2365);
nor U3993 (N_3993,N_1941,N_114);
nand U3994 (N_3994,N_1085,N_1468);
or U3995 (N_3995,N_1312,N_2260);
xor U3996 (N_3996,N_2211,N_1355);
xnor U3997 (N_3997,N_14,N_464);
nand U3998 (N_3998,N_40,N_2546);
nor U3999 (N_3999,N_1502,N_1586);
or U4000 (N_4000,N_707,N_1839);
nor U4001 (N_4001,N_2692,N_1188);
xnor U4002 (N_4002,N_2059,N_2108);
nand U4003 (N_4003,N_570,N_2334);
and U4004 (N_4004,N_1135,N_2447);
nand U4005 (N_4005,N_1695,N_894);
and U4006 (N_4006,N_884,N_1380);
nand U4007 (N_4007,N_2927,N_1081);
nor U4008 (N_4008,N_2525,N_1012);
nand U4009 (N_4009,N_1707,N_2067);
nand U4010 (N_4010,N_2032,N_2520);
or U4011 (N_4011,N_2972,N_1026);
nor U4012 (N_4012,N_1132,N_2427);
and U4013 (N_4013,N_1090,N_2584);
nor U4014 (N_4014,N_824,N_330);
xnor U4015 (N_4015,N_275,N_2600);
xor U4016 (N_4016,N_2371,N_20);
nand U4017 (N_4017,N_688,N_1838);
or U4018 (N_4018,N_797,N_1946);
nor U4019 (N_4019,N_416,N_514);
nand U4020 (N_4020,N_2919,N_939);
nand U4021 (N_4021,N_2400,N_1673);
nand U4022 (N_4022,N_2954,N_1911);
nand U4023 (N_4023,N_2800,N_2735);
nand U4024 (N_4024,N_1484,N_886);
xnor U4025 (N_4025,N_1162,N_2021);
or U4026 (N_4026,N_298,N_411);
xnor U4027 (N_4027,N_1124,N_1236);
nor U4028 (N_4028,N_995,N_630);
and U4029 (N_4029,N_1940,N_284);
nor U4030 (N_4030,N_2921,N_2565);
nor U4031 (N_4031,N_7,N_1133);
and U4032 (N_4032,N_213,N_772);
xnor U4033 (N_4033,N_515,N_2607);
xnor U4034 (N_4034,N_2699,N_528);
xor U4035 (N_4035,N_1573,N_369);
nor U4036 (N_4036,N_2257,N_2475);
xor U4037 (N_4037,N_461,N_2742);
or U4038 (N_4038,N_2798,N_988);
nor U4039 (N_4039,N_372,N_2237);
xnor U4040 (N_4040,N_2522,N_856);
nand U4041 (N_4041,N_2017,N_580);
or U4042 (N_4042,N_1981,N_1667);
or U4043 (N_4043,N_160,N_2982);
or U4044 (N_4044,N_1792,N_55);
xnor U4045 (N_4045,N_405,N_1098);
and U4046 (N_4046,N_2718,N_1579);
and U4047 (N_4047,N_46,N_215);
nor U4048 (N_4048,N_285,N_1016);
and U4049 (N_4049,N_978,N_1797);
or U4050 (N_4050,N_1650,N_794);
or U4051 (N_4051,N_2736,N_384);
or U4052 (N_4052,N_1415,N_449);
nor U4053 (N_4053,N_1515,N_337);
or U4054 (N_4054,N_920,N_917);
xor U4055 (N_4055,N_1471,N_2738);
or U4056 (N_4056,N_1232,N_80);
nand U4057 (N_4057,N_2074,N_305);
nand U4058 (N_4058,N_463,N_2935);
nor U4059 (N_4059,N_1048,N_2787);
and U4060 (N_4060,N_1131,N_6);
nor U4061 (N_4061,N_1802,N_1783);
and U4062 (N_4062,N_557,N_1491);
nand U4063 (N_4063,N_711,N_2777);
nand U4064 (N_4064,N_1051,N_67);
and U4065 (N_4065,N_786,N_2441);
nand U4066 (N_4066,N_694,N_373);
and U4067 (N_4067,N_1406,N_2374);
or U4068 (N_4068,N_2657,N_1381);
or U4069 (N_4069,N_1243,N_695);
and U4070 (N_4070,N_1954,N_2574);
xnor U4071 (N_4071,N_1244,N_1387);
nand U4072 (N_4072,N_1698,N_359);
xnor U4073 (N_4073,N_465,N_1768);
xnor U4074 (N_4074,N_2419,N_1062);
nand U4075 (N_4075,N_1582,N_2346);
and U4076 (N_4076,N_1310,N_1861);
nor U4077 (N_4077,N_1226,N_1399);
and U4078 (N_4078,N_2858,N_1482);
xnor U4079 (N_4079,N_1430,N_791);
and U4080 (N_4080,N_2691,N_611);
or U4081 (N_4081,N_1459,N_2971);
nand U4082 (N_4082,N_1271,N_243);
or U4083 (N_4083,N_2299,N_316);
nand U4084 (N_4084,N_858,N_1116);
nand U4085 (N_4085,N_477,N_1507);
and U4086 (N_4086,N_244,N_1501);
nand U4087 (N_4087,N_1714,N_199);
or U4088 (N_4088,N_588,N_1643);
and U4089 (N_4089,N_702,N_1979);
or U4090 (N_4090,N_1657,N_2947);
xnor U4091 (N_4091,N_1444,N_245);
xor U4092 (N_4092,N_214,N_1665);
or U4093 (N_4093,N_2903,N_2275);
and U4094 (N_4094,N_776,N_821);
or U4095 (N_4095,N_1248,N_2201);
xnor U4096 (N_4096,N_1458,N_1262);
nand U4097 (N_4097,N_1506,N_2713);
or U4098 (N_4098,N_1059,N_1824);
nor U4099 (N_4099,N_335,N_628);
xor U4100 (N_4100,N_2541,N_1848);
and U4101 (N_4101,N_183,N_2683);
and U4102 (N_4102,N_1704,N_880);
or U4103 (N_4103,N_1358,N_309);
nor U4104 (N_4104,N_1877,N_2560);
xnor U4105 (N_4105,N_1242,N_476);
or U4106 (N_4106,N_2039,N_2329);
xnor U4107 (N_4107,N_1626,N_2123);
or U4108 (N_4108,N_2153,N_1418);
and U4109 (N_4109,N_1354,N_811);
or U4110 (N_4110,N_1079,N_971);
nand U4111 (N_4111,N_546,N_1397);
and U4112 (N_4112,N_876,N_1356);
and U4113 (N_4113,N_1801,N_760);
nor U4114 (N_4114,N_2076,N_2324);
xor U4115 (N_4115,N_525,N_2926);
and U4116 (N_4116,N_895,N_336);
nor U4117 (N_4117,N_221,N_693);
or U4118 (N_4118,N_487,N_595);
and U4119 (N_4119,N_1916,N_784);
nor U4120 (N_4120,N_2444,N_442);
nand U4121 (N_4121,N_921,N_1884);
nand U4122 (N_4122,N_2236,N_2509);
nor U4123 (N_4123,N_2068,N_2579);
xor U4124 (N_4124,N_1937,N_2559);
and U4125 (N_4125,N_1045,N_300);
xor U4126 (N_4126,N_2740,N_1920);
nor U4127 (N_4127,N_1424,N_1385);
nand U4128 (N_4128,N_897,N_2502);
xnor U4129 (N_4129,N_2962,N_2197);
and U4130 (N_4130,N_1681,N_993);
nand U4131 (N_4131,N_1411,N_2797);
or U4132 (N_4132,N_1818,N_2277);
or U4133 (N_4133,N_1971,N_1155);
nor U4134 (N_4134,N_2221,N_1726);
or U4135 (N_4135,N_473,N_1893);
and U4136 (N_4136,N_1849,N_2900);
xnor U4137 (N_4137,N_177,N_1157);
or U4138 (N_4138,N_1874,N_1306);
nand U4139 (N_4139,N_1774,N_1303);
or U4140 (N_4140,N_2976,N_2852);
xor U4141 (N_4141,N_1879,N_2353);
nor U4142 (N_4142,N_1627,N_2748);
nand U4143 (N_4143,N_722,N_2312);
xor U4144 (N_4144,N_867,N_1963);
or U4145 (N_4145,N_1671,N_138);
and U4146 (N_4146,N_149,N_1436);
nor U4147 (N_4147,N_2180,N_207);
nor U4148 (N_4148,N_1396,N_1164);
or U4149 (N_4149,N_1898,N_1533);
nand U4150 (N_4150,N_102,N_100);
and U4151 (N_4151,N_2389,N_1728);
nor U4152 (N_4152,N_236,N_2366);
or U4153 (N_4153,N_2308,N_2397);
or U4154 (N_4154,N_2316,N_1209);
nor U4155 (N_4155,N_909,N_765);
nor U4156 (N_4156,N_2540,N_406);
nor U4157 (N_4157,N_2667,N_1055);
xnor U4158 (N_4158,N_2140,N_2022);
or U4159 (N_4159,N_1563,N_2040);
and U4160 (N_4160,N_2866,N_912);
xor U4161 (N_4161,N_1960,N_2170);
and U4162 (N_4162,N_48,N_2861);
and U4163 (N_4163,N_2923,N_2611);
and U4164 (N_4164,N_469,N_2178);
nor U4165 (N_4165,N_1166,N_2220);
or U4166 (N_4166,N_1063,N_2009);
or U4167 (N_4167,N_981,N_2254);
nor U4168 (N_4168,N_209,N_2386);
nor U4169 (N_4169,N_1605,N_537);
nor U4170 (N_4170,N_375,N_347);
nor U4171 (N_4171,N_2707,N_1091);
xnor U4172 (N_4172,N_388,N_184);
and U4173 (N_4173,N_1740,N_583);
nand U4174 (N_4174,N_1290,N_314);
xor U4175 (N_4175,N_1453,N_2809);
or U4176 (N_4176,N_196,N_400);
nor U4177 (N_4177,N_1061,N_137);
or U4178 (N_4178,N_1165,N_2985);
xnor U4179 (N_4179,N_19,N_472);
nor U4180 (N_4180,N_2879,N_2504);
xor U4181 (N_4181,N_2256,N_2737);
xor U4182 (N_4182,N_1495,N_454);
and U4183 (N_4183,N_1902,N_1220);
nand U4184 (N_4184,N_361,N_1793);
nor U4185 (N_4185,N_1351,N_340);
and U4186 (N_4186,N_1624,N_2033);
and U4187 (N_4187,N_1700,N_1352);
or U4188 (N_4188,N_532,N_1332);
nor U4189 (N_4189,N_1474,N_545);
nand U4190 (N_4190,N_1067,N_287);
nand U4191 (N_4191,N_2853,N_1095);
nand U4192 (N_4192,N_1706,N_891);
xor U4193 (N_4193,N_2234,N_2199);
and U4194 (N_4194,N_2654,N_66);
nand U4195 (N_4195,N_2979,N_1254);
or U4196 (N_4196,N_818,N_2655);
nor U4197 (N_4197,N_2700,N_1330);
nand U4198 (N_4198,N_2669,N_1005);
and U4199 (N_4199,N_253,N_2614);
nor U4200 (N_4200,N_1718,N_1193);
or U4201 (N_4201,N_563,N_977);
or U4202 (N_4202,N_293,N_2695);
nand U4203 (N_4203,N_1504,N_651);
xor U4204 (N_4204,N_2758,N_2136);
and U4205 (N_4205,N_2045,N_919);
nand U4206 (N_4206,N_460,N_2272);
nand U4207 (N_4207,N_1518,N_2634);
and U4208 (N_4208,N_2470,N_1175);
nor U4209 (N_4209,N_2387,N_133);
or U4210 (N_4210,N_2589,N_428);
nand U4211 (N_4211,N_1799,N_2970);
and U4212 (N_4212,N_2801,N_1525);
nand U4213 (N_4213,N_2571,N_2294);
nand U4214 (N_4214,N_961,N_2212);
or U4215 (N_4215,N_2974,N_2007);
nand U4216 (N_4216,N_265,N_523);
nand U4217 (N_4217,N_180,N_5);
nor U4218 (N_4218,N_448,N_1892);
nand U4219 (N_4219,N_553,N_2271);
nor U4220 (N_4220,N_2468,N_1654);
nand U4221 (N_4221,N_534,N_589);
xor U4222 (N_4222,N_703,N_1416);
nand U4223 (N_4223,N_730,N_202);
nor U4224 (N_4224,N_190,N_2557);
and U4225 (N_4225,N_2860,N_768);
nand U4226 (N_4226,N_2664,N_2726);
xor U4227 (N_4227,N_451,N_661);
xor U4228 (N_4228,N_1440,N_325);
and U4229 (N_4229,N_1926,N_657);
or U4230 (N_4230,N_785,N_945);
or U4231 (N_4231,N_2580,N_2474);
or U4232 (N_4232,N_1620,N_2453);
or U4233 (N_4233,N_1250,N_1696);
or U4234 (N_4234,N_1284,N_1782);
nand U4235 (N_4235,N_1100,N_800);
xor U4236 (N_4236,N_1729,N_1276);
or U4237 (N_4237,N_447,N_673);
nand U4238 (N_4238,N_985,N_2772);
nand U4239 (N_4239,N_2864,N_2466);
xor U4240 (N_4240,N_2701,N_887);
and U4241 (N_4241,N_192,N_2393);
nand U4242 (N_4242,N_2823,N_1298);
nand U4243 (N_4243,N_663,N_437);
and U4244 (N_4244,N_2172,N_896);
nor U4245 (N_4245,N_838,N_1143);
nor U4246 (N_4246,N_2036,N_560);
nand U4247 (N_4247,N_1072,N_2791);
nor U4248 (N_4248,N_28,N_2235);
and U4249 (N_4249,N_1680,N_1273);
xnor U4250 (N_4250,N_827,N_2345);
nand U4251 (N_4251,N_2767,N_937);
nor U4252 (N_4252,N_2310,N_2843);
nor U4253 (N_4253,N_2130,N_2773);
nand U4254 (N_4254,N_1934,N_1487);
and U4255 (N_4255,N_1407,N_2785);
nor U4256 (N_4256,N_1693,N_2515);
and U4257 (N_4257,N_98,N_2094);
nor U4258 (N_4258,N_2716,N_345);
and U4259 (N_4259,N_927,N_453);
or U4260 (N_4260,N_1456,N_2633);
or U4261 (N_4261,N_2030,N_2598);
nand U4262 (N_4262,N_2219,N_362);
nand U4263 (N_4263,N_2796,N_1906);
or U4264 (N_4264,N_2523,N_2120);
or U4265 (N_4265,N_1550,N_246);
nor U4266 (N_4266,N_269,N_2350);
or U4267 (N_4267,N_524,N_2025);
nor U4268 (N_4268,N_2063,N_2394);
nor U4269 (N_4269,N_2534,N_466);
xnor U4270 (N_4270,N_718,N_420);
xor U4271 (N_4271,N_2642,N_266);
or U4272 (N_4272,N_105,N_144);
nand U4273 (N_4273,N_1989,N_1891);
nor U4274 (N_4274,N_2448,N_2774);
or U4275 (N_4275,N_1701,N_210);
and U4276 (N_4276,N_1854,N_143);
or U4277 (N_4277,N_2625,N_2992);
or U4278 (N_4278,N_2549,N_294);
or U4279 (N_4279,N_482,N_1229);
and U4280 (N_4280,N_502,N_1052);
nand U4281 (N_4281,N_2093,N_1545);
and U4282 (N_4282,N_2833,N_2569);
and U4283 (N_4283,N_1214,N_2315);
and U4284 (N_4284,N_720,N_1000);
and U4285 (N_4285,N_736,N_1664);
or U4286 (N_4286,N_1371,N_1716);
nand U4287 (N_4287,N_1329,N_2544);
or U4288 (N_4288,N_2539,N_145);
nor U4289 (N_4289,N_2859,N_2376);
nand U4290 (N_4290,N_2582,N_1690);
or U4291 (N_4291,N_50,N_1826);
nand U4292 (N_4292,N_2817,N_631);
xor U4293 (N_4293,N_1771,N_434);
and U4294 (N_4294,N_2618,N_2283);
and U4295 (N_4295,N_1958,N_648);
or U4296 (N_4296,N_2012,N_2802);
and U4297 (N_4297,N_2189,N_677);
or U4298 (N_4298,N_968,N_1630);
and U4299 (N_4299,N_1194,N_1710);
nor U4300 (N_4300,N_2847,N_944);
or U4301 (N_4301,N_2128,N_2687);
xnor U4302 (N_4302,N_1530,N_151);
nand U4303 (N_4303,N_479,N_2537);
nor U4304 (N_4304,N_182,N_2503);
and U4305 (N_4305,N_115,N_370);
or U4306 (N_4306,N_84,N_698);
or U4307 (N_4307,N_1715,N_1955);
nor U4308 (N_4308,N_2621,N_439);
or U4309 (N_4309,N_2592,N_2980);
xor U4310 (N_4310,N_782,N_1687);
or U4311 (N_4311,N_2746,N_778);
and U4312 (N_4312,N_1403,N_1569);
xnor U4313 (N_4313,N_1779,N_2924);
and U4314 (N_4314,N_796,N_237);
xnor U4315 (N_4315,N_470,N_2727);
nand U4316 (N_4316,N_2994,N_2930);
nand U4317 (N_4317,N_2487,N_4);
xnor U4318 (N_4318,N_1230,N_111);
or U4319 (N_4319,N_1198,N_1846);
nor U4320 (N_4320,N_1822,N_1347);
or U4321 (N_4321,N_704,N_139);
nand U4322 (N_4322,N_2111,N_1017);
nor U4323 (N_4323,N_1749,N_2881);
and U4324 (N_4324,N_2134,N_291);
xor U4325 (N_4325,N_512,N_2564);
nand U4326 (N_4326,N_1466,N_462);
or U4327 (N_4327,N_639,N_1984);
nand U4328 (N_4328,N_2443,N_290);
nor U4329 (N_4329,N_2456,N_2156);
xnor U4330 (N_4330,N_2282,N_1274);
nor U4331 (N_4331,N_1952,N_15);
nand U4332 (N_4332,N_1318,N_566);
nand U4333 (N_4333,N_1841,N_343);
and U4334 (N_4334,N_973,N_1342);
and U4335 (N_4335,N_717,N_678);
and U4336 (N_4336,N_421,N_601);
xnor U4337 (N_4337,N_2890,N_2467);
or U4338 (N_4338,N_2931,N_1190);
and U4339 (N_4339,N_1365,N_2214);
or U4340 (N_4340,N_2558,N_2368);
xnor U4341 (N_4341,N_1590,N_1420);
nand U4342 (N_4342,N_2831,N_1912);
and U4343 (N_4343,N_508,N_2327);
and U4344 (N_4344,N_2300,N_2013);
nand U4345 (N_4345,N_1535,N_1776);
nand U4346 (N_4346,N_1574,N_1439);
and U4347 (N_4347,N_1039,N_733);
xor U4348 (N_4348,N_468,N_931);
nor U4349 (N_4349,N_2144,N_2296);
or U4350 (N_4350,N_2604,N_1832);
or U4351 (N_4351,N_175,N_1750);
or U4352 (N_4352,N_1842,N_2157);
nand U4353 (N_4353,N_2066,N_1367);
nand U4354 (N_4354,N_881,N_2887);
or U4355 (N_4355,N_1976,N_1688);
xor U4356 (N_4356,N_552,N_665);
nand U4357 (N_4357,N_1556,N_2771);
xor U4358 (N_4358,N_1544,N_1619);
xor U4359 (N_4359,N_54,N_683);
or U4360 (N_4360,N_1388,N_2173);
nand U4361 (N_4361,N_2762,N_792);
and U4362 (N_4362,N_1493,N_863);
xnor U4363 (N_4363,N_2961,N_223);
nor U4364 (N_4364,N_2501,N_1331);
or U4365 (N_4365,N_1158,N_1289);
and U4366 (N_4366,N_1908,N_1510);
and U4367 (N_4367,N_2003,N_1816);
or U4368 (N_4368,N_835,N_2896);
nand U4369 (N_4369,N_273,N_1037);
and U4370 (N_4370,N_274,N_1900);
and U4371 (N_4371,N_1737,N_1307);
xnor U4372 (N_4372,N_1073,N_1860);
nand U4373 (N_4373,N_2733,N_527);
or U4374 (N_4374,N_2776,N_2262);
xor U4375 (N_4375,N_2287,N_338);
nor U4376 (N_4376,N_715,N_504);
and U4377 (N_4377,N_2680,N_1527);
nand U4378 (N_4378,N_1269,N_789);
and U4379 (N_4379,N_2129,N_820);
nand U4380 (N_4380,N_2905,N_97);
nor U4381 (N_4381,N_1924,N_1314);
xnor U4382 (N_4382,N_2205,N_1253);
and U4383 (N_4383,N_10,N_89);
nand U4384 (N_4384,N_1003,N_1564);
or U4385 (N_4385,N_1994,N_2705);
or U4386 (N_4386,N_2828,N_2637);
and U4387 (N_4387,N_1827,N_2483);
or U4388 (N_4388,N_861,N_1153);
nor U4389 (N_4389,N_2952,N_32);
nor U4390 (N_4390,N_173,N_1999);
or U4391 (N_4391,N_823,N_2630);
nor U4392 (N_4392,N_857,N_1957);
or U4393 (N_4393,N_1694,N_1514);
nand U4394 (N_4394,N_1473,N_2168);
and U4395 (N_4395,N_2396,N_1997);
nand U4396 (N_4396,N_708,N_775);
xor U4397 (N_4397,N_994,N_2672);
or U4398 (N_4398,N_2384,N_238);
and U4399 (N_4399,N_2001,N_1361);
nor U4400 (N_4400,N_1206,N_2910);
nand U4401 (N_4401,N_2290,N_2318);
or U4402 (N_4402,N_1168,N_624);
nand U4403 (N_4403,N_1748,N_915);
and U4404 (N_4404,N_349,N_854);
nor U4405 (N_4405,N_1821,N_2395);
xor U4406 (N_4406,N_1956,N_2276);
nand U4407 (N_4407,N_1177,N_990);
or U4408 (N_4408,N_2730,N_2414);
nand U4409 (N_4409,N_2284,N_2554);
or U4410 (N_4410,N_936,N_150);
or U4411 (N_4411,N_2326,N_1735);
nor U4412 (N_4412,N_1001,N_2928);
nor U4413 (N_4413,N_2080,N_2533);
and U4414 (N_4414,N_2304,N_1853);
and U4415 (N_4415,N_869,N_2477);
nand U4416 (N_4416,N_2519,N_2838);
xnor U4417 (N_4417,N_2020,N_929);
nor U4418 (N_4418,N_2369,N_1888);
xnor U4419 (N_4419,N_2845,N_655);
or U4420 (N_4420,N_2062,N_401);
nand U4421 (N_4421,N_2292,N_1786);
or U4422 (N_4422,N_958,N_750);
or U4423 (N_4423,N_805,N_1998);
nor U4424 (N_4424,N_544,N_2135);
nor U4425 (N_4425,N_1674,N_93);
nand U4426 (N_4426,N_2535,N_2159);
and U4427 (N_4427,N_2250,N_1007);
nor U4428 (N_4428,N_1973,N_2241);
xnor U4429 (N_4429,N_1870,N_578);
nor U4430 (N_4430,N_2678,N_1315);
and U4431 (N_4431,N_646,N_1899);
xor U4432 (N_4432,N_1498,N_1478);
nand U4433 (N_4433,N_289,N_1636);
nand U4434 (N_4434,N_219,N_1936);
and U4435 (N_4435,N_1663,N_1614);
xor U4436 (N_4436,N_2317,N_2462);
or U4437 (N_4437,N_976,N_147);
or U4438 (N_4438,N_1757,N_1856);
nand U4439 (N_4439,N_913,N_2906);
nand U4440 (N_4440,N_1068,N_2096);
and U4441 (N_4441,N_2388,N_88);
xnor U4442 (N_4442,N_709,N_2472);
nand U4443 (N_4443,N_2202,N_2807);
and U4444 (N_4444,N_1951,N_1125);
xnor U4445 (N_4445,N_1977,N_1078);
or U4446 (N_4446,N_483,N_1319);
or U4447 (N_4447,N_1753,N_2133);
xor U4448 (N_4448,N_2361,N_1454);
or U4449 (N_4449,N_2880,N_422);
nand U4450 (N_4450,N_1559,N_914);
nand U4451 (N_4451,N_529,N_2206);
nor U4452 (N_4452,N_2638,N_1931);
or U4453 (N_4453,N_1011,N_112);
nor U4454 (N_4454,N_2047,N_1817);
nor U4455 (N_4455,N_1350,N_1182);
nand U4456 (N_4456,N_1752,N_2252);
nor U4457 (N_4457,N_2359,N_2689);
and U4458 (N_4458,N_2675,N_124);
and U4459 (N_4459,N_1186,N_1609);
xnor U4460 (N_4460,N_2102,N_1172);
xnor U4461 (N_4461,N_2567,N_418);
xor U4462 (N_4462,N_1293,N_1772);
nand U4463 (N_4463,N_1561,N_1056);
xnor U4464 (N_4464,N_930,N_82);
xnor U4465 (N_4465,N_1719,N_2240);
and U4466 (N_4466,N_2086,N_1857);
and U4467 (N_4467,N_2217,N_2884);
or U4468 (N_4468,N_1819,N_2583);
xor U4469 (N_4469,N_1985,N_2146);
nand U4470 (N_4470,N_2698,N_485);
nor U4471 (N_4471,N_2875,N_1283);
nand U4472 (N_4472,N_1809,N_2851);
xor U4473 (N_4473,N_1709,N_783);
and U4474 (N_4474,N_1450,N_817);
xnor U4475 (N_4475,N_1313,N_942);
and U4476 (N_4476,N_2127,N_804);
xor U4477 (N_4477,N_2273,N_2876);
nand U4478 (N_4478,N_2375,N_68);
nor U4479 (N_4479,N_1568,N_2336);
nand U4480 (N_4480,N_1596,N_1909);
nor U4481 (N_4481,N_1496,N_2196);
nand U4482 (N_4482,N_1139,N_2628);
xnor U4483 (N_4483,N_2547,N_845);
nand U4484 (N_4484,N_1445,N_2570);
or U4485 (N_4485,N_2907,N_2243);
nand U4486 (N_4486,N_1427,N_675);
xor U4487 (N_4487,N_2431,N_270);
nor U4488 (N_4488,N_1183,N_195);
xnor U4489 (N_4489,N_2684,N_76);
and U4490 (N_4490,N_1552,N_790);
nand U4491 (N_4491,N_367,N_701);
xnor U4492 (N_4492,N_2330,N_368);
nor U4493 (N_4493,N_2297,N_2999);
nand U4494 (N_4494,N_1255,N_377);
xor U4495 (N_4495,N_1398,N_2911);
xnor U4496 (N_4496,N_813,N_2488);
nor U4497 (N_4497,N_1622,N_2335);
nor U4498 (N_4498,N_516,N_608);
and U4499 (N_4499,N_781,N_1618);
and U4500 (N_4500,N_2274,N_2022);
and U4501 (N_4501,N_2153,N_675);
and U4502 (N_4502,N_1654,N_30);
and U4503 (N_4503,N_2613,N_2934);
xnor U4504 (N_4504,N_965,N_2273);
xnor U4505 (N_4505,N_99,N_156);
xor U4506 (N_4506,N_2649,N_1430);
or U4507 (N_4507,N_1909,N_562);
nor U4508 (N_4508,N_525,N_1141);
nor U4509 (N_4509,N_2234,N_1172);
and U4510 (N_4510,N_1426,N_2961);
nor U4511 (N_4511,N_898,N_2346);
and U4512 (N_4512,N_1285,N_1710);
xor U4513 (N_4513,N_332,N_1121);
nor U4514 (N_4514,N_1551,N_726);
and U4515 (N_4515,N_952,N_2211);
xnor U4516 (N_4516,N_164,N_973);
and U4517 (N_4517,N_1418,N_686);
nand U4518 (N_4518,N_1854,N_45);
or U4519 (N_4519,N_1013,N_424);
nand U4520 (N_4520,N_1413,N_2062);
or U4521 (N_4521,N_2165,N_1120);
and U4522 (N_4522,N_1331,N_1814);
nand U4523 (N_4523,N_2844,N_357);
nand U4524 (N_4524,N_2623,N_2084);
and U4525 (N_4525,N_809,N_188);
nor U4526 (N_4526,N_940,N_761);
or U4527 (N_4527,N_164,N_159);
nor U4528 (N_4528,N_2046,N_2189);
nand U4529 (N_4529,N_2591,N_1090);
and U4530 (N_4530,N_2063,N_2084);
xor U4531 (N_4531,N_1972,N_1197);
or U4532 (N_4532,N_459,N_129);
nor U4533 (N_4533,N_1799,N_1064);
xnor U4534 (N_4534,N_2992,N_43);
and U4535 (N_4535,N_2730,N_639);
xor U4536 (N_4536,N_2475,N_1501);
nand U4537 (N_4537,N_425,N_1244);
xor U4538 (N_4538,N_1886,N_572);
nand U4539 (N_4539,N_506,N_2203);
xnor U4540 (N_4540,N_563,N_100);
and U4541 (N_4541,N_1343,N_728);
xnor U4542 (N_4542,N_1408,N_39);
or U4543 (N_4543,N_335,N_592);
or U4544 (N_4544,N_2805,N_1156);
and U4545 (N_4545,N_123,N_1911);
nor U4546 (N_4546,N_2599,N_1538);
nor U4547 (N_4547,N_1567,N_805);
nand U4548 (N_4548,N_1801,N_211);
or U4549 (N_4549,N_2221,N_1619);
and U4550 (N_4550,N_346,N_2062);
nor U4551 (N_4551,N_2344,N_1866);
or U4552 (N_4552,N_260,N_2432);
xnor U4553 (N_4553,N_942,N_2049);
and U4554 (N_4554,N_2466,N_2352);
xor U4555 (N_4555,N_2626,N_2509);
nand U4556 (N_4556,N_2450,N_2416);
or U4557 (N_4557,N_349,N_2020);
nor U4558 (N_4558,N_2164,N_2178);
and U4559 (N_4559,N_375,N_2114);
nand U4560 (N_4560,N_53,N_2454);
and U4561 (N_4561,N_338,N_1450);
or U4562 (N_4562,N_1190,N_2259);
nand U4563 (N_4563,N_258,N_1503);
nor U4564 (N_4564,N_2603,N_1430);
xor U4565 (N_4565,N_2831,N_2869);
nand U4566 (N_4566,N_749,N_986);
nor U4567 (N_4567,N_1077,N_2501);
and U4568 (N_4568,N_215,N_1413);
nor U4569 (N_4569,N_52,N_1870);
or U4570 (N_4570,N_511,N_870);
or U4571 (N_4571,N_2667,N_1754);
and U4572 (N_4572,N_1447,N_2623);
nor U4573 (N_4573,N_1598,N_1970);
xor U4574 (N_4574,N_1349,N_1906);
nor U4575 (N_4575,N_1493,N_95);
or U4576 (N_4576,N_2197,N_1488);
xor U4577 (N_4577,N_2705,N_2362);
nand U4578 (N_4578,N_1424,N_2734);
xnor U4579 (N_4579,N_1933,N_2904);
and U4580 (N_4580,N_2337,N_1836);
and U4581 (N_4581,N_730,N_6);
xor U4582 (N_4582,N_1403,N_1787);
xnor U4583 (N_4583,N_1989,N_1472);
and U4584 (N_4584,N_1598,N_1681);
or U4585 (N_4585,N_2052,N_939);
or U4586 (N_4586,N_292,N_696);
xnor U4587 (N_4587,N_2454,N_939);
and U4588 (N_4588,N_1099,N_494);
nor U4589 (N_4589,N_2242,N_294);
and U4590 (N_4590,N_901,N_269);
nor U4591 (N_4591,N_2197,N_2277);
and U4592 (N_4592,N_2020,N_1283);
xor U4593 (N_4593,N_2025,N_2990);
nor U4594 (N_4594,N_802,N_2682);
nand U4595 (N_4595,N_2022,N_1201);
or U4596 (N_4596,N_2248,N_447);
and U4597 (N_4597,N_1207,N_189);
nor U4598 (N_4598,N_1316,N_1371);
and U4599 (N_4599,N_2836,N_541);
nor U4600 (N_4600,N_899,N_720);
xnor U4601 (N_4601,N_1442,N_1890);
nor U4602 (N_4602,N_293,N_2052);
nand U4603 (N_4603,N_2645,N_2307);
nor U4604 (N_4604,N_964,N_2167);
xor U4605 (N_4605,N_141,N_1842);
nor U4606 (N_4606,N_2052,N_438);
nand U4607 (N_4607,N_174,N_1141);
xor U4608 (N_4608,N_1057,N_463);
and U4609 (N_4609,N_2950,N_1562);
nand U4610 (N_4610,N_1455,N_1842);
xnor U4611 (N_4611,N_617,N_1357);
and U4612 (N_4612,N_1584,N_2487);
or U4613 (N_4613,N_1657,N_519);
and U4614 (N_4614,N_148,N_1230);
nor U4615 (N_4615,N_1581,N_707);
and U4616 (N_4616,N_2431,N_433);
or U4617 (N_4617,N_763,N_679);
or U4618 (N_4618,N_1857,N_2951);
nand U4619 (N_4619,N_1391,N_1121);
xnor U4620 (N_4620,N_2295,N_1569);
nand U4621 (N_4621,N_789,N_2864);
xnor U4622 (N_4622,N_2355,N_871);
xor U4623 (N_4623,N_2292,N_303);
xor U4624 (N_4624,N_2440,N_2588);
nor U4625 (N_4625,N_2293,N_2399);
xor U4626 (N_4626,N_993,N_2749);
nor U4627 (N_4627,N_2872,N_531);
nor U4628 (N_4628,N_1481,N_1999);
nor U4629 (N_4629,N_1110,N_219);
xnor U4630 (N_4630,N_2344,N_2658);
and U4631 (N_4631,N_1892,N_535);
nor U4632 (N_4632,N_893,N_1632);
xnor U4633 (N_4633,N_2885,N_534);
or U4634 (N_4634,N_2004,N_2849);
nand U4635 (N_4635,N_350,N_771);
or U4636 (N_4636,N_1747,N_1836);
or U4637 (N_4637,N_2963,N_718);
or U4638 (N_4638,N_2127,N_2345);
and U4639 (N_4639,N_2325,N_1355);
xor U4640 (N_4640,N_103,N_379);
nor U4641 (N_4641,N_338,N_2112);
xnor U4642 (N_4642,N_2375,N_1706);
or U4643 (N_4643,N_2624,N_737);
nor U4644 (N_4644,N_827,N_1649);
nand U4645 (N_4645,N_165,N_1197);
nor U4646 (N_4646,N_1501,N_2423);
xor U4647 (N_4647,N_1741,N_471);
xor U4648 (N_4648,N_799,N_2880);
xor U4649 (N_4649,N_309,N_222);
nand U4650 (N_4650,N_1197,N_1062);
nor U4651 (N_4651,N_320,N_258);
xnor U4652 (N_4652,N_792,N_473);
or U4653 (N_4653,N_363,N_2097);
nand U4654 (N_4654,N_1960,N_1821);
nand U4655 (N_4655,N_1070,N_2498);
nand U4656 (N_4656,N_2398,N_2965);
nor U4657 (N_4657,N_711,N_2461);
and U4658 (N_4658,N_527,N_1557);
and U4659 (N_4659,N_288,N_2960);
nand U4660 (N_4660,N_2397,N_741);
xnor U4661 (N_4661,N_1795,N_1059);
nand U4662 (N_4662,N_1007,N_1024);
nor U4663 (N_4663,N_2789,N_1081);
or U4664 (N_4664,N_1198,N_817);
nor U4665 (N_4665,N_2608,N_2434);
xnor U4666 (N_4666,N_416,N_1050);
and U4667 (N_4667,N_923,N_604);
nand U4668 (N_4668,N_1310,N_2858);
xnor U4669 (N_4669,N_1982,N_283);
xnor U4670 (N_4670,N_1084,N_1750);
nand U4671 (N_4671,N_903,N_88);
or U4672 (N_4672,N_1059,N_929);
and U4673 (N_4673,N_86,N_1773);
and U4674 (N_4674,N_1913,N_996);
and U4675 (N_4675,N_2895,N_2922);
xor U4676 (N_4676,N_2352,N_2428);
or U4677 (N_4677,N_1570,N_1588);
nand U4678 (N_4678,N_1558,N_1088);
nand U4679 (N_4679,N_219,N_2605);
nor U4680 (N_4680,N_2819,N_2510);
nand U4681 (N_4681,N_1486,N_2086);
nor U4682 (N_4682,N_342,N_2199);
or U4683 (N_4683,N_1508,N_2180);
and U4684 (N_4684,N_929,N_793);
nor U4685 (N_4685,N_2248,N_765);
and U4686 (N_4686,N_2157,N_2952);
xor U4687 (N_4687,N_1037,N_2339);
and U4688 (N_4688,N_2501,N_78);
xor U4689 (N_4689,N_1263,N_1852);
or U4690 (N_4690,N_1556,N_754);
or U4691 (N_4691,N_2617,N_2549);
or U4692 (N_4692,N_1854,N_813);
nor U4693 (N_4693,N_1112,N_2078);
nand U4694 (N_4694,N_2106,N_1993);
nor U4695 (N_4695,N_1991,N_1037);
or U4696 (N_4696,N_874,N_1864);
nor U4697 (N_4697,N_186,N_1734);
and U4698 (N_4698,N_2576,N_336);
and U4699 (N_4699,N_1154,N_678);
nor U4700 (N_4700,N_962,N_1731);
and U4701 (N_4701,N_1861,N_217);
and U4702 (N_4702,N_2391,N_1545);
nor U4703 (N_4703,N_2529,N_2035);
nand U4704 (N_4704,N_961,N_1230);
and U4705 (N_4705,N_1837,N_1985);
nand U4706 (N_4706,N_2428,N_2636);
nor U4707 (N_4707,N_265,N_901);
or U4708 (N_4708,N_2389,N_540);
or U4709 (N_4709,N_519,N_1020);
nor U4710 (N_4710,N_1452,N_1153);
or U4711 (N_4711,N_1952,N_1686);
and U4712 (N_4712,N_1139,N_2680);
nor U4713 (N_4713,N_909,N_2247);
or U4714 (N_4714,N_1682,N_2079);
xor U4715 (N_4715,N_1846,N_326);
or U4716 (N_4716,N_1517,N_1246);
or U4717 (N_4717,N_1487,N_2957);
xor U4718 (N_4718,N_826,N_2860);
or U4719 (N_4719,N_1139,N_1643);
nor U4720 (N_4720,N_664,N_2530);
or U4721 (N_4721,N_1676,N_637);
or U4722 (N_4722,N_2672,N_943);
nor U4723 (N_4723,N_1202,N_1400);
nand U4724 (N_4724,N_954,N_313);
and U4725 (N_4725,N_1095,N_2917);
or U4726 (N_4726,N_586,N_2404);
xor U4727 (N_4727,N_1965,N_1050);
and U4728 (N_4728,N_130,N_2875);
nor U4729 (N_4729,N_46,N_336);
nor U4730 (N_4730,N_2242,N_642);
xor U4731 (N_4731,N_1837,N_2091);
and U4732 (N_4732,N_423,N_2987);
nor U4733 (N_4733,N_977,N_1620);
and U4734 (N_4734,N_43,N_28);
nor U4735 (N_4735,N_65,N_2938);
or U4736 (N_4736,N_756,N_978);
xor U4737 (N_4737,N_1297,N_1154);
and U4738 (N_4738,N_718,N_2449);
nor U4739 (N_4739,N_570,N_1481);
and U4740 (N_4740,N_2657,N_2626);
nor U4741 (N_4741,N_313,N_1229);
or U4742 (N_4742,N_1217,N_2419);
xnor U4743 (N_4743,N_2812,N_427);
or U4744 (N_4744,N_2486,N_2861);
nor U4745 (N_4745,N_1585,N_1568);
nand U4746 (N_4746,N_849,N_2477);
nand U4747 (N_4747,N_2652,N_2921);
nand U4748 (N_4748,N_2231,N_1596);
xor U4749 (N_4749,N_2455,N_515);
and U4750 (N_4750,N_360,N_1375);
nor U4751 (N_4751,N_887,N_298);
nand U4752 (N_4752,N_1629,N_2273);
nor U4753 (N_4753,N_2619,N_469);
and U4754 (N_4754,N_1723,N_2425);
nor U4755 (N_4755,N_1001,N_2782);
nor U4756 (N_4756,N_145,N_278);
nor U4757 (N_4757,N_321,N_645);
nand U4758 (N_4758,N_745,N_2485);
or U4759 (N_4759,N_2664,N_70);
and U4760 (N_4760,N_1604,N_1729);
and U4761 (N_4761,N_113,N_1908);
nor U4762 (N_4762,N_279,N_2029);
xor U4763 (N_4763,N_2703,N_2643);
xor U4764 (N_4764,N_875,N_1359);
xnor U4765 (N_4765,N_2818,N_2055);
and U4766 (N_4766,N_2383,N_2386);
xnor U4767 (N_4767,N_2832,N_1939);
nand U4768 (N_4768,N_1330,N_2386);
nor U4769 (N_4769,N_1838,N_2054);
or U4770 (N_4770,N_1640,N_2815);
and U4771 (N_4771,N_1472,N_461);
nor U4772 (N_4772,N_892,N_0);
and U4773 (N_4773,N_572,N_936);
xnor U4774 (N_4774,N_2173,N_850);
nor U4775 (N_4775,N_1100,N_1533);
nor U4776 (N_4776,N_1837,N_1474);
or U4777 (N_4777,N_1710,N_1294);
nand U4778 (N_4778,N_2328,N_1842);
xor U4779 (N_4779,N_136,N_94);
or U4780 (N_4780,N_1057,N_12);
nand U4781 (N_4781,N_2787,N_452);
nand U4782 (N_4782,N_1637,N_2642);
nand U4783 (N_4783,N_2882,N_685);
or U4784 (N_4784,N_523,N_1040);
xor U4785 (N_4785,N_2880,N_770);
or U4786 (N_4786,N_2072,N_1855);
xor U4787 (N_4787,N_898,N_779);
and U4788 (N_4788,N_608,N_2859);
and U4789 (N_4789,N_771,N_2139);
or U4790 (N_4790,N_272,N_1627);
nand U4791 (N_4791,N_2010,N_1262);
nand U4792 (N_4792,N_545,N_2238);
nor U4793 (N_4793,N_1715,N_654);
nor U4794 (N_4794,N_2965,N_1294);
and U4795 (N_4795,N_2775,N_190);
nand U4796 (N_4796,N_474,N_1083);
and U4797 (N_4797,N_307,N_1396);
xor U4798 (N_4798,N_1694,N_1834);
and U4799 (N_4799,N_985,N_448);
or U4800 (N_4800,N_653,N_208);
and U4801 (N_4801,N_536,N_1496);
and U4802 (N_4802,N_1981,N_2959);
or U4803 (N_4803,N_2137,N_1434);
and U4804 (N_4804,N_1978,N_272);
nand U4805 (N_4805,N_2221,N_430);
or U4806 (N_4806,N_1816,N_1843);
xnor U4807 (N_4807,N_994,N_593);
and U4808 (N_4808,N_2080,N_2168);
nor U4809 (N_4809,N_580,N_2891);
nor U4810 (N_4810,N_2852,N_1149);
nand U4811 (N_4811,N_1851,N_2935);
nor U4812 (N_4812,N_1350,N_1261);
xor U4813 (N_4813,N_2958,N_2033);
nor U4814 (N_4814,N_1581,N_1585);
nand U4815 (N_4815,N_611,N_2484);
or U4816 (N_4816,N_2471,N_246);
nand U4817 (N_4817,N_1877,N_2186);
nand U4818 (N_4818,N_1372,N_2333);
or U4819 (N_4819,N_1917,N_1160);
or U4820 (N_4820,N_1600,N_2175);
or U4821 (N_4821,N_335,N_2465);
nand U4822 (N_4822,N_32,N_183);
or U4823 (N_4823,N_562,N_396);
or U4824 (N_4824,N_2599,N_2645);
and U4825 (N_4825,N_2798,N_2950);
or U4826 (N_4826,N_2849,N_578);
or U4827 (N_4827,N_1644,N_2749);
nor U4828 (N_4828,N_2364,N_2697);
xnor U4829 (N_4829,N_2991,N_333);
and U4830 (N_4830,N_1376,N_2707);
nand U4831 (N_4831,N_338,N_1928);
nand U4832 (N_4832,N_2710,N_2892);
and U4833 (N_4833,N_1182,N_471);
and U4834 (N_4834,N_2147,N_1878);
nand U4835 (N_4835,N_208,N_182);
xor U4836 (N_4836,N_2710,N_634);
nand U4837 (N_4837,N_1185,N_877);
xnor U4838 (N_4838,N_471,N_846);
nor U4839 (N_4839,N_2441,N_2762);
or U4840 (N_4840,N_2287,N_1523);
nand U4841 (N_4841,N_1543,N_2455);
nand U4842 (N_4842,N_416,N_1768);
nand U4843 (N_4843,N_630,N_389);
xnor U4844 (N_4844,N_123,N_1203);
and U4845 (N_4845,N_2815,N_2536);
and U4846 (N_4846,N_1537,N_151);
nor U4847 (N_4847,N_2788,N_2305);
xnor U4848 (N_4848,N_103,N_2742);
nand U4849 (N_4849,N_1662,N_888);
and U4850 (N_4850,N_1133,N_1356);
nand U4851 (N_4851,N_2795,N_2969);
nor U4852 (N_4852,N_1401,N_2982);
nor U4853 (N_4853,N_2302,N_665);
xor U4854 (N_4854,N_855,N_2829);
or U4855 (N_4855,N_580,N_2932);
nand U4856 (N_4856,N_2794,N_652);
nand U4857 (N_4857,N_2272,N_1937);
xnor U4858 (N_4858,N_1660,N_1255);
xor U4859 (N_4859,N_1395,N_1332);
nor U4860 (N_4860,N_2339,N_2552);
or U4861 (N_4861,N_1041,N_2546);
nand U4862 (N_4862,N_2675,N_1339);
and U4863 (N_4863,N_1080,N_306);
or U4864 (N_4864,N_214,N_352);
or U4865 (N_4865,N_1906,N_1286);
nand U4866 (N_4866,N_405,N_2748);
nand U4867 (N_4867,N_1067,N_726);
nor U4868 (N_4868,N_203,N_2561);
and U4869 (N_4869,N_1892,N_1015);
or U4870 (N_4870,N_1727,N_314);
nand U4871 (N_4871,N_2553,N_1095);
and U4872 (N_4872,N_2907,N_2055);
nand U4873 (N_4873,N_2678,N_2759);
nor U4874 (N_4874,N_2321,N_1768);
nand U4875 (N_4875,N_2427,N_443);
and U4876 (N_4876,N_2306,N_781);
or U4877 (N_4877,N_782,N_536);
or U4878 (N_4878,N_2622,N_2245);
xor U4879 (N_4879,N_1573,N_2569);
xor U4880 (N_4880,N_1910,N_1136);
nand U4881 (N_4881,N_310,N_2513);
and U4882 (N_4882,N_2017,N_1411);
xor U4883 (N_4883,N_1823,N_2905);
or U4884 (N_4884,N_486,N_9);
and U4885 (N_4885,N_2948,N_233);
xnor U4886 (N_4886,N_2272,N_1135);
xnor U4887 (N_4887,N_2011,N_2519);
nor U4888 (N_4888,N_2231,N_331);
and U4889 (N_4889,N_814,N_827);
nor U4890 (N_4890,N_1565,N_1683);
nand U4891 (N_4891,N_2673,N_1320);
nor U4892 (N_4892,N_733,N_2867);
or U4893 (N_4893,N_407,N_763);
nor U4894 (N_4894,N_2841,N_2315);
or U4895 (N_4895,N_253,N_2972);
and U4896 (N_4896,N_927,N_691);
and U4897 (N_4897,N_1621,N_1133);
nor U4898 (N_4898,N_1446,N_1648);
nand U4899 (N_4899,N_2296,N_1190);
or U4900 (N_4900,N_992,N_1182);
nand U4901 (N_4901,N_1657,N_1993);
nor U4902 (N_4902,N_1166,N_1542);
xnor U4903 (N_4903,N_2731,N_2641);
or U4904 (N_4904,N_918,N_2543);
or U4905 (N_4905,N_2940,N_365);
and U4906 (N_4906,N_988,N_506);
xor U4907 (N_4907,N_1104,N_960);
or U4908 (N_4908,N_2835,N_1772);
or U4909 (N_4909,N_148,N_130);
or U4910 (N_4910,N_361,N_2290);
and U4911 (N_4911,N_1983,N_335);
xnor U4912 (N_4912,N_1407,N_2622);
xnor U4913 (N_4913,N_2158,N_791);
nor U4914 (N_4914,N_616,N_2525);
nand U4915 (N_4915,N_2413,N_909);
xor U4916 (N_4916,N_2398,N_536);
or U4917 (N_4917,N_20,N_1370);
nor U4918 (N_4918,N_2424,N_702);
nor U4919 (N_4919,N_2628,N_2240);
nor U4920 (N_4920,N_2710,N_1417);
nand U4921 (N_4921,N_1032,N_2878);
and U4922 (N_4922,N_2019,N_622);
xnor U4923 (N_4923,N_2798,N_315);
nor U4924 (N_4924,N_2652,N_2624);
or U4925 (N_4925,N_890,N_180);
nor U4926 (N_4926,N_1730,N_694);
nand U4927 (N_4927,N_1439,N_2063);
or U4928 (N_4928,N_556,N_602);
nand U4929 (N_4929,N_1043,N_2157);
nor U4930 (N_4930,N_1657,N_556);
xnor U4931 (N_4931,N_2838,N_1818);
nand U4932 (N_4932,N_21,N_1635);
and U4933 (N_4933,N_2696,N_2056);
and U4934 (N_4934,N_626,N_2754);
nor U4935 (N_4935,N_2503,N_2818);
and U4936 (N_4936,N_1013,N_704);
or U4937 (N_4937,N_1812,N_815);
nand U4938 (N_4938,N_2948,N_1358);
nor U4939 (N_4939,N_63,N_2392);
nor U4940 (N_4940,N_1142,N_1176);
or U4941 (N_4941,N_335,N_1943);
nor U4942 (N_4942,N_1614,N_596);
nor U4943 (N_4943,N_2017,N_2419);
xnor U4944 (N_4944,N_567,N_1976);
or U4945 (N_4945,N_2541,N_253);
nand U4946 (N_4946,N_750,N_2763);
nor U4947 (N_4947,N_719,N_1524);
and U4948 (N_4948,N_1913,N_1584);
nor U4949 (N_4949,N_1186,N_2751);
xnor U4950 (N_4950,N_1612,N_1101);
or U4951 (N_4951,N_2127,N_1659);
or U4952 (N_4952,N_1619,N_1565);
nor U4953 (N_4953,N_1633,N_2916);
xnor U4954 (N_4954,N_99,N_2937);
nor U4955 (N_4955,N_197,N_974);
nand U4956 (N_4956,N_2702,N_1366);
nand U4957 (N_4957,N_1477,N_908);
nand U4958 (N_4958,N_1930,N_1299);
nand U4959 (N_4959,N_1151,N_983);
or U4960 (N_4960,N_2069,N_2606);
nor U4961 (N_4961,N_533,N_843);
nor U4962 (N_4962,N_2701,N_434);
nor U4963 (N_4963,N_421,N_2051);
nand U4964 (N_4964,N_759,N_1549);
nand U4965 (N_4965,N_2454,N_463);
and U4966 (N_4966,N_1526,N_1865);
xor U4967 (N_4967,N_2658,N_1002);
nor U4968 (N_4968,N_105,N_2021);
and U4969 (N_4969,N_293,N_1227);
nand U4970 (N_4970,N_440,N_2225);
nand U4971 (N_4971,N_1394,N_1180);
nor U4972 (N_4972,N_2217,N_1891);
or U4973 (N_4973,N_2081,N_2603);
and U4974 (N_4974,N_851,N_409);
nor U4975 (N_4975,N_456,N_994);
nand U4976 (N_4976,N_1885,N_2813);
nor U4977 (N_4977,N_2270,N_430);
or U4978 (N_4978,N_116,N_73);
or U4979 (N_4979,N_2412,N_2301);
and U4980 (N_4980,N_342,N_2571);
and U4981 (N_4981,N_2858,N_1460);
and U4982 (N_4982,N_2587,N_1880);
nand U4983 (N_4983,N_2554,N_2329);
and U4984 (N_4984,N_2938,N_152);
nand U4985 (N_4985,N_2611,N_2943);
or U4986 (N_4986,N_2514,N_2850);
nor U4987 (N_4987,N_192,N_735);
or U4988 (N_4988,N_881,N_290);
or U4989 (N_4989,N_2184,N_2520);
nand U4990 (N_4990,N_25,N_544);
xor U4991 (N_4991,N_2134,N_1103);
nand U4992 (N_4992,N_2014,N_2298);
nor U4993 (N_4993,N_453,N_1458);
nand U4994 (N_4994,N_75,N_557);
and U4995 (N_4995,N_1983,N_1974);
nand U4996 (N_4996,N_2083,N_762);
xor U4997 (N_4997,N_2341,N_2541);
xnor U4998 (N_4998,N_398,N_1389);
nand U4999 (N_4999,N_1294,N_1141);
nor U5000 (N_5000,N_2480,N_987);
nor U5001 (N_5001,N_574,N_2507);
or U5002 (N_5002,N_562,N_1224);
or U5003 (N_5003,N_212,N_2151);
nor U5004 (N_5004,N_938,N_89);
nor U5005 (N_5005,N_2320,N_927);
xor U5006 (N_5006,N_1479,N_1309);
and U5007 (N_5007,N_2436,N_2600);
nor U5008 (N_5008,N_761,N_2818);
and U5009 (N_5009,N_2369,N_2741);
nand U5010 (N_5010,N_2623,N_221);
nor U5011 (N_5011,N_2212,N_573);
nand U5012 (N_5012,N_973,N_1305);
nand U5013 (N_5013,N_1512,N_1075);
xnor U5014 (N_5014,N_1650,N_1858);
or U5015 (N_5015,N_2025,N_1335);
xor U5016 (N_5016,N_1159,N_2201);
nor U5017 (N_5017,N_2428,N_1308);
and U5018 (N_5018,N_524,N_1373);
nor U5019 (N_5019,N_1991,N_2585);
nor U5020 (N_5020,N_217,N_2689);
nand U5021 (N_5021,N_2486,N_1053);
nand U5022 (N_5022,N_2288,N_1079);
and U5023 (N_5023,N_326,N_1210);
and U5024 (N_5024,N_2025,N_1451);
or U5025 (N_5025,N_2816,N_2396);
nor U5026 (N_5026,N_2163,N_677);
xnor U5027 (N_5027,N_624,N_2239);
nor U5028 (N_5028,N_200,N_1385);
xnor U5029 (N_5029,N_2487,N_2916);
xor U5030 (N_5030,N_404,N_1074);
and U5031 (N_5031,N_431,N_2836);
or U5032 (N_5032,N_2320,N_850);
and U5033 (N_5033,N_2610,N_296);
nor U5034 (N_5034,N_1669,N_392);
and U5035 (N_5035,N_1504,N_2701);
xnor U5036 (N_5036,N_1695,N_2508);
xnor U5037 (N_5037,N_877,N_2387);
xnor U5038 (N_5038,N_647,N_1583);
nand U5039 (N_5039,N_360,N_1170);
or U5040 (N_5040,N_1062,N_882);
nand U5041 (N_5041,N_1839,N_1167);
and U5042 (N_5042,N_660,N_2256);
nand U5043 (N_5043,N_2767,N_2402);
xor U5044 (N_5044,N_1186,N_1251);
or U5045 (N_5045,N_1543,N_2146);
xor U5046 (N_5046,N_343,N_1417);
nand U5047 (N_5047,N_2812,N_2162);
xor U5048 (N_5048,N_733,N_722);
or U5049 (N_5049,N_1676,N_2959);
nand U5050 (N_5050,N_2349,N_1215);
and U5051 (N_5051,N_495,N_105);
or U5052 (N_5052,N_312,N_1760);
or U5053 (N_5053,N_464,N_1493);
xor U5054 (N_5054,N_261,N_2333);
xor U5055 (N_5055,N_271,N_2573);
xnor U5056 (N_5056,N_142,N_2760);
nor U5057 (N_5057,N_2800,N_1481);
xor U5058 (N_5058,N_989,N_2213);
nand U5059 (N_5059,N_1300,N_578);
nand U5060 (N_5060,N_1612,N_1073);
xor U5061 (N_5061,N_2271,N_98);
nor U5062 (N_5062,N_2874,N_1595);
xor U5063 (N_5063,N_152,N_800);
nand U5064 (N_5064,N_2620,N_2548);
nand U5065 (N_5065,N_2776,N_448);
nand U5066 (N_5066,N_257,N_2202);
or U5067 (N_5067,N_169,N_468);
and U5068 (N_5068,N_215,N_83);
or U5069 (N_5069,N_264,N_1725);
nand U5070 (N_5070,N_572,N_2280);
nand U5071 (N_5071,N_855,N_1980);
and U5072 (N_5072,N_1889,N_2713);
or U5073 (N_5073,N_2557,N_2379);
nor U5074 (N_5074,N_664,N_1920);
nand U5075 (N_5075,N_2734,N_1945);
and U5076 (N_5076,N_164,N_2461);
nand U5077 (N_5077,N_1840,N_79);
nand U5078 (N_5078,N_1541,N_1396);
xnor U5079 (N_5079,N_2853,N_1372);
or U5080 (N_5080,N_2419,N_2463);
or U5081 (N_5081,N_744,N_2307);
nor U5082 (N_5082,N_1100,N_1654);
nand U5083 (N_5083,N_1806,N_2954);
and U5084 (N_5084,N_120,N_2710);
nor U5085 (N_5085,N_442,N_1672);
nor U5086 (N_5086,N_2842,N_2336);
xor U5087 (N_5087,N_1964,N_2440);
nand U5088 (N_5088,N_1676,N_357);
xor U5089 (N_5089,N_879,N_1310);
nor U5090 (N_5090,N_1550,N_2357);
xor U5091 (N_5091,N_2436,N_533);
xor U5092 (N_5092,N_2932,N_2111);
nor U5093 (N_5093,N_117,N_2700);
xnor U5094 (N_5094,N_443,N_758);
nor U5095 (N_5095,N_471,N_914);
nor U5096 (N_5096,N_1962,N_546);
xnor U5097 (N_5097,N_1919,N_143);
nand U5098 (N_5098,N_1315,N_2958);
nor U5099 (N_5099,N_743,N_18);
and U5100 (N_5100,N_1939,N_230);
nor U5101 (N_5101,N_1964,N_1129);
or U5102 (N_5102,N_40,N_1900);
nor U5103 (N_5103,N_27,N_937);
and U5104 (N_5104,N_1955,N_1568);
or U5105 (N_5105,N_2251,N_752);
xor U5106 (N_5106,N_1431,N_1651);
nand U5107 (N_5107,N_720,N_2664);
or U5108 (N_5108,N_316,N_2394);
nor U5109 (N_5109,N_766,N_2150);
nor U5110 (N_5110,N_108,N_1668);
and U5111 (N_5111,N_1843,N_2389);
or U5112 (N_5112,N_2607,N_1493);
or U5113 (N_5113,N_1577,N_717);
nor U5114 (N_5114,N_979,N_1739);
nor U5115 (N_5115,N_1941,N_2850);
and U5116 (N_5116,N_2487,N_320);
nand U5117 (N_5117,N_1315,N_505);
or U5118 (N_5118,N_2242,N_2756);
and U5119 (N_5119,N_1006,N_2500);
nor U5120 (N_5120,N_1833,N_2566);
xnor U5121 (N_5121,N_2092,N_2244);
or U5122 (N_5122,N_1350,N_1316);
xnor U5123 (N_5123,N_2282,N_535);
xnor U5124 (N_5124,N_1242,N_2066);
or U5125 (N_5125,N_1271,N_1793);
or U5126 (N_5126,N_2799,N_2290);
nand U5127 (N_5127,N_1191,N_88);
or U5128 (N_5128,N_2605,N_2899);
nand U5129 (N_5129,N_1434,N_1061);
and U5130 (N_5130,N_1703,N_530);
nor U5131 (N_5131,N_145,N_108);
nand U5132 (N_5132,N_1077,N_1561);
nand U5133 (N_5133,N_954,N_1467);
xor U5134 (N_5134,N_2479,N_914);
nor U5135 (N_5135,N_1872,N_2215);
xor U5136 (N_5136,N_1176,N_339);
nor U5137 (N_5137,N_2475,N_2973);
xnor U5138 (N_5138,N_2119,N_858);
xor U5139 (N_5139,N_2726,N_2984);
nand U5140 (N_5140,N_1195,N_379);
xnor U5141 (N_5141,N_490,N_1162);
nand U5142 (N_5142,N_2544,N_2460);
or U5143 (N_5143,N_1495,N_1084);
or U5144 (N_5144,N_2259,N_1161);
and U5145 (N_5145,N_1315,N_237);
or U5146 (N_5146,N_1338,N_393);
nor U5147 (N_5147,N_2173,N_2473);
nor U5148 (N_5148,N_1971,N_1599);
nor U5149 (N_5149,N_1486,N_1339);
nand U5150 (N_5150,N_2974,N_2190);
xor U5151 (N_5151,N_1561,N_1587);
and U5152 (N_5152,N_473,N_1059);
nor U5153 (N_5153,N_1329,N_2086);
and U5154 (N_5154,N_554,N_1048);
nor U5155 (N_5155,N_2774,N_760);
or U5156 (N_5156,N_289,N_2618);
or U5157 (N_5157,N_2731,N_1264);
nor U5158 (N_5158,N_2120,N_44);
or U5159 (N_5159,N_2773,N_2226);
and U5160 (N_5160,N_1580,N_413);
and U5161 (N_5161,N_2380,N_938);
and U5162 (N_5162,N_1935,N_2000);
or U5163 (N_5163,N_2896,N_1322);
and U5164 (N_5164,N_2059,N_1874);
xnor U5165 (N_5165,N_2387,N_2023);
and U5166 (N_5166,N_1508,N_966);
xor U5167 (N_5167,N_1677,N_1487);
xnor U5168 (N_5168,N_775,N_1106);
xnor U5169 (N_5169,N_2096,N_2146);
nand U5170 (N_5170,N_2419,N_2415);
and U5171 (N_5171,N_1063,N_2972);
and U5172 (N_5172,N_1717,N_308);
xor U5173 (N_5173,N_1848,N_8);
nand U5174 (N_5174,N_533,N_1318);
and U5175 (N_5175,N_2582,N_1625);
nand U5176 (N_5176,N_2873,N_688);
nor U5177 (N_5177,N_1117,N_2691);
nor U5178 (N_5178,N_1022,N_1157);
nor U5179 (N_5179,N_1527,N_1961);
nor U5180 (N_5180,N_69,N_678);
nor U5181 (N_5181,N_2567,N_2588);
xor U5182 (N_5182,N_2188,N_1270);
and U5183 (N_5183,N_150,N_730);
and U5184 (N_5184,N_77,N_2972);
nor U5185 (N_5185,N_1950,N_2153);
nand U5186 (N_5186,N_566,N_593);
or U5187 (N_5187,N_1739,N_486);
nor U5188 (N_5188,N_2714,N_1758);
or U5189 (N_5189,N_2382,N_2087);
or U5190 (N_5190,N_2150,N_1304);
nand U5191 (N_5191,N_2935,N_2815);
or U5192 (N_5192,N_1080,N_2159);
and U5193 (N_5193,N_2589,N_914);
nor U5194 (N_5194,N_1221,N_1436);
nor U5195 (N_5195,N_880,N_787);
nor U5196 (N_5196,N_339,N_2639);
nor U5197 (N_5197,N_2363,N_1817);
xnor U5198 (N_5198,N_41,N_1608);
nor U5199 (N_5199,N_2941,N_2538);
xor U5200 (N_5200,N_1902,N_1777);
nor U5201 (N_5201,N_781,N_1844);
xnor U5202 (N_5202,N_2472,N_1211);
nor U5203 (N_5203,N_1713,N_602);
and U5204 (N_5204,N_588,N_916);
nand U5205 (N_5205,N_441,N_1492);
or U5206 (N_5206,N_566,N_424);
and U5207 (N_5207,N_2698,N_1496);
and U5208 (N_5208,N_331,N_475);
and U5209 (N_5209,N_859,N_622);
nor U5210 (N_5210,N_2504,N_2149);
nand U5211 (N_5211,N_1767,N_388);
and U5212 (N_5212,N_2992,N_2591);
and U5213 (N_5213,N_1610,N_866);
nor U5214 (N_5214,N_2020,N_2368);
nor U5215 (N_5215,N_2497,N_2040);
or U5216 (N_5216,N_1151,N_2579);
or U5217 (N_5217,N_2654,N_1205);
xnor U5218 (N_5218,N_1216,N_371);
nor U5219 (N_5219,N_2021,N_993);
xnor U5220 (N_5220,N_1883,N_1384);
nand U5221 (N_5221,N_2791,N_2701);
nor U5222 (N_5222,N_1419,N_228);
and U5223 (N_5223,N_1084,N_2361);
and U5224 (N_5224,N_464,N_1284);
xnor U5225 (N_5225,N_674,N_433);
nor U5226 (N_5226,N_1032,N_1728);
and U5227 (N_5227,N_2915,N_1844);
nand U5228 (N_5228,N_2007,N_2711);
or U5229 (N_5229,N_2635,N_119);
or U5230 (N_5230,N_2310,N_2478);
and U5231 (N_5231,N_2417,N_190);
nor U5232 (N_5232,N_1037,N_2737);
and U5233 (N_5233,N_1869,N_684);
nand U5234 (N_5234,N_1880,N_281);
nor U5235 (N_5235,N_1935,N_172);
nand U5236 (N_5236,N_1593,N_1646);
nor U5237 (N_5237,N_744,N_2795);
xnor U5238 (N_5238,N_940,N_1817);
nor U5239 (N_5239,N_2213,N_2124);
nand U5240 (N_5240,N_2418,N_2556);
nand U5241 (N_5241,N_665,N_2881);
nand U5242 (N_5242,N_408,N_1518);
nor U5243 (N_5243,N_590,N_2043);
or U5244 (N_5244,N_1395,N_1489);
xnor U5245 (N_5245,N_1703,N_213);
and U5246 (N_5246,N_2412,N_219);
nand U5247 (N_5247,N_2677,N_929);
and U5248 (N_5248,N_2984,N_309);
nor U5249 (N_5249,N_1258,N_2949);
and U5250 (N_5250,N_2114,N_862);
nand U5251 (N_5251,N_209,N_2157);
or U5252 (N_5252,N_1987,N_216);
and U5253 (N_5253,N_1476,N_1461);
nor U5254 (N_5254,N_1053,N_911);
and U5255 (N_5255,N_2568,N_588);
nor U5256 (N_5256,N_1852,N_2830);
xor U5257 (N_5257,N_1212,N_1140);
and U5258 (N_5258,N_1532,N_1167);
nand U5259 (N_5259,N_1086,N_576);
nand U5260 (N_5260,N_542,N_1090);
and U5261 (N_5261,N_2201,N_2020);
xor U5262 (N_5262,N_1107,N_2560);
or U5263 (N_5263,N_1322,N_64);
or U5264 (N_5264,N_2726,N_1363);
xnor U5265 (N_5265,N_2321,N_774);
or U5266 (N_5266,N_1547,N_2684);
nor U5267 (N_5267,N_2713,N_2514);
nand U5268 (N_5268,N_1206,N_1925);
nor U5269 (N_5269,N_2182,N_2396);
xnor U5270 (N_5270,N_2467,N_2829);
xor U5271 (N_5271,N_2851,N_629);
and U5272 (N_5272,N_1365,N_2370);
nor U5273 (N_5273,N_2736,N_2598);
nor U5274 (N_5274,N_1818,N_1602);
nand U5275 (N_5275,N_1657,N_2852);
nand U5276 (N_5276,N_1541,N_1383);
or U5277 (N_5277,N_179,N_978);
xor U5278 (N_5278,N_1996,N_582);
and U5279 (N_5279,N_2828,N_2445);
xor U5280 (N_5280,N_583,N_422);
nor U5281 (N_5281,N_2626,N_2243);
nand U5282 (N_5282,N_1446,N_1637);
nor U5283 (N_5283,N_2064,N_2275);
nor U5284 (N_5284,N_2716,N_231);
and U5285 (N_5285,N_1402,N_1959);
and U5286 (N_5286,N_291,N_2009);
xor U5287 (N_5287,N_232,N_194);
or U5288 (N_5288,N_1222,N_1186);
nor U5289 (N_5289,N_2925,N_469);
or U5290 (N_5290,N_1899,N_167);
nand U5291 (N_5291,N_203,N_1237);
or U5292 (N_5292,N_836,N_1689);
xnor U5293 (N_5293,N_2747,N_2819);
xor U5294 (N_5294,N_2261,N_1256);
nor U5295 (N_5295,N_378,N_1045);
nand U5296 (N_5296,N_896,N_1238);
and U5297 (N_5297,N_2828,N_1118);
xor U5298 (N_5298,N_1172,N_1929);
nand U5299 (N_5299,N_765,N_127);
xnor U5300 (N_5300,N_656,N_2866);
and U5301 (N_5301,N_2206,N_1929);
and U5302 (N_5302,N_1290,N_243);
xnor U5303 (N_5303,N_2975,N_1144);
nor U5304 (N_5304,N_625,N_59);
nor U5305 (N_5305,N_2327,N_2333);
xor U5306 (N_5306,N_1083,N_2542);
xor U5307 (N_5307,N_1704,N_155);
nand U5308 (N_5308,N_51,N_2941);
nor U5309 (N_5309,N_622,N_1187);
or U5310 (N_5310,N_2809,N_2567);
nand U5311 (N_5311,N_2993,N_928);
nand U5312 (N_5312,N_579,N_2692);
and U5313 (N_5313,N_1415,N_2011);
nand U5314 (N_5314,N_1666,N_822);
and U5315 (N_5315,N_2014,N_2906);
nor U5316 (N_5316,N_467,N_439);
nand U5317 (N_5317,N_254,N_1461);
or U5318 (N_5318,N_1884,N_360);
or U5319 (N_5319,N_1492,N_854);
nand U5320 (N_5320,N_2121,N_2346);
xor U5321 (N_5321,N_1290,N_2543);
xnor U5322 (N_5322,N_2094,N_290);
nor U5323 (N_5323,N_1897,N_1604);
nand U5324 (N_5324,N_1932,N_1474);
xnor U5325 (N_5325,N_1645,N_2374);
nand U5326 (N_5326,N_1209,N_1810);
xor U5327 (N_5327,N_2304,N_2745);
nor U5328 (N_5328,N_469,N_1954);
xnor U5329 (N_5329,N_2017,N_1156);
nor U5330 (N_5330,N_8,N_2669);
or U5331 (N_5331,N_1584,N_171);
xor U5332 (N_5332,N_1255,N_997);
or U5333 (N_5333,N_400,N_1992);
nor U5334 (N_5334,N_2909,N_1897);
xor U5335 (N_5335,N_2201,N_2630);
or U5336 (N_5336,N_323,N_901);
and U5337 (N_5337,N_389,N_258);
and U5338 (N_5338,N_512,N_27);
or U5339 (N_5339,N_2436,N_857);
xor U5340 (N_5340,N_925,N_857);
or U5341 (N_5341,N_895,N_798);
xor U5342 (N_5342,N_447,N_2486);
and U5343 (N_5343,N_1939,N_1948);
xor U5344 (N_5344,N_1132,N_2815);
and U5345 (N_5345,N_20,N_43);
nand U5346 (N_5346,N_370,N_565);
and U5347 (N_5347,N_768,N_2519);
nor U5348 (N_5348,N_1513,N_984);
and U5349 (N_5349,N_1355,N_2832);
xnor U5350 (N_5350,N_1018,N_2256);
xnor U5351 (N_5351,N_929,N_2821);
or U5352 (N_5352,N_288,N_320);
nor U5353 (N_5353,N_648,N_992);
or U5354 (N_5354,N_2654,N_1638);
nor U5355 (N_5355,N_767,N_1603);
and U5356 (N_5356,N_209,N_1892);
nor U5357 (N_5357,N_323,N_2863);
or U5358 (N_5358,N_2999,N_1505);
or U5359 (N_5359,N_339,N_1575);
or U5360 (N_5360,N_1635,N_205);
nor U5361 (N_5361,N_1030,N_1976);
xor U5362 (N_5362,N_553,N_142);
and U5363 (N_5363,N_975,N_553);
and U5364 (N_5364,N_2622,N_1182);
xnor U5365 (N_5365,N_781,N_2226);
xor U5366 (N_5366,N_2965,N_2365);
and U5367 (N_5367,N_1513,N_1437);
xor U5368 (N_5368,N_1891,N_1586);
xor U5369 (N_5369,N_1681,N_2416);
and U5370 (N_5370,N_2790,N_2025);
and U5371 (N_5371,N_1774,N_87);
xnor U5372 (N_5372,N_1348,N_2535);
nand U5373 (N_5373,N_2863,N_484);
and U5374 (N_5374,N_2169,N_1534);
nand U5375 (N_5375,N_351,N_2137);
nor U5376 (N_5376,N_315,N_1077);
or U5377 (N_5377,N_291,N_9);
or U5378 (N_5378,N_2890,N_683);
nand U5379 (N_5379,N_371,N_702);
or U5380 (N_5380,N_2581,N_2477);
nor U5381 (N_5381,N_1284,N_1804);
or U5382 (N_5382,N_962,N_2130);
nand U5383 (N_5383,N_1987,N_1194);
nor U5384 (N_5384,N_63,N_2461);
nand U5385 (N_5385,N_2724,N_1289);
xnor U5386 (N_5386,N_462,N_249);
xor U5387 (N_5387,N_1647,N_2815);
nor U5388 (N_5388,N_1203,N_2249);
or U5389 (N_5389,N_2016,N_1097);
xnor U5390 (N_5390,N_1132,N_1113);
or U5391 (N_5391,N_1829,N_516);
or U5392 (N_5392,N_54,N_1608);
nor U5393 (N_5393,N_28,N_461);
nor U5394 (N_5394,N_1832,N_315);
and U5395 (N_5395,N_633,N_2120);
or U5396 (N_5396,N_1936,N_2060);
nor U5397 (N_5397,N_115,N_2738);
xnor U5398 (N_5398,N_284,N_875);
and U5399 (N_5399,N_99,N_2386);
xor U5400 (N_5400,N_1550,N_2589);
or U5401 (N_5401,N_1081,N_1100);
nor U5402 (N_5402,N_1832,N_684);
nor U5403 (N_5403,N_759,N_81);
and U5404 (N_5404,N_478,N_277);
and U5405 (N_5405,N_1330,N_1454);
xnor U5406 (N_5406,N_2435,N_1582);
or U5407 (N_5407,N_1231,N_2540);
or U5408 (N_5408,N_1078,N_1187);
nor U5409 (N_5409,N_2620,N_2597);
xor U5410 (N_5410,N_1071,N_649);
xnor U5411 (N_5411,N_2574,N_1034);
nand U5412 (N_5412,N_727,N_433);
xnor U5413 (N_5413,N_1320,N_1819);
or U5414 (N_5414,N_611,N_358);
and U5415 (N_5415,N_1829,N_1593);
nand U5416 (N_5416,N_2963,N_1391);
nor U5417 (N_5417,N_1914,N_2406);
or U5418 (N_5418,N_2949,N_1132);
or U5419 (N_5419,N_243,N_233);
or U5420 (N_5420,N_553,N_1869);
and U5421 (N_5421,N_2826,N_1005);
xnor U5422 (N_5422,N_207,N_2262);
nor U5423 (N_5423,N_2911,N_1811);
nor U5424 (N_5424,N_1296,N_2632);
nand U5425 (N_5425,N_2426,N_2233);
xnor U5426 (N_5426,N_517,N_2528);
and U5427 (N_5427,N_504,N_2721);
or U5428 (N_5428,N_2038,N_1609);
or U5429 (N_5429,N_1846,N_2841);
xor U5430 (N_5430,N_2152,N_1517);
nand U5431 (N_5431,N_73,N_1283);
and U5432 (N_5432,N_315,N_2845);
nor U5433 (N_5433,N_437,N_2858);
and U5434 (N_5434,N_1412,N_459);
xor U5435 (N_5435,N_635,N_1454);
or U5436 (N_5436,N_1992,N_2814);
nand U5437 (N_5437,N_2429,N_241);
nor U5438 (N_5438,N_333,N_1790);
nor U5439 (N_5439,N_1242,N_455);
xnor U5440 (N_5440,N_2771,N_248);
xor U5441 (N_5441,N_1375,N_1864);
and U5442 (N_5442,N_783,N_1321);
nand U5443 (N_5443,N_267,N_94);
xor U5444 (N_5444,N_962,N_1654);
xor U5445 (N_5445,N_2729,N_1336);
xor U5446 (N_5446,N_1669,N_2595);
xor U5447 (N_5447,N_148,N_2671);
nand U5448 (N_5448,N_783,N_368);
nand U5449 (N_5449,N_2048,N_456);
nand U5450 (N_5450,N_1785,N_193);
and U5451 (N_5451,N_1816,N_2829);
or U5452 (N_5452,N_424,N_569);
and U5453 (N_5453,N_1530,N_1920);
nor U5454 (N_5454,N_186,N_1407);
and U5455 (N_5455,N_957,N_1424);
nor U5456 (N_5456,N_2805,N_996);
xor U5457 (N_5457,N_690,N_329);
nor U5458 (N_5458,N_1817,N_321);
nand U5459 (N_5459,N_141,N_2154);
or U5460 (N_5460,N_2890,N_1952);
nand U5461 (N_5461,N_2120,N_1407);
and U5462 (N_5462,N_640,N_74);
or U5463 (N_5463,N_1679,N_2266);
and U5464 (N_5464,N_2039,N_2889);
nand U5465 (N_5465,N_1990,N_1359);
nand U5466 (N_5466,N_356,N_2735);
or U5467 (N_5467,N_2173,N_2101);
nor U5468 (N_5468,N_2674,N_2727);
and U5469 (N_5469,N_2408,N_399);
and U5470 (N_5470,N_336,N_1200);
and U5471 (N_5471,N_2526,N_48);
nand U5472 (N_5472,N_1248,N_2818);
xnor U5473 (N_5473,N_1414,N_505);
nor U5474 (N_5474,N_2030,N_2842);
nand U5475 (N_5475,N_1299,N_422);
nor U5476 (N_5476,N_1859,N_1592);
xor U5477 (N_5477,N_2354,N_821);
nor U5478 (N_5478,N_1031,N_235);
nand U5479 (N_5479,N_515,N_777);
nor U5480 (N_5480,N_1795,N_1403);
nand U5481 (N_5481,N_565,N_1722);
xor U5482 (N_5482,N_2834,N_1879);
or U5483 (N_5483,N_2981,N_1087);
xnor U5484 (N_5484,N_2584,N_79);
and U5485 (N_5485,N_913,N_498);
nand U5486 (N_5486,N_2045,N_1643);
nand U5487 (N_5487,N_2915,N_2623);
or U5488 (N_5488,N_1289,N_776);
nor U5489 (N_5489,N_1426,N_2605);
and U5490 (N_5490,N_531,N_2906);
nand U5491 (N_5491,N_1667,N_1781);
or U5492 (N_5492,N_1097,N_2809);
nor U5493 (N_5493,N_2973,N_1278);
or U5494 (N_5494,N_1637,N_93);
or U5495 (N_5495,N_593,N_2552);
nor U5496 (N_5496,N_332,N_778);
nor U5497 (N_5497,N_1239,N_1236);
and U5498 (N_5498,N_2495,N_1447);
and U5499 (N_5499,N_1953,N_1014);
nor U5500 (N_5500,N_2323,N_1717);
nor U5501 (N_5501,N_149,N_468);
or U5502 (N_5502,N_1695,N_2272);
nand U5503 (N_5503,N_889,N_1575);
nor U5504 (N_5504,N_410,N_1700);
nor U5505 (N_5505,N_1911,N_62);
nand U5506 (N_5506,N_71,N_1614);
nor U5507 (N_5507,N_1747,N_2016);
nand U5508 (N_5508,N_2014,N_2266);
xor U5509 (N_5509,N_374,N_1275);
nor U5510 (N_5510,N_218,N_847);
nand U5511 (N_5511,N_809,N_413);
nand U5512 (N_5512,N_2396,N_696);
nand U5513 (N_5513,N_2855,N_1761);
or U5514 (N_5514,N_1079,N_2882);
or U5515 (N_5515,N_831,N_186);
nor U5516 (N_5516,N_2060,N_188);
xor U5517 (N_5517,N_37,N_1377);
or U5518 (N_5518,N_77,N_2080);
nor U5519 (N_5519,N_505,N_2306);
xnor U5520 (N_5520,N_858,N_767);
xor U5521 (N_5521,N_2932,N_223);
xnor U5522 (N_5522,N_250,N_1122);
and U5523 (N_5523,N_846,N_1701);
xnor U5524 (N_5524,N_2323,N_195);
nor U5525 (N_5525,N_2443,N_1667);
xnor U5526 (N_5526,N_1103,N_2700);
nand U5527 (N_5527,N_2489,N_2592);
nor U5528 (N_5528,N_833,N_1665);
xor U5529 (N_5529,N_1074,N_280);
or U5530 (N_5530,N_1347,N_718);
or U5531 (N_5531,N_831,N_1692);
nor U5532 (N_5532,N_159,N_916);
or U5533 (N_5533,N_509,N_972);
xor U5534 (N_5534,N_2773,N_971);
and U5535 (N_5535,N_2124,N_2324);
or U5536 (N_5536,N_1904,N_217);
and U5537 (N_5537,N_2546,N_2603);
xnor U5538 (N_5538,N_2469,N_455);
nor U5539 (N_5539,N_34,N_2474);
and U5540 (N_5540,N_1453,N_2485);
xnor U5541 (N_5541,N_1821,N_2077);
xnor U5542 (N_5542,N_1470,N_384);
nand U5543 (N_5543,N_188,N_843);
xnor U5544 (N_5544,N_272,N_2630);
and U5545 (N_5545,N_2314,N_2223);
nand U5546 (N_5546,N_1185,N_1083);
nand U5547 (N_5547,N_2772,N_10);
and U5548 (N_5548,N_2536,N_782);
or U5549 (N_5549,N_2222,N_1625);
and U5550 (N_5550,N_2814,N_2265);
or U5551 (N_5551,N_10,N_1060);
and U5552 (N_5552,N_1487,N_2384);
or U5553 (N_5553,N_2705,N_582);
nor U5554 (N_5554,N_1087,N_2906);
xnor U5555 (N_5555,N_2554,N_1087);
xor U5556 (N_5556,N_1548,N_1183);
nor U5557 (N_5557,N_837,N_637);
xnor U5558 (N_5558,N_2993,N_2761);
nand U5559 (N_5559,N_1074,N_1340);
nand U5560 (N_5560,N_2803,N_1738);
nand U5561 (N_5561,N_2397,N_1262);
nand U5562 (N_5562,N_837,N_2389);
and U5563 (N_5563,N_1461,N_81);
nand U5564 (N_5564,N_1475,N_2604);
or U5565 (N_5565,N_125,N_1319);
nor U5566 (N_5566,N_1221,N_804);
nor U5567 (N_5567,N_1119,N_688);
or U5568 (N_5568,N_377,N_215);
nand U5569 (N_5569,N_1684,N_28);
and U5570 (N_5570,N_2102,N_2189);
or U5571 (N_5571,N_2881,N_2788);
nor U5572 (N_5572,N_1050,N_1955);
and U5573 (N_5573,N_1400,N_2726);
or U5574 (N_5574,N_1496,N_229);
nand U5575 (N_5575,N_438,N_2508);
or U5576 (N_5576,N_2499,N_398);
and U5577 (N_5577,N_801,N_1999);
and U5578 (N_5578,N_2544,N_180);
nand U5579 (N_5579,N_1767,N_955);
xnor U5580 (N_5580,N_2068,N_1099);
or U5581 (N_5581,N_751,N_1602);
and U5582 (N_5582,N_14,N_618);
nand U5583 (N_5583,N_1547,N_427);
xnor U5584 (N_5584,N_1456,N_1003);
or U5585 (N_5585,N_716,N_1763);
or U5586 (N_5586,N_1117,N_1584);
nor U5587 (N_5587,N_2547,N_1120);
nand U5588 (N_5588,N_810,N_792);
or U5589 (N_5589,N_1680,N_844);
nor U5590 (N_5590,N_581,N_1868);
xnor U5591 (N_5591,N_1277,N_1519);
xor U5592 (N_5592,N_963,N_1733);
nor U5593 (N_5593,N_701,N_2933);
nand U5594 (N_5594,N_1665,N_2948);
nor U5595 (N_5595,N_1222,N_2103);
nand U5596 (N_5596,N_2334,N_1364);
and U5597 (N_5597,N_2012,N_1451);
or U5598 (N_5598,N_2117,N_2712);
and U5599 (N_5599,N_1317,N_1376);
and U5600 (N_5600,N_667,N_2685);
nor U5601 (N_5601,N_2619,N_2882);
and U5602 (N_5602,N_1113,N_474);
nor U5603 (N_5603,N_2300,N_675);
nand U5604 (N_5604,N_1854,N_2887);
xnor U5605 (N_5605,N_547,N_99);
and U5606 (N_5606,N_1921,N_2188);
xnor U5607 (N_5607,N_264,N_560);
and U5608 (N_5608,N_1238,N_1637);
xnor U5609 (N_5609,N_968,N_2352);
xor U5610 (N_5610,N_1068,N_1795);
and U5611 (N_5611,N_1213,N_314);
nor U5612 (N_5612,N_2778,N_1053);
nor U5613 (N_5613,N_2655,N_1984);
nor U5614 (N_5614,N_2086,N_1950);
nor U5615 (N_5615,N_2262,N_590);
nor U5616 (N_5616,N_1857,N_1736);
or U5617 (N_5617,N_1115,N_2272);
or U5618 (N_5618,N_1700,N_289);
nand U5619 (N_5619,N_2542,N_1538);
and U5620 (N_5620,N_285,N_2860);
nor U5621 (N_5621,N_359,N_170);
nand U5622 (N_5622,N_1221,N_2211);
or U5623 (N_5623,N_3,N_1353);
or U5624 (N_5624,N_2774,N_452);
and U5625 (N_5625,N_1379,N_585);
nor U5626 (N_5626,N_49,N_504);
or U5627 (N_5627,N_2921,N_1331);
nor U5628 (N_5628,N_2310,N_2204);
xnor U5629 (N_5629,N_1309,N_2404);
or U5630 (N_5630,N_93,N_1238);
xor U5631 (N_5631,N_2728,N_2709);
and U5632 (N_5632,N_1963,N_2493);
nor U5633 (N_5633,N_2202,N_2410);
nand U5634 (N_5634,N_411,N_717);
nor U5635 (N_5635,N_2513,N_906);
xnor U5636 (N_5636,N_2198,N_291);
xor U5637 (N_5637,N_1643,N_1886);
nor U5638 (N_5638,N_2580,N_1556);
xnor U5639 (N_5639,N_1090,N_785);
and U5640 (N_5640,N_2578,N_1948);
or U5641 (N_5641,N_1182,N_54);
and U5642 (N_5642,N_1974,N_721);
nor U5643 (N_5643,N_2617,N_526);
and U5644 (N_5644,N_2851,N_483);
or U5645 (N_5645,N_1438,N_340);
nor U5646 (N_5646,N_888,N_305);
xnor U5647 (N_5647,N_925,N_359);
or U5648 (N_5648,N_2784,N_296);
nor U5649 (N_5649,N_2626,N_2682);
or U5650 (N_5650,N_153,N_1726);
or U5651 (N_5651,N_1047,N_185);
nor U5652 (N_5652,N_1344,N_1752);
nand U5653 (N_5653,N_496,N_1548);
xor U5654 (N_5654,N_2340,N_2765);
and U5655 (N_5655,N_1431,N_734);
or U5656 (N_5656,N_311,N_1012);
or U5657 (N_5657,N_202,N_1292);
nand U5658 (N_5658,N_177,N_2504);
xor U5659 (N_5659,N_1016,N_920);
xor U5660 (N_5660,N_805,N_481);
xnor U5661 (N_5661,N_799,N_1102);
xor U5662 (N_5662,N_2677,N_1776);
nand U5663 (N_5663,N_2349,N_1008);
and U5664 (N_5664,N_1724,N_78);
nor U5665 (N_5665,N_1610,N_136);
nand U5666 (N_5666,N_496,N_304);
and U5667 (N_5667,N_39,N_741);
xor U5668 (N_5668,N_2775,N_311);
nand U5669 (N_5669,N_2953,N_2059);
xnor U5670 (N_5670,N_576,N_2464);
xor U5671 (N_5671,N_1125,N_582);
and U5672 (N_5672,N_865,N_29);
nand U5673 (N_5673,N_2285,N_2204);
xor U5674 (N_5674,N_421,N_1938);
and U5675 (N_5675,N_1376,N_415);
xor U5676 (N_5676,N_685,N_263);
xnor U5677 (N_5677,N_2192,N_1510);
xor U5678 (N_5678,N_1373,N_1184);
xnor U5679 (N_5679,N_1038,N_756);
xor U5680 (N_5680,N_1699,N_2536);
nand U5681 (N_5681,N_46,N_389);
xnor U5682 (N_5682,N_1516,N_63);
xor U5683 (N_5683,N_1670,N_204);
nand U5684 (N_5684,N_2609,N_1973);
nand U5685 (N_5685,N_2649,N_1662);
nand U5686 (N_5686,N_2765,N_1681);
xnor U5687 (N_5687,N_2498,N_2622);
or U5688 (N_5688,N_2080,N_21);
nand U5689 (N_5689,N_1523,N_277);
or U5690 (N_5690,N_15,N_2498);
xor U5691 (N_5691,N_1837,N_1827);
or U5692 (N_5692,N_1161,N_1055);
xor U5693 (N_5693,N_2551,N_1174);
or U5694 (N_5694,N_226,N_479);
and U5695 (N_5695,N_1026,N_1237);
nand U5696 (N_5696,N_1235,N_2287);
nor U5697 (N_5697,N_988,N_453);
nor U5698 (N_5698,N_791,N_2563);
and U5699 (N_5699,N_517,N_1275);
xnor U5700 (N_5700,N_1401,N_1640);
nor U5701 (N_5701,N_1925,N_1614);
and U5702 (N_5702,N_2760,N_825);
and U5703 (N_5703,N_177,N_480);
nand U5704 (N_5704,N_2500,N_939);
nand U5705 (N_5705,N_2025,N_834);
or U5706 (N_5706,N_2971,N_2635);
nor U5707 (N_5707,N_200,N_1175);
xnor U5708 (N_5708,N_1594,N_1197);
nand U5709 (N_5709,N_1723,N_286);
nand U5710 (N_5710,N_993,N_1209);
or U5711 (N_5711,N_1365,N_1873);
or U5712 (N_5712,N_2366,N_81);
nor U5713 (N_5713,N_185,N_2852);
nor U5714 (N_5714,N_2992,N_0);
nand U5715 (N_5715,N_294,N_2564);
or U5716 (N_5716,N_434,N_1887);
nor U5717 (N_5717,N_2921,N_954);
nand U5718 (N_5718,N_754,N_924);
and U5719 (N_5719,N_1394,N_291);
and U5720 (N_5720,N_755,N_2748);
and U5721 (N_5721,N_845,N_2472);
nor U5722 (N_5722,N_419,N_117);
or U5723 (N_5723,N_1178,N_2884);
nand U5724 (N_5724,N_2585,N_246);
nor U5725 (N_5725,N_2560,N_896);
nor U5726 (N_5726,N_229,N_1897);
and U5727 (N_5727,N_81,N_1688);
nor U5728 (N_5728,N_2706,N_2962);
and U5729 (N_5729,N_933,N_878);
xnor U5730 (N_5730,N_1881,N_2277);
xnor U5731 (N_5731,N_1386,N_2319);
nor U5732 (N_5732,N_46,N_2199);
or U5733 (N_5733,N_1243,N_2983);
xor U5734 (N_5734,N_1467,N_558);
and U5735 (N_5735,N_198,N_669);
nor U5736 (N_5736,N_1302,N_2330);
nand U5737 (N_5737,N_982,N_761);
nor U5738 (N_5738,N_2071,N_1777);
and U5739 (N_5739,N_1707,N_480);
nor U5740 (N_5740,N_1439,N_708);
xnor U5741 (N_5741,N_1796,N_720);
xor U5742 (N_5742,N_1789,N_2877);
nand U5743 (N_5743,N_47,N_1062);
nor U5744 (N_5744,N_488,N_440);
or U5745 (N_5745,N_2166,N_822);
or U5746 (N_5746,N_1806,N_2228);
nand U5747 (N_5747,N_1434,N_1189);
nor U5748 (N_5748,N_2796,N_1034);
xor U5749 (N_5749,N_2428,N_2795);
or U5750 (N_5750,N_1057,N_1942);
or U5751 (N_5751,N_1065,N_1301);
or U5752 (N_5752,N_1214,N_2565);
nor U5753 (N_5753,N_1191,N_2452);
and U5754 (N_5754,N_707,N_2080);
and U5755 (N_5755,N_1381,N_2812);
xor U5756 (N_5756,N_1499,N_1225);
nor U5757 (N_5757,N_2675,N_40);
nor U5758 (N_5758,N_2776,N_2890);
nand U5759 (N_5759,N_2720,N_2220);
xor U5760 (N_5760,N_1429,N_1141);
or U5761 (N_5761,N_1500,N_550);
xnor U5762 (N_5762,N_2812,N_1374);
nor U5763 (N_5763,N_1701,N_2812);
and U5764 (N_5764,N_2728,N_749);
xnor U5765 (N_5765,N_2961,N_716);
nand U5766 (N_5766,N_2185,N_591);
nor U5767 (N_5767,N_1939,N_2270);
nor U5768 (N_5768,N_2960,N_1881);
nor U5769 (N_5769,N_2244,N_452);
or U5770 (N_5770,N_485,N_1714);
nor U5771 (N_5771,N_2060,N_1438);
nand U5772 (N_5772,N_2368,N_2081);
or U5773 (N_5773,N_2609,N_1971);
xnor U5774 (N_5774,N_1493,N_2403);
nor U5775 (N_5775,N_908,N_949);
xnor U5776 (N_5776,N_2728,N_1617);
nor U5777 (N_5777,N_1220,N_737);
nor U5778 (N_5778,N_2344,N_2675);
nor U5779 (N_5779,N_851,N_386);
nor U5780 (N_5780,N_2628,N_514);
nor U5781 (N_5781,N_1368,N_1117);
nand U5782 (N_5782,N_2185,N_519);
nand U5783 (N_5783,N_645,N_2172);
and U5784 (N_5784,N_529,N_422);
nand U5785 (N_5785,N_409,N_322);
xnor U5786 (N_5786,N_1500,N_1142);
or U5787 (N_5787,N_625,N_1587);
and U5788 (N_5788,N_2958,N_2668);
nor U5789 (N_5789,N_1055,N_767);
or U5790 (N_5790,N_2128,N_2789);
or U5791 (N_5791,N_2866,N_1014);
or U5792 (N_5792,N_1891,N_2265);
or U5793 (N_5793,N_1677,N_563);
or U5794 (N_5794,N_1150,N_534);
and U5795 (N_5795,N_1034,N_2363);
nand U5796 (N_5796,N_1867,N_2646);
and U5797 (N_5797,N_2457,N_2549);
or U5798 (N_5798,N_2677,N_791);
xnor U5799 (N_5799,N_164,N_2234);
nor U5800 (N_5800,N_2229,N_114);
xnor U5801 (N_5801,N_1101,N_551);
xor U5802 (N_5802,N_1238,N_2946);
or U5803 (N_5803,N_2433,N_2143);
or U5804 (N_5804,N_2898,N_1178);
xor U5805 (N_5805,N_933,N_1131);
and U5806 (N_5806,N_720,N_1224);
or U5807 (N_5807,N_1193,N_2219);
and U5808 (N_5808,N_2919,N_1991);
nand U5809 (N_5809,N_1575,N_138);
xnor U5810 (N_5810,N_1093,N_608);
or U5811 (N_5811,N_1681,N_2605);
nand U5812 (N_5812,N_578,N_1033);
or U5813 (N_5813,N_904,N_2658);
nand U5814 (N_5814,N_1178,N_2171);
and U5815 (N_5815,N_146,N_777);
xnor U5816 (N_5816,N_427,N_291);
nor U5817 (N_5817,N_1021,N_314);
nor U5818 (N_5818,N_1205,N_1227);
and U5819 (N_5819,N_565,N_185);
nand U5820 (N_5820,N_2072,N_1584);
nand U5821 (N_5821,N_856,N_2808);
and U5822 (N_5822,N_1155,N_2866);
nor U5823 (N_5823,N_2205,N_2410);
xor U5824 (N_5824,N_2148,N_905);
nor U5825 (N_5825,N_2582,N_2658);
nor U5826 (N_5826,N_2470,N_2999);
nand U5827 (N_5827,N_1956,N_2763);
or U5828 (N_5828,N_1353,N_2950);
xor U5829 (N_5829,N_709,N_22);
or U5830 (N_5830,N_348,N_1224);
or U5831 (N_5831,N_2099,N_1531);
nand U5832 (N_5832,N_2470,N_1822);
xnor U5833 (N_5833,N_554,N_936);
nor U5834 (N_5834,N_1159,N_542);
nand U5835 (N_5835,N_57,N_1820);
and U5836 (N_5836,N_495,N_1149);
nand U5837 (N_5837,N_2393,N_2506);
or U5838 (N_5838,N_1443,N_2855);
nor U5839 (N_5839,N_116,N_628);
or U5840 (N_5840,N_970,N_353);
nand U5841 (N_5841,N_2771,N_793);
nand U5842 (N_5842,N_687,N_1041);
xnor U5843 (N_5843,N_2944,N_243);
nor U5844 (N_5844,N_854,N_2512);
nand U5845 (N_5845,N_2900,N_1660);
xnor U5846 (N_5846,N_637,N_1723);
and U5847 (N_5847,N_1091,N_197);
xnor U5848 (N_5848,N_434,N_803);
nor U5849 (N_5849,N_453,N_459);
nand U5850 (N_5850,N_1047,N_356);
or U5851 (N_5851,N_1556,N_1063);
xnor U5852 (N_5852,N_1060,N_40);
or U5853 (N_5853,N_345,N_211);
or U5854 (N_5854,N_2529,N_755);
xnor U5855 (N_5855,N_1999,N_299);
and U5856 (N_5856,N_294,N_1678);
and U5857 (N_5857,N_97,N_301);
or U5858 (N_5858,N_750,N_995);
or U5859 (N_5859,N_858,N_2277);
nand U5860 (N_5860,N_470,N_350);
and U5861 (N_5861,N_2232,N_2904);
and U5862 (N_5862,N_1550,N_2989);
nor U5863 (N_5863,N_2460,N_2728);
nor U5864 (N_5864,N_2134,N_2464);
or U5865 (N_5865,N_1605,N_225);
nand U5866 (N_5866,N_962,N_1882);
xnor U5867 (N_5867,N_1340,N_2880);
nor U5868 (N_5868,N_1326,N_2228);
or U5869 (N_5869,N_612,N_1380);
and U5870 (N_5870,N_833,N_471);
nand U5871 (N_5871,N_2443,N_445);
or U5872 (N_5872,N_1889,N_896);
nand U5873 (N_5873,N_1158,N_2536);
nand U5874 (N_5874,N_335,N_1535);
and U5875 (N_5875,N_2556,N_612);
and U5876 (N_5876,N_2590,N_1019);
nand U5877 (N_5877,N_428,N_1208);
or U5878 (N_5878,N_509,N_2620);
xor U5879 (N_5879,N_14,N_800);
or U5880 (N_5880,N_699,N_2732);
xnor U5881 (N_5881,N_2025,N_850);
nor U5882 (N_5882,N_2548,N_413);
and U5883 (N_5883,N_1605,N_2334);
and U5884 (N_5884,N_2614,N_1922);
nand U5885 (N_5885,N_980,N_1116);
nor U5886 (N_5886,N_1521,N_891);
xor U5887 (N_5887,N_2063,N_1759);
xor U5888 (N_5888,N_2897,N_2342);
and U5889 (N_5889,N_1527,N_458);
or U5890 (N_5890,N_1095,N_1512);
xor U5891 (N_5891,N_141,N_2133);
xor U5892 (N_5892,N_868,N_2468);
nor U5893 (N_5893,N_1260,N_932);
nand U5894 (N_5894,N_2886,N_853);
and U5895 (N_5895,N_495,N_563);
nand U5896 (N_5896,N_2019,N_610);
nor U5897 (N_5897,N_2479,N_1144);
or U5898 (N_5898,N_1295,N_922);
and U5899 (N_5899,N_2824,N_151);
or U5900 (N_5900,N_313,N_1303);
nor U5901 (N_5901,N_1527,N_2527);
nor U5902 (N_5902,N_74,N_2003);
or U5903 (N_5903,N_663,N_400);
nor U5904 (N_5904,N_2353,N_1869);
and U5905 (N_5905,N_2921,N_310);
nor U5906 (N_5906,N_402,N_2767);
and U5907 (N_5907,N_1985,N_2295);
and U5908 (N_5908,N_1485,N_1441);
nor U5909 (N_5909,N_2330,N_534);
nand U5910 (N_5910,N_1896,N_731);
or U5911 (N_5911,N_2625,N_293);
nand U5912 (N_5912,N_271,N_513);
nand U5913 (N_5913,N_2626,N_2322);
nand U5914 (N_5914,N_2181,N_2816);
nand U5915 (N_5915,N_122,N_1580);
nor U5916 (N_5916,N_19,N_2303);
and U5917 (N_5917,N_208,N_2091);
and U5918 (N_5918,N_1162,N_59);
or U5919 (N_5919,N_2821,N_2167);
and U5920 (N_5920,N_432,N_1540);
xnor U5921 (N_5921,N_37,N_1916);
nand U5922 (N_5922,N_340,N_1783);
xor U5923 (N_5923,N_807,N_255);
nand U5924 (N_5924,N_2209,N_1153);
or U5925 (N_5925,N_2343,N_1877);
nor U5926 (N_5926,N_2800,N_9);
nor U5927 (N_5927,N_2544,N_1984);
xor U5928 (N_5928,N_479,N_2449);
or U5929 (N_5929,N_1847,N_31);
xor U5930 (N_5930,N_1951,N_390);
or U5931 (N_5931,N_363,N_1689);
xnor U5932 (N_5932,N_2929,N_1429);
nand U5933 (N_5933,N_1583,N_1247);
nor U5934 (N_5934,N_2797,N_1044);
or U5935 (N_5935,N_2186,N_2947);
nor U5936 (N_5936,N_807,N_333);
and U5937 (N_5937,N_2560,N_678);
nand U5938 (N_5938,N_1958,N_188);
xnor U5939 (N_5939,N_2404,N_931);
or U5940 (N_5940,N_2457,N_2278);
and U5941 (N_5941,N_37,N_2830);
nor U5942 (N_5942,N_2239,N_2093);
xor U5943 (N_5943,N_2353,N_613);
nor U5944 (N_5944,N_644,N_1339);
xnor U5945 (N_5945,N_2105,N_2612);
nand U5946 (N_5946,N_138,N_2988);
and U5947 (N_5947,N_2575,N_1615);
nand U5948 (N_5948,N_1277,N_2894);
nand U5949 (N_5949,N_771,N_1727);
and U5950 (N_5950,N_479,N_670);
and U5951 (N_5951,N_666,N_1986);
nand U5952 (N_5952,N_1688,N_89);
xor U5953 (N_5953,N_1470,N_455);
xnor U5954 (N_5954,N_73,N_2421);
or U5955 (N_5955,N_1118,N_1316);
nand U5956 (N_5956,N_1258,N_958);
or U5957 (N_5957,N_2066,N_1512);
xnor U5958 (N_5958,N_1438,N_262);
nand U5959 (N_5959,N_1511,N_2457);
nand U5960 (N_5960,N_1472,N_2785);
nor U5961 (N_5961,N_663,N_2271);
nor U5962 (N_5962,N_338,N_2558);
nand U5963 (N_5963,N_1565,N_2491);
and U5964 (N_5964,N_2758,N_2505);
xor U5965 (N_5965,N_901,N_1594);
nand U5966 (N_5966,N_2640,N_2944);
nand U5967 (N_5967,N_1553,N_1087);
xor U5968 (N_5968,N_2046,N_1444);
or U5969 (N_5969,N_2257,N_141);
nand U5970 (N_5970,N_2480,N_1740);
nor U5971 (N_5971,N_1792,N_127);
and U5972 (N_5972,N_498,N_294);
xor U5973 (N_5973,N_1394,N_585);
or U5974 (N_5974,N_1187,N_2108);
nor U5975 (N_5975,N_2795,N_2807);
nor U5976 (N_5976,N_1163,N_986);
or U5977 (N_5977,N_351,N_1134);
xnor U5978 (N_5978,N_70,N_1564);
xor U5979 (N_5979,N_1844,N_510);
or U5980 (N_5980,N_1193,N_1203);
and U5981 (N_5981,N_577,N_2118);
nand U5982 (N_5982,N_1921,N_2435);
or U5983 (N_5983,N_2312,N_1917);
or U5984 (N_5984,N_2352,N_1499);
nand U5985 (N_5985,N_2213,N_2602);
nand U5986 (N_5986,N_288,N_2654);
xnor U5987 (N_5987,N_315,N_1880);
xor U5988 (N_5988,N_1218,N_1762);
nand U5989 (N_5989,N_917,N_2143);
nor U5990 (N_5990,N_2377,N_1422);
and U5991 (N_5991,N_2939,N_2058);
or U5992 (N_5992,N_1834,N_2559);
nor U5993 (N_5993,N_1782,N_2488);
and U5994 (N_5994,N_526,N_1878);
nand U5995 (N_5995,N_2504,N_121);
nand U5996 (N_5996,N_710,N_1687);
and U5997 (N_5997,N_12,N_1063);
nor U5998 (N_5998,N_2346,N_1606);
nor U5999 (N_5999,N_287,N_1433);
xor U6000 (N_6000,N_3070,N_5084);
xnor U6001 (N_6001,N_5832,N_4311);
nor U6002 (N_6002,N_4115,N_3220);
nand U6003 (N_6003,N_3773,N_3041);
nor U6004 (N_6004,N_4869,N_5901);
and U6005 (N_6005,N_5926,N_3861);
and U6006 (N_6006,N_3822,N_3718);
xor U6007 (N_6007,N_5667,N_3143);
and U6008 (N_6008,N_5765,N_4771);
or U6009 (N_6009,N_4479,N_4693);
or U6010 (N_6010,N_3442,N_5664);
or U6011 (N_6011,N_5899,N_5722);
or U6012 (N_6012,N_5592,N_4126);
nor U6013 (N_6013,N_3342,N_3825);
and U6014 (N_6014,N_4895,N_3841);
and U6015 (N_6015,N_5790,N_4466);
xnor U6016 (N_6016,N_4616,N_3438);
or U6017 (N_6017,N_4719,N_3267);
and U6018 (N_6018,N_3660,N_5986);
or U6019 (N_6019,N_4852,N_3658);
nor U6020 (N_6020,N_4442,N_4822);
nand U6021 (N_6021,N_5402,N_3521);
xnor U6022 (N_6022,N_3706,N_4413);
or U6023 (N_6023,N_5346,N_5611);
xnor U6024 (N_6024,N_4043,N_3894);
and U6025 (N_6025,N_4261,N_5065);
nor U6026 (N_6026,N_3454,N_5030);
nand U6027 (N_6027,N_4424,N_3077);
xnor U6028 (N_6028,N_4829,N_5264);
or U6029 (N_6029,N_4603,N_3761);
and U6030 (N_6030,N_3466,N_5078);
or U6031 (N_6031,N_5163,N_5048);
nand U6032 (N_6032,N_4241,N_4416);
xnor U6033 (N_6033,N_5513,N_4515);
or U6034 (N_6034,N_3348,N_3066);
nor U6035 (N_6035,N_5888,N_5424);
xor U6036 (N_6036,N_4856,N_4784);
xnor U6037 (N_6037,N_4123,N_4551);
xor U6038 (N_6038,N_4761,N_5735);
or U6039 (N_6039,N_4091,N_4872);
nor U6040 (N_6040,N_3393,N_3802);
nand U6041 (N_6041,N_5826,N_5374);
nor U6042 (N_6042,N_3698,N_4972);
or U6043 (N_6043,N_4046,N_4720);
xnor U6044 (N_6044,N_5041,N_3238);
xnor U6045 (N_6045,N_3370,N_3211);
and U6046 (N_6046,N_3257,N_3952);
nand U6047 (N_6047,N_5138,N_3282);
or U6048 (N_6048,N_5243,N_3541);
and U6049 (N_6049,N_5267,N_4238);
and U6050 (N_6050,N_3852,N_4282);
nor U6051 (N_6051,N_4791,N_3312);
nand U6052 (N_6052,N_4219,N_5794);
or U6053 (N_6053,N_5809,N_4568);
nand U6054 (N_6054,N_3672,N_3303);
nand U6055 (N_6055,N_3863,N_4073);
and U6056 (N_6056,N_5439,N_4580);
and U6057 (N_6057,N_5983,N_4069);
xor U6058 (N_6058,N_5185,N_3098);
or U6059 (N_6059,N_4525,N_4445);
or U6060 (N_6060,N_3969,N_3446);
xnor U6061 (N_6061,N_5963,N_4854);
and U6062 (N_6062,N_3757,N_3518);
nand U6063 (N_6063,N_4229,N_4454);
nand U6064 (N_6064,N_4393,N_4557);
nand U6065 (N_6065,N_3359,N_3310);
nand U6066 (N_6066,N_4254,N_4853);
nor U6067 (N_6067,N_5519,N_3690);
nand U6068 (N_6068,N_3300,N_4200);
or U6069 (N_6069,N_4528,N_4604);
and U6070 (N_6070,N_5134,N_5271);
nor U6071 (N_6071,N_5458,N_4918);
and U6072 (N_6072,N_5702,N_3531);
xnor U6073 (N_6073,N_3369,N_4710);
nor U6074 (N_6074,N_4266,N_3708);
or U6075 (N_6075,N_5507,N_3404);
and U6076 (N_6076,N_3017,N_4265);
and U6077 (N_6077,N_5736,N_3021);
nor U6078 (N_6078,N_4201,N_4991);
and U6079 (N_6079,N_5207,N_4347);
or U6080 (N_6080,N_5177,N_4045);
or U6081 (N_6081,N_4334,N_4510);
and U6082 (N_6082,N_4776,N_5102);
nor U6083 (N_6083,N_4076,N_5654);
xnor U6084 (N_6084,N_5072,N_3354);
and U6085 (N_6085,N_4615,N_5497);
nand U6086 (N_6086,N_3172,N_3721);
or U6087 (N_6087,N_5012,N_5687);
and U6088 (N_6088,N_3772,N_4176);
nand U6089 (N_6089,N_4731,N_4906);
and U6090 (N_6090,N_5292,N_3752);
or U6091 (N_6091,N_3948,N_4927);
xor U6092 (N_6092,N_3262,N_4730);
and U6093 (N_6093,N_3659,N_4026);
xnor U6094 (N_6094,N_3272,N_5136);
xnor U6095 (N_6095,N_5997,N_4517);
and U6096 (N_6096,N_4954,N_5036);
xor U6097 (N_6097,N_5238,N_4996);
xor U6098 (N_6098,N_5886,N_4717);
and U6099 (N_6099,N_5674,N_3168);
or U6100 (N_6100,N_5103,N_3318);
or U6101 (N_6101,N_3054,N_3942);
nor U6102 (N_6102,N_4231,N_3668);
or U6103 (N_6103,N_5896,N_3946);
or U6104 (N_6104,N_4670,N_3217);
or U6105 (N_6105,N_4496,N_3062);
xor U6106 (N_6106,N_4101,N_3855);
and U6107 (N_6107,N_5393,N_4021);
and U6108 (N_6108,N_5337,N_4699);
and U6109 (N_6109,N_3611,N_4754);
nor U6110 (N_6110,N_3298,N_3705);
nand U6111 (N_6111,N_5808,N_5583);
nand U6112 (N_6112,N_5298,N_3274);
and U6113 (N_6113,N_4156,N_3760);
nand U6114 (N_6114,N_5144,N_3295);
and U6115 (N_6115,N_4928,N_5389);
nand U6116 (N_6116,N_3067,N_3947);
xor U6117 (N_6117,N_4813,N_3880);
nand U6118 (N_6118,N_3108,N_4967);
and U6119 (N_6119,N_3122,N_3590);
or U6120 (N_6120,N_5092,N_4308);
nor U6121 (N_6121,N_4422,N_5459);
nand U6122 (N_6122,N_4121,N_3783);
and U6123 (N_6123,N_3378,N_5567);
nor U6124 (N_6124,N_3877,N_3222);
or U6125 (N_6125,N_5588,N_3101);
nor U6126 (N_6126,N_3431,N_5518);
or U6127 (N_6127,N_4032,N_4990);
or U6128 (N_6128,N_5936,N_5712);
and U6129 (N_6129,N_5319,N_4049);
nor U6130 (N_6130,N_4942,N_4098);
nor U6131 (N_6131,N_3767,N_3171);
or U6132 (N_6132,N_4785,N_5898);
xnor U6133 (N_6133,N_3539,N_4215);
nor U6134 (N_6134,N_3657,N_3701);
xor U6135 (N_6135,N_3644,N_4932);
xnor U6136 (N_6136,N_3421,N_3100);
nand U6137 (N_6137,N_3824,N_5925);
nor U6138 (N_6138,N_5863,N_4096);
nand U6139 (N_6139,N_4269,N_4104);
or U6140 (N_6140,N_3019,N_5805);
nor U6141 (N_6141,N_4493,N_5636);
xnor U6142 (N_6142,N_5490,N_4980);
or U6143 (N_6143,N_3014,N_3888);
nand U6144 (N_6144,N_5698,N_4662);
and U6145 (N_6145,N_3157,N_3675);
nand U6146 (N_6146,N_3973,N_3710);
xor U6147 (N_6147,N_4508,N_4148);
nor U6148 (N_6148,N_4110,N_3670);
and U6149 (N_6149,N_5186,N_5620);
nor U6150 (N_6150,N_4673,N_5501);
and U6151 (N_6151,N_5630,N_5961);
nor U6152 (N_6152,N_4373,N_5892);
nand U6153 (N_6153,N_3397,N_5212);
xnor U6154 (N_6154,N_5035,N_4407);
or U6155 (N_6155,N_3195,N_3736);
nand U6156 (N_6156,N_5766,N_5201);
xor U6157 (N_6157,N_4486,N_4594);
xnor U6158 (N_6158,N_3984,N_5245);
and U6159 (N_6159,N_4707,N_4939);
xor U6160 (N_6160,N_4157,N_4816);
nand U6161 (N_6161,N_5731,N_5803);
xor U6162 (N_6162,N_3304,N_5645);
and U6163 (N_6163,N_5474,N_4626);
nor U6164 (N_6164,N_4645,N_3409);
or U6165 (N_6165,N_3651,N_4258);
nand U6166 (N_6166,N_3583,N_4572);
and U6167 (N_6167,N_3368,N_5590);
xor U6168 (N_6168,N_5923,N_3391);
and U6169 (N_6169,N_5087,N_4408);
and U6170 (N_6170,N_4327,N_3846);
xnor U6171 (N_6171,N_3545,N_3927);
and U6172 (N_6172,N_3548,N_3897);
and U6173 (N_6173,N_5757,N_4970);
nor U6174 (N_6174,N_3754,N_4881);
xnor U6175 (N_6175,N_3104,N_4489);
xnor U6176 (N_6176,N_3130,N_4500);
xor U6177 (N_6177,N_3037,N_5344);
nand U6178 (N_6178,N_3661,N_4708);
or U6179 (N_6179,N_4085,N_4544);
nand U6180 (N_6180,N_3805,N_3970);
or U6181 (N_6181,N_5689,N_3331);
and U6182 (N_6182,N_5121,N_3870);
nand U6183 (N_6183,N_3874,N_5093);
and U6184 (N_6184,N_4301,N_4807);
nor U6185 (N_6185,N_5489,N_4204);
or U6186 (N_6186,N_3528,N_3856);
xor U6187 (N_6187,N_3994,N_4826);
and U6188 (N_6188,N_5555,N_4586);
nor U6189 (N_6189,N_4938,N_4611);
or U6190 (N_6190,N_5659,N_3572);
xor U6191 (N_6191,N_4162,N_3107);
xor U6192 (N_6192,N_5777,N_3127);
and U6193 (N_6193,N_3681,N_3589);
or U6194 (N_6194,N_5605,N_4067);
and U6195 (N_6195,N_5246,N_5976);
nor U6196 (N_6196,N_3703,N_5379);
xnor U6197 (N_6197,N_3292,N_5066);
and U6198 (N_6198,N_4302,N_4288);
nor U6199 (N_6199,N_3992,N_3938);
and U6200 (N_6200,N_3782,N_5804);
xnor U6201 (N_6201,N_3616,N_5563);
nor U6202 (N_6202,N_3993,N_3297);
nand U6203 (N_6203,N_4394,N_5694);
and U6204 (N_6204,N_3480,N_5668);
xor U6205 (N_6205,N_5989,N_5112);
nor U6206 (N_6206,N_4925,N_4563);
or U6207 (N_6207,N_4575,N_4455);
and U6208 (N_6208,N_5509,N_4420);
or U6209 (N_6209,N_5133,N_4599);
or U6210 (N_6210,N_4569,N_5293);
and U6211 (N_6211,N_5830,N_3356);
nand U6212 (N_6212,N_3951,N_3123);
and U6213 (N_6213,N_3812,N_3945);
nand U6214 (N_6214,N_5366,N_5797);
and U6215 (N_6215,N_5942,N_5747);
and U6216 (N_6216,N_5175,N_4690);
or U6217 (N_6217,N_5340,N_3384);
or U6218 (N_6218,N_3857,N_5530);
and U6219 (N_6219,N_4718,N_3096);
nand U6220 (N_6220,N_3392,N_5054);
or U6221 (N_6221,N_3511,N_3150);
or U6222 (N_6222,N_3631,N_4798);
xnor U6223 (N_6223,N_5342,N_3620);
and U6224 (N_6224,N_4593,N_5994);
xor U6225 (N_6225,N_4333,N_5498);
and U6226 (N_6226,N_4184,N_5428);
and U6227 (N_6227,N_3428,N_4988);
nand U6228 (N_6228,N_5755,N_3003);
xnor U6229 (N_6229,N_3309,N_3596);
xnor U6230 (N_6230,N_5917,N_4644);
or U6231 (N_6231,N_3519,N_3135);
xnor U6232 (N_6232,N_3141,N_4960);
and U6233 (N_6233,N_5003,N_3922);
or U6234 (N_6234,N_5650,N_5594);
nand U6235 (N_6235,N_3876,N_5924);
or U6236 (N_6236,N_4030,N_3200);
xnor U6237 (N_6237,N_5970,N_4535);
or U6238 (N_6238,N_4409,N_5656);
nand U6239 (N_6239,N_5921,N_5361);
and U6240 (N_6240,N_3402,N_5380);
and U6241 (N_6241,N_4300,N_4780);
or U6242 (N_6242,N_3450,N_4884);
nand U6243 (N_6243,N_3998,N_4653);
xnor U6244 (N_6244,N_3883,N_3678);
and U6245 (N_6245,N_4709,N_3580);
and U6246 (N_6246,N_5665,N_5104);
or U6247 (N_6247,N_3607,N_3591);
nand U6248 (N_6248,N_5398,N_5649);
nand U6249 (N_6249,N_4364,N_4371);
nor U6250 (N_6250,N_5939,N_4655);
nand U6251 (N_6251,N_3281,N_5524);
and U6252 (N_6252,N_4433,N_3854);
or U6253 (N_6253,N_3890,N_5106);
nand U6254 (N_6254,N_3686,N_4277);
xnor U6255 (N_6255,N_3677,N_4392);
xnor U6256 (N_6256,N_4609,N_5690);
and U6257 (N_6257,N_4472,N_4546);
or U6258 (N_6258,N_5758,N_5703);
and U6259 (N_6259,N_5284,N_3893);
nor U6260 (N_6260,N_3080,N_4223);
nand U6261 (N_6261,N_3711,N_4395);
or U6262 (N_6262,N_5161,N_4566);
and U6263 (N_6263,N_4237,N_5868);
nor U6264 (N_6264,N_4839,N_4272);
xor U6265 (N_6265,N_5934,N_3790);
nand U6266 (N_6266,N_5914,N_3878);
xor U6267 (N_6267,N_3405,N_4167);
or U6268 (N_6268,N_3155,N_5331);
or U6269 (N_6269,N_3273,N_4198);
nand U6270 (N_6270,N_4444,N_4908);
or U6271 (N_6271,N_4956,N_3940);
xnor U6272 (N_6272,N_3555,N_5079);
and U6273 (N_6273,N_4834,N_4811);
nor U6274 (N_6274,N_4959,N_4310);
nand U6275 (N_6275,N_4802,N_3972);
nor U6276 (N_6276,N_3406,N_3099);
nor U6277 (N_6277,N_3779,N_3799);
xnor U6278 (N_6278,N_3410,N_3546);
nor U6279 (N_6279,N_5154,N_3110);
and U6280 (N_6280,N_5508,N_3839);
or U6281 (N_6281,N_4052,N_3278);
and U6282 (N_6282,N_4628,N_5495);
and U6283 (N_6283,N_5172,N_4504);
xnor U6284 (N_6284,N_4646,N_4485);
nand U6285 (N_6285,N_3334,N_5675);
or U6286 (N_6286,N_3682,N_3694);
or U6287 (N_6287,N_5843,N_4830);
or U6288 (N_6288,N_5454,N_3720);
and U6289 (N_6289,N_4497,N_4692);
xnor U6290 (N_6290,N_3755,N_4250);
nor U6291 (N_6291,N_5954,N_3366);
xnor U6292 (N_6292,N_3321,N_3319);
or U6293 (N_6293,N_5360,N_3351);
or U6294 (N_6294,N_4380,N_3192);
or U6295 (N_6295,N_3565,N_4099);
or U6296 (N_6296,N_3902,N_4211);
nand U6297 (N_6297,N_5915,N_4913);
or U6298 (N_6298,N_3484,N_5666);
nand U6299 (N_6299,N_5810,N_3087);
or U6300 (N_6300,N_4765,N_4117);
nand U6301 (N_6301,N_4057,N_4994);
xnor U6302 (N_6302,N_4635,N_4304);
xor U6303 (N_6303,N_4916,N_5377);
and U6304 (N_6304,N_4965,N_5388);
xnor U6305 (N_6305,N_5480,N_5335);
or U6306 (N_6306,N_4298,N_3291);
and U6307 (N_6307,N_3551,N_4159);
or U6308 (N_6308,N_3093,N_4756);
xor U6309 (N_6309,N_3513,N_3203);
and U6310 (N_6310,N_3197,N_3345);
and U6311 (N_6311,N_4886,N_4501);
and U6312 (N_6312,N_3072,N_5683);
nor U6313 (N_6313,N_5764,N_5623);
nand U6314 (N_6314,N_3317,N_5171);
nor U6315 (N_6315,N_5629,N_3925);
nand U6316 (N_6316,N_3018,N_5083);
nand U6317 (N_6317,N_4948,N_5523);
nand U6318 (N_6318,N_5252,N_5363);
xnor U6319 (N_6319,N_4689,N_3362);
nand U6320 (N_6320,N_5510,N_4782);
nand U6321 (N_6321,N_4081,N_5985);
xnor U6322 (N_6322,N_5394,N_4034);
and U6323 (N_6323,N_3688,N_4256);
xnor U6324 (N_6324,N_4318,N_4090);
nor U6325 (N_6325,N_4390,N_5918);
nor U6326 (N_6326,N_3959,N_4031);
xor U6327 (N_6327,N_4362,N_4700);
xor U6328 (N_6328,N_5254,N_5981);
xor U6329 (N_6329,N_4010,N_4289);
and U6330 (N_6330,N_4677,N_5053);
xnor U6331 (N_6331,N_5145,N_3559);
nor U6332 (N_6332,N_5565,N_3592);
and U6333 (N_6333,N_4864,N_4545);
and U6334 (N_6334,N_3806,N_4158);
or U6335 (N_6335,N_3522,N_4825);
nor U6336 (N_6336,N_5557,N_4674);
nand U6337 (N_6337,N_5466,N_4694);
nor U6338 (N_6338,N_3829,N_5435);
nand U6339 (N_6339,N_3588,N_3464);
or U6340 (N_6340,N_4428,N_5176);
nand U6341 (N_6341,N_4606,N_3040);
nand U6342 (N_6342,N_3045,N_3777);
xor U6343 (N_6343,N_5806,N_5927);
xor U6344 (N_6344,N_4622,N_5960);
or U6345 (N_6345,N_5317,N_5835);
xnor U6346 (N_6346,N_5032,N_3626);
and U6347 (N_6347,N_4770,N_4867);
xor U6348 (N_6348,N_3769,N_5152);
or U6349 (N_6349,N_5858,N_3512);
or U6350 (N_6350,N_4165,N_4490);
and U6351 (N_6351,N_4388,N_3801);
xnor U6352 (N_6352,N_4634,N_4105);
xnor U6353 (N_6353,N_3656,N_4372);
and U6354 (N_6354,N_3185,N_5058);
and U6355 (N_6355,N_3407,N_4190);
and U6356 (N_6356,N_3000,N_3139);
or U6357 (N_6357,N_3357,N_3057);
nand U6358 (N_6358,N_3071,N_4402);
nor U6359 (N_6359,N_4335,N_3862);
nand U6360 (N_6360,N_5546,N_5333);
xnor U6361 (N_6361,N_4658,N_4194);
or U6362 (N_6362,N_3928,N_5191);
xor U6363 (N_6363,N_5677,N_4352);
and U6364 (N_6364,N_3152,N_4801);
nor U6365 (N_6365,N_4549,N_3941);
nor U6366 (N_6366,N_3269,N_5752);
and U6367 (N_6367,N_5948,N_4132);
nor U6368 (N_6368,N_5531,N_5431);
nor U6369 (N_6369,N_5427,N_5792);
nor U6370 (N_6370,N_5932,N_3765);
nor U6371 (N_6371,N_3237,N_5125);
xnor U6372 (N_6372,N_3447,N_4640);
or U6373 (N_6373,N_5351,N_4449);
nand U6374 (N_6374,N_3955,N_5446);
nand U6375 (N_6375,N_3898,N_5597);
xnor U6376 (N_6376,N_4779,N_5070);
and U6377 (N_6377,N_5911,N_3886);
nor U6378 (N_6378,N_4312,N_5306);
nor U6379 (N_6379,N_5483,N_3208);
xnor U6380 (N_6380,N_3741,N_4177);
or U6381 (N_6381,N_3165,N_4226);
and U6382 (N_6382,N_5268,N_5815);
and U6383 (N_6383,N_4212,N_3470);
or U6384 (N_6384,N_4130,N_3467);
nor U6385 (N_6385,N_4998,N_4656);
nand U6386 (N_6386,N_5403,N_4072);
xnor U6387 (N_6387,N_3349,N_5571);
xnor U6388 (N_6388,N_5525,N_3056);
or U6389 (N_6389,N_4136,N_5006);
nor U6390 (N_6390,N_4592,N_4075);
nor U6391 (N_6391,N_4239,N_4411);
nor U6392 (N_6392,N_5094,N_3717);
and U6393 (N_6393,N_5204,N_4800);
xnor U6394 (N_6394,N_3674,N_5956);
nand U6395 (N_6395,N_3634,N_3284);
xnor U6396 (N_6396,N_4235,N_4792);
or U6397 (N_6397,N_4589,N_5085);
nor U6398 (N_6398,N_3229,N_4650);
or U6399 (N_6399,N_4147,N_5648);
or U6400 (N_6400,N_4435,N_4940);
or U6401 (N_6401,N_5718,N_4080);
nand U6402 (N_6402,N_3089,N_4897);
xnor U6403 (N_6403,N_5464,N_4011);
nand U6404 (N_6404,N_4915,N_5408);
nor U6405 (N_6405,N_4513,N_3495);
nand U6406 (N_6406,N_5206,N_5641);
and U6407 (N_6407,N_3859,N_5946);
xor U6408 (N_6408,N_5553,N_5734);
or U6409 (N_6409,N_5281,N_4170);
nand U6410 (N_6410,N_3383,N_4933);
and U6411 (N_6411,N_4866,N_4964);
nand U6412 (N_6412,N_3290,N_5062);
or U6413 (N_6413,N_3847,N_4732);
xnor U6414 (N_6414,N_3212,N_3361);
nand U6415 (N_6415,N_4815,N_4452);
nand U6416 (N_6416,N_4637,N_5912);
xor U6417 (N_6417,N_3215,N_4838);
and U6418 (N_6418,N_5568,N_4767);
xnor U6419 (N_6419,N_3882,N_5045);
or U6420 (N_6420,N_3140,N_5415);
nand U6421 (N_6421,N_3871,N_3568);
xor U6422 (N_6422,N_4614,N_3696);
and U6423 (N_6423,N_4541,N_5325);
xnor U6424 (N_6424,N_5199,N_4590);
and U6425 (N_6425,N_5330,N_4273);
nand U6426 (N_6426,N_3137,N_3027);
xnor U6427 (N_6427,N_3618,N_3709);
or U6428 (N_6428,N_3554,N_3786);
and U6429 (N_6429,N_5682,N_3896);
nor U6430 (N_6430,N_4507,N_3243);
or U6431 (N_6431,N_3923,N_4337);
or U6432 (N_6432,N_4654,N_4381);
and U6433 (N_6433,N_5552,N_4672);
and U6434 (N_6434,N_4214,N_5442);
nor U6435 (N_6435,N_5479,N_4898);
xor U6436 (N_6436,N_3427,N_5535);
and U6437 (N_6437,N_3451,N_4671);
and U6438 (N_6438,N_5762,N_3216);
nor U6439 (N_6439,N_5405,N_4303);
or U6440 (N_6440,N_3194,N_5320);
xnor U6441 (N_6441,N_5478,N_5990);
xnor U6442 (N_6442,N_3094,N_4003);
or U6443 (N_6443,N_3493,N_4721);
and U6444 (N_6444,N_5732,N_4876);
xnor U6445 (N_6445,N_3933,N_4934);
nor U6446 (N_6446,N_5140,N_4284);
xor U6447 (N_6447,N_3732,N_4931);
nand U6448 (N_6448,N_4025,N_4358);
or U6449 (N_6449,N_5496,N_4112);
and U6450 (N_6450,N_5108,N_5467);
nor U6451 (N_6451,N_4195,N_4062);
or U6452 (N_6452,N_3619,N_4977);
nor U6453 (N_6453,N_5862,N_5365);
nor U6454 (N_6454,N_5716,N_3266);
nor U6455 (N_6455,N_5748,N_4216);
or U6456 (N_6456,N_4855,N_5561);
or U6457 (N_6457,N_3248,N_4753);
or U6458 (N_6458,N_3601,N_4747);
xnor U6459 (N_6459,N_3912,N_3420);
xor U6460 (N_6460,N_4179,N_5704);
or U6461 (N_6461,N_4877,N_5075);
or U6462 (N_6462,N_4363,N_3417);
nand U6463 (N_6463,N_5647,N_5321);
nor U6464 (N_6464,N_5705,N_5135);
or U6465 (N_6465,N_4841,N_3202);
or U6466 (N_6466,N_5780,N_5433);
xnor U6467 (N_6467,N_3977,N_3884);
nor U6468 (N_6468,N_5681,N_5827);
or U6469 (N_6469,N_3434,N_5957);
or U6470 (N_6470,N_3652,N_5782);
or U6471 (N_6471,N_4728,N_4385);
or U6472 (N_6472,N_4506,N_4679);
nor U6473 (N_6473,N_3347,N_5534);
and U6474 (N_6474,N_5795,N_3489);
nor U6475 (N_6475,N_5151,N_3225);
nor U6476 (N_6476,N_3198,N_4332);
or U6477 (N_6477,N_5944,N_3307);
xnor U6478 (N_6478,N_3116,N_5099);
and U6479 (N_6479,N_3996,N_3508);
nor U6480 (N_6480,N_3774,N_5639);
nand U6481 (N_6481,N_5038,N_3939);
or U6482 (N_6482,N_4518,N_3460);
nor U6483 (N_6483,N_5548,N_4271);
or U6484 (N_6484,N_3990,N_5584);
or U6485 (N_6485,N_5369,N_3214);
and U6486 (N_6486,N_4168,N_3158);
xnor U6487 (N_6487,N_4232,N_5850);
nor U6488 (N_6488,N_3264,N_3693);
and U6489 (N_6489,N_5027,N_5071);
nand U6490 (N_6490,N_3569,N_5481);
and U6491 (N_6491,N_5975,N_3575);
or U6492 (N_6492,N_3147,N_4209);
xor U6493 (N_6493,N_4114,N_3289);
and U6494 (N_6494,N_4491,N_4750);
or U6495 (N_6495,N_4008,N_4896);
and U6496 (N_6496,N_3989,N_4446);
nor U6497 (N_6497,N_3453,N_4639);
xnor U6498 (N_6498,N_3429,N_3835);
xor U6499 (N_6499,N_5364,N_5796);
nand U6500 (N_6500,N_3544,N_4818);
nor U6501 (N_6501,N_4532,N_4343);
nand U6502 (N_6502,N_4066,N_4585);
xnor U6503 (N_6503,N_3265,N_4949);
nand U6504 (N_6504,N_3924,N_5110);
and U6505 (N_6505,N_3663,N_3504);
and U6506 (N_6506,N_3937,N_3556);
and U6507 (N_6507,N_5357,N_4421);
nand U6508 (N_6508,N_3179,N_3456);
xor U6509 (N_6509,N_3006,N_4118);
xor U6510 (N_6510,N_5273,N_5349);
nand U6511 (N_6511,N_4976,N_3075);
or U6512 (N_6512,N_4113,N_4329);
nand U6513 (N_6513,N_5156,N_5001);
nor U6514 (N_6514,N_3932,N_4181);
and U6515 (N_6515,N_4892,N_3314);
nand U6516 (N_6516,N_4503,N_4427);
nand U6517 (N_6517,N_3794,N_3604);
and U6518 (N_6518,N_5385,N_4068);
nor U6519 (N_6519,N_5695,N_3105);
and U6520 (N_6520,N_3031,N_5715);
nor U6521 (N_6521,N_4039,N_5680);
xor U6522 (N_6522,N_3136,N_3388);
or U6523 (N_6523,N_5516,N_4744);
or U6524 (N_6524,N_5223,N_5148);
or U6525 (N_6525,N_4262,N_3043);
xnor U6526 (N_6526,N_5746,N_5906);
nand U6527 (N_6527,N_5322,N_3308);
xnor U6528 (N_6528,N_3224,N_5878);
or U6529 (N_6529,N_5033,N_5599);
or U6530 (N_6530,N_5801,N_4533);
and U6531 (N_6531,N_5816,N_3443);
xnor U6532 (N_6532,N_4142,N_4840);
nand U6533 (N_6533,N_4937,N_4955);
and U6534 (N_6534,N_5067,N_5520);
nand U6535 (N_6535,N_3520,N_5618);
or U6536 (N_6536,N_4641,N_4505);
nand U6537 (N_6537,N_5115,N_3471);
nand U6538 (N_6538,N_3869,N_4257);
nor U6539 (N_6539,N_3302,N_5726);
nand U6540 (N_6540,N_4981,N_4597);
and U6541 (N_6541,N_4773,N_4849);
nor U6542 (N_6542,N_5010,N_3412);
and U6543 (N_6543,N_5697,N_4553);
nor U6544 (N_6544,N_5100,N_3594);
nor U6545 (N_6545,N_3086,N_5974);
xnor U6546 (N_6546,N_3069,N_3377);
or U6547 (N_6547,N_5371,N_4993);
nand U6548 (N_6548,N_5005,N_3895);
nor U6549 (N_6549,N_5776,N_4017);
nand U6550 (N_6550,N_5971,N_4768);
xor U6551 (N_6551,N_4322,N_4923);
and U6552 (N_6552,N_4281,N_3844);
nand U6553 (N_6553,N_4100,N_4244);
and U6554 (N_6554,N_4468,N_3971);
xor U6555 (N_6555,N_3461,N_3436);
or U6556 (N_6556,N_4094,N_5933);
xnor U6557 (N_6557,N_5308,N_5761);
and U6558 (N_6558,N_5713,N_5595);
and U6559 (N_6559,N_5484,N_3650);
nand U6560 (N_6560,N_5547,N_4848);
nand U6561 (N_6561,N_4704,N_3403);
nand U6562 (N_6562,N_5725,N_3763);
nand U6563 (N_6563,N_3360,N_3578);
and U6564 (N_6564,N_4169,N_4548);
nand U6565 (N_6565,N_4199,N_5631);
and U6566 (N_6566,N_5708,N_3126);
and U6567 (N_6567,N_3804,N_5591);
or U6568 (N_6568,N_3787,N_3133);
or U6569 (N_6569,N_5802,N_5673);
xor U6570 (N_6570,N_4396,N_5536);
nand U6571 (N_6571,N_3142,N_5515);
xnor U6572 (N_6572,N_3444,N_3227);
or U6573 (N_6573,N_5632,N_4680);
nor U6574 (N_6574,N_3485,N_5754);
nor U6575 (N_6575,N_3577,N_4401);
and U6576 (N_6576,N_3770,N_5891);
xor U6577 (N_6577,N_4082,N_5300);
or U6578 (N_6578,N_3324,N_3007);
nand U6579 (N_6579,N_3481,N_5875);
and U6580 (N_6580,N_5019,N_4038);
nor U6581 (N_6581,N_4920,N_3584);
or U6582 (N_6582,N_4120,N_5026);
nand U6583 (N_6583,N_5635,N_4643);
xnor U6584 (N_6584,N_5719,N_5126);
nand U6585 (N_6585,N_3389,N_3159);
xor U6586 (N_6586,N_3365,N_4014);
and U6587 (N_6587,N_3991,N_5096);
xnor U6588 (N_6588,N_3465,N_5662);
nand U6589 (N_6589,N_5608,N_5336);
and U6590 (N_6590,N_4474,N_4828);
or U6591 (N_6591,N_5313,N_3279);
nor U6592 (N_6592,N_3603,N_4758);
xnor U6593 (N_6593,N_4419,N_5159);
and U6594 (N_6594,N_4050,N_5544);
nor U6595 (N_6595,N_4279,N_3654);
nand U6596 (N_6596,N_5854,N_5375);
nand U6597 (N_6597,N_5485,N_4796);
nand U6598 (N_6598,N_5910,N_5562);
and U6599 (N_6599,N_4527,N_3160);
nor U6600 (N_6600,N_4607,N_4040);
nand U6601 (N_6601,N_3593,N_3561);
nand U6602 (N_6602,N_3490,N_3015);
nand U6603 (N_6603,N_5132,N_3585);
or U6604 (N_6604,N_4097,N_4664);
and U6605 (N_6605,N_5270,N_3088);
or U6606 (N_6606,N_4370,N_5461);
and U6607 (N_6607,N_5029,N_4880);
nand U6608 (N_6608,N_5416,N_4885);
nor U6609 (N_6609,N_5289,N_4820);
nor U6610 (N_6610,N_5737,N_4889);
nand U6611 (N_6611,N_3424,N_4957);
or U6612 (N_6612,N_4192,N_5147);
nor U6613 (N_6613,N_5160,N_3497);
nor U6614 (N_6614,N_5105,N_5966);
nor U6615 (N_6615,N_4509,N_4495);
or U6616 (N_6616,N_4145,N_3299);
nor U6617 (N_6617,N_5000,N_5052);
nor U6618 (N_6618,N_3949,N_3496);
and U6619 (N_6619,N_5170,N_5685);
and U6620 (N_6620,N_5107,N_4726);
or U6621 (N_6621,N_4969,N_5696);
or U6622 (N_6622,N_3386,N_3207);
and U6623 (N_6623,N_5291,N_4781);
or U6624 (N_6624,N_4883,N_3413);
xor U6625 (N_6625,N_5114,N_4354);
and U6626 (N_6626,N_3364,N_3113);
nand U6627 (N_6627,N_3375,N_4425);
xor U6628 (N_6628,N_3506,N_4974);
or U6629 (N_6629,N_3293,N_3363);
nor U6630 (N_6630,N_3146,N_4458);
or U6631 (N_6631,N_3549,N_5222);
xnor U6632 (N_6632,N_4160,N_5768);
nand U6633 (N_6633,N_4412,N_5076);
nand U6634 (N_6634,N_5141,N_4405);
or U6635 (N_6635,N_5157,N_4738);
xor U6636 (N_6636,N_3542,N_3191);
nor U6637 (N_6637,N_3457,N_5443);
nor U6638 (N_6638,N_3352,N_4598);
xor U6639 (N_6639,N_5573,N_5541);
and U6640 (N_6640,N_3891,N_5242);
or U6641 (N_6641,N_4398,N_5769);
xnor U6642 (N_6642,N_4795,N_5049);
or U6643 (N_6643,N_3673,N_3621);
xnor U6644 (N_6644,N_4835,N_5823);
or U6645 (N_6645,N_5771,N_3624);
nand U6646 (N_6646,N_3502,N_4002);
or U6647 (N_6647,N_5168,N_5150);
nor U6648 (N_6648,N_5845,N_3550);
nor U6649 (N_6649,N_5277,N_3962);
xnor U6650 (N_6650,N_5538,N_3726);
nor U6651 (N_6651,N_5717,N_5303);
nor U6652 (N_6652,N_3538,N_5286);
and U6653 (N_6653,N_5384,N_4763);
and U6654 (N_6654,N_3011,N_5015);
nand U6655 (N_6655,N_4360,N_4429);
or U6656 (N_6656,N_5213,N_3605);
and U6657 (N_6657,N_3335,N_4384);
nand U6658 (N_6658,N_5569,N_5211);
and U6659 (N_6659,N_5865,N_5158);
and U6660 (N_6660,N_3735,N_5128);
nor U6661 (N_6661,N_3441,N_3132);
nand U6662 (N_6662,N_4755,N_4986);
and U6663 (N_6663,N_5414,N_4171);
nor U6664 (N_6664,N_5542,N_3232);
nand U6665 (N_6665,N_4806,N_5074);
xor U6666 (N_6666,N_4962,N_3756);
and U6667 (N_6667,N_5676,N_4536);
and U6668 (N_6668,N_4382,N_4788);
xnor U6669 (N_6669,N_4483,N_4297);
or U6670 (N_6670,N_3048,N_3380);
nor U6671 (N_6671,N_5625,N_3954);
nand U6672 (N_6672,N_3164,N_4847);
or U6673 (N_6673,N_5169,N_3983);
nand U6674 (N_6674,N_5884,N_3630);
nor U6675 (N_6675,N_5039,N_5280);
and U6676 (N_6676,N_5355,N_5821);
nor U6677 (N_6677,N_5486,N_4456);
nand U6678 (N_6678,N_4374,N_5869);
xor U6679 (N_6679,N_5503,N_3781);
or U6680 (N_6680,N_4636,N_5740);
xor U6681 (N_6681,N_3401,N_4175);
xor U6682 (N_6682,N_4582,N_4183);
nor U6683 (N_6683,N_5226,N_4642);
nor U6684 (N_6684,N_4579,N_5476);
xnor U6685 (N_6685,N_3814,N_3817);
xor U6686 (N_6686,N_4074,N_5009);
nor U6687 (N_6687,N_4817,N_5642);
or U6688 (N_6688,N_5130,N_5205);
xor U6689 (N_6689,N_5274,N_5903);
xnor U6690 (N_6690,N_4437,N_5860);
and U6691 (N_6691,N_4982,N_5413);
nand U6692 (N_6692,N_3843,N_3190);
or U6693 (N_6693,N_4270,N_4059);
nand U6694 (N_6694,N_4185,N_5842);
and U6695 (N_6695,N_3529,N_3109);
nand U6696 (N_6696,N_4228,N_4448);
nor U6697 (N_6697,N_4748,N_5312);
nand U6698 (N_6698,N_4851,N_3287);
or U6699 (N_6699,N_4447,N_5822);
nor U6700 (N_6700,N_3714,N_3653);
nor U6701 (N_6701,N_4953,N_3785);
or U6702 (N_6702,N_3476,N_3022);
and U6703 (N_6703,N_5958,N_5447);
nand U6704 (N_6704,N_3739,N_3798);
nor U6705 (N_6705,N_4751,N_3636);
or U6706 (N_6706,N_3333,N_3134);
or U6707 (N_6707,N_5334,N_5596);
nor U6708 (N_6708,N_3976,N_3042);
nor U6709 (N_6709,N_3501,N_3263);
or U6710 (N_6710,N_4542,N_3235);
nor U6711 (N_6711,N_4345,N_5800);
xor U6712 (N_6712,N_5578,N_3762);
and U6713 (N_6713,N_5352,N_4294);
nand U6714 (N_6714,N_4328,N_5091);
and U6715 (N_6715,N_4789,N_3813);
nor U6716 (N_6716,N_4743,N_5068);
nand U6717 (N_6717,N_4109,N_4905);
nor U6718 (N_6718,N_3012,N_3646);
xor U6719 (N_6719,N_5056,N_4164);
and U6720 (N_6720,N_4295,N_3887);
or U6721 (N_6721,N_4152,N_4899);
or U6722 (N_6722,N_5962,N_3381);
and U6723 (N_6723,N_5577,N_4020);
nor U6724 (N_6724,N_4338,N_3306);
xor U6725 (N_6725,N_4365,N_4777);
and U6726 (N_6726,N_5462,N_3599);
nor U6727 (N_6727,N_5376,N_4574);
and U6728 (N_6728,N_5082,N_4987);
and U6729 (N_6729,N_5095,N_5880);
nand U6730 (N_6730,N_5772,N_5283);
and U6731 (N_6731,N_4227,N_3967);
nand U6732 (N_6732,N_5907,N_4827);
xnor U6733 (N_6733,N_5572,N_5955);
and U6734 (N_6734,N_5233,N_5438);
or U6735 (N_6735,N_3068,N_4375);
or U6736 (N_6736,N_5855,N_3753);
or U6737 (N_6737,N_5877,N_3968);
or U6738 (N_6738,N_4695,N_5602);
and U6739 (N_6739,N_4879,N_4457);
nor U6740 (N_6740,N_3323,N_5028);
xor U6741 (N_6741,N_4676,N_3904);
nand U6742 (N_6742,N_3074,N_4711);
nand U6743 (N_6743,N_4477,N_4725);
nor U6744 (N_6744,N_3622,N_3341);
nor U6745 (N_6745,N_4467,N_3058);
or U6746 (N_6746,N_4403,N_3979);
nor U6747 (N_6747,N_5370,N_3713);
nand U6748 (N_6748,N_5814,N_3499);
or U6749 (N_6749,N_5833,N_3664);
or U6750 (N_6750,N_3908,N_4203);
or U6751 (N_6751,N_3910,N_5904);
or U6752 (N_6752,N_5400,N_5190);
nand U6753 (N_6753,N_4106,N_5988);
or U6754 (N_6754,N_5208,N_5470);
and U6755 (N_6755,N_3564,N_5220);
nor U6756 (N_6756,N_3879,N_5350);
and U6757 (N_6757,N_5440,N_5943);
or U6758 (N_6758,N_3004,N_4317);
or U6759 (N_6759,N_5753,N_3514);
nand U6760 (N_6760,N_3469,N_4914);
and U6761 (N_6761,N_3242,N_5214);
or U6762 (N_6762,N_5016,N_5853);
xnor U6763 (N_6763,N_3246,N_5282);
nor U6764 (N_6764,N_4037,N_3328);
or U6765 (N_6765,N_4910,N_5276);
nor U6766 (N_6766,N_3486,N_5228);
or U6767 (N_6767,N_4028,N_5069);
or U6768 (N_6768,N_3842,N_4919);
nor U6769 (N_6769,N_3326,N_5077);
or U6770 (N_6770,N_5652,N_3055);
or U6771 (N_6771,N_4024,N_4805);
nor U6772 (N_6772,N_5143,N_5051);
and U6773 (N_6773,N_4907,N_4029);
nor U6774 (N_6774,N_5219,N_5589);
or U6775 (N_6775,N_5165,N_5897);
xor U6776 (N_6776,N_4882,N_4722);
nor U6777 (N_6777,N_5720,N_4961);
nor U6778 (N_6778,N_4376,N_5672);
or U6779 (N_6779,N_3254,N_4863);
or U6780 (N_6780,N_5908,N_3026);
nand U6781 (N_6781,N_5837,N_4570);
or U6782 (N_6782,N_4617,N_5728);
or U6783 (N_6783,N_4344,N_5013);
or U6784 (N_6784,N_4772,N_4033);
and U6785 (N_6785,N_3953,N_4543);
nand U6786 (N_6786,N_5874,N_5494);
and U6787 (N_6787,N_3926,N_3964);
nor U6788 (N_6788,N_5644,N_4259);
nand U6789 (N_6789,N_4296,N_4610);
nor U6790 (N_6790,N_3111,N_5297);
and U6791 (N_6791,N_5353,N_4391);
nand U6792 (N_6792,N_3166,N_4512);
nor U6793 (N_6793,N_3745,N_5521);
or U6794 (N_6794,N_5550,N_5811);
nor U6795 (N_6795,N_3515,N_4249);
nand U6796 (N_6796,N_5679,N_3228);
and U6797 (N_6797,N_3655,N_3353);
or U6798 (N_6798,N_4688,N_4652);
nor U6799 (N_6799,N_4742,N_3818);
nand U6800 (N_6800,N_4584,N_5315);
xnor U6801 (N_6801,N_4891,N_4006);
and U6802 (N_6802,N_4946,N_5081);
xnor U6803 (N_6803,N_4494,N_3598);
or U6804 (N_6804,N_5870,N_3563);
nand U6805 (N_6805,N_5166,N_3029);
xnor U6806 (N_6806,N_5972,N_4036);
nor U6807 (N_6807,N_3256,N_4070);
or U6808 (N_6808,N_4735,N_4698);
and U6809 (N_6809,N_5579,N_3828);
or U6810 (N_6810,N_5258,N_3680);
or U6811 (N_6811,N_5272,N_5059);
nand U6812 (N_6812,N_5527,N_5603);
xor U6813 (N_6813,N_4012,N_4760);
xnor U6814 (N_6814,N_4291,N_4958);
nor U6815 (N_6815,N_4736,N_4859);
or U6816 (N_6816,N_4389,N_5146);
or U6817 (N_6817,N_5612,N_3800);
xor U6818 (N_6818,N_4154,N_5316);
or U6819 (N_6819,N_3503,N_5537);
or U6820 (N_6820,N_5751,N_5127);
or U6821 (N_6821,N_3250,N_5749);
or U6822 (N_6822,N_4669,N_4438);
nand U6823 (N_6823,N_3199,N_4578);
and U6824 (N_6824,N_4865,N_5343);
or U6825 (N_6825,N_3860,N_3500);
and U6826 (N_6826,N_5299,N_5025);
and U6827 (N_6827,N_3667,N_3468);
nand U6828 (N_6828,N_4522,N_3305);
nand U6829 (N_6829,N_3396,N_4464);
nor U6830 (N_6830,N_5050,N_5216);
xnor U6831 (N_6831,N_3557,N_4992);
nand U6832 (N_6832,N_5008,N_3864);
and U6833 (N_6833,N_5564,N_4018);
or U6834 (N_6834,N_3076,N_4230);
or U6835 (N_6835,N_4724,N_5407);
or U6836 (N_6836,N_4292,N_5381);
nand U6837 (N_6837,N_5118,N_5354);
or U6838 (N_6838,N_5022,N_3586);
nor U6839 (N_6839,N_3913,N_3083);
xor U6840 (N_6840,N_5469,N_3437);
nor U6841 (N_6841,N_5999,N_3722);
nor U6842 (N_6842,N_5200,N_5818);
or U6843 (N_6843,N_4146,N_5194);
and U6844 (N_6844,N_5930,N_4555);
nand U6845 (N_6845,N_4022,N_4151);
nand U6846 (N_6846,N_3373,N_5634);
nand U6847 (N_6847,N_5181,N_3627);
nand U6848 (N_6848,N_3452,N_5857);
nand U6849 (N_6849,N_4186,N_5953);
xnor U6850 (N_6850,N_4979,N_5931);
nor U6851 (N_6851,N_4044,N_4079);
and U6852 (N_6852,N_5250,N_3867);
nand U6853 (N_6853,N_3112,N_5372);
and U6854 (N_6854,N_5998,N_3178);
nor U6855 (N_6855,N_3697,N_5453);
or U6856 (N_6856,N_3230,N_4797);
nand U6857 (N_6857,N_3176,N_5653);
nor U6858 (N_6858,N_5455,N_5345);
nand U6859 (N_6859,N_5700,N_3810);
nor U6860 (N_6860,N_5477,N_4783);
nor U6861 (N_6861,N_4926,N_3374);
or U6862 (N_6862,N_5788,N_5192);
xnor U6863 (N_6863,N_3051,N_5445);
xnor U6864 (N_6864,N_3005,N_5909);
and U6865 (N_6865,N_3400,N_3449);
nor U6866 (N_6866,N_3775,N_5411);
nor U6867 (N_6867,N_4122,N_4824);
nor U6868 (N_6868,N_4874,N_5444);
and U6869 (N_6869,N_3316,N_4499);
nand U6870 (N_6870,N_3629,N_3795);
and U6871 (N_6871,N_5506,N_3186);
and U6872 (N_6872,N_4850,N_3523);
or U6873 (N_6873,N_5265,N_3371);
and U6874 (N_6874,N_4150,N_5002);
nor U6875 (N_6875,N_4245,N_3759);
nand U6876 (N_6876,N_5784,N_4417);
xor U6877 (N_6877,N_4685,N_3776);
or U6878 (N_6878,N_5585,N_4093);
xor U6879 (N_6879,N_5873,N_3858);
nor U6880 (N_6880,N_4729,N_5617);
xnor U6881 (N_6881,N_5318,N_5155);
xnor U6882 (N_6882,N_5037,N_5063);
nor U6883 (N_6883,N_3725,N_3665);
nor U6884 (N_6884,N_4141,N_3793);
and U6885 (N_6885,N_4793,N_3095);
nor U6886 (N_6886,N_5744,N_5060);
nor U6887 (N_6887,N_4247,N_5783);
or U6888 (N_6888,N_3286,N_4902);
xor U6889 (N_6889,N_4305,N_3766);
nand U6890 (N_6890,N_3106,N_5324);
and U6891 (N_6891,N_5116,N_4149);
nor U6892 (N_6892,N_3034,N_4095);
nand U6893 (N_6893,N_3524,N_3065);
or U6894 (N_6894,N_5378,N_4552);
nand U6895 (N_6895,N_5890,N_3566);
or U6896 (N_6896,N_3830,N_5861);
or U6897 (N_6897,N_5951,N_3899);
nand U6898 (N_6898,N_4023,N_3445);
xnor U6899 (N_6899,N_5020,N_4538);
or U6900 (N_6900,N_3944,N_4930);
nand U6901 (N_6901,N_5928,N_3648);
and U6902 (N_6902,N_3695,N_3414);
and U6903 (N_6903,N_3277,N_3322);
or U6904 (N_6904,N_5073,N_5179);
xnor U6905 (N_6905,N_5120,N_3865);
xor U6906 (N_6906,N_3615,N_4526);
nand U6907 (N_6907,N_5109,N_3900);
or U6908 (N_6908,N_5401,N_5153);
and U6909 (N_6909,N_5604,N_5841);
nor U6910 (N_6910,N_4042,N_5269);
nor U6911 (N_6911,N_5261,N_5847);
xnor U6912 (N_6912,N_4737,N_4523);
xnor U6913 (N_6913,N_3534,N_4188);
xor U6914 (N_6914,N_3073,N_3398);
xnor U6915 (N_6915,N_5610,N_3156);
xor U6916 (N_6916,N_3980,N_3382);
xor U6917 (N_6917,N_3009,N_5643);
and U6918 (N_6918,N_3301,N_4524);
or U6919 (N_6919,N_5449,N_3905);
and U6920 (N_6920,N_3987,N_4224);
or U6921 (N_6921,N_3997,N_5097);
or U6922 (N_6922,N_5566,N_3025);
nand U6923 (N_6923,N_3320,N_5706);
or U6924 (N_6924,N_5294,N_5502);
and U6925 (N_6925,N_3740,N_4921);
or U6926 (N_6926,N_4723,N_5042);
and U6927 (N_6927,N_5367,N_4285);
or U6928 (N_6928,N_4947,N_5851);
xnor U6929 (N_6929,N_3909,N_5859);
xnor U6930 (N_6930,N_4336,N_4716);
nand U6931 (N_6931,N_3102,N_3986);
and U6932 (N_6932,N_3676,N_5193);
and U6933 (N_6933,N_5978,N_4173);
nor U6934 (N_6934,N_5973,N_4516);
xnor U6935 (N_6935,N_5721,N_4351);
nor U6936 (N_6936,N_3270,N_5473);
nor U6937 (N_6937,N_3571,N_3833);
nor U6938 (N_6938,N_5812,N_5164);
and U6939 (N_6939,N_4197,N_3016);
or U6940 (N_6940,N_5437,N_3091);
xnor U6941 (N_6941,N_4220,N_3999);
nand U6942 (N_6942,N_5867,N_5257);
xnor U6943 (N_6943,N_4618,N_5624);
or U6944 (N_6944,N_4207,N_4912);
xor U6945 (N_6945,N_3163,N_5262);
nand U6946 (N_6946,N_3789,N_5348);
xnor U6947 (N_6947,N_4727,N_4868);
nor U6948 (N_6948,N_3671,N_5249);
and U6949 (N_6949,N_3840,N_5301);
or U6950 (N_6950,N_3850,N_5807);
nor U6951 (N_6951,N_3749,N_3498);
nand U6952 (N_6952,N_5993,N_4514);
nand U6953 (N_6953,N_5730,N_3809);
nand U6954 (N_6954,N_4196,N_5663);
nand U6955 (N_6955,N_3081,N_3535);
or U6956 (N_6956,N_3866,N_4206);
nor U6957 (N_6957,N_3119,N_5491);
xor U6958 (N_6958,N_5789,N_4809);
nor U6959 (N_6959,N_3567,N_5131);
xor U6960 (N_6960,N_5236,N_5023);
nor U6961 (N_6961,N_4556,N_4144);
or U6962 (N_6962,N_5895,N_3811);
nand U6963 (N_6963,N_3613,N_5991);
nand U6964 (N_6964,N_5329,N_3643);
or U6965 (N_6965,N_3685,N_3647);
and U6966 (N_6966,N_5256,N_4260);
and U6967 (N_6967,N_5326,N_5390);
nor U6968 (N_6968,N_5938,N_4134);
nor U6969 (N_6969,N_3275,N_3838);
and U6970 (N_6970,N_3553,N_5323);
xor U6971 (N_6971,N_5900,N_3587);
xor U6972 (N_6972,N_3313,N_3716);
nand U6973 (N_6973,N_5710,N_3372);
nand U6974 (N_6974,N_3052,N_3687);
nor U6975 (N_6975,N_4346,N_5089);
nor U6976 (N_6976,N_4463,N_4234);
nor U6977 (N_6977,N_3418,N_4276);
and U6978 (N_6978,N_5871,N_5139);
xnor U6979 (N_6979,N_5678,N_5441);
nor U6980 (N_6980,N_5180,N_3816);
and U6981 (N_6981,N_4682,N_5406);
and U6982 (N_6982,N_3509,N_3482);
nor U6983 (N_6983,N_4129,N_3796);
xor U6984 (N_6984,N_5196,N_3344);
xnor U6985 (N_6985,N_5472,N_5819);
and U6986 (N_6986,N_3148,N_4187);
xor U6987 (N_6987,N_5633,N_4786);
xnor U6988 (N_6988,N_4857,N_4377);
nor U6989 (N_6989,N_4092,N_3574);
nand U6990 (N_6990,N_4691,N_3526);
and U6991 (N_6991,N_5043,N_3315);
xnor U6992 (N_6992,N_4832,N_3117);
nor U6993 (N_6993,N_4651,N_5533);
nor U6994 (N_6994,N_3712,N_5399);
nor U6995 (N_6995,N_5729,N_4667);
nor U6996 (N_6996,N_4127,N_4350);
xnor U6997 (N_6997,N_5215,N_3336);
xnor U6998 (N_6998,N_4875,N_4478);
nand U6999 (N_6999,N_4053,N_4339);
nor U7000 (N_7000,N_4116,N_3930);
nor U7001 (N_7001,N_4290,N_4415);
or U7002 (N_7002,N_3174,N_4701);
xnor U7003 (N_7003,N_3579,N_4087);
nor U7004 (N_7004,N_4687,N_3934);
and U7005 (N_7005,N_4842,N_4629);
nand U7006 (N_7006,N_3188,N_4661);
and U7007 (N_7007,N_4316,N_5558);
or U7008 (N_7008,N_4769,N_4462);
and U7009 (N_7009,N_4191,N_4357);
nand U7010 (N_7010,N_3573,N_5123);
nand U7011 (N_7011,N_4814,N_5601);
and U7012 (N_7012,N_5373,N_4089);
xnor U7013 (N_7013,N_5017,N_4621);
or U7014 (N_7014,N_4222,N_3339);
and U7015 (N_7015,N_4470,N_5593);
and U7016 (N_7016,N_4366,N_5434);
xor U7017 (N_7017,N_4476,N_4903);
or U7018 (N_7018,N_3064,N_4973);
xor U7019 (N_7019,N_3525,N_5040);
xor U7020 (N_7020,N_3516,N_4471);
xor U7021 (N_7021,N_5787,N_3649);
and U7022 (N_7022,N_3296,N_3346);
nor U7023 (N_7023,N_4323,N_4812);
nor U7024 (N_7024,N_4684,N_3778);
xor U7025 (N_7025,N_3731,N_3387);
nand U7026 (N_7026,N_4665,N_3259);
nor U7027 (N_7027,N_5707,N_3035);
nand U7028 (N_7028,N_4440,N_5395);
nor U7029 (N_7029,N_5436,N_3053);
and U7030 (N_7030,N_3260,N_4844);
and U7031 (N_7031,N_4612,N_4340);
or U7032 (N_7032,N_5798,N_4107);
nand U7033 (N_7033,N_3780,N_4619);
or U7034 (N_7034,N_4561,N_5980);
or U7035 (N_7035,N_5137,N_4166);
and U7036 (N_7036,N_5007,N_5984);
nor U7037 (N_7037,N_4697,N_5111);
and U7038 (N_7038,N_4571,N_4410);
nor U7039 (N_7039,N_4143,N_4054);
nor U7040 (N_7040,N_4632,N_4379);
nor U7041 (N_7041,N_4041,N_3684);
nor U7042 (N_7042,N_5450,N_3689);
or U7043 (N_7043,N_4058,N_4624);
xor U7044 (N_7044,N_3196,N_5420);
xnor U7045 (N_7045,N_4633,N_5429);
or U7046 (N_7046,N_3921,N_4821);
nand U7047 (N_7047,N_3981,N_3807);
nor U7048 (N_7048,N_5221,N_3435);
and U7049 (N_7049,N_5251,N_3985);
nor U7050 (N_7050,N_5688,N_3737);
nand U7051 (N_7051,N_4035,N_5198);
xnor U7052 (N_7052,N_4950,N_3911);
nand U7053 (N_7053,N_5034,N_5119);
xnor U7054 (N_7054,N_5724,N_4935);
and U7055 (N_7055,N_3826,N_5014);
nor U7056 (N_7056,N_4833,N_4746);
xnor U7057 (N_7057,N_3875,N_4803);
xnor U7058 (N_7058,N_5739,N_3358);
nor U7059 (N_7059,N_4657,N_3919);
and U7060 (N_7060,N_5129,N_3038);
and U7061 (N_7061,N_3283,N_3124);
nand U7062 (N_7062,N_3084,N_3023);
xor U7063 (N_7063,N_5799,N_3961);
xor U7064 (N_7064,N_4369,N_5259);
and U7065 (N_7065,N_4860,N_4901);
nor U7066 (N_7066,N_5122,N_4924);
nor U7067 (N_7067,N_5266,N_5263);
and U7068 (N_7068,N_5575,N_3803);
nand U7069 (N_7069,N_4752,N_3558);
nand U7070 (N_7070,N_5426,N_3920);
xor U7071 (N_7071,N_4917,N_5451);
nor U7072 (N_7072,N_5763,N_3249);
nor U7073 (N_7073,N_5511,N_3638);
or U7074 (N_7074,N_3245,N_4172);
xor U7075 (N_7075,N_5432,N_3533);
and U7076 (N_7076,N_5723,N_4348);
nand U7077 (N_7077,N_3595,N_3046);
xor U7078 (N_7078,N_5358,N_3151);
and U7079 (N_7079,N_4086,N_3576);
and U7080 (N_7080,N_3848,N_3343);
or U7081 (N_7081,N_3540,N_5504);
nor U7082 (N_7082,N_5825,N_5658);
nand U7083 (N_7083,N_4989,N_5813);
and U7084 (N_7084,N_3666,N_5968);
or U7085 (N_7085,N_4502,N_3459);
nand U7086 (N_7086,N_5711,N_5500);
xor U7087 (N_7087,N_3885,N_5482);
nand U7088 (N_7088,N_5229,N_3115);
and U7089 (N_7089,N_5661,N_4182);
or U7090 (N_7090,N_3845,N_5493);
or U7091 (N_7091,N_3002,N_5781);
or U7092 (N_7092,N_4706,N_3221);
nor U7093 (N_7093,N_5785,N_5613);
nor U7094 (N_7094,N_4155,N_4627);
and U7095 (N_7095,N_4858,N_3271);
and U7096 (N_7096,N_3187,N_5866);
nor U7097 (N_7097,N_5031,N_5660);
or U7098 (N_7098,N_4306,N_5505);
nor U7099 (N_7099,N_5225,N_4246);
or U7100 (N_7100,N_5686,N_3881);
nand U7101 (N_7101,N_5759,N_5760);
and U7102 (N_7102,N_4359,N_4430);
nor U7103 (N_7103,N_3285,N_5386);
and U7104 (N_7104,N_3063,N_4498);
or U7105 (N_7105,N_4135,N_5295);
xor U7106 (N_7106,N_4349,N_3614);
nand U7107 (N_7107,N_3892,N_5064);
or U7108 (N_7108,N_4368,N_5995);
nor U7109 (N_7109,N_5829,N_5992);
xor U7110 (N_7110,N_4064,N_5305);
xor U7111 (N_7111,N_5549,N_5756);
xor U7112 (N_7112,N_5964,N_3915);
or U7113 (N_7113,N_4210,N_5969);
or U7114 (N_7114,N_4480,N_4367);
and U7115 (N_7115,N_3536,N_3917);
and U7116 (N_7116,N_3820,N_3837);
and U7117 (N_7117,N_3422,N_3743);
nor U7118 (N_7118,N_3472,N_3832);
nand U7119 (N_7119,N_3600,N_3532);
nor U7120 (N_7120,N_5627,N_4577);
nand U7121 (N_7121,N_3943,N_3728);
nor U7122 (N_7122,N_5582,N_3975);
or U7123 (N_7123,N_5404,N_3543);
and U7124 (N_7124,N_4764,N_5362);
nand U7125 (N_7125,N_5098,N_5430);
xnor U7126 (N_7126,N_5727,N_4999);
or U7127 (N_7127,N_4620,N_4267);
nor U7128 (N_7128,N_5916,N_4941);
or U7129 (N_7129,N_3177,N_5307);
nor U7130 (N_7130,N_3487,N_3423);
nor U7131 (N_7131,N_5580,N_3868);
nand U7132 (N_7132,N_3792,N_4713);
nand U7133 (N_7133,N_3213,N_5905);
and U7134 (N_7134,N_5392,N_5227);
or U7135 (N_7135,N_3704,N_4587);
or U7136 (N_7136,N_4278,N_5061);
and U7137 (N_7137,N_5770,N_5743);
nand U7138 (N_7138,N_3764,N_5465);
xor U7139 (N_7139,N_3411,N_4406);
and U7140 (N_7140,N_5691,N_5275);
and U7141 (N_7141,N_4757,N_5849);
or U7142 (N_7142,N_3114,N_5628);
nor U7143 (N_7143,N_5701,N_4361);
xnor U7144 (N_7144,N_3827,N_5457);
or U7145 (N_7145,N_4605,N_3276);
nand U7146 (N_7146,N_5397,N_5622);
and U7147 (N_7147,N_5396,N_3153);
nand U7148 (N_7148,N_3201,N_4383);
and U7149 (N_7149,N_4414,N_4890);
xnor U7150 (N_7150,N_4236,N_4125);
nand U7151 (N_7151,N_3399,N_5619);
or U7152 (N_7152,N_5260,N_5197);
and U7153 (N_7153,N_4263,N_4558);
and U7154 (N_7154,N_4766,N_4831);
nand U7155 (N_7155,N_3090,N_5836);
xnor U7156 (N_7156,N_5738,N_3145);
and U7157 (N_7157,N_3719,N_3982);
nand U7158 (N_7158,N_3608,N_4944);
or U7159 (N_7159,N_3252,N_5965);
or U7160 (N_7160,N_3560,N_3853);
and U7161 (N_7161,N_3623,N_4307);
or U7162 (N_7162,N_4775,N_5383);
or U7163 (N_7163,N_4174,N_3639);
or U7164 (N_7164,N_3103,N_4660);
or U7165 (N_7165,N_4137,N_5793);
and U7166 (N_7166,N_4124,N_3692);
or U7167 (N_7167,N_5218,N_3036);
nand U7168 (N_7168,N_4423,N_4696);
nand U7169 (N_7169,N_5714,N_5425);
or U7170 (N_7170,N_4686,N_5902);
or U7171 (N_7171,N_5671,N_4314);
nand U7172 (N_7172,N_5838,N_4180);
and U7173 (N_7173,N_3432,N_5279);
nor U7174 (N_7174,N_5586,N_3247);
and U7175 (N_7175,N_3478,N_4404);
nand U7176 (N_7176,N_5311,N_3416);
xor U7177 (N_7177,N_3582,N_3030);
xor U7178 (N_7178,N_4591,N_4459);
xnor U7179 (N_7179,N_3965,N_5919);
or U7180 (N_7180,N_5733,N_3206);
xor U7181 (N_7181,N_4630,N_5609);
or U7182 (N_7182,N_4862,N_4397);
or U7183 (N_7183,N_4911,N_3872);
nor U7184 (N_7184,N_5339,N_5290);
nand U7185 (N_7185,N_5241,N_5047);
and U7186 (N_7186,N_4233,N_5203);
xnor U7187 (N_7187,N_5876,N_3612);
and U7188 (N_7188,N_4519,N_4922);
xor U7189 (N_7189,N_3625,N_4596);
and U7190 (N_7190,N_5574,N_3258);
nand U7191 (N_7191,N_4243,N_3390);
and U7192 (N_7192,N_4019,N_3797);
or U7193 (N_7193,N_5210,N_4681);
xnor U7194 (N_7194,N_5741,N_4888);
nor U7195 (N_7195,N_5230,N_4683);
xor U7196 (N_7196,N_4108,N_5996);
or U7197 (N_7197,N_3958,N_3209);
xor U7198 (N_7198,N_3226,N_5670);
and U7199 (N_7199,N_3032,N_5209);
and U7200 (N_7200,N_5856,N_5745);
xor U7201 (N_7201,N_5894,N_5621);
or U7202 (N_7202,N_3294,N_5839);
and U7203 (N_7203,N_4450,N_3610);
and U7204 (N_7204,N_4319,N_4705);
or U7205 (N_7205,N_3552,N_5699);
xor U7206 (N_7206,N_5545,N_3823);
xor U7207 (N_7207,N_5952,N_4061);
xnor U7208 (N_7208,N_4997,N_4894);
nor U7209 (N_7209,N_4559,N_3458);
nor U7210 (N_7210,N_5778,N_3426);
nor U7211 (N_7211,N_5234,N_3873);
nor U7212 (N_7212,N_3415,N_3385);
nor U7213 (N_7213,N_5824,N_4588);
and U7214 (N_7214,N_3079,N_4225);
xor U7215 (N_7215,N_4666,N_3916);
or U7216 (N_7216,N_5775,N_4819);
nand U7217 (N_7217,N_3218,N_3729);
or U7218 (N_7218,N_5247,N_5600);
and U7219 (N_7219,N_3483,N_5184);
xor U7220 (N_7220,N_3606,N_5412);
xnor U7221 (N_7221,N_4004,N_4749);
nor U7222 (N_7222,N_3233,N_4252);
or U7223 (N_7223,N_3261,N_3988);
or U7224 (N_7224,N_3517,N_5487);
nor U7225 (N_7225,N_4161,N_3950);
nand U7226 (N_7226,N_4208,N_5285);
xor U7227 (N_7227,N_3748,N_5640);
or U7228 (N_7228,N_4530,N_4461);
nand U7229 (N_7229,N_3477,N_3433);
nand U7230 (N_7230,N_5419,N_4475);
xor U7231 (N_7231,N_3505,N_5011);
nor U7232 (N_7232,N_5872,N_4315);
nand U7233 (N_7233,N_4119,N_4878);
nand U7234 (N_7234,N_4027,N_3849);
and U7235 (N_7235,N_4283,N_4016);
nor U7236 (N_7236,N_5391,N_3907);
or U7237 (N_7237,N_3047,N_3700);
or U7238 (N_7238,N_5576,N_3008);
nor U7239 (N_7239,N_5646,N_4945);
xnor U7240 (N_7240,N_4534,N_3617);
nand U7241 (N_7241,N_5879,N_4712);
nand U7242 (N_7242,N_4560,N_4521);
xnor U7243 (N_7243,N_4808,N_5657);
and U7244 (N_7244,N_3597,N_4648);
and U7245 (N_7245,N_5356,N_3699);
xor U7246 (N_7246,N_3231,N_4217);
nand U7247 (N_7247,N_5080,N_4103);
or U7248 (N_7248,N_5288,N_3376);
nand U7249 (N_7249,N_3162,N_3138);
and U7250 (N_7250,N_3244,N_5195);
xor U7251 (N_7251,N_3641,N_3581);
xnor U7252 (N_7252,N_5468,N_5309);
or U7253 (N_7253,N_5174,N_5651);
or U7254 (N_7254,N_4469,N_4268);
nand U7255 (N_7255,N_4904,N_3788);
nor U7256 (N_7256,N_3831,N_5341);
nand U7257 (N_7257,N_5581,N_3730);
nor U7258 (N_7258,N_3268,N_3020);
and U7259 (N_7259,N_4386,N_3635);
nor U7260 (N_7260,N_4734,N_3632);
and U7261 (N_7261,N_4492,N_4326);
or U7262 (N_7262,N_3758,N_3430);
nor U7263 (N_7263,N_5224,N_3889);
or U7264 (N_7264,N_3669,N_4715);
or U7265 (N_7265,N_4321,N_5499);
xor U7266 (N_7266,N_4251,N_4529);
nand U7267 (N_7267,N_3028,N_4060);
or U7268 (N_7268,N_3903,N_4520);
or U7269 (N_7269,N_4583,N_3723);
xnor U7270 (N_7270,N_3183,N_3929);
and U7271 (N_7271,N_3747,N_4900);
nand U7272 (N_7272,N_5044,N_4565);
nor U7273 (N_7273,N_5940,N_4287);
nor U7274 (N_7274,N_5327,N_5638);
nand U7275 (N_7275,N_5844,N_5086);
and U7276 (N_7276,N_4601,N_4567);
nor U7277 (N_7277,N_3240,N_4274);
xor U7278 (N_7278,N_5421,N_5554);
xor U7279 (N_7279,N_5979,N_4077);
nor U7280 (N_7280,N_4963,N_4595);
or U7281 (N_7281,N_3024,N_3746);
nor U7282 (N_7282,N_3205,N_3311);
or U7283 (N_7283,N_4088,N_3974);
xor U7284 (N_7284,N_5551,N_3475);
nor U7285 (N_7285,N_5882,N_3120);
nand U7286 (N_7286,N_4426,N_4436);
xor U7287 (N_7287,N_4845,N_4140);
or U7288 (N_7288,N_5183,N_3819);
nor U7289 (N_7289,N_4078,N_5922);
and U7290 (N_7290,N_3180,N_5941);
and U7291 (N_7291,N_5117,N_3914);
and U7292 (N_7292,N_4983,N_5248);
nor U7293 (N_7293,N_5239,N_4837);
xor U7294 (N_7294,N_5021,N_4733);
xor U7295 (N_7295,N_4564,N_4065);
xnor U7296 (N_7296,N_3050,N_5471);
nand U7297 (N_7297,N_4465,N_5314);
nand U7298 (N_7298,N_4714,N_3121);
or U7299 (N_7299,N_5231,N_4759);
and U7300 (N_7300,N_3118,N_4309);
or U7301 (N_7301,N_5057,N_3255);
or U7302 (N_7302,N_4739,N_3645);
and U7303 (N_7303,N_4804,N_4511);
and U7304 (N_7304,N_3125,N_4487);
and U7305 (N_7305,N_4399,N_3901);
and U7306 (N_7306,N_3488,N_3181);
and U7307 (N_7307,N_4051,N_5742);
nor U7308 (N_7308,N_3474,N_5347);
xor U7309 (N_7309,N_4810,N_3170);
nor U7310 (N_7310,N_5570,N_4400);
nor U7311 (N_7311,N_4131,N_5615);
or U7312 (N_7312,N_5359,N_4573);
and U7313 (N_7313,N_3082,N_3957);
nor U7314 (N_7314,N_4678,N_4623);
and U7315 (N_7315,N_4951,N_4659);
and U7316 (N_7316,N_5492,N_5834);
xnor U7317 (N_7317,N_3144,N_5302);
or U7318 (N_7318,N_4608,N_5460);
or U7319 (N_7319,N_5945,N_5101);
or U7320 (N_7320,N_3492,N_3161);
xor U7321 (N_7321,N_4778,N_4929);
xor U7322 (N_7322,N_5750,N_4631);
or U7323 (N_7323,N_4015,N_4331);
nor U7324 (N_7324,N_3189,N_5187);
or U7325 (N_7325,N_3039,N_4213);
nand U7326 (N_7326,N_3060,N_5779);
and U7327 (N_7327,N_5189,N_3061);
xnor U7328 (N_7328,N_4048,N_4013);
nor U7329 (N_7329,N_3223,N_5217);
or U7330 (N_7330,N_4133,N_3408);
xor U7331 (N_7331,N_4005,N_4846);
nand U7332 (N_7332,N_4794,N_3236);
and U7333 (N_7333,N_5967,N_3049);
nor U7334 (N_7334,N_5409,N_3078);
or U7335 (N_7335,N_3332,N_5423);
and U7336 (N_7336,N_5840,N_4330);
xnor U7337 (N_7337,N_5935,N_4001);
and U7338 (N_7338,N_3547,N_4995);
and U7339 (N_7339,N_3173,N_5514);
nand U7340 (N_7340,N_3808,N_4264);
nand U7341 (N_7341,N_4275,N_5607);
xor U7342 (N_7342,N_4355,N_3479);
or U7343 (N_7343,N_4341,N_4320);
xor U7344 (N_7344,N_5684,N_5529);
nand U7345 (N_7345,N_4083,N_3637);
or U7346 (N_7346,N_5817,N_5848);
xor U7347 (N_7347,N_5913,N_3727);
and U7348 (N_7348,N_5018,N_3491);
xor U7349 (N_7349,N_3013,N_4378);
or U7350 (N_7350,N_3425,N_4102);
nand U7351 (N_7351,N_3204,N_5709);
or U7352 (N_7352,N_4887,N_3906);
or U7353 (N_7353,N_4299,N_3288);
nand U7354 (N_7354,N_3815,N_4056);
nand U7355 (N_7355,N_3234,N_4649);
and U7356 (N_7356,N_3253,N_3738);
or U7357 (N_7357,N_4787,N_4009);
and U7358 (N_7358,N_3527,N_3239);
nor U7359 (N_7359,N_4823,N_4952);
nor U7360 (N_7360,N_4971,N_5368);
nand U7361 (N_7361,N_4218,N_4286);
nand U7362 (N_7362,N_5410,N_3044);
or U7363 (N_7363,N_5864,N_4451);
xor U7364 (N_7364,N_3836,N_3448);
xor U7365 (N_7365,N_4481,N_4745);
nor U7366 (N_7366,N_3707,N_5528);
and U7367 (N_7367,N_3175,N_3001);
nand U7368 (N_7368,N_3733,N_4562);
nand U7369 (N_7369,N_4434,N_3330);
nor U7370 (N_7370,N_5598,N_3978);
xor U7371 (N_7371,N_4178,N_5977);
and U7372 (N_7372,N_3918,N_4539);
and U7373 (N_7373,N_5088,N_4153);
and U7374 (N_7374,N_3149,N_4313);
xnor U7375 (N_7375,N_3097,N_3325);
and U7376 (N_7376,N_4873,N_3935);
nor U7377 (N_7377,N_3768,N_4625);
xnor U7378 (N_7378,N_3210,N_4554);
or U7379 (N_7379,N_5920,N_5947);
xnor U7380 (N_7380,N_3340,N_3562);
or U7381 (N_7381,N_5113,N_3131);
and U7382 (N_7382,N_4985,N_5448);
and U7383 (N_7383,N_5587,N_5655);
and U7384 (N_7384,N_5182,N_4488);
xnor U7385 (N_7385,N_4790,N_3750);
nor U7386 (N_7386,N_4531,N_4240);
and U7387 (N_7387,N_4071,N_3936);
nand U7388 (N_7388,N_5767,N_5539);
and U7389 (N_7389,N_5637,N_4253);
xor U7390 (N_7390,N_3537,N_5173);
or U7391 (N_7391,N_3167,N_5887);
xor U7392 (N_7392,N_5142,N_5310);
xor U7393 (N_7393,N_5328,N_5950);
and U7394 (N_7394,N_5881,N_5162);
nand U7395 (N_7395,N_4221,N_4638);
nor U7396 (N_7396,N_3394,N_4431);
or U7397 (N_7397,N_5774,N_5614);
xnor U7398 (N_7398,N_3338,N_4441);
nor U7399 (N_7399,N_5949,N_4163);
or U7400 (N_7400,N_5846,N_3010);
nand U7401 (N_7401,N_4537,N_5332);
xor U7402 (N_7402,N_5982,N_4007);
nor U7403 (N_7403,N_4280,N_4600);
nand U7404 (N_7404,N_5090,N_4893);
nor U7405 (N_7405,N_5202,N_3724);
or U7406 (N_7406,N_5237,N_4581);
nand U7407 (N_7407,N_5543,N_3280);
xnor U7408 (N_7408,N_5512,N_3463);
nor U7409 (N_7409,N_3751,N_3251);
xnor U7410 (N_7410,N_3379,N_4000);
or U7411 (N_7411,N_3337,N_4861);
and U7412 (N_7412,N_5422,N_4439);
and U7413 (N_7413,N_4975,N_4843);
nand U7414 (N_7414,N_4613,N_3455);
or U7415 (N_7415,N_3960,N_3570);
nand U7416 (N_7416,N_5893,N_3821);
and U7417 (N_7417,N_5606,N_4293);
xor U7418 (N_7418,N_3182,N_3742);
and U7419 (N_7419,N_3715,N_3956);
or U7420 (N_7420,N_3633,N_3642);
or U7421 (N_7421,N_4205,N_4647);
xnor U7422 (N_7422,N_3995,N_5831);
xnor U7423 (N_7423,N_3085,N_4128);
nand U7424 (N_7424,N_5517,N_4774);
and U7425 (N_7425,N_3350,N_3931);
and U7426 (N_7426,N_4675,N_4460);
nor U7427 (N_7427,N_4602,N_3473);
and U7428 (N_7428,N_4255,N_5559);
nand U7429 (N_7429,N_4193,N_4189);
xnor U7430 (N_7430,N_4909,N_5456);
nor U7431 (N_7431,N_5452,N_3219);
xnor U7432 (N_7432,N_4540,N_4111);
and U7433 (N_7433,N_3851,N_3744);
xor U7434 (N_7434,N_4387,N_4242);
and U7435 (N_7435,N_3834,N_4740);
xor U7436 (N_7436,N_5852,N_5987);
nand U7437 (N_7437,N_4943,N_3169);
xnor U7438 (N_7438,N_5820,N_4342);
or U7439 (N_7439,N_5149,N_5255);
or U7440 (N_7440,N_5287,N_5055);
or U7441 (N_7441,N_3609,N_5616);
and U7442 (N_7442,N_3184,N_4443);
nand U7443 (N_7443,N_5828,N_3128);
and U7444 (N_7444,N_5540,N_5387);
nor U7445 (N_7445,N_5418,N_5240);
nand U7446 (N_7446,N_3033,N_4055);
nor U7447 (N_7447,N_3510,N_4473);
xor U7448 (N_7448,N_5773,N_3602);
nand U7449 (N_7449,N_3129,N_4984);
nand U7450 (N_7450,N_5488,N_3966);
or U7451 (N_7451,N_5167,N_5046);
nand U7452 (N_7452,N_4484,N_4482);
nor U7453 (N_7453,N_5959,N_5475);
and U7454 (N_7454,N_4138,N_5791);
and U7455 (N_7455,N_3494,N_3355);
and U7456 (N_7456,N_4836,N_5417);
nand U7457 (N_7457,N_3640,N_3691);
nand U7458 (N_7458,N_3059,N_3327);
nor U7459 (N_7459,N_4248,N_3419);
and U7460 (N_7460,N_3507,N_3784);
nor U7461 (N_7461,N_5929,N_5560);
nor U7462 (N_7462,N_4741,N_3734);
nand U7463 (N_7463,N_5669,N_4762);
or U7464 (N_7464,N_5786,N_5278);
and U7465 (N_7465,N_5296,N_4063);
or U7466 (N_7466,N_4432,N_5244);
xnor U7467 (N_7467,N_3241,N_5338);
and U7468 (N_7468,N_5188,N_4547);
and U7469 (N_7469,N_5304,N_3440);
or U7470 (N_7470,N_4325,N_3662);
and U7471 (N_7471,N_5178,N_5526);
and U7472 (N_7472,N_3683,N_3367);
and U7473 (N_7473,N_3439,N_3679);
xor U7474 (N_7474,N_4978,N_4139);
nor U7475 (N_7475,N_4799,N_4576);
nor U7476 (N_7476,N_5522,N_4202);
and U7477 (N_7477,N_4084,N_3092);
nand U7478 (N_7478,N_5692,N_3530);
nand U7479 (N_7479,N_5885,N_5124);
and U7480 (N_7480,N_4353,N_3963);
xor U7481 (N_7481,N_3791,N_4871);
xnor U7482 (N_7482,N_3628,N_4936);
xor U7483 (N_7483,N_4324,N_3395);
xnor U7484 (N_7484,N_3771,N_3154);
nand U7485 (N_7485,N_5232,N_4968);
nor U7486 (N_7486,N_5253,N_5235);
and U7487 (N_7487,N_5693,N_4703);
nor U7488 (N_7488,N_5024,N_4356);
nor U7489 (N_7489,N_5382,N_5463);
or U7490 (N_7490,N_4550,N_3462);
or U7491 (N_7491,N_4702,N_5532);
nor U7492 (N_7492,N_4870,N_4453);
and U7493 (N_7493,N_4663,N_4047);
nor U7494 (N_7494,N_5004,N_5889);
and U7495 (N_7495,N_5937,N_3193);
or U7496 (N_7496,N_3329,N_4668);
xnor U7497 (N_7497,N_4418,N_5556);
nand U7498 (N_7498,N_5626,N_4966);
xor U7499 (N_7499,N_3702,N_5883);
xnor U7500 (N_7500,N_5060,N_5082);
nor U7501 (N_7501,N_4243,N_5889);
and U7502 (N_7502,N_4189,N_3431);
and U7503 (N_7503,N_5898,N_3832);
nor U7504 (N_7504,N_4300,N_3148);
nand U7505 (N_7505,N_4529,N_3590);
and U7506 (N_7506,N_4980,N_4678);
xnor U7507 (N_7507,N_4443,N_3549);
nand U7508 (N_7508,N_4526,N_4317);
and U7509 (N_7509,N_3169,N_3082);
or U7510 (N_7510,N_3363,N_5137);
or U7511 (N_7511,N_5370,N_5547);
nand U7512 (N_7512,N_3754,N_4518);
xnor U7513 (N_7513,N_5183,N_3014);
nand U7514 (N_7514,N_3199,N_5036);
nand U7515 (N_7515,N_3082,N_5879);
nor U7516 (N_7516,N_4676,N_3308);
nand U7517 (N_7517,N_5706,N_4616);
nand U7518 (N_7518,N_3071,N_4179);
nor U7519 (N_7519,N_3898,N_3713);
nor U7520 (N_7520,N_3868,N_3819);
or U7521 (N_7521,N_4371,N_4098);
xnor U7522 (N_7522,N_3690,N_3343);
and U7523 (N_7523,N_4962,N_4471);
xnor U7524 (N_7524,N_4218,N_4101);
nand U7525 (N_7525,N_3673,N_5889);
nor U7526 (N_7526,N_4671,N_3914);
and U7527 (N_7527,N_4286,N_5434);
xor U7528 (N_7528,N_4156,N_4417);
nand U7529 (N_7529,N_3508,N_5636);
xnor U7530 (N_7530,N_5102,N_3898);
nor U7531 (N_7531,N_3981,N_3702);
or U7532 (N_7532,N_4117,N_5599);
nand U7533 (N_7533,N_4218,N_4198);
and U7534 (N_7534,N_4670,N_5759);
or U7535 (N_7535,N_3480,N_3385);
or U7536 (N_7536,N_4945,N_4207);
or U7537 (N_7537,N_4414,N_5570);
nand U7538 (N_7538,N_3265,N_5154);
and U7539 (N_7539,N_4693,N_3058);
xnor U7540 (N_7540,N_4643,N_3193);
xnor U7541 (N_7541,N_4536,N_3476);
nor U7542 (N_7542,N_3556,N_5856);
and U7543 (N_7543,N_5366,N_3293);
nor U7544 (N_7544,N_4999,N_5974);
xor U7545 (N_7545,N_5282,N_3337);
nor U7546 (N_7546,N_3641,N_4361);
xor U7547 (N_7547,N_3929,N_4196);
and U7548 (N_7548,N_5127,N_3495);
and U7549 (N_7549,N_3823,N_4021);
xor U7550 (N_7550,N_4985,N_5374);
and U7551 (N_7551,N_5063,N_5497);
nor U7552 (N_7552,N_5208,N_3518);
nand U7553 (N_7553,N_5865,N_5829);
or U7554 (N_7554,N_3352,N_4861);
and U7555 (N_7555,N_3059,N_3348);
and U7556 (N_7556,N_4446,N_4968);
nor U7557 (N_7557,N_5571,N_4808);
nand U7558 (N_7558,N_4546,N_5870);
xnor U7559 (N_7559,N_4871,N_4043);
nand U7560 (N_7560,N_5618,N_3031);
or U7561 (N_7561,N_3173,N_3220);
xor U7562 (N_7562,N_3403,N_5685);
nand U7563 (N_7563,N_4731,N_4761);
and U7564 (N_7564,N_3719,N_4329);
nand U7565 (N_7565,N_4636,N_3490);
and U7566 (N_7566,N_5319,N_3577);
nor U7567 (N_7567,N_4288,N_5850);
and U7568 (N_7568,N_5156,N_3587);
or U7569 (N_7569,N_4384,N_4238);
and U7570 (N_7570,N_4902,N_4888);
xnor U7571 (N_7571,N_5005,N_4083);
or U7572 (N_7572,N_4179,N_3649);
nor U7573 (N_7573,N_3004,N_4728);
nand U7574 (N_7574,N_4095,N_4702);
and U7575 (N_7575,N_5208,N_4246);
xnor U7576 (N_7576,N_3930,N_4273);
xor U7577 (N_7577,N_3551,N_4543);
and U7578 (N_7578,N_3219,N_3276);
nand U7579 (N_7579,N_3610,N_4678);
xnor U7580 (N_7580,N_3794,N_3374);
or U7581 (N_7581,N_4128,N_5488);
or U7582 (N_7582,N_4074,N_3827);
and U7583 (N_7583,N_4795,N_5211);
and U7584 (N_7584,N_3631,N_4276);
and U7585 (N_7585,N_5120,N_4684);
nand U7586 (N_7586,N_5713,N_5611);
or U7587 (N_7587,N_3553,N_5717);
or U7588 (N_7588,N_3244,N_3717);
nor U7589 (N_7589,N_3844,N_4853);
or U7590 (N_7590,N_5209,N_3955);
xor U7591 (N_7591,N_3779,N_5628);
nand U7592 (N_7592,N_5329,N_5143);
xnor U7593 (N_7593,N_3347,N_5021);
and U7594 (N_7594,N_3212,N_4891);
nand U7595 (N_7595,N_3320,N_3615);
and U7596 (N_7596,N_4025,N_5817);
xor U7597 (N_7597,N_4239,N_5910);
xnor U7598 (N_7598,N_5728,N_3500);
xor U7599 (N_7599,N_5015,N_5439);
and U7600 (N_7600,N_4102,N_4638);
or U7601 (N_7601,N_3555,N_4737);
xnor U7602 (N_7602,N_4130,N_5443);
xor U7603 (N_7603,N_5999,N_4844);
nor U7604 (N_7604,N_4995,N_5149);
nand U7605 (N_7605,N_5758,N_5028);
xnor U7606 (N_7606,N_3569,N_3945);
xor U7607 (N_7607,N_3783,N_3417);
nor U7608 (N_7608,N_4653,N_4501);
nor U7609 (N_7609,N_5225,N_5383);
and U7610 (N_7610,N_3283,N_5476);
and U7611 (N_7611,N_4927,N_4809);
or U7612 (N_7612,N_3376,N_3420);
nand U7613 (N_7613,N_4786,N_3668);
or U7614 (N_7614,N_3375,N_4696);
nor U7615 (N_7615,N_3639,N_3345);
nor U7616 (N_7616,N_4583,N_5748);
or U7617 (N_7617,N_4113,N_5433);
xnor U7618 (N_7618,N_4207,N_3065);
xnor U7619 (N_7619,N_5963,N_3432);
and U7620 (N_7620,N_4007,N_5249);
xor U7621 (N_7621,N_5826,N_5544);
or U7622 (N_7622,N_5436,N_3018);
and U7623 (N_7623,N_5583,N_5174);
nor U7624 (N_7624,N_5761,N_4673);
xor U7625 (N_7625,N_5650,N_4772);
and U7626 (N_7626,N_4285,N_3853);
or U7627 (N_7627,N_4614,N_3338);
or U7628 (N_7628,N_5312,N_5212);
and U7629 (N_7629,N_4458,N_5119);
nand U7630 (N_7630,N_5815,N_4252);
nand U7631 (N_7631,N_4290,N_4972);
xor U7632 (N_7632,N_5446,N_4656);
xnor U7633 (N_7633,N_3936,N_5323);
xor U7634 (N_7634,N_4242,N_4085);
or U7635 (N_7635,N_5317,N_5947);
and U7636 (N_7636,N_4065,N_5226);
and U7637 (N_7637,N_3320,N_3561);
xnor U7638 (N_7638,N_4586,N_4902);
xor U7639 (N_7639,N_5008,N_5673);
nor U7640 (N_7640,N_3475,N_3752);
nand U7641 (N_7641,N_3539,N_5375);
xnor U7642 (N_7642,N_4375,N_4208);
nand U7643 (N_7643,N_3384,N_5153);
nor U7644 (N_7644,N_4916,N_5596);
nand U7645 (N_7645,N_5411,N_3528);
nor U7646 (N_7646,N_3262,N_4009);
or U7647 (N_7647,N_3304,N_4510);
nand U7648 (N_7648,N_4458,N_4331);
xnor U7649 (N_7649,N_3405,N_4441);
nor U7650 (N_7650,N_5202,N_3540);
xor U7651 (N_7651,N_4551,N_3981);
xnor U7652 (N_7652,N_4018,N_5204);
nand U7653 (N_7653,N_4808,N_4968);
and U7654 (N_7654,N_5680,N_4412);
xnor U7655 (N_7655,N_3777,N_5894);
and U7656 (N_7656,N_3223,N_4885);
and U7657 (N_7657,N_4024,N_3946);
and U7658 (N_7658,N_3813,N_3593);
nand U7659 (N_7659,N_5762,N_4617);
nand U7660 (N_7660,N_5599,N_3797);
xor U7661 (N_7661,N_4619,N_4708);
or U7662 (N_7662,N_4039,N_3863);
xnor U7663 (N_7663,N_3767,N_3299);
nor U7664 (N_7664,N_4817,N_5041);
and U7665 (N_7665,N_5086,N_3799);
or U7666 (N_7666,N_4991,N_3815);
nand U7667 (N_7667,N_5844,N_4462);
or U7668 (N_7668,N_3298,N_5571);
and U7669 (N_7669,N_4471,N_4161);
or U7670 (N_7670,N_5936,N_5632);
xnor U7671 (N_7671,N_4844,N_5344);
nand U7672 (N_7672,N_5604,N_5223);
nor U7673 (N_7673,N_5042,N_5672);
and U7674 (N_7674,N_5530,N_5219);
and U7675 (N_7675,N_5269,N_3984);
or U7676 (N_7676,N_4740,N_5982);
nand U7677 (N_7677,N_5703,N_4573);
or U7678 (N_7678,N_4518,N_4520);
nor U7679 (N_7679,N_4427,N_3836);
nor U7680 (N_7680,N_3269,N_3455);
and U7681 (N_7681,N_3267,N_5063);
nor U7682 (N_7682,N_3806,N_5006);
nand U7683 (N_7683,N_4344,N_4700);
or U7684 (N_7684,N_5003,N_3218);
or U7685 (N_7685,N_3331,N_3614);
xor U7686 (N_7686,N_3318,N_4344);
xnor U7687 (N_7687,N_4935,N_3523);
and U7688 (N_7688,N_5594,N_4686);
xor U7689 (N_7689,N_5653,N_5039);
or U7690 (N_7690,N_5460,N_3180);
xor U7691 (N_7691,N_3328,N_3341);
xnor U7692 (N_7692,N_5027,N_5861);
nand U7693 (N_7693,N_5382,N_3197);
xnor U7694 (N_7694,N_4322,N_4260);
nand U7695 (N_7695,N_3537,N_4673);
xor U7696 (N_7696,N_3526,N_3205);
xor U7697 (N_7697,N_5974,N_5280);
nor U7698 (N_7698,N_5103,N_4413);
xor U7699 (N_7699,N_3984,N_3746);
or U7700 (N_7700,N_5355,N_3947);
or U7701 (N_7701,N_4216,N_4474);
and U7702 (N_7702,N_4485,N_3432);
or U7703 (N_7703,N_4751,N_5455);
nand U7704 (N_7704,N_5553,N_3348);
or U7705 (N_7705,N_4509,N_3835);
nor U7706 (N_7706,N_5025,N_4907);
nand U7707 (N_7707,N_3905,N_5626);
xnor U7708 (N_7708,N_5209,N_4033);
nor U7709 (N_7709,N_4618,N_4226);
nand U7710 (N_7710,N_4466,N_5636);
and U7711 (N_7711,N_4421,N_5175);
xor U7712 (N_7712,N_5723,N_3544);
nor U7713 (N_7713,N_5605,N_5323);
nand U7714 (N_7714,N_4293,N_4382);
and U7715 (N_7715,N_3427,N_4843);
or U7716 (N_7716,N_4494,N_4625);
nor U7717 (N_7717,N_5064,N_3829);
and U7718 (N_7718,N_4232,N_5867);
or U7719 (N_7719,N_4485,N_5763);
or U7720 (N_7720,N_3990,N_3965);
xnor U7721 (N_7721,N_5968,N_5221);
or U7722 (N_7722,N_4531,N_4644);
nor U7723 (N_7723,N_3197,N_4814);
nor U7724 (N_7724,N_4803,N_3553);
xnor U7725 (N_7725,N_4193,N_5329);
nand U7726 (N_7726,N_5755,N_5014);
nand U7727 (N_7727,N_4504,N_4495);
nor U7728 (N_7728,N_3597,N_5297);
and U7729 (N_7729,N_4837,N_4578);
xnor U7730 (N_7730,N_3911,N_4869);
nand U7731 (N_7731,N_3273,N_4285);
and U7732 (N_7732,N_4618,N_4066);
nor U7733 (N_7733,N_5990,N_5802);
xnor U7734 (N_7734,N_5098,N_3927);
nor U7735 (N_7735,N_3094,N_5391);
and U7736 (N_7736,N_3783,N_5514);
nand U7737 (N_7737,N_5429,N_5144);
nor U7738 (N_7738,N_3504,N_4696);
xor U7739 (N_7739,N_4114,N_5180);
nand U7740 (N_7740,N_4048,N_3735);
xor U7741 (N_7741,N_4070,N_4687);
nand U7742 (N_7742,N_3256,N_5184);
and U7743 (N_7743,N_5996,N_3458);
nand U7744 (N_7744,N_5707,N_5950);
or U7745 (N_7745,N_5466,N_5113);
xnor U7746 (N_7746,N_5620,N_5744);
nor U7747 (N_7747,N_4492,N_3797);
and U7748 (N_7748,N_5621,N_4050);
and U7749 (N_7749,N_4184,N_4878);
nand U7750 (N_7750,N_4058,N_5053);
xor U7751 (N_7751,N_5590,N_5611);
nand U7752 (N_7752,N_4021,N_5375);
nor U7753 (N_7753,N_4730,N_4977);
xnor U7754 (N_7754,N_4526,N_5254);
and U7755 (N_7755,N_3967,N_3881);
xor U7756 (N_7756,N_4393,N_3362);
and U7757 (N_7757,N_4663,N_3264);
nor U7758 (N_7758,N_5069,N_3642);
or U7759 (N_7759,N_5812,N_4308);
nor U7760 (N_7760,N_5498,N_3283);
nand U7761 (N_7761,N_4469,N_3643);
and U7762 (N_7762,N_4252,N_4223);
and U7763 (N_7763,N_5531,N_5443);
nor U7764 (N_7764,N_3909,N_4091);
or U7765 (N_7765,N_3951,N_3897);
nor U7766 (N_7766,N_4883,N_4742);
or U7767 (N_7767,N_4522,N_4436);
nand U7768 (N_7768,N_4292,N_4425);
and U7769 (N_7769,N_5828,N_5975);
xor U7770 (N_7770,N_4698,N_4589);
or U7771 (N_7771,N_5266,N_4925);
nand U7772 (N_7772,N_3035,N_5901);
nand U7773 (N_7773,N_5316,N_3591);
nor U7774 (N_7774,N_3552,N_4588);
nand U7775 (N_7775,N_3720,N_3051);
xnor U7776 (N_7776,N_3328,N_5268);
xor U7777 (N_7777,N_5883,N_5052);
xor U7778 (N_7778,N_4877,N_5486);
nand U7779 (N_7779,N_4317,N_5010);
xor U7780 (N_7780,N_3747,N_5302);
nand U7781 (N_7781,N_3863,N_3306);
nand U7782 (N_7782,N_5937,N_5042);
xor U7783 (N_7783,N_5312,N_4070);
xnor U7784 (N_7784,N_4253,N_3165);
xor U7785 (N_7785,N_3808,N_3795);
and U7786 (N_7786,N_5355,N_4628);
xor U7787 (N_7787,N_5977,N_4211);
xor U7788 (N_7788,N_5101,N_3244);
nor U7789 (N_7789,N_3587,N_4471);
and U7790 (N_7790,N_3164,N_3512);
nor U7791 (N_7791,N_4378,N_4939);
nor U7792 (N_7792,N_4902,N_3515);
xor U7793 (N_7793,N_3989,N_4173);
and U7794 (N_7794,N_3761,N_4484);
or U7795 (N_7795,N_3966,N_5756);
xor U7796 (N_7796,N_3657,N_4990);
or U7797 (N_7797,N_4130,N_4321);
nand U7798 (N_7798,N_3186,N_5425);
nor U7799 (N_7799,N_4783,N_3116);
xnor U7800 (N_7800,N_5614,N_4786);
and U7801 (N_7801,N_4089,N_4594);
and U7802 (N_7802,N_4706,N_3450);
and U7803 (N_7803,N_4713,N_4060);
nand U7804 (N_7804,N_5897,N_5027);
nand U7805 (N_7805,N_4423,N_5537);
nand U7806 (N_7806,N_3910,N_3738);
and U7807 (N_7807,N_5026,N_3565);
or U7808 (N_7808,N_5880,N_5785);
nor U7809 (N_7809,N_5024,N_4451);
xnor U7810 (N_7810,N_5389,N_4441);
or U7811 (N_7811,N_4758,N_5377);
and U7812 (N_7812,N_5386,N_5376);
nand U7813 (N_7813,N_4401,N_5872);
nor U7814 (N_7814,N_3196,N_5047);
and U7815 (N_7815,N_4915,N_5521);
or U7816 (N_7816,N_3426,N_5048);
nor U7817 (N_7817,N_3208,N_3393);
or U7818 (N_7818,N_5940,N_5963);
nor U7819 (N_7819,N_4601,N_4096);
xor U7820 (N_7820,N_4223,N_5457);
or U7821 (N_7821,N_5586,N_4459);
and U7822 (N_7822,N_4651,N_3990);
or U7823 (N_7823,N_3589,N_4804);
xor U7824 (N_7824,N_4375,N_3628);
nand U7825 (N_7825,N_4108,N_4576);
or U7826 (N_7826,N_5423,N_3979);
xnor U7827 (N_7827,N_4811,N_4729);
nand U7828 (N_7828,N_5783,N_5882);
nor U7829 (N_7829,N_3675,N_3035);
and U7830 (N_7830,N_5962,N_4821);
and U7831 (N_7831,N_5964,N_4968);
xnor U7832 (N_7832,N_3444,N_4804);
xnor U7833 (N_7833,N_5004,N_3450);
xnor U7834 (N_7834,N_4112,N_4918);
or U7835 (N_7835,N_3702,N_5590);
nand U7836 (N_7836,N_3655,N_3729);
nor U7837 (N_7837,N_3502,N_5115);
xnor U7838 (N_7838,N_3371,N_3120);
nor U7839 (N_7839,N_4399,N_3025);
nor U7840 (N_7840,N_3572,N_3834);
nor U7841 (N_7841,N_5197,N_4621);
nor U7842 (N_7842,N_4812,N_4701);
nor U7843 (N_7843,N_4106,N_3803);
nor U7844 (N_7844,N_5028,N_5243);
nand U7845 (N_7845,N_3399,N_4839);
or U7846 (N_7846,N_4265,N_3527);
nand U7847 (N_7847,N_5894,N_3099);
or U7848 (N_7848,N_5405,N_4519);
and U7849 (N_7849,N_3964,N_4442);
nor U7850 (N_7850,N_3022,N_5021);
and U7851 (N_7851,N_3549,N_5566);
or U7852 (N_7852,N_4814,N_4712);
xnor U7853 (N_7853,N_4471,N_4917);
nor U7854 (N_7854,N_4062,N_5651);
and U7855 (N_7855,N_5635,N_5249);
xor U7856 (N_7856,N_5381,N_5561);
or U7857 (N_7857,N_5492,N_5470);
nand U7858 (N_7858,N_5390,N_5785);
xnor U7859 (N_7859,N_3404,N_5864);
nand U7860 (N_7860,N_5267,N_3723);
nand U7861 (N_7861,N_3238,N_3568);
xor U7862 (N_7862,N_3454,N_5600);
or U7863 (N_7863,N_5300,N_3816);
and U7864 (N_7864,N_4090,N_4321);
and U7865 (N_7865,N_3044,N_4650);
or U7866 (N_7866,N_4712,N_5018);
and U7867 (N_7867,N_4951,N_5476);
nand U7868 (N_7868,N_5115,N_4020);
nor U7869 (N_7869,N_4476,N_5197);
nor U7870 (N_7870,N_5298,N_5867);
or U7871 (N_7871,N_3666,N_4145);
nand U7872 (N_7872,N_5524,N_4833);
or U7873 (N_7873,N_4883,N_4255);
or U7874 (N_7874,N_3327,N_5419);
and U7875 (N_7875,N_5251,N_5312);
nor U7876 (N_7876,N_3039,N_5195);
xnor U7877 (N_7877,N_3421,N_3728);
or U7878 (N_7878,N_3313,N_5922);
or U7879 (N_7879,N_4101,N_4476);
nor U7880 (N_7880,N_4669,N_3707);
nand U7881 (N_7881,N_4103,N_4016);
nor U7882 (N_7882,N_5512,N_3435);
and U7883 (N_7883,N_3299,N_5366);
or U7884 (N_7884,N_3065,N_3428);
nor U7885 (N_7885,N_3589,N_3592);
nand U7886 (N_7886,N_3202,N_4484);
and U7887 (N_7887,N_5855,N_4506);
nand U7888 (N_7888,N_3782,N_3579);
and U7889 (N_7889,N_4191,N_5151);
or U7890 (N_7890,N_4792,N_4832);
nand U7891 (N_7891,N_5587,N_4949);
xnor U7892 (N_7892,N_4910,N_3740);
nor U7893 (N_7893,N_4088,N_3139);
nand U7894 (N_7894,N_4699,N_5644);
nand U7895 (N_7895,N_3295,N_3558);
nor U7896 (N_7896,N_3625,N_4270);
and U7897 (N_7897,N_4214,N_3039);
xnor U7898 (N_7898,N_3659,N_5940);
xor U7899 (N_7899,N_3674,N_5202);
nor U7900 (N_7900,N_3366,N_3587);
nor U7901 (N_7901,N_5019,N_4503);
nand U7902 (N_7902,N_4083,N_3544);
nor U7903 (N_7903,N_3281,N_5958);
nand U7904 (N_7904,N_3926,N_4083);
nor U7905 (N_7905,N_4419,N_5414);
xnor U7906 (N_7906,N_4552,N_4435);
nand U7907 (N_7907,N_3958,N_5329);
nor U7908 (N_7908,N_4838,N_5570);
xor U7909 (N_7909,N_4425,N_4812);
xnor U7910 (N_7910,N_3559,N_4818);
or U7911 (N_7911,N_4236,N_3132);
and U7912 (N_7912,N_4166,N_4581);
or U7913 (N_7913,N_5690,N_5696);
nor U7914 (N_7914,N_3863,N_4036);
nor U7915 (N_7915,N_3739,N_4269);
xor U7916 (N_7916,N_3672,N_5164);
nand U7917 (N_7917,N_4657,N_4519);
nor U7918 (N_7918,N_4322,N_3809);
or U7919 (N_7919,N_3301,N_3354);
and U7920 (N_7920,N_3737,N_4749);
xnor U7921 (N_7921,N_5109,N_4734);
xor U7922 (N_7922,N_4957,N_4866);
or U7923 (N_7923,N_4583,N_3054);
xor U7924 (N_7924,N_3116,N_5275);
and U7925 (N_7925,N_3952,N_3571);
nand U7926 (N_7926,N_3626,N_5422);
nand U7927 (N_7927,N_3958,N_5232);
nor U7928 (N_7928,N_5274,N_5846);
and U7929 (N_7929,N_5330,N_3548);
nor U7930 (N_7930,N_5062,N_5008);
or U7931 (N_7931,N_3167,N_5022);
nand U7932 (N_7932,N_3579,N_4064);
nor U7933 (N_7933,N_5568,N_3365);
nor U7934 (N_7934,N_3470,N_5401);
and U7935 (N_7935,N_5579,N_3692);
or U7936 (N_7936,N_4066,N_3221);
nor U7937 (N_7937,N_5678,N_3086);
nand U7938 (N_7938,N_3072,N_5916);
nand U7939 (N_7939,N_4236,N_5678);
and U7940 (N_7940,N_3072,N_5726);
and U7941 (N_7941,N_4097,N_4501);
or U7942 (N_7942,N_4047,N_5269);
nor U7943 (N_7943,N_4275,N_5508);
nor U7944 (N_7944,N_4344,N_4488);
or U7945 (N_7945,N_5742,N_5462);
xor U7946 (N_7946,N_3845,N_5524);
xnor U7947 (N_7947,N_5288,N_5873);
and U7948 (N_7948,N_3003,N_4780);
xor U7949 (N_7949,N_4003,N_5121);
nand U7950 (N_7950,N_3527,N_5299);
and U7951 (N_7951,N_4921,N_3788);
nand U7952 (N_7952,N_5730,N_5337);
or U7953 (N_7953,N_3956,N_3709);
xor U7954 (N_7954,N_3658,N_5000);
nand U7955 (N_7955,N_5589,N_5575);
or U7956 (N_7956,N_5987,N_3697);
and U7957 (N_7957,N_5890,N_4060);
nand U7958 (N_7958,N_4789,N_4291);
nor U7959 (N_7959,N_3966,N_4620);
or U7960 (N_7960,N_4317,N_3147);
nor U7961 (N_7961,N_5390,N_4356);
nor U7962 (N_7962,N_5693,N_5367);
nor U7963 (N_7963,N_4496,N_4058);
xor U7964 (N_7964,N_4879,N_4511);
nand U7965 (N_7965,N_3394,N_5312);
nor U7966 (N_7966,N_4008,N_5764);
nor U7967 (N_7967,N_5348,N_3794);
nor U7968 (N_7968,N_3099,N_4716);
and U7969 (N_7969,N_5834,N_5641);
or U7970 (N_7970,N_4485,N_3226);
xnor U7971 (N_7971,N_4805,N_5923);
or U7972 (N_7972,N_5117,N_4272);
and U7973 (N_7973,N_5018,N_4902);
or U7974 (N_7974,N_3060,N_4336);
and U7975 (N_7975,N_5476,N_3799);
xnor U7976 (N_7976,N_3325,N_4158);
nor U7977 (N_7977,N_4512,N_5447);
or U7978 (N_7978,N_3397,N_5208);
xor U7979 (N_7979,N_4893,N_5685);
and U7980 (N_7980,N_3481,N_3892);
and U7981 (N_7981,N_3066,N_3106);
xnor U7982 (N_7982,N_5810,N_3353);
or U7983 (N_7983,N_3288,N_5747);
nand U7984 (N_7984,N_5234,N_4754);
nor U7985 (N_7985,N_3986,N_4522);
and U7986 (N_7986,N_5653,N_5179);
nand U7987 (N_7987,N_5699,N_4071);
nand U7988 (N_7988,N_3998,N_3178);
or U7989 (N_7989,N_3399,N_4922);
and U7990 (N_7990,N_4622,N_3095);
or U7991 (N_7991,N_4083,N_5430);
or U7992 (N_7992,N_3066,N_4617);
and U7993 (N_7993,N_3038,N_5856);
nand U7994 (N_7994,N_3775,N_5756);
nor U7995 (N_7995,N_3361,N_3580);
and U7996 (N_7996,N_3024,N_4974);
and U7997 (N_7997,N_5932,N_5438);
or U7998 (N_7998,N_5280,N_4156);
xor U7999 (N_7999,N_4790,N_5289);
xor U8000 (N_8000,N_5640,N_5450);
and U8001 (N_8001,N_3797,N_4907);
and U8002 (N_8002,N_4842,N_4715);
nand U8003 (N_8003,N_4066,N_4699);
xor U8004 (N_8004,N_4334,N_4670);
or U8005 (N_8005,N_4193,N_4751);
nand U8006 (N_8006,N_4057,N_4943);
xor U8007 (N_8007,N_3814,N_4035);
nand U8008 (N_8008,N_4234,N_5224);
and U8009 (N_8009,N_3922,N_3363);
nand U8010 (N_8010,N_5062,N_5492);
nor U8011 (N_8011,N_5153,N_4358);
nand U8012 (N_8012,N_5017,N_4267);
nor U8013 (N_8013,N_3036,N_5437);
nand U8014 (N_8014,N_3851,N_4610);
xor U8015 (N_8015,N_4260,N_5968);
and U8016 (N_8016,N_4384,N_4296);
or U8017 (N_8017,N_3803,N_3333);
or U8018 (N_8018,N_5343,N_4446);
and U8019 (N_8019,N_3102,N_5673);
and U8020 (N_8020,N_5766,N_5490);
or U8021 (N_8021,N_4881,N_3030);
xnor U8022 (N_8022,N_4494,N_3187);
or U8023 (N_8023,N_4679,N_3107);
or U8024 (N_8024,N_5630,N_4730);
nand U8025 (N_8025,N_5247,N_5113);
nor U8026 (N_8026,N_4380,N_5349);
and U8027 (N_8027,N_4906,N_4310);
xnor U8028 (N_8028,N_5538,N_5199);
nor U8029 (N_8029,N_5933,N_3664);
nand U8030 (N_8030,N_5067,N_5404);
or U8031 (N_8031,N_3608,N_5773);
nand U8032 (N_8032,N_5913,N_3732);
xor U8033 (N_8033,N_4541,N_5059);
xor U8034 (N_8034,N_3047,N_3451);
nor U8035 (N_8035,N_4134,N_5090);
and U8036 (N_8036,N_3543,N_4160);
xor U8037 (N_8037,N_3087,N_4356);
nand U8038 (N_8038,N_5201,N_5842);
xnor U8039 (N_8039,N_4177,N_5928);
nand U8040 (N_8040,N_5098,N_4257);
nand U8041 (N_8041,N_4309,N_4004);
and U8042 (N_8042,N_4879,N_4213);
and U8043 (N_8043,N_3347,N_3879);
xnor U8044 (N_8044,N_4441,N_3044);
and U8045 (N_8045,N_5758,N_4692);
or U8046 (N_8046,N_3416,N_3101);
or U8047 (N_8047,N_4970,N_3985);
nand U8048 (N_8048,N_5064,N_5176);
nor U8049 (N_8049,N_5598,N_3511);
nor U8050 (N_8050,N_4955,N_4609);
xor U8051 (N_8051,N_4699,N_4777);
nor U8052 (N_8052,N_4585,N_5274);
or U8053 (N_8053,N_4925,N_3383);
xor U8054 (N_8054,N_3094,N_3205);
nor U8055 (N_8055,N_4446,N_3052);
or U8056 (N_8056,N_5498,N_3538);
xor U8057 (N_8057,N_4905,N_4259);
xnor U8058 (N_8058,N_3476,N_4801);
and U8059 (N_8059,N_5022,N_5252);
xor U8060 (N_8060,N_5855,N_5332);
nor U8061 (N_8061,N_4783,N_5457);
and U8062 (N_8062,N_3605,N_4709);
nand U8063 (N_8063,N_4952,N_5568);
nand U8064 (N_8064,N_5900,N_5370);
and U8065 (N_8065,N_3865,N_5468);
or U8066 (N_8066,N_3490,N_4048);
and U8067 (N_8067,N_4588,N_4519);
nand U8068 (N_8068,N_3592,N_4037);
and U8069 (N_8069,N_5852,N_4479);
or U8070 (N_8070,N_4768,N_5611);
nand U8071 (N_8071,N_5966,N_4061);
nor U8072 (N_8072,N_3590,N_3730);
nor U8073 (N_8073,N_5477,N_4338);
xnor U8074 (N_8074,N_5882,N_5460);
xor U8075 (N_8075,N_5380,N_5482);
nor U8076 (N_8076,N_4152,N_3658);
nand U8077 (N_8077,N_5060,N_5417);
and U8078 (N_8078,N_3140,N_5785);
and U8079 (N_8079,N_3891,N_3872);
nor U8080 (N_8080,N_5857,N_5288);
nand U8081 (N_8081,N_4860,N_5354);
nor U8082 (N_8082,N_3205,N_3609);
nor U8083 (N_8083,N_5664,N_5613);
and U8084 (N_8084,N_3783,N_5454);
xor U8085 (N_8085,N_4132,N_3314);
xor U8086 (N_8086,N_3553,N_4938);
nor U8087 (N_8087,N_3818,N_4920);
or U8088 (N_8088,N_3225,N_3084);
or U8089 (N_8089,N_5679,N_4951);
nand U8090 (N_8090,N_3514,N_3757);
or U8091 (N_8091,N_5923,N_3580);
and U8092 (N_8092,N_5438,N_5268);
nor U8093 (N_8093,N_4429,N_3676);
and U8094 (N_8094,N_3494,N_5133);
nand U8095 (N_8095,N_5492,N_5187);
xor U8096 (N_8096,N_3800,N_3970);
and U8097 (N_8097,N_4486,N_4166);
nor U8098 (N_8098,N_5347,N_5130);
xor U8099 (N_8099,N_5478,N_5826);
nor U8100 (N_8100,N_4691,N_4268);
or U8101 (N_8101,N_4075,N_3041);
and U8102 (N_8102,N_3961,N_4864);
xor U8103 (N_8103,N_4544,N_5816);
or U8104 (N_8104,N_5169,N_3138);
nor U8105 (N_8105,N_5239,N_3386);
and U8106 (N_8106,N_5353,N_3837);
or U8107 (N_8107,N_3430,N_4791);
or U8108 (N_8108,N_5127,N_3790);
and U8109 (N_8109,N_5399,N_4052);
xnor U8110 (N_8110,N_4636,N_3412);
xnor U8111 (N_8111,N_3752,N_4883);
nor U8112 (N_8112,N_5546,N_3632);
nand U8113 (N_8113,N_5810,N_5172);
nor U8114 (N_8114,N_4340,N_5135);
or U8115 (N_8115,N_5992,N_4679);
or U8116 (N_8116,N_3448,N_4374);
xnor U8117 (N_8117,N_4702,N_3225);
and U8118 (N_8118,N_3349,N_3161);
xnor U8119 (N_8119,N_4585,N_4724);
xnor U8120 (N_8120,N_4760,N_3112);
nand U8121 (N_8121,N_3393,N_5608);
nor U8122 (N_8122,N_3673,N_3026);
or U8123 (N_8123,N_5867,N_3199);
nor U8124 (N_8124,N_3296,N_3365);
and U8125 (N_8125,N_4797,N_4603);
xnor U8126 (N_8126,N_3193,N_5175);
or U8127 (N_8127,N_4009,N_3048);
xnor U8128 (N_8128,N_4508,N_5217);
nand U8129 (N_8129,N_3614,N_4702);
or U8130 (N_8130,N_4640,N_4612);
or U8131 (N_8131,N_5273,N_4337);
nor U8132 (N_8132,N_4824,N_3625);
nor U8133 (N_8133,N_3928,N_4745);
nor U8134 (N_8134,N_4492,N_4452);
or U8135 (N_8135,N_3039,N_5567);
nor U8136 (N_8136,N_5247,N_4401);
nor U8137 (N_8137,N_3454,N_5085);
or U8138 (N_8138,N_4990,N_3293);
or U8139 (N_8139,N_5111,N_5635);
xor U8140 (N_8140,N_4728,N_4041);
nor U8141 (N_8141,N_4860,N_3530);
xor U8142 (N_8142,N_3929,N_5523);
nor U8143 (N_8143,N_3807,N_5752);
nand U8144 (N_8144,N_5984,N_5933);
and U8145 (N_8145,N_4368,N_5884);
xor U8146 (N_8146,N_4671,N_4852);
or U8147 (N_8147,N_3489,N_5258);
and U8148 (N_8148,N_3466,N_4961);
xnor U8149 (N_8149,N_3377,N_5074);
and U8150 (N_8150,N_5366,N_5886);
xor U8151 (N_8151,N_3879,N_3793);
or U8152 (N_8152,N_4909,N_4957);
and U8153 (N_8153,N_3816,N_5657);
xnor U8154 (N_8154,N_5605,N_3323);
or U8155 (N_8155,N_3326,N_3870);
or U8156 (N_8156,N_3150,N_4299);
xor U8157 (N_8157,N_5781,N_5794);
and U8158 (N_8158,N_5624,N_4822);
or U8159 (N_8159,N_3306,N_5871);
or U8160 (N_8160,N_3462,N_3304);
nand U8161 (N_8161,N_4237,N_3671);
and U8162 (N_8162,N_4901,N_5664);
and U8163 (N_8163,N_5744,N_3309);
nor U8164 (N_8164,N_5746,N_5011);
nand U8165 (N_8165,N_4883,N_5794);
xor U8166 (N_8166,N_3467,N_5013);
or U8167 (N_8167,N_3062,N_3933);
or U8168 (N_8168,N_4063,N_5235);
or U8169 (N_8169,N_3164,N_3607);
and U8170 (N_8170,N_5559,N_3689);
nand U8171 (N_8171,N_4782,N_4978);
or U8172 (N_8172,N_3930,N_4140);
xor U8173 (N_8173,N_3672,N_5449);
or U8174 (N_8174,N_3737,N_4087);
or U8175 (N_8175,N_5932,N_5461);
or U8176 (N_8176,N_3346,N_3455);
and U8177 (N_8177,N_3715,N_4907);
and U8178 (N_8178,N_5108,N_5978);
nor U8179 (N_8179,N_4301,N_5724);
nor U8180 (N_8180,N_5654,N_5079);
xnor U8181 (N_8181,N_5051,N_4120);
xnor U8182 (N_8182,N_4039,N_3978);
nor U8183 (N_8183,N_5711,N_5442);
and U8184 (N_8184,N_3353,N_3259);
and U8185 (N_8185,N_5808,N_3610);
or U8186 (N_8186,N_5110,N_3745);
xnor U8187 (N_8187,N_3719,N_4952);
or U8188 (N_8188,N_4128,N_3204);
or U8189 (N_8189,N_5046,N_4182);
and U8190 (N_8190,N_5663,N_3955);
nand U8191 (N_8191,N_5458,N_4262);
nand U8192 (N_8192,N_5837,N_4080);
and U8193 (N_8193,N_4172,N_5648);
xnor U8194 (N_8194,N_3510,N_4678);
nand U8195 (N_8195,N_3575,N_3914);
xnor U8196 (N_8196,N_4150,N_3774);
and U8197 (N_8197,N_5532,N_4460);
and U8198 (N_8198,N_5209,N_4048);
nor U8199 (N_8199,N_5949,N_3442);
xor U8200 (N_8200,N_5438,N_3159);
nor U8201 (N_8201,N_5688,N_4876);
nor U8202 (N_8202,N_3402,N_3403);
nor U8203 (N_8203,N_3935,N_4609);
or U8204 (N_8204,N_3913,N_5122);
nor U8205 (N_8205,N_3613,N_4934);
nor U8206 (N_8206,N_4743,N_4368);
nor U8207 (N_8207,N_3941,N_4649);
xnor U8208 (N_8208,N_5993,N_5682);
nand U8209 (N_8209,N_4750,N_3004);
and U8210 (N_8210,N_5227,N_4912);
or U8211 (N_8211,N_4500,N_4371);
and U8212 (N_8212,N_5513,N_4888);
nand U8213 (N_8213,N_5102,N_5434);
and U8214 (N_8214,N_5983,N_4918);
and U8215 (N_8215,N_4644,N_4368);
nor U8216 (N_8216,N_4299,N_5590);
xnor U8217 (N_8217,N_3378,N_5607);
nand U8218 (N_8218,N_3630,N_3239);
or U8219 (N_8219,N_5841,N_5064);
and U8220 (N_8220,N_3752,N_4059);
nand U8221 (N_8221,N_5929,N_3400);
nor U8222 (N_8222,N_4932,N_4806);
or U8223 (N_8223,N_3343,N_4383);
nor U8224 (N_8224,N_4528,N_4537);
nand U8225 (N_8225,N_4410,N_3411);
or U8226 (N_8226,N_3183,N_3129);
nor U8227 (N_8227,N_4176,N_5508);
xnor U8228 (N_8228,N_4817,N_4693);
or U8229 (N_8229,N_5859,N_5464);
or U8230 (N_8230,N_4932,N_4997);
nor U8231 (N_8231,N_5220,N_3601);
or U8232 (N_8232,N_4545,N_3481);
nand U8233 (N_8233,N_5728,N_5296);
nor U8234 (N_8234,N_5111,N_4067);
nor U8235 (N_8235,N_4466,N_3465);
and U8236 (N_8236,N_4579,N_3860);
nor U8237 (N_8237,N_3563,N_5341);
and U8238 (N_8238,N_5226,N_4122);
or U8239 (N_8239,N_3632,N_3169);
nand U8240 (N_8240,N_5095,N_3305);
nor U8241 (N_8241,N_3239,N_3774);
or U8242 (N_8242,N_5215,N_5982);
or U8243 (N_8243,N_3674,N_3231);
and U8244 (N_8244,N_4695,N_3997);
nand U8245 (N_8245,N_4499,N_3832);
and U8246 (N_8246,N_3275,N_4229);
nand U8247 (N_8247,N_4762,N_4765);
and U8248 (N_8248,N_5184,N_3981);
xor U8249 (N_8249,N_4755,N_4675);
xnor U8250 (N_8250,N_4095,N_3060);
or U8251 (N_8251,N_3460,N_4256);
xor U8252 (N_8252,N_3546,N_4967);
nand U8253 (N_8253,N_5621,N_5586);
and U8254 (N_8254,N_5355,N_4437);
or U8255 (N_8255,N_3979,N_3906);
xnor U8256 (N_8256,N_4005,N_3909);
and U8257 (N_8257,N_3861,N_4667);
nand U8258 (N_8258,N_4779,N_4201);
or U8259 (N_8259,N_5107,N_4786);
and U8260 (N_8260,N_4926,N_3742);
nor U8261 (N_8261,N_4610,N_3338);
xor U8262 (N_8262,N_3243,N_5366);
nand U8263 (N_8263,N_3361,N_3480);
or U8264 (N_8264,N_5005,N_4937);
xnor U8265 (N_8265,N_3741,N_4367);
and U8266 (N_8266,N_5908,N_5423);
or U8267 (N_8267,N_5790,N_4987);
xnor U8268 (N_8268,N_5276,N_4884);
xnor U8269 (N_8269,N_3019,N_5747);
xor U8270 (N_8270,N_3407,N_4219);
and U8271 (N_8271,N_4928,N_4826);
xnor U8272 (N_8272,N_3954,N_5294);
nor U8273 (N_8273,N_3896,N_5476);
or U8274 (N_8274,N_4700,N_4849);
or U8275 (N_8275,N_5217,N_4771);
nand U8276 (N_8276,N_5890,N_4126);
nor U8277 (N_8277,N_5749,N_4845);
or U8278 (N_8278,N_3518,N_5188);
nand U8279 (N_8279,N_3677,N_3446);
or U8280 (N_8280,N_3219,N_5888);
xor U8281 (N_8281,N_5847,N_5364);
xor U8282 (N_8282,N_3975,N_4302);
nand U8283 (N_8283,N_4921,N_4172);
xnor U8284 (N_8284,N_3055,N_3929);
nand U8285 (N_8285,N_5599,N_3129);
or U8286 (N_8286,N_5239,N_5137);
nand U8287 (N_8287,N_5230,N_5752);
nand U8288 (N_8288,N_4384,N_3317);
or U8289 (N_8289,N_3620,N_5244);
xor U8290 (N_8290,N_3055,N_3451);
nand U8291 (N_8291,N_4128,N_5282);
xor U8292 (N_8292,N_5193,N_4615);
or U8293 (N_8293,N_5733,N_3777);
nand U8294 (N_8294,N_4129,N_4808);
and U8295 (N_8295,N_5547,N_5962);
xnor U8296 (N_8296,N_4913,N_5882);
nand U8297 (N_8297,N_5063,N_5831);
nor U8298 (N_8298,N_5337,N_4854);
or U8299 (N_8299,N_5339,N_5404);
xnor U8300 (N_8300,N_4176,N_5356);
nand U8301 (N_8301,N_4205,N_3679);
nand U8302 (N_8302,N_5476,N_3338);
nor U8303 (N_8303,N_5776,N_4561);
or U8304 (N_8304,N_5818,N_3352);
and U8305 (N_8305,N_4539,N_3226);
or U8306 (N_8306,N_5145,N_4941);
nand U8307 (N_8307,N_5109,N_4151);
nand U8308 (N_8308,N_5096,N_3333);
or U8309 (N_8309,N_3375,N_4472);
nand U8310 (N_8310,N_3582,N_5849);
and U8311 (N_8311,N_4940,N_4051);
xnor U8312 (N_8312,N_5591,N_5223);
and U8313 (N_8313,N_5068,N_4949);
or U8314 (N_8314,N_4173,N_3582);
nand U8315 (N_8315,N_3292,N_5083);
nand U8316 (N_8316,N_3786,N_3587);
and U8317 (N_8317,N_4078,N_4872);
or U8318 (N_8318,N_3508,N_3375);
and U8319 (N_8319,N_3255,N_4251);
or U8320 (N_8320,N_4063,N_4024);
xor U8321 (N_8321,N_3658,N_4793);
nor U8322 (N_8322,N_5378,N_3572);
or U8323 (N_8323,N_4667,N_3143);
or U8324 (N_8324,N_5766,N_4136);
nand U8325 (N_8325,N_3042,N_3454);
nand U8326 (N_8326,N_4005,N_3656);
nand U8327 (N_8327,N_4875,N_5696);
and U8328 (N_8328,N_3971,N_3013);
nand U8329 (N_8329,N_5469,N_3034);
nor U8330 (N_8330,N_3206,N_5412);
xor U8331 (N_8331,N_3415,N_4648);
and U8332 (N_8332,N_5924,N_5816);
nand U8333 (N_8333,N_4008,N_5293);
xnor U8334 (N_8334,N_5007,N_5445);
xor U8335 (N_8335,N_4631,N_5314);
nor U8336 (N_8336,N_5229,N_5270);
or U8337 (N_8337,N_4442,N_4322);
xnor U8338 (N_8338,N_5143,N_5373);
and U8339 (N_8339,N_3904,N_3981);
xor U8340 (N_8340,N_4948,N_4710);
nor U8341 (N_8341,N_5459,N_5607);
or U8342 (N_8342,N_5336,N_5822);
and U8343 (N_8343,N_4371,N_4618);
nand U8344 (N_8344,N_5610,N_4424);
or U8345 (N_8345,N_5430,N_4695);
nand U8346 (N_8346,N_4041,N_4363);
or U8347 (N_8347,N_3278,N_5783);
nand U8348 (N_8348,N_5866,N_3286);
and U8349 (N_8349,N_3220,N_3035);
nand U8350 (N_8350,N_4650,N_4405);
and U8351 (N_8351,N_4008,N_5863);
nand U8352 (N_8352,N_5280,N_3545);
xnor U8353 (N_8353,N_3726,N_4184);
nand U8354 (N_8354,N_3234,N_5505);
xnor U8355 (N_8355,N_3057,N_3939);
or U8356 (N_8356,N_5297,N_3318);
nor U8357 (N_8357,N_4896,N_5423);
and U8358 (N_8358,N_5245,N_5301);
nor U8359 (N_8359,N_5022,N_3752);
or U8360 (N_8360,N_4227,N_5773);
and U8361 (N_8361,N_5504,N_5353);
or U8362 (N_8362,N_4669,N_5194);
nand U8363 (N_8363,N_5927,N_4277);
and U8364 (N_8364,N_3539,N_4757);
xor U8365 (N_8365,N_3761,N_4018);
nor U8366 (N_8366,N_3409,N_5277);
xor U8367 (N_8367,N_3302,N_5065);
nor U8368 (N_8368,N_5493,N_4209);
nand U8369 (N_8369,N_3170,N_3356);
or U8370 (N_8370,N_5385,N_5998);
or U8371 (N_8371,N_5249,N_4079);
or U8372 (N_8372,N_3964,N_5316);
nand U8373 (N_8373,N_3493,N_5215);
or U8374 (N_8374,N_4879,N_5897);
xnor U8375 (N_8375,N_5034,N_3043);
xor U8376 (N_8376,N_4403,N_3841);
nand U8377 (N_8377,N_3320,N_5338);
nand U8378 (N_8378,N_4176,N_3632);
nand U8379 (N_8379,N_4719,N_3150);
and U8380 (N_8380,N_3698,N_5738);
and U8381 (N_8381,N_3693,N_4060);
nor U8382 (N_8382,N_5800,N_3279);
xnor U8383 (N_8383,N_5188,N_3374);
and U8384 (N_8384,N_3216,N_5000);
nor U8385 (N_8385,N_4119,N_3333);
xor U8386 (N_8386,N_4628,N_3552);
xor U8387 (N_8387,N_5592,N_5480);
nand U8388 (N_8388,N_3791,N_5345);
nor U8389 (N_8389,N_4126,N_5007);
nor U8390 (N_8390,N_4094,N_3460);
or U8391 (N_8391,N_3903,N_5593);
nor U8392 (N_8392,N_3818,N_4969);
or U8393 (N_8393,N_4208,N_5266);
nand U8394 (N_8394,N_4295,N_3253);
or U8395 (N_8395,N_4231,N_4565);
nor U8396 (N_8396,N_4038,N_4408);
xnor U8397 (N_8397,N_4870,N_5439);
or U8398 (N_8398,N_5703,N_5355);
nand U8399 (N_8399,N_5641,N_5946);
nand U8400 (N_8400,N_4576,N_3468);
nand U8401 (N_8401,N_5019,N_4718);
and U8402 (N_8402,N_3982,N_5005);
or U8403 (N_8403,N_5797,N_5267);
and U8404 (N_8404,N_3309,N_3007);
nand U8405 (N_8405,N_5677,N_4653);
xor U8406 (N_8406,N_4458,N_5640);
and U8407 (N_8407,N_3352,N_4508);
nor U8408 (N_8408,N_4261,N_4398);
and U8409 (N_8409,N_3121,N_5244);
nor U8410 (N_8410,N_3775,N_4941);
nand U8411 (N_8411,N_3316,N_4394);
nand U8412 (N_8412,N_5333,N_5526);
xor U8413 (N_8413,N_3198,N_5580);
nor U8414 (N_8414,N_5349,N_5473);
nor U8415 (N_8415,N_5654,N_4226);
xor U8416 (N_8416,N_5632,N_5582);
or U8417 (N_8417,N_3964,N_3902);
and U8418 (N_8418,N_5458,N_3924);
or U8419 (N_8419,N_4142,N_3112);
and U8420 (N_8420,N_4795,N_3635);
or U8421 (N_8421,N_3259,N_3735);
xor U8422 (N_8422,N_4822,N_3422);
xnor U8423 (N_8423,N_3495,N_3211);
or U8424 (N_8424,N_3543,N_5249);
nand U8425 (N_8425,N_4120,N_3210);
and U8426 (N_8426,N_4680,N_3596);
or U8427 (N_8427,N_4491,N_3427);
nand U8428 (N_8428,N_3715,N_5858);
or U8429 (N_8429,N_3944,N_5997);
and U8430 (N_8430,N_4222,N_3982);
and U8431 (N_8431,N_3282,N_3313);
xnor U8432 (N_8432,N_4161,N_5758);
nor U8433 (N_8433,N_5902,N_4901);
or U8434 (N_8434,N_4272,N_3335);
and U8435 (N_8435,N_4349,N_3935);
nor U8436 (N_8436,N_5442,N_4984);
and U8437 (N_8437,N_4924,N_3460);
xnor U8438 (N_8438,N_4186,N_5261);
or U8439 (N_8439,N_4998,N_5871);
xor U8440 (N_8440,N_5931,N_5023);
nand U8441 (N_8441,N_5512,N_5240);
or U8442 (N_8442,N_4858,N_4468);
nand U8443 (N_8443,N_3077,N_5851);
and U8444 (N_8444,N_5694,N_3532);
and U8445 (N_8445,N_3776,N_5658);
or U8446 (N_8446,N_3471,N_4260);
nand U8447 (N_8447,N_3701,N_3214);
xnor U8448 (N_8448,N_4579,N_5829);
xor U8449 (N_8449,N_5909,N_5336);
and U8450 (N_8450,N_4827,N_4371);
xnor U8451 (N_8451,N_3380,N_3148);
and U8452 (N_8452,N_4522,N_5184);
or U8453 (N_8453,N_5443,N_4771);
nand U8454 (N_8454,N_4658,N_5536);
nor U8455 (N_8455,N_5989,N_3124);
nor U8456 (N_8456,N_5050,N_4962);
nand U8457 (N_8457,N_4951,N_4896);
and U8458 (N_8458,N_5450,N_4536);
or U8459 (N_8459,N_4359,N_4607);
or U8460 (N_8460,N_5335,N_4398);
or U8461 (N_8461,N_5310,N_3319);
xnor U8462 (N_8462,N_5390,N_4123);
and U8463 (N_8463,N_5219,N_4347);
and U8464 (N_8464,N_5646,N_3222);
and U8465 (N_8465,N_4515,N_4157);
nor U8466 (N_8466,N_5504,N_5890);
and U8467 (N_8467,N_4598,N_5572);
xnor U8468 (N_8468,N_4558,N_4043);
and U8469 (N_8469,N_3393,N_3483);
and U8470 (N_8470,N_3147,N_4661);
or U8471 (N_8471,N_5395,N_3699);
and U8472 (N_8472,N_5106,N_4533);
and U8473 (N_8473,N_4384,N_4312);
or U8474 (N_8474,N_4257,N_5243);
nand U8475 (N_8475,N_3208,N_5195);
and U8476 (N_8476,N_5646,N_5784);
nand U8477 (N_8477,N_5153,N_5248);
and U8478 (N_8478,N_4314,N_5191);
nand U8479 (N_8479,N_4027,N_3918);
and U8480 (N_8480,N_5282,N_3330);
nand U8481 (N_8481,N_5462,N_5791);
or U8482 (N_8482,N_4080,N_5678);
nand U8483 (N_8483,N_5409,N_5544);
xnor U8484 (N_8484,N_4083,N_4193);
nor U8485 (N_8485,N_3280,N_4156);
nor U8486 (N_8486,N_3507,N_5141);
and U8487 (N_8487,N_4441,N_4556);
and U8488 (N_8488,N_3528,N_3671);
or U8489 (N_8489,N_3896,N_3732);
xnor U8490 (N_8490,N_5433,N_3843);
and U8491 (N_8491,N_5962,N_4810);
nand U8492 (N_8492,N_4575,N_4042);
xor U8493 (N_8493,N_5374,N_5560);
nor U8494 (N_8494,N_3633,N_5940);
and U8495 (N_8495,N_3008,N_3323);
or U8496 (N_8496,N_3297,N_4921);
and U8497 (N_8497,N_3112,N_5263);
and U8498 (N_8498,N_3701,N_4323);
nor U8499 (N_8499,N_4394,N_3217);
nor U8500 (N_8500,N_4142,N_5730);
or U8501 (N_8501,N_3991,N_4428);
nor U8502 (N_8502,N_4139,N_5793);
nand U8503 (N_8503,N_3995,N_5467);
nand U8504 (N_8504,N_3633,N_3206);
xor U8505 (N_8505,N_4625,N_3026);
or U8506 (N_8506,N_3895,N_5735);
xor U8507 (N_8507,N_4718,N_3639);
nor U8508 (N_8508,N_3609,N_5417);
nand U8509 (N_8509,N_5541,N_5929);
nor U8510 (N_8510,N_5795,N_4742);
xor U8511 (N_8511,N_3683,N_5712);
nor U8512 (N_8512,N_3073,N_3572);
or U8513 (N_8513,N_4925,N_4431);
or U8514 (N_8514,N_5884,N_3317);
nand U8515 (N_8515,N_4769,N_5815);
nor U8516 (N_8516,N_5805,N_5385);
and U8517 (N_8517,N_3597,N_4960);
or U8518 (N_8518,N_3972,N_5239);
or U8519 (N_8519,N_3518,N_5448);
and U8520 (N_8520,N_5986,N_5309);
and U8521 (N_8521,N_4748,N_3307);
xnor U8522 (N_8522,N_3448,N_3510);
or U8523 (N_8523,N_4656,N_4391);
nor U8524 (N_8524,N_5057,N_3534);
xor U8525 (N_8525,N_5813,N_3441);
or U8526 (N_8526,N_5016,N_5261);
and U8527 (N_8527,N_3626,N_5806);
xnor U8528 (N_8528,N_5586,N_4053);
and U8529 (N_8529,N_3368,N_4366);
nor U8530 (N_8530,N_3150,N_5932);
xnor U8531 (N_8531,N_5577,N_3577);
and U8532 (N_8532,N_5220,N_3842);
or U8533 (N_8533,N_4586,N_4746);
and U8534 (N_8534,N_5972,N_5874);
xor U8535 (N_8535,N_5510,N_4353);
or U8536 (N_8536,N_4214,N_5481);
and U8537 (N_8537,N_4239,N_4443);
nand U8538 (N_8538,N_5409,N_3761);
xor U8539 (N_8539,N_3357,N_4697);
nand U8540 (N_8540,N_5143,N_5475);
or U8541 (N_8541,N_5049,N_4959);
and U8542 (N_8542,N_4806,N_5035);
xnor U8543 (N_8543,N_5090,N_3705);
or U8544 (N_8544,N_5778,N_5298);
or U8545 (N_8545,N_3681,N_4139);
or U8546 (N_8546,N_5642,N_5080);
xnor U8547 (N_8547,N_4199,N_5222);
nor U8548 (N_8548,N_4397,N_5738);
nand U8549 (N_8549,N_3595,N_3660);
xor U8550 (N_8550,N_5629,N_4994);
xor U8551 (N_8551,N_4848,N_4474);
and U8552 (N_8552,N_3987,N_4715);
and U8553 (N_8553,N_4923,N_5782);
or U8554 (N_8554,N_5324,N_4844);
and U8555 (N_8555,N_4394,N_5925);
nand U8556 (N_8556,N_5846,N_3970);
or U8557 (N_8557,N_4880,N_3983);
xnor U8558 (N_8558,N_4463,N_5624);
nor U8559 (N_8559,N_4998,N_5522);
nor U8560 (N_8560,N_3780,N_4234);
xnor U8561 (N_8561,N_4229,N_5762);
and U8562 (N_8562,N_5777,N_4149);
xor U8563 (N_8563,N_3552,N_4611);
nor U8564 (N_8564,N_3762,N_3396);
nor U8565 (N_8565,N_5490,N_4694);
xor U8566 (N_8566,N_3872,N_4954);
or U8567 (N_8567,N_4434,N_3521);
nand U8568 (N_8568,N_3403,N_3746);
xor U8569 (N_8569,N_4715,N_4963);
nand U8570 (N_8570,N_3232,N_3589);
nand U8571 (N_8571,N_5709,N_5332);
nand U8572 (N_8572,N_3791,N_3120);
or U8573 (N_8573,N_4380,N_5873);
or U8574 (N_8574,N_4114,N_5544);
nor U8575 (N_8575,N_4807,N_4996);
nor U8576 (N_8576,N_3196,N_5106);
xnor U8577 (N_8577,N_4653,N_5944);
nand U8578 (N_8578,N_4518,N_4342);
or U8579 (N_8579,N_3611,N_5668);
xor U8580 (N_8580,N_3143,N_4030);
nand U8581 (N_8581,N_3044,N_4642);
xnor U8582 (N_8582,N_4465,N_5599);
and U8583 (N_8583,N_4450,N_5027);
nor U8584 (N_8584,N_3905,N_5232);
nor U8585 (N_8585,N_3731,N_5842);
and U8586 (N_8586,N_3227,N_5896);
nor U8587 (N_8587,N_5940,N_4234);
nand U8588 (N_8588,N_4116,N_3777);
or U8589 (N_8589,N_3758,N_3792);
nand U8590 (N_8590,N_5529,N_3946);
nand U8591 (N_8591,N_3617,N_4323);
and U8592 (N_8592,N_4540,N_3081);
nor U8593 (N_8593,N_5653,N_5500);
or U8594 (N_8594,N_4418,N_5793);
nor U8595 (N_8595,N_4521,N_5945);
nand U8596 (N_8596,N_3597,N_5558);
or U8597 (N_8597,N_4139,N_4127);
nand U8598 (N_8598,N_3443,N_3037);
nor U8599 (N_8599,N_5406,N_4423);
nor U8600 (N_8600,N_3677,N_3600);
or U8601 (N_8601,N_5545,N_3443);
xnor U8602 (N_8602,N_3697,N_5340);
nand U8603 (N_8603,N_4131,N_5617);
and U8604 (N_8604,N_5401,N_5864);
nor U8605 (N_8605,N_5138,N_5425);
xor U8606 (N_8606,N_3634,N_3074);
nand U8607 (N_8607,N_4992,N_4761);
nand U8608 (N_8608,N_5219,N_4092);
xnor U8609 (N_8609,N_4438,N_4834);
xor U8610 (N_8610,N_5247,N_4509);
or U8611 (N_8611,N_4054,N_3323);
nor U8612 (N_8612,N_3292,N_3259);
xnor U8613 (N_8613,N_4841,N_3489);
or U8614 (N_8614,N_3280,N_3081);
and U8615 (N_8615,N_3186,N_4330);
nand U8616 (N_8616,N_3443,N_3989);
xor U8617 (N_8617,N_4446,N_5255);
and U8618 (N_8618,N_3622,N_4229);
or U8619 (N_8619,N_3330,N_3939);
xnor U8620 (N_8620,N_4167,N_3380);
nand U8621 (N_8621,N_4507,N_3547);
or U8622 (N_8622,N_3640,N_5388);
nor U8623 (N_8623,N_5938,N_3223);
or U8624 (N_8624,N_4368,N_3798);
xnor U8625 (N_8625,N_4634,N_3841);
or U8626 (N_8626,N_5250,N_4068);
nor U8627 (N_8627,N_5424,N_4422);
nor U8628 (N_8628,N_4916,N_3018);
or U8629 (N_8629,N_5958,N_5495);
and U8630 (N_8630,N_5699,N_4400);
xor U8631 (N_8631,N_4885,N_5206);
nand U8632 (N_8632,N_4944,N_5944);
xor U8633 (N_8633,N_4669,N_3901);
nor U8634 (N_8634,N_5885,N_4226);
nand U8635 (N_8635,N_5707,N_5160);
nand U8636 (N_8636,N_4924,N_3515);
nand U8637 (N_8637,N_5607,N_5720);
nand U8638 (N_8638,N_4858,N_4130);
nor U8639 (N_8639,N_3266,N_5961);
nor U8640 (N_8640,N_5216,N_4855);
or U8641 (N_8641,N_4690,N_5067);
nor U8642 (N_8642,N_5478,N_5696);
and U8643 (N_8643,N_3470,N_5533);
nor U8644 (N_8644,N_5029,N_5053);
or U8645 (N_8645,N_3996,N_4285);
nor U8646 (N_8646,N_5528,N_3133);
and U8647 (N_8647,N_5426,N_4960);
and U8648 (N_8648,N_5259,N_3535);
and U8649 (N_8649,N_4941,N_3713);
xor U8650 (N_8650,N_4211,N_4834);
nor U8651 (N_8651,N_3515,N_4283);
or U8652 (N_8652,N_3188,N_3203);
nand U8653 (N_8653,N_3144,N_4183);
nand U8654 (N_8654,N_4647,N_4287);
nor U8655 (N_8655,N_5494,N_5283);
nor U8656 (N_8656,N_5645,N_4296);
and U8657 (N_8657,N_5129,N_3977);
or U8658 (N_8658,N_5954,N_5084);
or U8659 (N_8659,N_3377,N_4138);
nor U8660 (N_8660,N_5655,N_5897);
xnor U8661 (N_8661,N_3898,N_4159);
xnor U8662 (N_8662,N_5667,N_4014);
nand U8663 (N_8663,N_3624,N_3886);
xor U8664 (N_8664,N_4806,N_4703);
and U8665 (N_8665,N_4610,N_4145);
nor U8666 (N_8666,N_4417,N_4980);
nand U8667 (N_8667,N_5000,N_4969);
or U8668 (N_8668,N_5714,N_3569);
xnor U8669 (N_8669,N_5650,N_4973);
nor U8670 (N_8670,N_3900,N_5276);
and U8671 (N_8671,N_4541,N_5259);
and U8672 (N_8672,N_5302,N_4208);
xor U8673 (N_8673,N_3992,N_5842);
and U8674 (N_8674,N_4172,N_5133);
nand U8675 (N_8675,N_3004,N_3799);
nor U8676 (N_8676,N_5099,N_4278);
nand U8677 (N_8677,N_3838,N_4695);
or U8678 (N_8678,N_3324,N_4114);
nor U8679 (N_8679,N_3259,N_3699);
nand U8680 (N_8680,N_3483,N_3234);
and U8681 (N_8681,N_4472,N_4455);
nand U8682 (N_8682,N_5156,N_4024);
nor U8683 (N_8683,N_5713,N_3951);
xnor U8684 (N_8684,N_3669,N_4156);
xnor U8685 (N_8685,N_3017,N_3372);
or U8686 (N_8686,N_3978,N_3175);
nand U8687 (N_8687,N_3731,N_5087);
or U8688 (N_8688,N_3703,N_4150);
or U8689 (N_8689,N_3534,N_4084);
or U8690 (N_8690,N_3390,N_3413);
or U8691 (N_8691,N_4290,N_5619);
and U8692 (N_8692,N_4065,N_5434);
or U8693 (N_8693,N_4628,N_5604);
xor U8694 (N_8694,N_4905,N_4260);
and U8695 (N_8695,N_4369,N_3316);
nor U8696 (N_8696,N_5504,N_5320);
nand U8697 (N_8697,N_3436,N_3976);
nor U8698 (N_8698,N_4506,N_4989);
nor U8699 (N_8699,N_4653,N_4517);
or U8700 (N_8700,N_5948,N_3746);
nor U8701 (N_8701,N_4246,N_5670);
or U8702 (N_8702,N_4321,N_4305);
and U8703 (N_8703,N_5168,N_4547);
nor U8704 (N_8704,N_5743,N_3782);
xnor U8705 (N_8705,N_3147,N_4552);
nor U8706 (N_8706,N_5317,N_4962);
or U8707 (N_8707,N_3797,N_5226);
nor U8708 (N_8708,N_5680,N_3155);
or U8709 (N_8709,N_3957,N_3996);
nor U8710 (N_8710,N_4057,N_3724);
nor U8711 (N_8711,N_3122,N_4146);
nor U8712 (N_8712,N_3120,N_3260);
nor U8713 (N_8713,N_4563,N_5807);
xor U8714 (N_8714,N_4912,N_3398);
xor U8715 (N_8715,N_5544,N_5429);
or U8716 (N_8716,N_3955,N_5317);
or U8717 (N_8717,N_4115,N_5710);
nor U8718 (N_8718,N_3439,N_3358);
and U8719 (N_8719,N_3788,N_5873);
and U8720 (N_8720,N_3527,N_3248);
xnor U8721 (N_8721,N_5112,N_4422);
and U8722 (N_8722,N_4836,N_5686);
xnor U8723 (N_8723,N_5218,N_4889);
or U8724 (N_8724,N_3172,N_4176);
and U8725 (N_8725,N_5797,N_4339);
nor U8726 (N_8726,N_4105,N_4411);
xor U8727 (N_8727,N_5812,N_3099);
or U8728 (N_8728,N_5803,N_5225);
xnor U8729 (N_8729,N_5254,N_3825);
nand U8730 (N_8730,N_4664,N_3075);
or U8731 (N_8731,N_4871,N_5486);
or U8732 (N_8732,N_5316,N_5624);
or U8733 (N_8733,N_5589,N_5152);
or U8734 (N_8734,N_4622,N_4462);
or U8735 (N_8735,N_5705,N_3197);
nor U8736 (N_8736,N_5098,N_4759);
and U8737 (N_8737,N_3381,N_5484);
nand U8738 (N_8738,N_4493,N_3046);
xnor U8739 (N_8739,N_3276,N_4688);
or U8740 (N_8740,N_3517,N_3669);
and U8741 (N_8741,N_3322,N_3364);
xor U8742 (N_8742,N_3015,N_4312);
and U8743 (N_8743,N_4082,N_3191);
nand U8744 (N_8744,N_4090,N_4381);
nand U8745 (N_8745,N_4509,N_5113);
or U8746 (N_8746,N_4093,N_5932);
nand U8747 (N_8747,N_4829,N_5991);
nor U8748 (N_8748,N_4102,N_5695);
or U8749 (N_8749,N_5886,N_3839);
nor U8750 (N_8750,N_3367,N_4534);
or U8751 (N_8751,N_5443,N_5275);
or U8752 (N_8752,N_4241,N_3896);
xor U8753 (N_8753,N_3629,N_5255);
xor U8754 (N_8754,N_3557,N_3195);
xnor U8755 (N_8755,N_4348,N_4753);
xor U8756 (N_8756,N_3317,N_3377);
or U8757 (N_8757,N_5666,N_4977);
or U8758 (N_8758,N_3128,N_5304);
nor U8759 (N_8759,N_5754,N_5057);
nand U8760 (N_8760,N_3124,N_3314);
nor U8761 (N_8761,N_4337,N_4613);
or U8762 (N_8762,N_5287,N_4055);
and U8763 (N_8763,N_3005,N_4724);
nand U8764 (N_8764,N_3054,N_5508);
nor U8765 (N_8765,N_3379,N_3862);
or U8766 (N_8766,N_4439,N_4831);
or U8767 (N_8767,N_3847,N_4703);
and U8768 (N_8768,N_4821,N_5562);
and U8769 (N_8769,N_4777,N_4579);
nor U8770 (N_8770,N_4382,N_4385);
nand U8771 (N_8771,N_3327,N_5345);
nor U8772 (N_8772,N_3987,N_5076);
xnor U8773 (N_8773,N_4645,N_5831);
or U8774 (N_8774,N_5845,N_4677);
xor U8775 (N_8775,N_3985,N_4313);
or U8776 (N_8776,N_3394,N_4840);
xor U8777 (N_8777,N_3827,N_5089);
nor U8778 (N_8778,N_3256,N_3320);
or U8779 (N_8779,N_5947,N_4651);
nor U8780 (N_8780,N_3605,N_4885);
nor U8781 (N_8781,N_4674,N_4493);
nor U8782 (N_8782,N_4770,N_4166);
nor U8783 (N_8783,N_4148,N_3407);
xor U8784 (N_8784,N_3393,N_4657);
and U8785 (N_8785,N_5105,N_4441);
or U8786 (N_8786,N_3141,N_5203);
nor U8787 (N_8787,N_4538,N_4310);
nand U8788 (N_8788,N_5668,N_3249);
nor U8789 (N_8789,N_5094,N_5043);
xor U8790 (N_8790,N_5479,N_3498);
xor U8791 (N_8791,N_3457,N_5836);
and U8792 (N_8792,N_4711,N_5475);
or U8793 (N_8793,N_3284,N_3809);
nor U8794 (N_8794,N_4184,N_3604);
and U8795 (N_8795,N_3010,N_3372);
nand U8796 (N_8796,N_4893,N_3547);
nand U8797 (N_8797,N_3252,N_5349);
nor U8798 (N_8798,N_4965,N_5317);
xnor U8799 (N_8799,N_5757,N_4357);
nand U8800 (N_8800,N_3368,N_4583);
and U8801 (N_8801,N_5681,N_3092);
xnor U8802 (N_8802,N_5293,N_3379);
and U8803 (N_8803,N_4165,N_4354);
nor U8804 (N_8804,N_5700,N_3605);
and U8805 (N_8805,N_5661,N_3676);
and U8806 (N_8806,N_3489,N_3055);
xnor U8807 (N_8807,N_4836,N_4559);
nand U8808 (N_8808,N_3264,N_5257);
or U8809 (N_8809,N_5317,N_3531);
nor U8810 (N_8810,N_5083,N_3435);
xnor U8811 (N_8811,N_5603,N_3555);
nor U8812 (N_8812,N_5576,N_3027);
or U8813 (N_8813,N_5190,N_3950);
nand U8814 (N_8814,N_4925,N_4751);
xnor U8815 (N_8815,N_4158,N_5045);
nand U8816 (N_8816,N_3096,N_4675);
xnor U8817 (N_8817,N_3315,N_4400);
nand U8818 (N_8818,N_5734,N_3634);
nor U8819 (N_8819,N_5502,N_3909);
nand U8820 (N_8820,N_4449,N_4486);
and U8821 (N_8821,N_5464,N_4548);
nor U8822 (N_8822,N_3928,N_5044);
and U8823 (N_8823,N_5305,N_4368);
and U8824 (N_8824,N_5501,N_5723);
and U8825 (N_8825,N_5798,N_5922);
nand U8826 (N_8826,N_5712,N_4916);
or U8827 (N_8827,N_5250,N_3640);
and U8828 (N_8828,N_4359,N_5716);
and U8829 (N_8829,N_5340,N_3332);
xnor U8830 (N_8830,N_3575,N_5722);
nor U8831 (N_8831,N_4425,N_5850);
and U8832 (N_8832,N_4140,N_3328);
nor U8833 (N_8833,N_5999,N_5075);
or U8834 (N_8834,N_4561,N_5531);
nor U8835 (N_8835,N_4950,N_4716);
nor U8836 (N_8836,N_5993,N_3906);
or U8837 (N_8837,N_5146,N_3061);
xnor U8838 (N_8838,N_4126,N_5343);
or U8839 (N_8839,N_3305,N_4297);
nor U8840 (N_8840,N_5306,N_3447);
and U8841 (N_8841,N_5334,N_5731);
nand U8842 (N_8842,N_3678,N_3151);
xor U8843 (N_8843,N_3118,N_5048);
or U8844 (N_8844,N_5556,N_3468);
nand U8845 (N_8845,N_3130,N_5773);
or U8846 (N_8846,N_3076,N_5536);
and U8847 (N_8847,N_3051,N_5513);
nand U8848 (N_8848,N_5025,N_5194);
xor U8849 (N_8849,N_3722,N_4253);
xnor U8850 (N_8850,N_4507,N_3886);
xnor U8851 (N_8851,N_4225,N_4149);
nand U8852 (N_8852,N_4319,N_5265);
or U8853 (N_8853,N_3205,N_3632);
and U8854 (N_8854,N_4806,N_3514);
and U8855 (N_8855,N_4798,N_4369);
nand U8856 (N_8856,N_4322,N_3454);
xor U8857 (N_8857,N_5827,N_5849);
xnor U8858 (N_8858,N_3722,N_3034);
nor U8859 (N_8859,N_3375,N_4984);
xor U8860 (N_8860,N_4992,N_4598);
nor U8861 (N_8861,N_3058,N_3284);
or U8862 (N_8862,N_4598,N_4513);
nand U8863 (N_8863,N_4388,N_4153);
and U8864 (N_8864,N_3741,N_5328);
nand U8865 (N_8865,N_5128,N_5883);
or U8866 (N_8866,N_3055,N_4445);
nor U8867 (N_8867,N_5373,N_3113);
nor U8868 (N_8868,N_4694,N_3573);
nor U8869 (N_8869,N_3682,N_4652);
nor U8870 (N_8870,N_4915,N_5637);
nand U8871 (N_8871,N_4597,N_3742);
nand U8872 (N_8872,N_4105,N_4426);
or U8873 (N_8873,N_3447,N_3521);
nor U8874 (N_8874,N_4748,N_4388);
and U8875 (N_8875,N_3484,N_5056);
and U8876 (N_8876,N_3382,N_4050);
and U8877 (N_8877,N_5036,N_3309);
and U8878 (N_8878,N_4785,N_3020);
or U8879 (N_8879,N_4401,N_5046);
nand U8880 (N_8880,N_5490,N_3092);
nand U8881 (N_8881,N_3606,N_5550);
nor U8882 (N_8882,N_4821,N_5943);
nand U8883 (N_8883,N_5080,N_5387);
nor U8884 (N_8884,N_5514,N_4225);
and U8885 (N_8885,N_5859,N_5263);
nand U8886 (N_8886,N_5013,N_4225);
nand U8887 (N_8887,N_5146,N_4655);
or U8888 (N_8888,N_5503,N_4468);
xnor U8889 (N_8889,N_4904,N_3121);
or U8890 (N_8890,N_5752,N_3458);
xnor U8891 (N_8891,N_4273,N_3955);
or U8892 (N_8892,N_5231,N_4337);
xor U8893 (N_8893,N_3718,N_3602);
or U8894 (N_8894,N_4705,N_3464);
nand U8895 (N_8895,N_4744,N_5232);
nand U8896 (N_8896,N_5695,N_5968);
xnor U8897 (N_8897,N_3471,N_5657);
xor U8898 (N_8898,N_5443,N_3615);
xnor U8899 (N_8899,N_3609,N_3422);
and U8900 (N_8900,N_3594,N_3244);
nor U8901 (N_8901,N_4294,N_4673);
or U8902 (N_8902,N_4876,N_3781);
nor U8903 (N_8903,N_3481,N_5993);
or U8904 (N_8904,N_4656,N_3465);
nand U8905 (N_8905,N_5408,N_5667);
nor U8906 (N_8906,N_5491,N_3789);
and U8907 (N_8907,N_4528,N_5976);
nor U8908 (N_8908,N_3417,N_5708);
nor U8909 (N_8909,N_4198,N_4030);
xor U8910 (N_8910,N_5071,N_3757);
and U8911 (N_8911,N_3327,N_3344);
or U8912 (N_8912,N_4769,N_5481);
nor U8913 (N_8913,N_3997,N_3871);
and U8914 (N_8914,N_5233,N_4082);
nand U8915 (N_8915,N_3492,N_3182);
xor U8916 (N_8916,N_5338,N_4801);
nand U8917 (N_8917,N_4836,N_5373);
nand U8918 (N_8918,N_4560,N_5116);
and U8919 (N_8919,N_3239,N_4090);
or U8920 (N_8920,N_3924,N_4750);
nand U8921 (N_8921,N_3228,N_4631);
nand U8922 (N_8922,N_5768,N_3409);
nand U8923 (N_8923,N_4582,N_4305);
or U8924 (N_8924,N_5896,N_5937);
nand U8925 (N_8925,N_4897,N_5741);
nor U8926 (N_8926,N_4000,N_5279);
xor U8927 (N_8927,N_5089,N_3719);
nor U8928 (N_8928,N_3732,N_5383);
nor U8929 (N_8929,N_5709,N_4273);
nor U8930 (N_8930,N_3058,N_5846);
xnor U8931 (N_8931,N_4222,N_4010);
or U8932 (N_8932,N_3967,N_5512);
or U8933 (N_8933,N_3154,N_5216);
and U8934 (N_8934,N_5563,N_3452);
nor U8935 (N_8935,N_3326,N_3689);
nor U8936 (N_8936,N_5542,N_5197);
nor U8937 (N_8937,N_5561,N_5168);
nand U8938 (N_8938,N_4987,N_5636);
xnor U8939 (N_8939,N_3760,N_3751);
nor U8940 (N_8940,N_4053,N_3260);
nand U8941 (N_8941,N_4473,N_3543);
nor U8942 (N_8942,N_5638,N_5340);
nand U8943 (N_8943,N_4409,N_4372);
nand U8944 (N_8944,N_5725,N_4369);
and U8945 (N_8945,N_4304,N_4019);
or U8946 (N_8946,N_3075,N_5121);
xnor U8947 (N_8947,N_5303,N_3663);
nor U8948 (N_8948,N_5764,N_3737);
nor U8949 (N_8949,N_3158,N_4696);
nand U8950 (N_8950,N_3893,N_4304);
xor U8951 (N_8951,N_3018,N_3492);
and U8952 (N_8952,N_4779,N_5420);
nor U8953 (N_8953,N_4621,N_4537);
nand U8954 (N_8954,N_4369,N_5472);
nor U8955 (N_8955,N_5734,N_5510);
xor U8956 (N_8956,N_3169,N_5645);
or U8957 (N_8957,N_3050,N_3348);
nand U8958 (N_8958,N_5784,N_3163);
or U8959 (N_8959,N_5816,N_4649);
and U8960 (N_8960,N_5121,N_5026);
and U8961 (N_8961,N_5801,N_3084);
or U8962 (N_8962,N_4838,N_3379);
or U8963 (N_8963,N_4245,N_3539);
and U8964 (N_8964,N_5602,N_3018);
and U8965 (N_8965,N_3118,N_4348);
or U8966 (N_8966,N_5366,N_4931);
nand U8967 (N_8967,N_3841,N_5772);
or U8968 (N_8968,N_3687,N_3547);
xor U8969 (N_8969,N_4087,N_3648);
and U8970 (N_8970,N_5986,N_4168);
nor U8971 (N_8971,N_4034,N_3806);
or U8972 (N_8972,N_3602,N_3192);
nand U8973 (N_8973,N_3684,N_5210);
and U8974 (N_8974,N_4965,N_5158);
nor U8975 (N_8975,N_5268,N_5147);
nor U8976 (N_8976,N_4719,N_3812);
nand U8977 (N_8977,N_4757,N_3042);
nand U8978 (N_8978,N_4884,N_5709);
nand U8979 (N_8979,N_5168,N_3532);
nand U8980 (N_8980,N_4453,N_5245);
xor U8981 (N_8981,N_3226,N_5771);
and U8982 (N_8982,N_3088,N_5564);
or U8983 (N_8983,N_4850,N_5459);
and U8984 (N_8984,N_5437,N_4173);
nand U8985 (N_8985,N_4816,N_5829);
xnor U8986 (N_8986,N_4782,N_5327);
nand U8987 (N_8987,N_3196,N_5500);
nor U8988 (N_8988,N_3556,N_4653);
or U8989 (N_8989,N_3880,N_3132);
and U8990 (N_8990,N_4214,N_5137);
nand U8991 (N_8991,N_5209,N_5376);
xor U8992 (N_8992,N_4620,N_4095);
or U8993 (N_8993,N_5409,N_4244);
or U8994 (N_8994,N_5601,N_4142);
nand U8995 (N_8995,N_3328,N_5233);
and U8996 (N_8996,N_3274,N_3122);
or U8997 (N_8997,N_3384,N_5908);
nor U8998 (N_8998,N_3541,N_5930);
nor U8999 (N_8999,N_4605,N_4643);
or U9000 (N_9000,N_6733,N_8612);
nand U9001 (N_9001,N_6946,N_8472);
or U9002 (N_9002,N_7414,N_8462);
xor U9003 (N_9003,N_8961,N_6283);
and U9004 (N_9004,N_8769,N_7224);
nor U9005 (N_9005,N_7928,N_7062);
nand U9006 (N_9006,N_8082,N_8992);
xnor U9007 (N_9007,N_7831,N_8118);
and U9008 (N_9008,N_6561,N_8302);
nor U9009 (N_9009,N_7233,N_6851);
or U9010 (N_9010,N_6228,N_8407);
xnor U9011 (N_9011,N_7871,N_8734);
nand U9012 (N_9012,N_7097,N_8062);
xnor U9013 (N_9013,N_8964,N_8994);
and U9014 (N_9014,N_7323,N_8575);
nand U9015 (N_9015,N_8367,N_7113);
nand U9016 (N_9016,N_8516,N_6813);
or U9017 (N_9017,N_6142,N_8751);
xnor U9018 (N_9018,N_7412,N_8726);
and U9019 (N_9019,N_8607,N_7713);
or U9020 (N_9020,N_7168,N_6651);
and U9021 (N_9021,N_8598,N_6490);
or U9022 (N_9022,N_7760,N_6601);
xor U9023 (N_9023,N_6973,N_6747);
nor U9024 (N_9024,N_6670,N_7196);
or U9025 (N_9025,N_7806,N_8117);
nor U9026 (N_9026,N_8145,N_7725);
or U9027 (N_9027,N_8599,N_7158);
and U9028 (N_9028,N_6237,N_8323);
or U9029 (N_9029,N_6047,N_7704);
nor U9030 (N_9030,N_8121,N_6684);
or U9031 (N_9031,N_8949,N_7161);
xnor U9032 (N_9032,N_8907,N_6693);
or U9033 (N_9033,N_7345,N_6333);
nor U9034 (N_9034,N_8996,N_7883);
nor U9035 (N_9035,N_6661,N_8287);
nor U9036 (N_9036,N_7121,N_7467);
nor U9037 (N_9037,N_6307,N_6203);
nand U9038 (N_9038,N_6274,N_8748);
nand U9039 (N_9039,N_6359,N_6809);
or U9040 (N_9040,N_7696,N_6939);
or U9041 (N_9041,N_6550,N_8700);
or U9042 (N_9042,N_8661,N_7302);
nand U9043 (N_9043,N_7108,N_7423);
xor U9044 (N_9044,N_8356,N_7321);
or U9045 (N_9045,N_7261,N_8016);
nand U9046 (N_9046,N_8552,N_8417);
nor U9047 (N_9047,N_6450,N_6887);
nand U9048 (N_9048,N_7024,N_7583);
and U9049 (N_9049,N_8034,N_6064);
and U9050 (N_9050,N_8923,N_7661);
nand U9051 (N_9051,N_7201,N_7951);
nand U9052 (N_9052,N_6463,N_6816);
xnor U9053 (N_9053,N_8251,N_6572);
nor U9054 (N_9054,N_7660,N_8317);
and U9055 (N_9055,N_7053,N_8878);
and U9056 (N_9056,N_6111,N_8547);
nand U9057 (N_9057,N_6563,N_6583);
and U9058 (N_9058,N_7734,N_6381);
nor U9059 (N_9059,N_7172,N_8132);
or U9060 (N_9060,N_6270,N_8150);
and U9061 (N_9061,N_7350,N_6850);
and U9062 (N_9062,N_8384,N_6522);
and U9063 (N_9063,N_7156,N_6830);
xor U9064 (N_9064,N_6368,N_7629);
xor U9065 (N_9065,N_6995,N_7563);
xnor U9066 (N_9066,N_6054,N_8203);
nand U9067 (N_9067,N_7356,N_7052);
nand U9068 (N_9068,N_6180,N_7538);
xnor U9069 (N_9069,N_8095,N_8777);
nor U9070 (N_9070,N_6714,N_6039);
xor U9071 (N_9071,N_6652,N_7343);
or U9072 (N_9072,N_8479,N_7422);
and U9073 (N_9073,N_7564,N_7372);
and U9074 (N_9074,N_8913,N_8678);
nor U9075 (N_9075,N_8187,N_6502);
nand U9076 (N_9076,N_8020,N_8890);
or U9077 (N_9077,N_7145,N_7726);
and U9078 (N_9078,N_8089,N_6048);
nand U9079 (N_9079,N_6428,N_8693);
nor U9080 (N_9080,N_8432,N_6750);
xnor U9081 (N_9081,N_8279,N_6390);
xnor U9082 (N_9082,N_8378,N_6051);
nand U9083 (N_9083,N_7642,N_6314);
nor U9084 (N_9084,N_6781,N_6343);
or U9085 (N_9085,N_7243,N_6771);
or U9086 (N_9086,N_8563,N_7665);
xor U9087 (N_9087,N_6788,N_8894);
nand U9088 (N_9088,N_7087,N_6501);
xor U9089 (N_9089,N_8393,N_6569);
nand U9090 (N_9090,N_7293,N_7600);
xor U9091 (N_9091,N_7494,N_6627);
or U9092 (N_9092,N_8053,N_7995);
and U9093 (N_9093,N_7747,N_8795);
nor U9094 (N_9094,N_7718,N_6593);
xnor U9095 (N_9095,N_6863,N_7681);
nand U9096 (N_9096,N_7502,N_6199);
or U9097 (N_9097,N_8239,N_8242);
nor U9098 (N_9098,N_8540,N_7046);
nor U9099 (N_9099,N_7832,N_7673);
and U9100 (N_9100,N_6742,N_7917);
and U9101 (N_9101,N_7477,N_7756);
nor U9102 (N_9102,N_6188,N_7662);
and U9103 (N_9103,N_8589,N_6053);
or U9104 (N_9104,N_6177,N_7728);
xor U9105 (N_9105,N_8667,N_7389);
nor U9106 (N_9106,N_7214,N_6003);
or U9107 (N_9107,N_6857,N_8762);
nor U9108 (N_9108,N_7096,N_6056);
or U9109 (N_9109,N_8106,N_8899);
or U9110 (N_9110,N_6751,N_7391);
nor U9111 (N_9111,N_7587,N_8206);
nand U9112 (N_9112,N_8229,N_7171);
nor U9113 (N_9113,N_8997,N_8880);
or U9114 (N_9114,N_6447,N_7887);
nand U9115 (N_9115,N_6535,N_6908);
and U9116 (N_9116,N_6746,N_6941);
or U9117 (N_9117,N_7899,N_8136);
and U9118 (N_9118,N_8647,N_7792);
or U9119 (N_9119,N_7915,N_8860);
nand U9120 (N_9120,N_6193,N_8993);
nand U9121 (N_9121,N_6358,N_7855);
xnor U9122 (N_9122,N_7004,N_8398);
nor U9123 (N_9123,N_6831,N_6139);
and U9124 (N_9124,N_6155,N_7309);
xor U9125 (N_9125,N_6372,N_6801);
and U9126 (N_9126,N_7842,N_8405);
nor U9127 (N_9127,N_8837,N_8070);
nand U9128 (N_9128,N_8278,N_7187);
nand U9129 (N_9129,N_6235,N_8525);
and U9130 (N_9130,N_8389,N_8138);
nor U9131 (N_9131,N_6564,N_7548);
xor U9132 (N_9132,N_8725,N_8652);
nand U9133 (N_9133,N_6391,N_6726);
and U9134 (N_9134,N_7940,N_7688);
and U9135 (N_9135,N_8243,N_7257);
nor U9136 (N_9136,N_7297,N_6917);
and U9137 (N_9137,N_8987,N_6800);
nand U9138 (N_9138,N_6758,N_7900);
nor U9139 (N_9139,N_6578,N_6660);
and U9140 (N_9140,N_8654,N_7455);
xor U9141 (N_9141,N_6271,N_8827);
and U9142 (N_9142,N_7997,N_7485);
or U9143 (N_9143,N_7955,N_6414);
nand U9144 (N_9144,N_7542,N_8212);
and U9145 (N_9145,N_8934,N_6434);
nand U9146 (N_9146,N_6062,N_6439);
or U9147 (N_9147,N_7784,N_7326);
xnor U9148 (N_9148,N_7875,N_7432);
or U9149 (N_9149,N_6192,N_6632);
xnor U9150 (N_9150,N_6157,N_8511);
nor U9151 (N_9151,N_7579,N_8971);
and U9152 (N_9152,N_6256,N_7212);
and U9153 (N_9153,N_8705,N_7625);
nand U9154 (N_9154,N_6443,N_6398);
xnor U9155 (N_9155,N_7802,N_8608);
and U9156 (N_9156,N_8901,N_7801);
nor U9157 (N_9157,N_6138,N_7393);
and U9158 (N_9158,N_6663,N_7264);
or U9159 (N_9159,N_8979,N_6201);
nor U9160 (N_9160,N_7607,N_6027);
or U9161 (N_9161,N_8784,N_8530);
or U9162 (N_9162,N_6979,N_7516);
nand U9163 (N_9163,N_7762,N_6957);
nand U9164 (N_9164,N_7410,N_6770);
nor U9165 (N_9165,N_7666,N_6913);
or U9166 (N_9166,N_8597,N_6776);
and U9167 (N_9167,N_8768,N_7394);
and U9168 (N_9168,N_6392,N_6609);
nor U9169 (N_9169,N_8090,N_8675);
nor U9170 (N_9170,N_6621,N_7973);
or U9171 (N_9171,N_8110,N_8583);
xnor U9172 (N_9172,N_7618,N_6150);
nor U9173 (N_9173,N_6253,N_8859);
nand U9174 (N_9174,N_7653,N_8969);
and U9175 (N_9175,N_6864,N_7054);
xor U9176 (N_9176,N_8353,N_6233);
or U9177 (N_9177,N_8260,N_8303);
and U9178 (N_9178,N_7633,N_7898);
and U9179 (N_9179,N_7225,N_6956);
xnor U9180 (N_9180,N_7813,N_7631);
nor U9181 (N_9181,N_6264,N_8368);
and U9182 (N_9182,N_6539,N_8579);
nand U9183 (N_9183,N_6037,N_8096);
nor U9184 (N_9184,N_6260,N_8346);
and U9185 (N_9185,N_7700,N_7519);
xor U9186 (N_9186,N_8263,N_7687);
xnor U9187 (N_9187,N_8402,N_8126);
or U9188 (N_9188,N_7064,N_7032);
and U9189 (N_9189,N_7836,N_8708);
nand U9190 (N_9190,N_8764,N_7169);
or U9191 (N_9191,N_8253,N_7619);
xor U9192 (N_9192,N_8486,N_8600);
or U9193 (N_9193,N_8871,N_7329);
nor U9194 (N_9194,N_8195,N_6635);
nand U9195 (N_9195,N_6006,N_8141);
xor U9196 (N_9196,N_8103,N_6702);
xor U9197 (N_9197,N_6504,N_8876);
nand U9198 (N_9198,N_6616,N_6907);
or U9199 (N_9199,N_6473,N_8753);
or U9200 (N_9200,N_7162,N_8033);
or U9201 (N_9201,N_7180,N_8325);
and U9202 (N_9202,N_6029,N_6404);
xor U9203 (N_9203,N_7082,N_6206);
nor U9204 (N_9204,N_7884,N_8989);
or U9205 (N_9205,N_6239,N_6774);
and U9206 (N_9206,N_8856,N_8201);
nand U9207 (N_9207,N_6780,N_8478);
and U9208 (N_9208,N_8666,N_7199);
and U9209 (N_9209,N_8444,N_8151);
xnor U9210 (N_9210,N_7528,N_7349);
xnor U9211 (N_9211,N_6495,N_6075);
nor U9212 (N_9212,N_8464,N_8018);
nor U9213 (N_9213,N_8925,N_8177);
and U9214 (N_9214,N_7965,N_6181);
or U9215 (N_9215,N_7308,N_6148);
nand U9216 (N_9216,N_7002,N_7868);
xor U9217 (N_9217,N_7818,N_7193);
nor U9218 (N_9218,N_6292,N_8165);
nand U9219 (N_9219,N_8382,N_8646);
nand U9220 (N_9220,N_7525,N_7550);
and U9221 (N_9221,N_6184,N_7846);
nand U9222 (N_9222,N_8208,N_6007);
nor U9223 (N_9223,N_8483,N_8637);
or U9224 (N_9224,N_7263,N_7289);
nand U9225 (N_9225,N_8749,N_8928);
nand U9226 (N_9226,N_7649,N_7545);
nor U9227 (N_9227,N_7654,N_6527);
or U9228 (N_9228,N_6306,N_7421);
xor U9229 (N_9229,N_6113,N_8143);
or U9230 (N_9230,N_7408,N_8746);
xor U9231 (N_9231,N_7879,N_7111);
xor U9232 (N_9232,N_6920,N_6068);
nor U9233 (N_9233,N_8766,N_8869);
and U9234 (N_9234,N_8079,N_6044);
or U9235 (N_9235,N_6089,N_7668);
and U9236 (N_9236,N_8670,N_6735);
or U9237 (N_9237,N_7292,N_6402);
and U9238 (N_9238,N_7512,N_8805);
and U9239 (N_9239,N_6134,N_7778);
and U9240 (N_9240,N_8972,N_6244);
and U9241 (N_9241,N_8192,N_7042);
nand U9242 (N_9242,N_8350,N_7626);
xnor U9243 (N_9243,N_7106,N_6592);
or U9244 (N_9244,N_8945,N_6509);
nor U9245 (N_9245,N_6168,N_8280);
and U9246 (N_9246,N_6553,N_7300);
xor U9247 (N_9247,N_8509,N_6005);
and U9248 (N_9248,N_8456,N_7347);
xor U9249 (N_9249,N_8175,N_7979);
nand U9250 (N_9250,N_8737,N_8801);
or U9251 (N_9251,N_6794,N_7585);
nor U9252 (N_9252,N_8178,N_7067);
nor U9253 (N_9253,N_7615,N_7014);
or U9254 (N_9254,N_8198,N_8065);
nand U9255 (N_9255,N_7999,N_6699);
nor U9256 (N_9256,N_7849,N_8386);
nor U9257 (N_9257,N_7694,N_8204);
nor U9258 (N_9258,N_7524,N_8852);
nand U9259 (N_9259,N_7731,N_7645);
nand U9260 (N_9260,N_6485,N_7796);
or U9261 (N_9261,N_7902,N_7234);
and U9262 (N_9262,N_8290,N_7707);
and U9263 (N_9263,N_8450,N_6654);
nand U9264 (N_9264,N_6667,N_8381);
nor U9265 (N_9265,N_8691,N_8824);
or U9266 (N_9266,N_6665,N_6812);
xnor U9267 (N_9267,N_6369,N_6845);
nor U9268 (N_9268,N_6680,N_7730);
nand U9269 (N_9269,N_6551,N_8793);
nand U9270 (N_9270,N_6508,N_7904);
nor U9271 (N_9271,N_8301,N_7367);
xnor U9272 (N_9272,N_6933,N_8221);
or U9273 (N_9273,N_6940,N_8735);
nand U9274 (N_9274,N_6634,N_6230);
and U9275 (N_9275,N_8093,N_7606);
nand U9276 (N_9276,N_7251,N_8501);
nor U9277 (N_9277,N_7683,N_8976);
xor U9278 (N_9278,N_6859,N_8534);
xnor U9279 (N_9279,N_7094,N_7692);
xor U9280 (N_9280,N_7711,N_8505);
and U9281 (N_9281,N_7213,N_7110);
and U9282 (N_9282,N_7338,N_8409);
and U9283 (N_9283,N_7019,N_6300);
or U9284 (N_9284,N_6642,N_8754);
or U9285 (N_9285,N_6376,N_7434);
nand U9286 (N_9286,N_6886,N_8051);
nor U9287 (N_9287,N_6722,N_6612);
nand U9288 (N_9288,N_7510,N_6420);
nor U9289 (N_9289,N_8767,N_6034);
xor U9290 (N_9290,N_6133,N_7775);
nand U9291 (N_9291,N_6412,N_6308);
and U9292 (N_9292,N_7107,N_7152);
nand U9293 (N_9293,N_7958,N_6810);
or U9294 (N_9294,N_6069,N_7670);
xor U9295 (N_9295,N_8621,N_8397);
xnor U9296 (N_9296,N_6879,N_8538);
or U9297 (N_9297,N_7444,N_6968);
nand U9298 (N_9298,N_8508,N_7648);
nand U9299 (N_9299,N_7624,N_7745);
nor U9300 (N_9300,N_7878,N_7268);
nand U9301 (N_9301,N_6744,N_6768);
xnor U9302 (N_9302,N_7889,N_7613);
xor U9303 (N_9303,N_7920,N_6442);
nor U9304 (N_9304,N_7943,N_8731);
xnor U9305 (N_9305,N_7777,N_8673);
and U9306 (N_9306,N_7266,N_6513);
or U9307 (N_9307,N_8650,N_7829);
and U9308 (N_9308,N_8888,N_8980);
xor U9309 (N_9309,N_8237,N_6936);
nor U9310 (N_9310,N_7810,N_7558);
or U9311 (N_9311,N_7119,N_6440);
and U9312 (N_9312,N_8312,N_7208);
nand U9313 (N_9313,N_8938,N_7129);
nand U9314 (N_9314,N_7771,N_8028);
xnor U9315 (N_9315,N_6025,N_8196);
xor U9316 (N_9316,N_7581,N_8788);
or U9317 (N_9317,N_7870,N_6147);
or U9318 (N_9318,N_7667,N_6524);
nor U9319 (N_9319,N_7727,N_6659);
or U9320 (N_9320,N_6738,N_6694);
xnor U9321 (N_9321,N_6273,N_6072);
xnor U9322 (N_9322,N_6295,N_8335);
nor U9323 (N_9323,N_6938,N_8797);
and U9324 (N_9324,N_8539,N_6488);
nor U9325 (N_9325,N_7809,N_8811);
nor U9326 (N_9326,N_6585,N_8222);
xor U9327 (N_9327,N_7690,N_6017);
or U9328 (N_9328,N_7919,N_7739);
or U9329 (N_9329,N_7102,N_6163);
nor U9330 (N_9330,N_8180,N_7176);
xnor U9331 (N_9331,N_6900,N_7114);
or U9332 (N_9332,N_8403,N_8513);
nor U9333 (N_9333,N_6437,N_8703);
nor U9334 (N_9334,N_6481,N_8931);
or U9335 (N_9335,N_7737,N_7761);
or U9336 (N_9336,N_8413,N_7010);
and U9337 (N_9337,N_7281,N_6586);
nand U9338 (N_9338,N_7228,N_7783);
or U9339 (N_9339,N_6647,N_7449);
and U9340 (N_9340,N_7975,N_7886);
nand U9341 (N_9341,N_7142,N_8102);
nor U9342 (N_9342,N_8850,N_6266);
and U9343 (N_9343,N_7573,N_7250);
or U9344 (N_9344,N_8952,N_6397);
nor U9345 (N_9345,N_8401,N_7722);
and U9346 (N_9346,N_6178,N_6753);
and U9347 (N_9347,N_7079,N_8744);
or U9348 (N_9348,N_6807,N_6000);
or U9349 (N_9349,N_8581,N_7947);
nor U9350 (N_9350,N_6249,N_8819);
or U9351 (N_9351,N_6918,N_6221);
xor U9352 (N_9352,N_6602,N_7369);
and U9353 (N_9353,N_7523,N_6453);
nand U9354 (N_9354,N_8254,N_6227);
nand U9355 (N_9355,N_8499,N_6669);
xor U9356 (N_9356,N_8215,N_6759);
nor U9357 (N_9357,N_7776,N_7075);
xor U9358 (N_9358,N_6389,N_8156);
or U9359 (N_9359,N_8271,N_6196);
nor U9360 (N_9360,N_8715,N_8814);
nand U9361 (N_9361,N_7273,N_7479);
xor U9362 (N_9362,N_8828,N_8921);
nor U9363 (N_9363,N_6015,N_6004);
nor U9364 (N_9364,N_7593,N_7377);
and U9365 (N_9365,N_6324,N_6873);
xor U9366 (N_9366,N_8101,N_6289);
or U9367 (N_9367,N_8171,N_6937);
nor U9368 (N_9368,N_7639,N_6534);
and U9369 (N_9369,N_7003,N_8959);
or U9370 (N_9370,N_8585,N_8718);
and U9371 (N_9371,N_7560,N_7604);
xnor U9372 (N_9372,N_7252,N_7521);
nor U9373 (N_9373,N_7402,N_7427);
nor U9374 (N_9374,N_7513,N_8474);
and U9375 (N_9375,N_8269,N_8849);
nor U9376 (N_9376,N_6761,N_6330);
nor U9377 (N_9377,N_6243,N_7353);
nand U9378 (N_9378,N_6876,N_7463);
and U9379 (N_9379,N_7209,N_6896);
xnor U9380 (N_9380,N_7008,N_7395);
nor U9381 (N_9381,N_7993,N_7277);
nand U9382 (N_9382,N_6791,N_6158);
xnor U9383 (N_9383,N_6286,N_7183);
nand U9384 (N_9384,N_7246,N_6408);
nor U9385 (N_9385,N_6421,N_7122);
xnor U9386 (N_9386,N_7500,N_7013);
or U9387 (N_9387,N_6285,N_7317);
nand U9388 (N_9388,N_7984,N_6950);
nand U9389 (N_9389,N_7921,N_6949);
or U9390 (N_9390,N_6341,N_8041);
and U9391 (N_9391,N_8365,N_6600);
nand U9392 (N_9392,N_8742,N_7627);
xnor U9393 (N_9393,N_6154,N_8297);
and U9394 (N_9394,N_7443,N_7016);
and U9395 (N_9395,N_8832,N_8477);
or U9396 (N_9396,N_8685,N_8895);
or U9397 (N_9397,N_8634,N_8296);
nand U9398 (N_9398,N_8798,N_8022);
nand U9399 (N_9399,N_7532,N_8304);
xnor U9400 (N_9400,N_7074,N_8231);
or U9401 (N_9401,N_7888,N_8146);
or U9402 (N_9402,N_6028,N_8546);
xnor U9403 (N_9403,N_7753,N_8991);
xnor U9404 (N_9404,N_6380,N_6451);
or U9405 (N_9405,N_7167,N_7229);
and U9406 (N_9406,N_6644,N_7344);
nand U9407 (N_9407,N_7651,N_6340);
nand U9408 (N_9408,N_7354,N_8185);
xnor U9409 (N_9409,N_8241,N_7848);
or U9410 (N_9410,N_8990,N_7379);
and U9411 (N_9411,N_7045,N_6388);
xor U9412 (N_9412,N_7346,N_6518);
nor U9413 (N_9413,N_6162,N_6444);
or U9414 (N_9414,N_7569,N_8752);
and U9415 (N_9415,N_7636,N_8283);
nor U9416 (N_9416,N_7695,N_7570);
nand U9417 (N_9417,N_8882,N_8506);
xnor U9418 (N_9418,N_8439,N_8435);
xor U9419 (N_9419,N_7612,N_8536);
nor U9420 (N_9420,N_8580,N_6383);
nor U9421 (N_9421,N_8821,N_7816);
xor U9422 (N_9422,N_6290,N_8848);
or U9423 (N_9423,N_6337,N_6231);
nand U9424 (N_9424,N_7088,N_6410);
or U9425 (N_9425,N_8707,N_6349);
and U9426 (N_9426,N_6756,N_8702);
xnor U9427 (N_9427,N_6570,N_6784);
and U9428 (N_9428,N_7361,N_8037);
and U9429 (N_9429,N_6861,N_7307);
xor U9430 (N_9430,N_8298,N_8168);
or U9431 (N_9431,N_6361,N_6709);
xor U9432 (N_9432,N_8069,N_6910);
or U9433 (N_9433,N_8729,N_8080);
xnor U9434 (N_9434,N_8388,N_6697);
xnor U9435 (N_9435,N_6474,N_6821);
or U9436 (N_9436,N_6705,N_6893);
nor U9437 (N_9437,N_6581,N_8940);
nand U9438 (N_9438,N_7961,N_6707);
or U9439 (N_9439,N_6066,N_7862);
nand U9440 (N_9440,N_8174,N_6107);
nor U9441 (N_9441,N_6675,N_6731);
nand U9442 (N_9442,N_6890,N_7603);
and U9443 (N_9443,N_8706,N_6186);
nand U9444 (N_9444,N_7769,N_6772);
xor U9445 (N_9445,N_7314,N_8182);
or U9446 (N_9446,N_7034,N_7048);
or U9447 (N_9447,N_7078,N_6038);
nand U9448 (N_9448,N_6467,N_6208);
nor U9449 (N_9449,N_7520,N_6603);
nand U9450 (N_9450,N_7280,N_7589);
xnor U9451 (N_9451,N_6220,N_8105);
nor U9452 (N_9452,N_6441,N_6422);
nor U9453 (N_9453,N_7478,N_6288);
xnor U9454 (N_9454,N_8152,N_7702);
xor U9455 (N_9455,N_7123,N_6310);
or U9456 (N_9456,N_8234,N_7499);
xor U9457 (N_9457,N_7766,N_8591);
nor U9458 (N_9458,N_7441,N_6123);
nor U9459 (N_9459,N_6322,N_6523);
nand U9460 (N_9460,N_7466,N_8502);
and U9461 (N_9461,N_6649,N_8326);
and U9462 (N_9462,N_8383,N_8434);
nand U9463 (N_9463,N_6338,N_8316);
xnor U9464 (N_9464,N_8111,N_8363);
and U9465 (N_9465,N_7927,N_7908);
xnor U9466 (N_9466,N_8039,N_8288);
xor U9467 (N_9467,N_7650,N_6921);
nand U9468 (N_9468,N_6137,N_6385);
nand U9469 (N_9469,N_8379,N_6429);
xor U9470 (N_9470,N_8445,N_6826);
nor U9471 (N_9471,N_6386,N_6091);
xnor U9472 (N_9472,N_8676,N_8906);
xor U9473 (N_9473,N_7039,N_6131);
or U9474 (N_9474,N_8484,N_8864);
nand U9475 (N_9475,N_8497,N_7789);
or U9476 (N_9476,N_6083,N_6655);
nor U9477 (N_9477,N_6245,N_8338);
nand U9478 (N_9478,N_8252,N_7911);
and U9479 (N_9479,N_6374,N_7677);
nand U9480 (N_9480,N_8681,N_7556);
and U9481 (N_9481,N_8305,N_7946);
nor U9482 (N_9482,N_7155,N_7216);
or U9483 (N_9483,N_8515,N_8528);
nand U9484 (N_9484,N_7204,N_8962);
nor U9485 (N_9485,N_7741,N_8314);
and U9486 (N_9486,N_8319,N_8336);
nand U9487 (N_9487,N_7638,N_7752);
nand U9488 (N_9488,N_7854,N_6172);
and U9489 (N_9489,N_7241,N_6345);
and U9490 (N_9490,N_6842,N_7203);
xor U9491 (N_9491,N_8815,N_7207);
and U9492 (N_9492,N_7254,N_6713);
nand U9493 (N_9493,N_7348,N_6323);
nor U9494 (N_9494,N_7924,N_6505);
or U9495 (N_9495,N_6828,N_6118);
or U9496 (N_9496,N_7419,N_7006);
or U9497 (N_9497,N_6448,N_6078);
or U9498 (N_9498,N_6418,N_6868);
nand U9499 (N_9499,N_8163,N_6318);
xor U9500 (N_9500,N_6461,N_8765);
xnor U9501 (N_9501,N_6811,N_6363);
nand U9502 (N_9502,N_7127,N_8123);
xor U9503 (N_9503,N_7844,N_8449);
and U9504 (N_9504,N_8559,N_7227);
or U9505 (N_9505,N_6901,N_7033);
xnor U9506 (N_9506,N_6765,N_8331);
xnor U9507 (N_9507,N_6943,N_8442);
nor U9508 (N_9508,N_8113,N_7577);
or U9509 (N_9509,N_7023,N_8340);
or U9510 (N_9510,N_6460,N_7630);
nand U9511 (N_9511,N_8355,N_6269);
nand U9512 (N_9512,N_6378,N_7529);
and U9513 (N_9513,N_7489,N_7027);
and U9514 (N_9514,N_6964,N_7426);
nand U9515 (N_9515,N_8507,N_6135);
and U9516 (N_9516,N_7452,N_8321);
and U9517 (N_9517,N_8602,N_6413);
and U9518 (N_9518,N_8043,N_8429);
nor U9519 (N_9519,N_7882,N_8745);
nand U9520 (N_9520,N_8264,N_8722);
or U9521 (N_9521,N_8176,N_7117);
xor U9522 (N_9522,N_6605,N_6970);
and U9523 (N_9523,N_8937,N_8838);
or U9524 (N_9524,N_8709,N_6074);
nor U9525 (N_9525,N_7566,N_6202);
xnor U9526 (N_9526,N_8169,N_7235);
nand U9527 (N_9527,N_6835,N_7793);
or U9528 (N_9528,N_8818,N_7336);
nand U9529 (N_9529,N_7405,N_7276);
xnor U9530 (N_9530,N_8481,N_8569);
and U9531 (N_9531,N_7460,N_8724);
and U9532 (N_9532,N_7283,N_6112);
xnor U9533 (N_9533,N_6588,N_6959);
or U9534 (N_9534,N_6140,N_8306);
or U9535 (N_9535,N_7351,N_6519);
nor U9536 (N_9536,N_6631,N_7853);
and U9537 (N_9537,N_6980,N_8473);
nand U9538 (N_9538,N_8930,N_7530);
nor U9539 (N_9539,N_6255,N_7001);
xnor U9540 (N_9540,N_7290,N_7931);
xor U9541 (N_9541,N_6119,N_7893);
and U9542 (N_9542,N_7397,N_8299);
xnor U9543 (N_9543,N_8698,N_6001);
nor U9544 (N_9544,N_6483,N_6435);
nand U9545 (N_9545,N_8226,N_7480);
xor U9546 (N_9546,N_8714,N_6127);
nand U9547 (N_9547,N_6217,N_8307);
and U9548 (N_9548,N_6197,N_8912);
and U9549 (N_9549,N_6617,N_7749);
xor U9550 (N_9550,N_7782,N_7781);
nor U9551 (N_9551,N_8328,N_8390);
xnor U9552 (N_9552,N_6677,N_7120);
and U9553 (N_9553,N_8119,N_7856);
nand U9554 (N_9554,N_6057,N_8233);
and U9555 (N_9555,N_8266,N_8656);
or U9556 (N_9556,N_6546,N_7964);
xnor U9557 (N_9557,N_8716,N_7706);
nand U9558 (N_9558,N_8071,N_8300);
nor U9559 (N_9559,N_8200,N_6817);
or U9560 (N_9560,N_7905,N_8642);
nand U9561 (N_9561,N_6101,N_7980);
or U9562 (N_9562,N_6303,N_7959);
xor U9563 (N_9563,N_6082,N_6613);
xor U9564 (N_9564,N_7584,N_8343);
nand U9565 (N_9565,N_6824,N_8427);
nor U9566 (N_9566,N_8900,N_7837);
xor U9567 (N_9567,N_7680,N_6486);
or U9568 (N_9568,N_7318,N_8437);
xnor U9569 (N_9569,N_7051,N_8274);
or U9570 (N_9570,N_7486,N_6880);
nor U9571 (N_9571,N_7599,N_8448);
nand U9572 (N_9572,N_6580,N_8669);
nand U9573 (N_9573,N_6061,N_8626);
or U9574 (N_9574,N_8172,N_6844);
nor U9575 (N_9575,N_6382,N_6106);
and U9576 (N_9576,N_7179,N_8216);
or U9577 (N_9577,N_8935,N_7515);
nand U9578 (N_9578,N_8561,N_6790);
nor U9579 (N_9579,N_8728,N_8825);
nor U9580 (N_9580,N_8672,N_7953);
or U9581 (N_9581,N_7440,N_6167);
or U9582 (N_9582,N_6419,N_6405);
and U9583 (N_9583,N_6478,N_8470);
nor U9584 (N_9584,N_7025,N_8362);
or U9585 (N_9585,N_7798,N_8339);
xor U9586 (N_9586,N_8738,N_8076);
or U9587 (N_9587,N_7143,N_8806);
or U9588 (N_9588,N_8419,N_8066);
xnor U9589 (N_9589,N_8526,N_7366);
nor U9590 (N_9590,N_7664,N_6806);
and U9591 (N_9591,N_7989,N_8808);
and U9592 (N_9592,N_6222,N_6843);
nor U9593 (N_9593,N_8002,N_7238);
and U9594 (N_9594,N_8618,N_6117);
nor U9595 (N_9595,N_8845,N_8686);
nand U9596 (N_9596,N_6805,N_7833);
xnor U9597 (N_9597,N_7828,N_8866);
and U9598 (N_9598,N_7190,N_7977);
nor U9599 (N_9599,N_8813,N_8455);
and U9600 (N_9600,N_7269,N_7331);
and U9601 (N_9601,N_6792,N_6657);
xnor U9602 (N_9602,N_7963,N_6803);
nand U9603 (N_9603,N_7549,N_8730);
and U9604 (N_9604,N_8835,N_8988);
xor U9605 (N_9605,N_8587,N_6628);
or U9606 (N_9606,N_7719,N_7622);
nand U9607 (N_9607,N_8857,N_7948);
or U9608 (N_9608,N_7253,N_8190);
nor U9609 (N_9609,N_6297,N_6326);
and U9610 (N_9610,N_6454,N_8466);
xor U9611 (N_9611,N_6436,N_6275);
and U9612 (N_9612,N_7086,N_6302);
or U9613 (N_9613,N_6898,N_8829);
nor U9614 (N_9614,N_8574,N_7493);
nor U9615 (N_9615,N_7077,N_6575);
and U9616 (N_9616,N_6915,N_8914);
or U9617 (N_9617,N_8493,N_8567);
nand U9618 (N_9618,N_8732,N_6576);
nand U9619 (N_9619,N_7018,N_7823);
nand U9620 (N_9620,N_8476,N_7655);
nor U9621 (N_9621,N_6475,N_7970);
nand U9622 (N_9622,N_7557,N_7357);
or U9623 (N_9623,N_6798,N_6019);
nand U9624 (N_9624,N_7750,N_7551);
nand U9625 (N_9625,N_6591,N_7141);
and U9626 (N_9626,N_7211,N_8446);
xor U9627 (N_9627,N_7194,N_8088);
and U9628 (N_9628,N_7457,N_6105);
xnor U9629 (N_9629,N_7996,N_7721);
and U9630 (N_9630,N_7978,N_6988);
xor U9631 (N_9631,N_6594,N_7804);
or U9632 (N_9632,N_7249,N_7101);
and U9633 (N_9633,N_8556,N_6717);
nand U9634 (N_9634,N_7501,N_6254);
xnor U9635 (N_9635,N_8351,N_6611);
nor U9636 (N_9636,N_8711,N_7388);
nand U9637 (N_9637,N_6216,N_6406);
xnor U9638 (N_9638,N_8024,N_7890);
or U9639 (N_9639,N_7215,N_6493);
or U9640 (N_9640,N_6741,N_8202);
and U9641 (N_9641,N_6179,N_7578);
xnor U9642 (N_9642,N_6793,N_8130);
and U9643 (N_9643,N_7104,N_7260);
or U9644 (N_9644,N_6639,N_8144);
nand U9645 (N_9645,N_8684,N_6926);
or U9646 (N_9646,N_6689,N_6084);
xnor U9647 (N_9647,N_8903,N_6251);
nand U9648 (N_9648,N_8469,N_7689);
xnor U9649 (N_9649,N_6268,N_6415);
and U9650 (N_9650,N_6598,N_6279);
xnor U9651 (N_9651,N_6558,N_6121);
and U9652 (N_9652,N_6232,N_8440);
or U9653 (N_9653,N_7819,N_8853);
xor U9654 (N_9654,N_8048,N_6566);
and U9655 (N_9655,N_6482,N_7710);
nor U9656 (N_9656,N_8776,N_6909);
nand U9657 (N_9657,N_6520,N_7795);
nand U9658 (N_9658,N_8104,N_8782);
nor U9659 (N_9659,N_7223,N_7424);
or U9660 (N_9660,N_7658,N_6449);
nand U9661 (N_9661,N_6262,N_8697);
and U9662 (N_9662,N_6965,N_7863);
xor U9663 (N_9663,N_8046,N_6721);
nor U9664 (N_9664,N_6205,N_8527);
or U9665 (N_9665,N_8858,N_6969);
nor U9666 (N_9666,N_7055,N_7697);
nand U9667 (N_9667,N_8733,N_6394);
xor U9668 (N_9668,N_8713,N_8453);
and U9669 (N_9669,N_8131,N_6225);
nand U9670 (N_9670,N_6762,N_7780);
xnor U9671 (N_9671,N_8761,N_6783);
and U9672 (N_9672,N_8503,N_8757);
and U9673 (N_9673,N_7592,N_6510);
or U9674 (N_9674,N_8087,N_7450);
nand U9675 (N_9675,N_6532,N_8865);
and U9676 (N_9676,N_7267,N_7678);
xor U9677 (N_9677,N_8426,N_6452);
xor U9678 (N_9678,N_7272,N_6189);
or U9679 (N_9679,N_6755,N_7872);
nand U9680 (N_9680,N_7284,N_7417);
nor U9681 (N_9681,N_8885,N_6008);
and U9682 (N_9682,N_6736,N_6097);
and U9683 (N_9683,N_8512,N_8488);
or U9684 (N_9684,N_7845,N_6769);
and U9685 (N_9685,N_7305,N_8061);
or U9686 (N_9686,N_8613,N_8490);
or U9687 (N_9687,N_6894,N_8884);
xnor U9688 (N_9688,N_8327,N_6610);
or U9689 (N_9689,N_8167,N_6766);
nand U9690 (N_9690,N_8915,N_8441);
or U9691 (N_9691,N_6676,N_6931);
xor U9692 (N_9692,N_8586,N_6209);
xnor U9693 (N_9693,N_6777,N_7239);
nor U9694 (N_9694,N_6854,N_8594);
and U9695 (N_9695,N_8982,N_8292);
xor U9696 (N_9696,N_6280,N_7376);
and U9697 (N_9697,N_8369,N_7504);
nand U9698 (N_9698,N_7746,N_7825);
and U9699 (N_9699,N_8674,N_7288);
nand U9700 (N_9700,N_8614,N_7939);
xnor U9701 (N_9701,N_8542,N_7400);
or U9702 (N_9702,N_8376,N_8960);
nor U9703 (N_9703,N_7543,N_6212);
and U9704 (N_9704,N_6737,N_7647);
and U9705 (N_9705,N_8875,N_6869);
nor U9706 (N_9706,N_8116,N_8219);
xnor U9707 (N_9707,N_6629,N_7474);
nand U9708 (N_9708,N_7571,N_8360);
and U9709 (N_9709,N_6267,N_8480);
and U9710 (N_9710,N_8529,N_7906);
or U9711 (N_9711,N_6104,N_6346);
nor U9712 (N_9712,N_7069,N_6529);
or U9713 (N_9713,N_8334,N_7210);
nand U9714 (N_9714,N_7922,N_8710);
or U9715 (N_9715,N_8644,N_7954);
or U9716 (N_9716,N_7195,N_6571);
or U9717 (N_9717,N_8758,N_6424);
or U9718 (N_9718,N_6176,N_8843);
xor U9719 (N_9719,N_8522,N_6971);
or U9720 (N_9720,N_7436,N_8008);
nand U9721 (N_9721,N_8005,N_6013);
nor U9722 (N_9722,N_8064,N_6263);
nor U9723 (N_9723,N_6497,N_6014);
xnor U9724 (N_9724,N_7160,N_7095);
nand U9725 (N_9725,N_8179,N_8332);
xnor U9726 (N_9726,N_7852,N_6589);
or U9727 (N_9727,N_6210,N_8791);
and U9728 (N_9728,N_8910,N_8412);
and U9729 (N_9729,N_7859,N_7236);
or U9730 (N_9730,N_7803,N_8348);
xor U9731 (N_9731,N_7539,N_6818);
and U9732 (N_9732,N_7759,N_8091);
nor U9733 (N_9733,N_7313,N_8973);
nand U9734 (N_9734,N_7858,N_8354);
xnor U9735 (N_9735,N_6226,N_6582);
or U9736 (N_9736,N_7497,N_6955);
nand U9737 (N_9737,N_7574,N_8524);
xnor U9738 (N_9738,N_7546,N_8653);
nor U9739 (N_9739,N_6377,N_8025);
nand U9740 (N_9740,N_7131,N_8966);
nor U9741 (N_9741,N_7286,N_8606);
nor U9742 (N_9742,N_8322,N_8235);
nand U9743 (N_9743,N_6132,N_6547);
or U9744 (N_9744,N_6948,N_8454);
or U9745 (N_9745,N_6981,N_8347);
nand U9746 (N_9746,N_6549,N_6035);
and U9747 (N_9747,N_7262,N_6674);
xor U9748 (N_9748,N_8747,N_8873);
xor U9749 (N_9749,N_6214,N_8663);
nand U9750 (N_9750,N_8166,N_8755);
and U9751 (N_9751,N_8773,N_7682);
nor U9752 (N_9752,N_7867,N_7580);
nor U9753 (N_9753,N_7540,N_8861);
xnor U9754 (N_9754,N_6740,N_7065);
or U9755 (N_9755,N_7118,N_6364);
and U9756 (N_9756,N_7866,N_6311);
or U9757 (N_9757,N_6599,N_6904);
xor U9758 (N_9758,N_6952,N_8680);
and U9759 (N_9759,N_7221,N_8953);
and U9760 (N_9760,N_7751,N_7640);
nand U9761 (N_9761,N_7219,N_6745);
nand U9762 (N_9762,N_6018,N_6141);
nor U9763 (N_9763,N_7137,N_6344);
xor U9764 (N_9764,N_7465,N_8073);
nor U9765 (N_9765,N_7838,N_8475);
nor U9766 (N_9766,N_8671,N_6977);
xnor U9767 (N_9767,N_8623,N_7693);
nand U9768 (N_9768,N_6839,N_6387);
and U9769 (N_9769,N_7072,N_6992);
and U9770 (N_9770,N_7185,N_6384);
or U9771 (N_9771,N_6194,N_7154);
xor U9772 (N_9772,N_6716,N_8485);
nor U9773 (N_9773,N_7470,N_6650);
xor U9774 (N_9774,N_6871,N_6814);
nor U9775 (N_9775,N_6373,N_7509);
nand U9776 (N_9776,N_8139,N_6897);
and U9777 (N_9777,N_8545,N_8164);
and U9778 (N_9778,N_6077,N_8003);
or U9779 (N_9779,N_7617,N_7547);
and U9780 (N_9780,N_7881,N_8975);
xnor U9781 (N_9781,N_7797,N_7386);
nor U9782 (N_9782,N_8616,N_7503);
and U9783 (N_9783,N_7830,N_7983);
or U9784 (N_9784,N_7365,N_6799);
nand U9785 (N_9785,N_8521,N_6704);
xnor U9786 (N_9786,N_6425,N_8750);
nor U9787 (N_9787,N_6278,N_6515);
nor U9788 (N_9788,N_7035,N_6469);
or U9789 (N_9789,N_7496,N_8425);
or U9790 (N_9790,N_6562,N_8147);
xor U9791 (N_9791,N_8891,N_8756);
nand U9792 (N_9792,N_7126,N_6881);
xnor U9793 (N_9793,N_7258,N_6129);
and U9794 (N_9794,N_7597,N_8963);
or U9795 (N_9795,N_6494,N_7605);
nor U9796 (N_9796,N_6618,N_7632);
and U9797 (N_9797,N_7488,N_7876);
nand U9798 (N_9798,N_6982,N_6983);
xnor U9799 (N_9799,N_7009,N_8687);
nor U9800 (N_9800,N_7643,N_8240);
nor U9801 (N_9801,N_8690,N_8739);
xnor U9802 (N_9802,N_6749,N_7770);
nor U9803 (N_9803,N_7826,N_8236);
nor U9804 (N_9804,N_8892,N_6067);
xor U9805 (N_9805,N_7582,N_7610);
and U9806 (N_9806,N_7271,N_7807);
or U9807 (N_9807,N_6304,N_7976);
nand U9808 (N_9808,N_6808,N_7602);
xnor U9809 (N_9809,N_7705,N_7135);
nor U9810 (N_9810,N_6984,N_7971);
nand U9811 (N_9811,N_8097,N_8985);
xnor U9812 (N_9812,N_6711,N_7732);
and U9813 (N_9813,N_8630,N_7950);
nand U9814 (N_9814,N_7659,N_6489);
xor U9815 (N_9815,N_8199,N_8918);
or U9816 (N_9816,N_6503,N_8640);
or U9817 (N_9817,N_8406,N_7812);
nand U9818 (N_9818,N_7646,N_6321);
nand U9819 (N_9819,N_7186,N_8799);
xnor U9820 (N_9820,N_6417,N_8631);
xnor U9821 (N_9821,N_6685,N_6020);
or U9822 (N_9822,N_8566,N_7220);
nor U9823 (N_9823,N_8584,N_6185);
xor U9824 (N_9824,N_8197,N_6573);
nor U9825 (N_9825,N_8225,N_6870);
and U9826 (N_9826,N_8840,N_8210);
or U9827 (N_9827,N_7843,N_6187);
nor U9828 (N_9828,N_8911,N_6533);
or U9829 (N_9829,N_6109,N_7050);
and U9830 (N_9830,N_7330,N_6395);
and U9831 (N_9831,N_6692,N_6682);
and U9832 (N_9832,N_7568,N_6615);
xor U9833 (N_9833,N_8627,N_7860);
and U9834 (N_9834,N_6401,N_7740);
xor U9835 (N_9835,N_6875,N_6954);
nor U9836 (N_9836,N_6156,N_7428);
nor U9837 (N_9837,N_7047,N_6079);
or U9838 (N_9838,N_8086,N_7382);
xor U9839 (N_9839,N_8807,N_8100);
xor U9840 (N_9840,N_8084,N_6085);
xnor U9841 (N_9841,N_8603,N_8781);
xnor U9842 (N_9842,N_6545,N_7912);
nor U9843 (N_9843,N_7371,N_7327);
nand U9844 (N_9844,N_7720,N_6802);
xor U9845 (N_9845,N_6614,N_7758);
xnor U9846 (N_9846,N_8601,N_8659);
nand U9847 (N_9847,N_7601,N_8785);
and U9848 (N_9848,N_6700,N_8047);
and U9849 (N_9849,N_6922,N_7063);
nand U9850 (N_9850,N_6191,N_7081);
nand U9851 (N_9851,N_6362,N_8217);
or U9852 (N_9852,N_8984,N_6011);
nor U9853 (N_9853,N_7611,N_7116);
nor U9854 (N_9854,N_7998,N_8696);
xnor U9855 (N_9855,N_6604,N_7287);
nor U9856 (N_9856,N_7941,N_6862);
xnor U9857 (N_9857,N_6479,N_7401);
nor U9858 (N_9858,N_7672,N_8433);
or U9859 (N_9859,N_6867,N_8780);
nand U9860 (N_9860,N_8518,N_6767);
nor U9861 (N_9861,N_6329,N_7788);
nand U9862 (N_9862,N_8056,N_6748);
xnor U9863 (N_9863,N_7319,N_6258);
and U9864 (N_9864,N_8794,N_8135);
or U9865 (N_9865,N_8075,N_6276);
xor U9866 (N_9866,N_6153,N_7709);
and U9867 (N_9867,N_6645,N_8057);
or U9868 (N_9868,N_6720,N_6899);
or U9869 (N_9869,N_8418,N_7461);
or U9870 (N_9870,N_8438,N_8759);
xor U9871 (N_9871,N_7473,N_6099);
xnor U9872 (N_9872,N_8926,N_8974);
nor U9873 (N_9873,N_6284,N_6877);
nor U9874 (N_9874,N_6924,N_6606);
and U9875 (N_9875,N_6853,N_6081);
nor U9876 (N_9876,N_8609,N_6261);
and U9877 (N_9877,N_6446,N_8820);
nand U9878 (N_9878,N_6822,N_8112);
or U9879 (N_9879,N_6120,N_7370);
nor U9880 (N_9880,N_7935,N_8373);
and U9881 (N_9881,N_8120,N_8308);
nand U9882 (N_9882,N_8683,N_8967);
and U9883 (N_9883,N_7595,N_6365);
nand U9884 (N_9884,N_7821,N_8344);
or U9885 (N_9885,N_6125,N_8588);
and U9886 (N_9886,N_7555,N_6691);
nor U9887 (N_9887,N_7933,N_6891);
and U9888 (N_9888,N_8268,N_7385);
and U9889 (N_9889,N_7469,N_8500);
nand U9890 (N_9890,N_7458,N_6498);
and U9891 (N_9891,N_7945,N_8995);
nor U9892 (N_9892,N_8148,N_7960);
xor U9893 (N_9893,N_6686,N_7429);
nand U9894 (N_9894,N_6108,N_6568);
xor U9895 (N_9895,N_6895,N_7471);
xnor U9896 (N_9896,N_8465,N_6248);
nand U9897 (N_9897,N_8137,N_8699);
nand U9898 (N_9898,N_7894,N_7028);
nor U9899 (N_9899,N_8230,N_6538);
xnor U9900 (N_9900,N_8294,N_6433);
nor U9901 (N_9901,N_7743,N_6071);
xnor U9902 (N_9902,N_7572,N_8611);
and U9903 (N_9903,N_6315,N_7840);
xor U9904 (N_9904,N_8564,N_8568);
or U9905 (N_9905,N_7518,N_7005);
nand U9906 (N_9906,N_6164,N_6466);
or U9907 (N_9907,N_8181,N_8560);
or U9908 (N_9908,N_7132,N_7085);
xnor U9909 (N_9909,N_8717,N_8459);
or U9910 (N_9910,N_8886,N_7712);
and U9911 (N_9911,N_6919,N_8183);
nor U9912 (N_9912,N_8723,N_6916);
nor U9913 (N_9913,N_6653,N_6171);
nand U9914 (N_9914,N_8648,N_6190);
and U9915 (N_9915,N_6521,N_7544);
or U9916 (N_9916,N_7942,N_7841);
nand U9917 (N_9917,N_7609,N_6010);
xor U9918 (N_9918,N_7178,N_7808);
nor U9919 (N_9919,N_7827,N_8932);
nor U9920 (N_9920,N_6122,N_7641);
nand U9921 (N_9921,N_7533,N_7418);
and U9922 (N_9922,N_8170,N_8514);
nor U9923 (N_9923,N_6002,N_7166);
or U9924 (N_9924,N_8660,N_7565);
and U9925 (N_9925,N_6114,N_7916);
and U9926 (N_9926,N_8471,N_7614);
or U9927 (N_9927,N_8107,N_7433);
or U9928 (N_9928,N_7298,N_7378);
nand U9929 (N_9929,N_8817,N_7124);
xor U9930 (N_9930,N_7134,N_8114);
xor U9931 (N_9931,N_6668,N_8320);
nand U9932 (N_9932,N_8443,N_7060);
or U9933 (N_9933,N_6856,N_7988);
nand U9934 (N_9934,N_7552,N_7880);
or U9935 (N_9935,N_7691,N_6215);
xnor U9936 (N_9936,N_6294,N_8549);
and U9937 (N_9937,N_8573,N_7409);
xnor U9938 (N_9938,N_8592,N_7275);
xor U9939 (N_9939,N_8083,N_7021);
and U9940 (N_9940,N_7495,N_7222);
or U9941 (N_9941,N_8374,N_7952);
and U9942 (N_9942,N_6499,N_8803);
nand U9943 (N_9943,N_7058,N_7957);
or U9944 (N_9944,N_8007,N_7679);
xnor U9945 (N_9945,N_8689,N_6590);
xor U9946 (N_9946,N_7192,N_7676);
or U9947 (N_9947,N_6942,N_6953);
xnor U9948 (N_9948,N_6760,N_7150);
or U9949 (N_9949,N_8533,N_7398);
nor U9950 (N_9950,N_8127,N_7218);
nor U9951 (N_9951,N_8329,N_8638);
nand U9952 (N_9952,N_7381,N_8846);
nor U9953 (N_9953,N_8129,N_7015);
nor U9954 (N_9954,N_7406,N_8295);
xnor U9955 (N_9955,N_6009,N_8955);
xnor U9956 (N_9956,N_7184,N_7068);
or U9957 (N_9957,N_6063,N_8027);
or U9958 (N_9958,N_7644,N_8617);
or U9959 (N_9959,N_8870,N_7322);
and U9960 (N_9960,N_6690,N_8565);
and U9961 (N_9961,N_8380,N_7453);
xor U9962 (N_9962,N_7559,N_8615);
nand U9963 (N_9963,N_6170,N_7869);
nand U9964 (N_9964,N_7851,N_7907);
and U9965 (N_9965,N_7029,N_6462);
and U9966 (N_9966,N_7669,N_8628);
and U9967 (N_9967,N_7017,N_8679);
xor U9968 (N_9968,N_8941,N_8247);
and U9969 (N_9969,N_7320,N_6804);
or U9970 (N_9970,N_6033,N_6218);
xnor U9971 (N_9971,N_6043,N_6174);
nor U9972 (N_9972,N_8154,N_6785);
and U9973 (N_9973,N_6507,N_7411);
or U9974 (N_9974,N_6730,N_8044);
or U9975 (N_9975,N_7699,N_6432);
xnor U9976 (N_9976,N_7787,N_8063);
xnor U9977 (N_9977,N_6065,N_7754);
nand U9978 (N_9978,N_6997,N_6152);
xnor U9979 (N_9979,N_7043,N_8281);
nor U9980 (N_9980,N_6012,N_7399);
xnor U9981 (N_9981,N_6985,N_7454);
nor U9982 (N_9982,N_6471,N_6087);
xnor U9983 (N_9983,N_7476,N_6673);
nand U9984 (N_9984,N_6656,N_8917);
and U9985 (N_9985,N_7360,N_6128);
and U9986 (N_9986,N_7736,N_6030);
and U9987 (N_9987,N_6366,N_8833);
xor U9988 (N_9988,N_6130,N_7755);
or U9989 (N_9989,N_7484,N_6641);
xor U9990 (N_9990,N_6175,N_6967);
xor U9991 (N_9991,N_6637,N_7439);
xor U9992 (N_9992,N_6866,N_7413);
xor U9993 (N_9993,N_7765,N_8223);
and U9994 (N_9994,N_8361,N_7066);
and U9995 (N_9995,N_6336,N_6914);
nand U9996 (N_9996,N_7561,N_8364);
and U9997 (N_9997,N_6902,N_8872);
nor U9998 (N_9998,N_8358,N_6219);
xor U9999 (N_9999,N_6696,N_7089);
nand U10000 (N_10000,N_6815,N_8482);
or U10001 (N_10001,N_7182,N_8898);
nor U10002 (N_10002,N_6124,N_8986);
and U10003 (N_10003,N_7531,N_7442);
and U10004 (N_10004,N_7177,N_6929);
xor U10005 (N_10005,N_7786,N_8520);
nor U10006 (N_10006,N_7191,N_7767);
nand U10007 (N_10007,N_6257,N_6559);
and U10008 (N_10008,N_7608,N_6246);
or U10009 (N_10009,N_7596,N_8207);
nor U10010 (N_10010,N_6928,N_6698);
nand U10011 (N_10011,N_7456,N_8188);
or U10012 (N_10012,N_8839,N_6317);
xor U10013 (N_10013,N_8720,N_8701);
nor U10014 (N_10014,N_7312,N_7968);
and U10015 (N_10015,N_8619,N_6312);
nand U10016 (N_10016,N_6636,N_6543);
and U10017 (N_10017,N_8804,N_8191);
or U10018 (N_10018,N_6795,N_8030);
nand U10019 (N_10019,N_7635,N_7598);
xnor U10020 (N_10020,N_6247,N_8017);
nor U10021 (N_10021,N_8140,N_6796);
or U10022 (N_10022,N_7929,N_8544);
or U10023 (N_10023,N_8704,N_8255);
xnor U10024 (N_10024,N_6183,N_6357);
and U10025 (N_10025,N_8834,N_6718);
or U10026 (N_10026,N_7811,N_6238);
and U10027 (N_10027,N_8430,N_6883);
and U10028 (N_10028,N_6960,N_6182);
nand U10029 (N_10029,N_7535,N_7041);
xor U10030 (N_10030,N_8489,N_8468);
or U10031 (N_10031,N_8719,N_7656);
and U10032 (N_10032,N_6240,N_6360);
nand U10033 (N_10033,N_8011,N_6282);
nor U10034 (N_10034,N_8889,N_6633);
and U10035 (N_10035,N_6477,N_6042);
nor U10036 (N_10036,N_7462,N_8655);
or U10037 (N_10037,N_7334,N_8399);
nor U10038 (N_10038,N_7061,N_6430);
or U10039 (N_10039,N_8404,N_8457);
nor U10040 (N_10040,N_6608,N_6169);
nor U10041 (N_10041,N_6379,N_8554);
or U10042 (N_10042,N_7768,N_8593);
nor U10043 (N_10043,N_7715,N_6906);
nor U10044 (N_10044,N_7159,N_6468);
or U10045 (N_10045,N_8249,N_8330);
and U10046 (N_10046,N_7451,N_7139);
xor U10047 (N_10047,N_7040,N_7575);
and U10048 (N_10048,N_8012,N_6165);
and U10049 (N_10049,N_8194,N_8411);
xor U10050 (N_10050,N_6710,N_8277);
or U10051 (N_10051,N_8965,N_6403);
nand U10052 (N_10052,N_8948,N_6102);
or U10053 (N_10053,N_7822,N_8826);
and U10054 (N_10054,N_7256,N_7628);
nor U10055 (N_10055,N_8149,N_7146);
xor U10056 (N_10056,N_8658,N_8262);
nand U10057 (N_10057,N_6350,N_8387);
nor U10058 (N_10058,N_8001,N_6658);
xnor U10059 (N_10059,N_8855,N_6849);
xor U10060 (N_10060,N_7527,N_6517);
or U10061 (N_10061,N_7895,N_8031);
nor U10062 (N_10062,N_6565,N_7967);
or U10063 (N_10063,N_8059,N_8023);
nand U10064 (N_10064,N_8916,N_6234);
nand U10065 (N_10065,N_6024,N_8125);
xor U10066 (N_10066,N_7994,N_7652);
and U10067 (N_10067,N_7763,N_6577);
nor U10068 (N_10068,N_8740,N_6754);
nand U10069 (N_10069,N_6021,N_6841);
nor U10070 (N_10070,N_7153,N_8774);
nor U10071 (N_10071,N_6829,N_7198);
xnor U10072 (N_10072,N_7425,N_8887);
xor U10073 (N_10073,N_8391,N_8313);
nand U10074 (N_10074,N_8015,N_7310);
or U10075 (N_10075,N_8157,N_7774);
and U10076 (N_10076,N_6242,N_6500);
or U10077 (N_10077,N_8787,N_8779);
nand U10078 (N_10078,N_8424,N_6059);
xnor U10079 (N_10079,N_7517,N_7733);
nand U10080 (N_10080,N_6166,N_7173);
or U10081 (N_10081,N_7105,N_6996);
and U10082 (N_10082,N_7011,N_6241);
xor U10083 (N_10083,N_7165,N_8492);
and U10084 (N_10084,N_7491,N_8595);
nand U10085 (N_10085,N_8877,N_7487);
nor U10086 (N_10086,N_6878,N_7084);
or U10087 (N_10087,N_8414,N_7303);
nand U10088 (N_10088,N_7717,N_7729);
or U10089 (N_10089,N_6472,N_8458);
nand U10090 (N_10090,N_8108,N_8881);
xnor U10091 (N_10091,N_6512,N_8293);
or U10092 (N_10092,N_8371,N_6396);
nor U10093 (N_10093,N_8357,N_6287);
nand U10094 (N_10094,N_8919,N_7447);
and U10095 (N_10095,N_8385,N_6342);
or U10096 (N_10096,N_6537,N_7337);
and U10097 (N_10097,N_6778,N_6506);
nor U10098 (N_10098,N_7125,N_7316);
nand U10099 (N_10099,N_7294,N_7620);
nor U10100 (N_10100,N_7567,N_6149);
or U10101 (N_10101,N_8625,N_8420);
and U10102 (N_10102,N_8649,N_6136);
or U10103 (N_10103,N_7364,N_6325);
nor U10104 (N_10104,N_8908,N_6250);
or U10105 (N_10105,N_7324,N_6678);
and U10106 (N_10106,N_7663,N_7764);
and U10107 (N_10107,N_6492,N_7468);
nand U10108 (N_10108,N_6525,N_7675);
nand U10109 (N_10109,N_6464,N_8802);
or U10110 (N_10110,N_6595,N_8286);
nor U10111 (N_10111,N_6719,N_7701);
nor U10112 (N_10112,N_8778,N_8922);
xnor U10113 (N_10113,N_8159,N_7232);
or U10114 (N_10114,N_6832,N_6672);
nor U10115 (N_10115,N_8842,N_6993);
or U10116 (N_10116,N_8267,N_6516);
nor U10117 (N_10117,N_8109,N_6200);
and U10118 (N_10118,N_6291,N_8999);
nor U10119 (N_10119,N_7415,N_7987);
nand U10120 (N_10120,N_8491,N_7092);
nand U10121 (N_10121,N_7202,N_6734);
and U10122 (N_10122,N_6093,N_7355);
nand U10123 (N_10123,N_7794,N_8897);
nor U10124 (N_10124,N_7188,N_7835);
xor U10125 (N_10125,N_7403,N_8248);
nand U10126 (N_10126,N_6407,N_6476);
and U10127 (N_10127,N_6046,N_7026);
xor U10128 (N_10128,N_6540,N_8553);
and U10129 (N_10129,N_7136,N_8836);
nand U10130 (N_10130,N_6144,N_7164);
or U10131 (N_10131,N_7735,N_8712);
xor U10132 (N_10132,N_6820,N_6145);
or U10133 (N_10133,N_6757,N_7864);
or U10134 (N_10134,N_6426,N_7044);
and U10135 (N_10135,N_7420,N_8036);
or U10136 (N_10136,N_6840,N_8841);
or U10137 (N_10137,N_7071,N_8645);
nor U10138 (N_10138,N_7392,N_6945);
xor U10139 (N_10139,N_7340,N_7514);
nor U10140 (N_10140,N_7616,N_6779);
nand U10141 (N_10141,N_8978,N_7247);
and U10142 (N_10142,N_7295,N_8193);
and U10143 (N_10143,N_6966,N_7472);
nor U10144 (N_10144,N_7839,N_8352);
or U10145 (N_10145,N_8596,N_8019);
nand U10146 (N_10146,N_6367,N_6624);
nand U10147 (N_10147,N_6470,N_7637);
nand U10148 (N_10148,N_8431,N_8496);
nand U10149 (N_10149,N_8851,N_6872);
xor U10150 (N_10150,N_7339,N_7363);
xor U10151 (N_10151,N_8844,N_8548);
xor U10152 (N_10152,N_7000,N_6252);
xor U10153 (N_10153,N_6852,N_6487);
xor U10154 (N_10154,N_6836,N_7772);
nand U10155 (N_10155,N_7070,N_8173);
nor U10156 (N_10156,N_8944,N_7708);
nor U10157 (N_10157,N_8232,N_7541);
xor U10158 (N_10158,N_6789,N_6838);
xor U10159 (N_10159,N_8610,N_6541);
and U10160 (N_10160,N_6456,N_7359);
nor U10161 (N_10161,N_7594,N_7157);
or U10162 (N_10162,N_6630,N_8863);
xor U10163 (N_10163,N_6356,N_6671);
nand U10164 (N_10164,N_8867,N_8311);
nor U10165 (N_10165,N_8142,N_8400);
nand U10166 (N_10166,N_7657,N_6110);
or U10167 (N_10167,N_8289,N_8265);
nor U10168 (N_10168,N_6947,N_7901);
nand U10169 (N_10169,N_6903,N_6882);
xor U10170 (N_10170,N_6098,N_6160);
nand U10171 (N_10171,N_7022,N_7990);
or U10172 (N_10172,N_6978,N_8771);
nand U10173 (N_10173,N_6328,N_6313);
or U10174 (N_10174,N_6305,N_6552);
xor U10175 (N_10175,N_8081,N_8160);
or U10176 (N_10176,N_6480,N_7748);
nor U10177 (N_10177,N_7799,N_7328);
or U10178 (N_10178,N_6912,N_7255);
xor U10179 (N_10179,N_8032,N_6281);
nor U10180 (N_10180,N_6773,N_6173);
nand U10181 (N_10181,N_8158,N_8537);
and U10182 (N_10182,N_6625,N_7128);
nand U10183 (N_10183,N_8098,N_6556);
or U10184 (N_10184,N_7291,N_6775);
or U10185 (N_10185,N_7446,N_8000);
or U10186 (N_10186,N_8341,N_7438);
and U10187 (N_10187,N_7483,N_8282);
xnor U10188 (N_10188,N_6732,N_7785);
or U10189 (N_10189,N_6986,N_8639);
nor U10190 (N_10190,N_6623,N_8092);
or U10191 (N_10191,N_8085,N_6393);
and U10192 (N_10192,N_6319,N_6060);
nor U10193 (N_10193,N_6664,N_7237);
nor U10194 (N_10194,N_7181,N_8463);
and U10195 (N_10195,N_6646,N_8372);
or U10196 (N_10196,N_6375,N_8133);
and U10197 (N_10197,N_8677,N_6560);
xnor U10198 (N_10198,N_7537,N_8721);
nand U10199 (N_10199,N_6272,N_7985);
xnor U10200 (N_10200,N_6352,N_7897);
and U10201 (N_10201,N_7554,N_8009);
nand U10202 (N_10202,N_7197,N_8220);
xnor U10203 (N_10203,N_8227,N_8629);
and U10204 (N_10204,N_6884,N_6207);
xor U10205 (N_10205,N_8415,N_8428);
and U10206 (N_10206,N_6837,N_7773);
xnor U10207 (N_10207,N_7861,N_6331);
nor U10208 (N_10208,N_7304,N_6348);
and U10209 (N_10209,N_8970,N_6662);
or U10210 (N_10210,N_6683,N_6092);
and U10211 (N_10211,N_7992,N_6548);
nor U10212 (N_10212,N_8950,N_6701);
and U10213 (N_10213,N_8816,N_8049);
xor U10214 (N_10214,N_8743,N_8318);
nor U10215 (N_10215,N_6787,N_8324);
xnor U10216 (N_10216,N_7779,N_8519);
or U10217 (N_10217,N_7974,N_8055);
nand U10218 (N_10218,N_7464,N_7492);
or U10219 (N_10219,N_6036,N_7374);
or U10220 (N_10220,N_8946,N_6855);
nand U10221 (N_10221,N_8228,N_8416);
and U10222 (N_10222,N_8968,N_7534);
and U10223 (N_10223,N_7151,N_7698);
nand U10224 (N_10224,N_6905,N_7384);
and U10225 (N_10225,N_6999,N_8688);
or U10226 (N_10226,N_8261,N_7138);
nor U10227 (N_10227,N_8770,N_8909);
xor U10228 (N_10228,N_7368,N_7245);
and U10229 (N_10229,N_7674,N_6301);
and U10230 (N_10230,N_8186,N_6347);
nor U10231 (N_10231,N_7685,N_8582);
xor U10232 (N_10232,N_7972,N_7431);
and U10233 (N_10233,N_8823,N_7744);
and U10234 (N_10234,N_7536,N_6076);
nand U10235 (N_10235,N_7850,N_6729);
xor U10236 (N_10236,N_7100,N_6458);
xnor U10237 (N_10237,N_6335,N_8211);
and U10238 (N_10238,N_8924,N_6400);
xnor U10239 (N_10239,N_8981,N_6052);
xnor U10240 (N_10240,N_8577,N_7815);
and U10241 (N_10241,N_7944,N_8523);
nand U10242 (N_10242,N_7325,N_7938);
xor U10243 (N_10243,N_8929,N_7877);
or U10244 (N_10244,N_7270,N_8451);
and U10245 (N_10245,N_6848,N_7703);
xor U10246 (N_10246,N_6116,N_8487);
nand U10247 (N_10247,N_7130,N_6725);
nor U10248 (N_10248,N_6782,N_6115);
or U10249 (N_10249,N_7576,N_6620);
xnor U10250 (N_10250,N_8532,N_8783);
or U10251 (N_10251,N_7914,N_8570);
nand U10252 (N_10252,N_8238,N_8270);
or U10253 (N_10253,N_7030,N_7590);
nand U10254 (N_10254,N_8256,N_7057);
or U10255 (N_10255,N_7522,N_6058);
and U10256 (N_10256,N_7248,N_6459);
nor U10257 (N_10257,N_8275,N_8883);
or U10258 (N_10258,N_8040,N_7857);
or U10259 (N_10259,N_6320,N_8665);
or U10260 (N_10260,N_8342,N_8452);
xnor U10261 (N_10261,N_7073,N_8285);
nor U10262 (N_10262,N_7723,N_8624);
nand U10263 (N_10263,N_7634,N_7562);
or U10264 (N_10264,N_7416,N_6073);
xnor U10265 (N_10265,N_7170,N_8736);
and U10266 (N_10266,N_6211,N_8571);
nand U10267 (N_10267,N_8535,N_7684);
nor U10268 (N_10268,N_8460,N_7149);
or U10269 (N_10269,N_6596,N_8983);
nor U10270 (N_10270,N_8224,N_6159);
or U10271 (N_10271,N_8620,N_7482);
and U10272 (N_10272,N_7982,N_8695);
nand U10273 (N_10273,N_6224,N_8014);
nand U10274 (N_10274,N_7956,N_7091);
nand U10275 (N_10275,N_7274,N_8622);
xnor U10276 (N_10276,N_8006,N_6706);
or U10277 (N_10277,N_7140,N_8447);
or U10278 (N_10278,N_8760,N_7342);
nor U10279 (N_10279,N_8209,N_8244);
or U10280 (N_10280,N_6688,N_7430);
xor U10281 (N_10281,N_6935,N_6026);
or U10282 (N_10282,N_8377,N_7936);
nand U10283 (N_10283,N_6679,N_6484);
and U10284 (N_10284,N_6465,N_6445);
or U10285 (N_10285,N_8862,N_6991);
nor U10286 (N_10286,N_8184,N_7407);
xor U10287 (N_10287,N_8467,N_8578);
xor U10288 (N_10288,N_7259,N_8957);
and U10289 (N_10289,N_8396,N_7588);
or U10290 (N_10290,N_7037,N_7790);
nor U10291 (N_10291,N_8421,N_8359);
and U10292 (N_10292,N_6259,N_8422);
xnor U10293 (N_10293,N_8042,N_8920);
nand U10294 (N_10294,N_7873,N_8531);
and U10295 (N_10295,N_7333,N_8392);
xnor U10296 (N_10296,N_6743,N_6198);
xnor U10297 (N_10297,N_7038,N_6370);
nor U10298 (N_10298,N_8309,N_8026);
nand U10299 (N_10299,N_8035,N_8517);
nor U10300 (N_10300,N_8874,N_6457);
nand U10301 (N_10301,N_8099,N_8605);
nor U10302 (N_10302,N_6739,N_6554);
nand U10303 (N_10303,N_6293,N_7049);
nand U10304 (N_10304,N_7285,N_6090);
nand U10305 (N_10305,N_8436,N_8790);
nand U10306 (N_10306,N_7686,N_8060);
nand U10307 (N_10307,N_8879,N_8205);
nand U10308 (N_10308,N_6161,N_6764);
xor U10309 (N_10309,N_6334,N_8831);
and U10310 (N_10310,N_8657,N_8074);
and U10311 (N_10311,N_8635,N_6146);
or U10312 (N_10312,N_6797,N_8812);
or U10313 (N_10313,N_7020,N_7435);
nor U10314 (N_10314,N_6846,N_6987);
nand U10315 (N_10315,N_7724,N_8050);
or U10316 (N_10316,N_7098,N_7910);
nand U10317 (N_10317,N_8189,N_7981);
xnor U10318 (N_10318,N_6687,N_7820);
or U10319 (N_10319,N_6351,N_6975);
or U10320 (N_10320,N_6934,N_8366);
or U10321 (N_10321,N_6994,N_7189);
and U10322 (N_10322,N_6536,N_8800);
and U10323 (N_10323,N_6195,N_6088);
and U10324 (N_10324,N_7115,N_6544);
xor U10325 (N_10325,N_7090,N_6724);
nor U10326 (N_10326,N_8847,N_8796);
xor U10327 (N_10327,N_7390,N_8077);
nand U10328 (N_10328,N_6355,N_8029);
and U10329 (N_10329,N_7144,N_8830);
or U10330 (N_10330,N_8557,N_6622);
nand U10331 (N_10331,N_6825,N_8951);
xor U10332 (N_10332,N_6951,N_7380);
and U10333 (N_10333,N_8694,N_6607);
nor U10334 (N_10334,N_8643,N_7373);
nand U10335 (N_10335,N_6597,N_7109);
nor U10336 (N_10336,N_7200,N_7874);
xnor U10337 (N_10337,N_8541,N_6023);
or U10338 (N_10338,N_8010,N_7966);
xor U10339 (N_10339,N_6874,N_8943);
nor U10340 (N_10340,N_8245,N_7332);
xnor U10341 (N_10341,N_7553,N_7059);
nor U10342 (N_10342,N_6666,N_6223);
nor U10343 (N_10343,N_8636,N_7885);
nor U10344 (N_10344,N_6096,N_7031);
nand U10345 (N_10345,N_7244,N_6958);
xnor U10346 (N_10346,N_8124,N_6889);
nand U10347 (N_10347,N_7511,N_7949);
nand U10348 (N_10348,N_8904,N_6332);
xnor U10349 (N_10349,N_6786,N_6643);
nor U10350 (N_10350,N_8498,N_7080);
nor U10351 (N_10351,N_7716,N_7913);
and U10352 (N_10352,N_6126,N_8905);
and U10353 (N_10353,N_8664,N_6531);
and U10354 (N_10354,N_6574,N_8162);
or U10355 (N_10355,N_7437,N_8868);
nand U10356 (N_10356,N_6944,N_8927);
nor U10357 (N_10357,N_6858,N_8013);
and U10358 (N_10358,N_7834,N_7791);
xnor U10359 (N_10359,N_8273,N_6213);
nor U10360 (N_10360,N_6961,N_7671);
xnor U10361 (N_10361,N_8933,N_6555);
and U10362 (N_10362,N_8977,N_7586);
nor U10363 (N_10363,N_8161,N_8021);
xnor U10364 (N_10364,N_7481,N_7459);
or U10365 (N_10365,N_8054,N_8956);
or U10366 (N_10366,N_7932,N_6976);
nor U10367 (N_10367,N_7896,N_6299);
and U10368 (N_10368,N_8250,N_8315);
xor U10369 (N_10369,N_8058,N_8510);
or U10370 (N_10370,N_7358,N_6409);
nand U10371 (N_10371,N_7362,N_8122);
nand U10372 (N_10372,N_7163,N_8333);
xor U10373 (N_10373,N_7112,N_6695);
nand U10374 (N_10374,N_8558,N_8822);
xor U10375 (N_10375,N_6055,N_6892);
or U10376 (N_10376,N_6371,N_8786);
xnor U10377 (N_10377,N_6514,N_6427);
and U10378 (N_10378,N_7926,N_6963);
and U10379 (N_10379,N_6530,N_8410);
and U10380 (N_10380,N_6860,N_7865);
xnor U10381 (N_10381,N_6041,N_6455);
or U10382 (N_10382,N_7230,N_7279);
or U10383 (N_10383,N_7282,N_8763);
nand U10384 (N_10384,N_6703,N_7036);
nand U10385 (N_10385,N_6925,N_8741);
nand U10386 (N_10386,N_6032,N_7396);
and U10387 (N_10387,N_8128,N_6411);
and U10388 (N_10388,N_8078,N_8772);
and U10389 (N_10389,N_6022,N_8551);
nand U10390 (N_10390,N_6587,N_8896);
nand U10391 (N_10391,N_8094,N_8947);
nor U10392 (N_10392,N_6998,N_7301);
nand U10393 (N_10393,N_6990,N_6277);
xnor U10394 (N_10394,N_8310,N_7306);
or U10395 (N_10395,N_7205,N_6962);
xor U10396 (N_10396,N_8633,N_7498);
nand U10397 (N_10397,N_7937,N_7824);
or U10398 (N_10398,N_7738,N_7526);
nor U10399 (N_10399,N_6819,N_6728);
nor U10400 (N_10400,N_7265,N_8562);
and U10401 (N_10401,N_6151,N_6727);
and U10402 (N_10402,N_6103,N_8543);
and U10403 (N_10403,N_7445,N_8809);
and U10404 (N_10404,N_6265,N_6031);
nor U10405 (N_10405,N_7174,N_8052);
and U10406 (N_10406,N_6491,N_8272);
and U10407 (N_10407,N_8692,N_8682);
nand U10408 (N_10408,N_7083,N_8954);
and U10409 (N_10409,N_6681,N_6712);
nor U10410 (N_10410,N_8349,N_6708);
nor U10411 (N_10411,N_7296,N_7231);
or U10412 (N_10412,N_6296,N_8155);
nor U10413 (N_10413,N_7133,N_6752);
nor U10414 (N_10414,N_8134,N_8727);
xnor U10415 (N_10415,N_7805,N_8115);
nand U10416 (N_10416,N_8257,N_7962);
xnor U10417 (N_10417,N_8038,N_8576);
or U10418 (N_10418,N_6236,N_7148);
nand U10419 (N_10419,N_8218,N_8590);
nand U10420 (N_10420,N_7311,N_7891);
nand U10421 (N_10421,N_6833,N_7918);
nand U10422 (N_10422,N_7969,N_7909);
or U10423 (N_10423,N_6885,N_8572);
xnor U10424 (N_10424,N_7923,N_6040);
nand U10425 (N_10425,N_7591,N_7507);
nor U10426 (N_10426,N_6827,N_6989);
nor U10427 (N_10427,N_7934,N_7621);
xnor U10428 (N_10428,N_7240,N_7448);
xor U10429 (N_10429,N_6354,N_6327);
and U10430 (N_10430,N_6648,N_6567);
or U10431 (N_10431,N_8792,N_6888);
nand U10432 (N_10432,N_8641,N_8461);
nor U10433 (N_10433,N_8375,N_7242);
and U10434 (N_10434,N_6911,N_8651);
nand U10435 (N_10435,N_6763,N_8998);
nand U10436 (N_10436,N_6823,N_8555);
or U10437 (N_10437,N_8004,N_6100);
nor U10438 (N_10438,N_7315,N_8902);
and U10439 (N_10439,N_7012,N_8408);
nor U10440 (N_10440,N_8246,N_7076);
nor U10441 (N_10441,N_7341,N_7278);
nor U10442 (N_10442,N_8423,N_6086);
nor U10443 (N_10443,N_8662,N_7103);
or U10444 (N_10444,N_6095,N_7007);
or U10445 (N_10445,N_7991,N_6847);
xor U10446 (N_10446,N_6865,N_7404);
and U10447 (N_10447,N_8604,N_7800);
or U10448 (N_10448,N_7475,N_8067);
nor U10449 (N_10449,N_6204,N_6416);
nand U10450 (N_10450,N_7335,N_6526);
nand U10451 (N_10451,N_6050,N_6626);
nor U10452 (N_10452,N_6049,N_8632);
and U10453 (N_10453,N_6723,N_7892);
and U10454 (N_10454,N_8775,N_8893);
nand U10455 (N_10455,N_6339,N_8494);
and U10456 (N_10456,N_6927,N_8072);
and U10457 (N_10457,N_8258,N_8854);
nand U10458 (N_10458,N_7623,N_7986);
or U10459 (N_10459,N_6619,N_7375);
nand U10460 (N_10460,N_6438,N_7175);
or U10461 (N_10461,N_7817,N_6298);
nor U10462 (N_10462,N_6399,N_8276);
or U10463 (N_10463,N_8345,N_6143);
xnor U10464 (N_10464,N_6496,N_8370);
or U10465 (N_10465,N_6542,N_7925);
or U10466 (N_10466,N_6972,N_6080);
nor U10467 (N_10467,N_7930,N_8284);
nand U10468 (N_10468,N_6930,N_8495);
or U10469 (N_10469,N_7147,N_7099);
and U10470 (N_10470,N_6638,N_8789);
nand U10471 (N_10471,N_7383,N_7757);
or U10472 (N_10472,N_6431,N_8942);
and U10473 (N_10473,N_6923,N_6932);
and U10474 (N_10474,N_7508,N_8213);
nor U10475 (N_10475,N_8153,N_7206);
nand U10476 (N_10476,N_6584,N_8045);
or U10477 (N_10477,N_8214,N_8395);
or U10478 (N_10478,N_7352,N_7226);
and U10479 (N_10479,N_6528,N_7903);
xor U10480 (N_10480,N_7387,N_6715);
nor U10481 (N_10481,N_6640,N_8394);
xnor U10482 (N_10482,N_8939,N_6309);
and U10483 (N_10483,N_7093,N_6016);
and U10484 (N_10484,N_8504,N_7742);
and U10485 (N_10485,N_6070,N_7814);
or U10486 (N_10486,N_6316,N_6423);
xnor U10487 (N_10487,N_6557,N_6353);
or U10488 (N_10488,N_7505,N_8068);
nand U10489 (N_10489,N_8668,N_6579);
or U10490 (N_10490,N_7847,N_8291);
and U10491 (N_10491,N_7714,N_6094);
and U10492 (N_10492,N_8337,N_8958);
or U10493 (N_10493,N_6974,N_6834);
or U10494 (N_10494,N_7056,N_8550);
and U10495 (N_10495,N_7217,N_8936);
xnor U10496 (N_10496,N_6229,N_6511);
nand U10497 (N_10497,N_6045,N_7506);
xnor U10498 (N_10498,N_7299,N_8810);
xor U10499 (N_10499,N_7490,N_8259);
nand U10500 (N_10500,N_6581,N_8165);
or U10501 (N_10501,N_8267,N_8420);
nor U10502 (N_10502,N_6813,N_7304);
xor U10503 (N_10503,N_8935,N_8548);
nor U10504 (N_10504,N_6270,N_8787);
or U10505 (N_10505,N_7313,N_6676);
and U10506 (N_10506,N_6422,N_6915);
xor U10507 (N_10507,N_6495,N_6546);
nand U10508 (N_10508,N_6145,N_7051);
nand U10509 (N_10509,N_8282,N_7954);
and U10510 (N_10510,N_6352,N_6228);
xor U10511 (N_10511,N_6140,N_8227);
and U10512 (N_10512,N_8652,N_6241);
nand U10513 (N_10513,N_6647,N_8321);
and U10514 (N_10514,N_8601,N_6542);
xnor U10515 (N_10515,N_8375,N_8845);
xor U10516 (N_10516,N_8325,N_7580);
xor U10517 (N_10517,N_8546,N_6855);
xnor U10518 (N_10518,N_6838,N_6998);
and U10519 (N_10519,N_6560,N_8863);
or U10520 (N_10520,N_7105,N_7725);
and U10521 (N_10521,N_7864,N_6970);
nand U10522 (N_10522,N_6864,N_7195);
nor U10523 (N_10523,N_8235,N_8344);
nor U10524 (N_10524,N_8907,N_6818);
and U10525 (N_10525,N_8214,N_7559);
xor U10526 (N_10526,N_7830,N_8601);
xnor U10527 (N_10527,N_7471,N_8940);
xor U10528 (N_10528,N_7317,N_6874);
nand U10529 (N_10529,N_8338,N_8834);
nand U10530 (N_10530,N_8021,N_6095);
or U10531 (N_10531,N_8881,N_8348);
and U10532 (N_10532,N_6305,N_6509);
nor U10533 (N_10533,N_8097,N_7187);
nor U10534 (N_10534,N_8754,N_7164);
nand U10535 (N_10535,N_8470,N_7615);
xor U10536 (N_10536,N_8750,N_7931);
xnor U10537 (N_10537,N_6955,N_8957);
nor U10538 (N_10538,N_6224,N_8938);
nand U10539 (N_10539,N_6112,N_8440);
nand U10540 (N_10540,N_8502,N_7411);
and U10541 (N_10541,N_7275,N_8900);
and U10542 (N_10542,N_6139,N_8492);
or U10543 (N_10543,N_6798,N_6864);
nor U10544 (N_10544,N_8000,N_6763);
or U10545 (N_10545,N_7239,N_8159);
nor U10546 (N_10546,N_8818,N_8315);
nand U10547 (N_10547,N_8653,N_6766);
nand U10548 (N_10548,N_7594,N_6792);
and U10549 (N_10549,N_6730,N_7455);
or U10550 (N_10550,N_8441,N_8601);
xnor U10551 (N_10551,N_6225,N_6860);
nor U10552 (N_10552,N_6666,N_8913);
nand U10553 (N_10553,N_6950,N_8388);
nand U10554 (N_10554,N_7913,N_7859);
nor U10555 (N_10555,N_6658,N_8329);
nand U10556 (N_10556,N_7991,N_6121);
or U10557 (N_10557,N_6225,N_7153);
or U10558 (N_10558,N_8448,N_8513);
nor U10559 (N_10559,N_6627,N_7208);
nand U10560 (N_10560,N_8692,N_7333);
or U10561 (N_10561,N_8096,N_7405);
or U10562 (N_10562,N_7909,N_7986);
or U10563 (N_10563,N_6234,N_7805);
xnor U10564 (N_10564,N_8641,N_8597);
nor U10565 (N_10565,N_7261,N_6198);
nor U10566 (N_10566,N_6614,N_7729);
xor U10567 (N_10567,N_6836,N_7650);
or U10568 (N_10568,N_7568,N_6143);
or U10569 (N_10569,N_7966,N_8420);
or U10570 (N_10570,N_6045,N_8574);
or U10571 (N_10571,N_8991,N_6371);
and U10572 (N_10572,N_8459,N_8656);
xnor U10573 (N_10573,N_7103,N_6216);
and U10574 (N_10574,N_7107,N_8816);
xor U10575 (N_10575,N_8351,N_7948);
xnor U10576 (N_10576,N_8360,N_8759);
and U10577 (N_10577,N_7150,N_6847);
and U10578 (N_10578,N_7239,N_7730);
nand U10579 (N_10579,N_8102,N_6659);
xor U10580 (N_10580,N_6883,N_8149);
and U10581 (N_10581,N_6421,N_7836);
and U10582 (N_10582,N_6828,N_7709);
and U10583 (N_10583,N_7436,N_8610);
xnor U10584 (N_10584,N_6009,N_6168);
xnor U10585 (N_10585,N_8291,N_6443);
xor U10586 (N_10586,N_8847,N_8457);
or U10587 (N_10587,N_6893,N_7444);
and U10588 (N_10588,N_7187,N_8208);
xor U10589 (N_10589,N_6848,N_7437);
nor U10590 (N_10590,N_6772,N_8683);
nand U10591 (N_10591,N_6629,N_7056);
nand U10592 (N_10592,N_7037,N_6541);
or U10593 (N_10593,N_8840,N_7318);
xnor U10594 (N_10594,N_7005,N_6619);
nor U10595 (N_10595,N_7426,N_7447);
and U10596 (N_10596,N_8801,N_6828);
nor U10597 (N_10597,N_7415,N_7797);
or U10598 (N_10598,N_7049,N_7558);
nand U10599 (N_10599,N_6080,N_6441);
or U10600 (N_10600,N_7254,N_7979);
xor U10601 (N_10601,N_6721,N_8584);
xor U10602 (N_10602,N_7645,N_8879);
xor U10603 (N_10603,N_7771,N_6908);
xor U10604 (N_10604,N_7146,N_6104);
nor U10605 (N_10605,N_7241,N_8614);
and U10606 (N_10606,N_6180,N_7640);
xor U10607 (N_10607,N_6819,N_8632);
or U10608 (N_10608,N_7081,N_7773);
and U10609 (N_10609,N_8574,N_8754);
xnor U10610 (N_10610,N_7106,N_6152);
or U10611 (N_10611,N_6538,N_7590);
xor U10612 (N_10612,N_7188,N_8797);
or U10613 (N_10613,N_7835,N_7655);
nand U10614 (N_10614,N_8229,N_6509);
nor U10615 (N_10615,N_8613,N_6848);
nor U10616 (N_10616,N_6049,N_8991);
nand U10617 (N_10617,N_7747,N_6886);
and U10618 (N_10618,N_6861,N_7021);
and U10619 (N_10619,N_6634,N_6705);
nor U10620 (N_10620,N_8211,N_7758);
xnor U10621 (N_10621,N_6875,N_7387);
and U10622 (N_10622,N_7923,N_8172);
or U10623 (N_10623,N_8272,N_7649);
nor U10624 (N_10624,N_8852,N_8554);
nor U10625 (N_10625,N_8454,N_7470);
or U10626 (N_10626,N_7978,N_8074);
or U10627 (N_10627,N_8799,N_6317);
nor U10628 (N_10628,N_6460,N_6244);
nor U10629 (N_10629,N_6827,N_8455);
and U10630 (N_10630,N_7172,N_8131);
or U10631 (N_10631,N_7363,N_6737);
and U10632 (N_10632,N_7126,N_7076);
and U10633 (N_10633,N_6147,N_7063);
or U10634 (N_10634,N_6339,N_7057);
xnor U10635 (N_10635,N_8843,N_8320);
nand U10636 (N_10636,N_8665,N_7118);
xnor U10637 (N_10637,N_8995,N_8969);
and U10638 (N_10638,N_7426,N_8044);
or U10639 (N_10639,N_7336,N_8163);
and U10640 (N_10640,N_8219,N_7065);
nand U10641 (N_10641,N_7205,N_7920);
nand U10642 (N_10642,N_7467,N_7925);
xor U10643 (N_10643,N_7930,N_7448);
and U10644 (N_10644,N_6738,N_6929);
nor U10645 (N_10645,N_6464,N_6963);
and U10646 (N_10646,N_8602,N_6520);
xnor U10647 (N_10647,N_8498,N_8949);
or U10648 (N_10648,N_7217,N_7676);
or U10649 (N_10649,N_6870,N_8601);
nor U10650 (N_10650,N_6362,N_8604);
or U10651 (N_10651,N_8536,N_7715);
and U10652 (N_10652,N_7630,N_7724);
or U10653 (N_10653,N_8535,N_6837);
and U10654 (N_10654,N_7360,N_7188);
nand U10655 (N_10655,N_7284,N_6787);
nor U10656 (N_10656,N_7267,N_7193);
or U10657 (N_10657,N_8362,N_7122);
xnor U10658 (N_10658,N_8765,N_8940);
and U10659 (N_10659,N_6359,N_6642);
or U10660 (N_10660,N_8976,N_6948);
and U10661 (N_10661,N_6334,N_7751);
nand U10662 (N_10662,N_8380,N_7519);
and U10663 (N_10663,N_7790,N_7518);
xor U10664 (N_10664,N_8279,N_8155);
and U10665 (N_10665,N_6773,N_8585);
and U10666 (N_10666,N_7560,N_6891);
and U10667 (N_10667,N_7162,N_8848);
or U10668 (N_10668,N_7101,N_8153);
or U10669 (N_10669,N_7323,N_7215);
nand U10670 (N_10670,N_8207,N_7591);
nor U10671 (N_10671,N_8411,N_6931);
nand U10672 (N_10672,N_7459,N_8138);
or U10673 (N_10673,N_8252,N_7071);
nand U10674 (N_10674,N_6370,N_6260);
nand U10675 (N_10675,N_8526,N_8342);
and U10676 (N_10676,N_8182,N_6915);
nor U10677 (N_10677,N_8030,N_6714);
and U10678 (N_10678,N_7136,N_7633);
and U10679 (N_10679,N_7139,N_6925);
xnor U10680 (N_10680,N_8118,N_8237);
or U10681 (N_10681,N_7121,N_7832);
nor U10682 (N_10682,N_6734,N_6992);
nor U10683 (N_10683,N_6181,N_7154);
xor U10684 (N_10684,N_8668,N_6364);
or U10685 (N_10685,N_6103,N_8130);
and U10686 (N_10686,N_7161,N_7677);
nand U10687 (N_10687,N_6989,N_8652);
nor U10688 (N_10688,N_7556,N_8441);
and U10689 (N_10689,N_8345,N_6428);
nor U10690 (N_10690,N_8591,N_8063);
nor U10691 (N_10691,N_8192,N_6884);
nor U10692 (N_10692,N_6179,N_7501);
nand U10693 (N_10693,N_8916,N_8827);
xnor U10694 (N_10694,N_6789,N_8843);
nor U10695 (N_10695,N_7035,N_8419);
nor U10696 (N_10696,N_6897,N_8757);
nand U10697 (N_10697,N_6885,N_8943);
nor U10698 (N_10698,N_8223,N_7656);
xor U10699 (N_10699,N_6923,N_7102);
and U10700 (N_10700,N_6379,N_8498);
or U10701 (N_10701,N_8424,N_6550);
or U10702 (N_10702,N_7401,N_7021);
xor U10703 (N_10703,N_7486,N_8724);
or U10704 (N_10704,N_6613,N_8688);
and U10705 (N_10705,N_8751,N_7105);
nor U10706 (N_10706,N_6779,N_7525);
nand U10707 (N_10707,N_6440,N_7747);
or U10708 (N_10708,N_7568,N_8678);
xor U10709 (N_10709,N_8286,N_7686);
or U10710 (N_10710,N_6811,N_8633);
nand U10711 (N_10711,N_7926,N_6184);
nor U10712 (N_10712,N_7182,N_8175);
or U10713 (N_10713,N_6218,N_8731);
or U10714 (N_10714,N_6022,N_7716);
nand U10715 (N_10715,N_7887,N_8886);
and U10716 (N_10716,N_8364,N_6503);
nor U10717 (N_10717,N_7246,N_6759);
xnor U10718 (N_10718,N_8233,N_8449);
or U10719 (N_10719,N_6179,N_6263);
nor U10720 (N_10720,N_6721,N_6592);
and U10721 (N_10721,N_7731,N_6564);
nand U10722 (N_10722,N_7041,N_8404);
or U10723 (N_10723,N_8906,N_7043);
xnor U10724 (N_10724,N_7281,N_6172);
and U10725 (N_10725,N_7384,N_6490);
and U10726 (N_10726,N_6773,N_7655);
xnor U10727 (N_10727,N_7303,N_8433);
and U10728 (N_10728,N_6773,N_8291);
nand U10729 (N_10729,N_8237,N_6861);
or U10730 (N_10730,N_8293,N_8168);
nor U10731 (N_10731,N_6157,N_7778);
nand U10732 (N_10732,N_8226,N_7488);
nor U10733 (N_10733,N_6787,N_6574);
xor U10734 (N_10734,N_6612,N_7997);
and U10735 (N_10735,N_7034,N_6735);
and U10736 (N_10736,N_7301,N_8744);
xor U10737 (N_10737,N_8147,N_8241);
and U10738 (N_10738,N_6299,N_6724);
and U10739 (N_10739,N_6242,N_6211);
or U10740 (N_10740,N_8153,N_7237);
and U10741 (N_10741,N_8248,N_7405);
or U10742 (N_10742,N_7406,N_6874);
or U10743 (N_10743,N_7138,N_7924);
and U10744 (N_10744,N_7750,N_6732);
nor U10745 (N_10745,N_7533,N_7669);
or U10746 (N_10746,N_6730,N_7957);
or U10747 (N_10747,N_6861,N_6517);
or U10748 (N_10748,N_8839,N_8564);
xor U10749 (N_10749,N_7684,N_7043);
and U10750 (N_10750,N_7359,N_8916);
nand U10751 (N_10751,N_6706,N_8418);
xnor U10752 (N_10752,N_8365,N_8103);
nand U10753 (N_10753,N_6878,N_6041);
xnor U10754 (N_10754,N_7297,N_8511);
xor U10755 (N_10755,N_8109,N_7851);
nor U10756 (N_10756,N_7118,N_7944);
nor U10757 (N_10757,N_6529,N_8970);
and U10758 (N_10758,N_8790,N_7883);
nand U10759 (N_10759,N_7228,N_7234);
nand U10760 (N_10760,N_8937,N_7210);
xnor U10761 (N_10761,N_6508,N_8560);
and U10762 (N_10762,N_7748,N_7899);
nand U10763 (N_10763,N_7362,N_7688);
xnor U10764 (N_10764,N_8189,N_6965);
and U10765 (N_10765,N_8884,N_6891);
xor U10766 (N_10766,N_7945,N_8908);
xnor U10767 (N_10767,N_8743,N_8700);
or U10768 (N_10768,N_8633,N_6441);
nand U10769 (N_10769,N_8639,N_7101);
and U10770 (N_10770,N_7258,N_8108);
xnor U10771 (N_10771,N_7907,N_6850);
xor U10772 (N_10772,N_8158,N_6799);
nand U10773 (N_10773,N_6784,N_8248);
xnor U10774 (N_10774,N_8605,N_7852);
nand U10775 (N_10775,N_6877,N_8421);
xnor U10776 (N_10776,N_8650,N_6095);
xnor U10777 (N_10777,N_7117,N_6008);
nor U10778 (N_10778,N_7216,N_6503);
nor U10779 (N_10779,N_6751,N_8517);
and U10780 (N_10780,N_6083,N_6985);
and U10781 (N_10781,N_7363,N_8908);
xnor U10782 (N_10782,N_8529,N_6613);
nand U10783 (N_10783,N_7555,N_8481);
nand U10784 (N_10784,N_8940,N_7881);
and U10785 (N_10785,N_7469,N_7682);
nand U10786 (N_10786,N_6127,N_8506);
or U10787 (N_10787,N_8739,N_6977);
nor U10788 (N_10788,N_7590,N_7713);
or U10789 (N_10789,N_8356,N_7326);
xnor U10790 (N_10790,N_8994,N_7116);
nand U10791 (N_10791,N_7571,N_7474);
nand U10792 (N_10792,N_8129,N_8351);
nand U10793 (N_10793,N_6492,N_7588);
nand U10794 (N_10794,N_8290,N_8489);
nand U10795 (N_10795,N_6873,N_7352);
nor U10796 (N_10796,N_6975,N_7684);
nand U10797 (N_10797,N_8519,N_8564);
nand U10798 (N_10798,N_6894,N_8629);
nor U10799 (N_10799,N_8799,N_6732);
nor U10800 (N_10800,N_8261,N_8977);
or U10801 (N_10801,N_7916,N_6214);
and U10802 (N_10802,N_6829,N_6748);
nor U10803 (N_10803,N_6745,N_7394);
or U10804 (N_10804,N_8362,N_7007);
xnor U10805 (N_10805,N_6288,N_6292);
xnor U10806 (N_10806,N_8360,N_7980);
and U10807 (N_10807,N_6213,N_8418);
xor U10808 (N_10808,N_7330,N_6945);
nor U10809 (N_10809,N_6084,N_6970);
and U10810 (N_10810,N_7042,N_7068);
nor U10811 (N_10811,N_7353,N_6507);
nor U10812 (N_10812,N_6942,N_8490);
nand U10813 (N_10813,N_7764,N_6396);
and U10814 (N_10814,N_6056,N_7180);
or U10815 (N_10815,N_6135,N_6827);
xnor U10816 (N_10816,N_6296,N_8974);
xor U10817 (N_10817,N_7888,N_7874);
nand U10818 (N_10818,N_6416,N_7447);
or U10819 (N_10819,N_6430,N_6890);
or U10820 (N_10820,N_8872,N_8610);
xor U10821 (N_10821,N_6251,N_7167);
or U10822 (N_10822,N_7983,N_6915);
nand U10823 (N_10823,N_7660,N_8530);
or U10824 (N_10824,N_8560,N_8994);
or U10825 (N_10825,N_6108,N_7144);
and U10826 (N_10826,N_8303,N_8820);
nand U10827 (N_10827,N_8571,N_8017);
nor U10828 (N_10828,N_6845,N_6996);
and U10829 (N_10829,N_6745,N_8984);
and U10830 (N_10830,N_8476,N_7369);
or U10831 (N_10831,N_6960,N_6587);
or U10832 (N_10832,N_7687,N_7854);
and U10833 (N_10833,N_6127,N_8801);
nor U10834 (N_10834,N_8814,N_7318);
nor U10835 (N_10835,N_7162,N_7386);
or U10836 (N_10836,N_6371,N_6481);
nand U10837 (N_10837,N_7362,N_6868);
nor U10838 (N_10838,N_7099,N_6522);
nor U10839 (N_10839,N_8526,N_7221);
or U10840 (N_10840,N_8389,N_7562);
xor U10841 (N_10841,N_7954,N_7723);
or U10842 (N_10842,N_8744,N_6730);
or U10843 (N_10843,N_6216,N_6636);
and U10844 (N_10844,N_6483,N_7580);
xor U10845 (N_10845,N_7381,N_7316);
nor U10846 (N_10846,N_6319,N_8043);
xor U10847 (N_10847,N_7192,N_7891);
nor U10848 (N_10848,N_6395,N_7080);
nand U10849 (N_10849,N_6353,N_6926);
or U10850 (N_10850,N_6058,N_7790);
nand U10851 (N_10851,N_8610,N_8726);
nor U10852 (N_10852,N_7868,N_7670);
or U10853 (N_10853,N_7184,N_8247);
nor U10854 (N_10854,N_6953,N_6807);
xor U10855 (N_10855,N_7351,N_6109);
nor U10856 (N_10856,N_8870,N_8758);
nand U10857 (N_10857,N_7819,N_7066);
and U10858 (N_10858,N_8984,N_8238);
or U10859 (N_10859,N_7984,N_6328);
nand U10860 (N_10860,N_8842,N_7143);
xor U10861 (N_10861,N_8626,N_8428);
xor U10862 (N_10862,N_8914,N_6560);
nand U10863 (N_10863,N_7292,N_8033);
or U10864 (N_10864,N_8137,N_6155);
nor U10865 (N_10865,N_6254,N_7389);
and U10866 (N_10866,N_7432,N_7591);
xnor U10867 (N_10867,N_8920,N_6336);
nand U10868 (N_10868,N_6686,N_6513);
xor U10869 (N_10869,N_8657,N_7775);
and U10870 (N_10870,N_6584,N_8397);
and U10871 (N_10871,N_7761,N_7701);
nand U10872 (N_10872,N_7100,N_8215);
and U10873 (N_10873,N_7382,N_7659);
and U10874 (N_10874,N_7180,N_6567);
nand U10875 (N_10875,N_6533,N_7678);
or U10876 (N_10876,N_6913,N_7742);
or U10877 (N_10877,N_8265,N_7841);
nor U10878 (N_10878,N_6058,N_7189);
nor U10879 (N_10879,N_8791,N_7552);
and U10880 (N_10880,N_6773,N_7739);
nand U10881 (N_10881,N_6446,N_6691);
nor U10882 (N_10882,N_8248,N_7870);
nor U10883 (N_10883,N_8637,N_8097);
nand U10884 (N_10884,N_7427,N_6790);
nor U10885 (N_10885,N_8811,N_6432);
xnor U10886 (N_10886,N_7572,N_7387);
or U10887 (N_10887,N_8659,N_8529);
nor U10888 (N_10888,N_6798,N_6673);
nand U10889 (N_10889,N_6638,N_6469);
nor U10890 (N_10890,N_6430,N_6987);
xnor U10891 (N_10891,N_8367,N_6032);
xnor U10892 (N_10892,N_6349,N_7793);
or U10893 (N_10893,N_7594,N_6851);
or U10894 (N_10894,N_8796,N_8372);
nor U10895 (N_10895,N_8789,N_6613);
xor U10896 (N_10896,N_7408,N_6947);
nor U10897 (N_10897,N_7546,N_6168);
nor U10898 (N_10898,N_7610,N_7633);
xor U10899 (N_10899,N_7012,N_8410);
and U10900 (N_10900,N_6846,N_6574);
or U10901 (N_10901,N_6340,N_6240);
nand U10902 (N_10902,N_6348,N_8177);
xnor U10903 (N_10903,N_8611,N_6073);
xor U10904 (N_10904,N_6555,N_7270);
nand U10905 (N_10905,N_8805,N_8210);
and U10906 (N_10906,N_7954,N_7238);
and U10907 (N_10907,N_6257,N_6186);
or U10908 (N_10908,N_8686,N_7651);
or U10909 (N_10909,N_7087,N_7632);
nor U10910 (N_10910,N_8220,N_8406);
nor U10911 (N_10911,N_7927,N_6699);
or U10912 (N_10912,N_8029,N_6057);
and U10913 (N_10913,N_8931,N_7580);
nor U10914 (N_10914,N_7943,N_8228);
nand U10915 (N_10915,N_6145,N_8961);
and U10916 (N_10916,N_6827,N_6748);
or U10917 (N_10917,N_7138,N_8872);
nor U10918 (N_10918,N_6684,N_6465);
nand U10919 (N_10919,N_8092,N_8412);
xnor U10920 (N_10920,N_7511,N_7239);
nor U10921 (N_10921,N_6168,N_7753);
xor U10922 (N_10922,N_7891,N_8853);
nand U10923 (N_10923,N_7714,N_7711);
or U10924 (N_10924,N_8864,N_6015);
and U10925 (N_10925,N_7094,N_6295);
or U10926 (N_10926,N_7090,N_8932);
or U10927 (N_10927,N_6121,N_7539);
xnor U10928 (N_10928,N_6632,N_6916);
nor U10929 (N_10929,N_8554,N_6411);
and U10930 (N_10930,N_7319,N_6922);
and U10931 (N_10931,N_8159,N_6356);
and U10932 (N_10932,N_8862,N_6567);
xnor U10933 (N_10933,N_7641,N_7962);
and U10934 (N_10934,N_6291,N_7192);
or U10935 (N_10935,N_8145,N_6506);
or U10936 (N_10936,N_8306,N_7449);
xnor U10937 (N_10937,N_8812,N_6291);
xor U10938 (N_10938,N_8425,N_7628);
nor U10939 (N_10939,N_8753,N_8185);
xor U10940 (N_10940,N_7644,N_7088);
and U10941 (N_10941,N_8701,N_6456);
xor U10942 (N_10942,N_7486,N_7852);
and U10943 (N_10943,N_7964,N_7242);
or U10944 (N_10944,N_8829,N_6331);
nand U10945 (N_10945,N_8669,N_7875);
nor U10946 (N_10946,N_6135,N_8726);
nand U10947 (N_10947,N_8511,N_8930);
and U10948 (N_10948,N_7040,N_8536);
nor U10949 (N_10949,N_8555,N_6328);
nor U10950 (N_10950,N_8757,N_8684);
nand U10951 (N_10951,N_8258,N_7258);
or U10952 (N_10952,N_6614,N_8076);
and U10953 (N_10953,N_6544,N_6182);
xor U10954 (N_10954,N_7026,N_7709);
nor U10955 (N_10955,N_8548,N_6121);
nor U10956 (N_10956,N_6175,N_6646);
xor U10957 (N_10957,N_8264,N_6990);
xor U10958 (N_10958,N_8669,N_7780);
nand U10959 (N_10959,N_6467,N_6419);
nor U10960 (N_10960,N_7533,N_6113);
or U10961 (N_10961,N_7615,N_6104);
and U10962 (N_10962,N_6087,N_7769);
nor U10963 (N_10963,N_7564,N_6938);
nor U10964 (N_10964,N_6126,N_7775);
and U10965 (N_10965,N_7422,N_6085);
or U10966 (N_10966,N_8797,N_6618);
or U10967 (N_10967,N_8473,N_8250);
and U10968 (N_10968,N_6556,N_7973);
nand U10969 (N_10969,N_6286,N_6493);
and U10970 (N_10970,N_8054,N_8608);
nor U10971 (N_10971,N_6053,N_7321);
and U10972 (N_10972,N_6940,N_7759);
or U10973 (N_10973,N_6767,N_6233);
and U10974 (N_10974,N_6652,N_7423);
or U10975 (N_10975,N_8112,N_7695);
and U10976 (N_10976,N_6635,N_7384);
and U10977 (N_10977,N_8881,N_6404);
xor U10978 (N_10978,N_8659,N_8974);
xor U10979 (N_10979,N_8839,N_8535);
or U10980 (N_10980,N_6188,N_7093);
nor U10981 (N_10981,N_6603,N_7912);
and U10982 (N_10982,N_8230,N_6739);
or U10983 (N_10983,N_6711,N_7328);
nor U10984 (N_10984,N_7741,N_7263);
or U10985 (N_10985,N_7170,N_7141);
xnor U10986 (N_10986,N_7039,N_7484);
and U10987 (N_10987,N_6094,N_6726);
nor U10988 (N_10988,N_7127,N_7612);
nand U10989 (N_10989,N_7227,N_6469);
nor U10990 (N_10990,N_6068,N_8756);
and U10991 (N_10991,N_7351,N_8545);
xor U10992 (N_10992,N_6459,N_8721);
or U10993 (N_10993,N_6015,N_6121);
or U10994 (N_10994,N_6123,N_7602);
xor U10995 (N_10995,N_7206,N_8328);
nor U10996 (N_10996,N_6648,N_6403);
xor U10997 (N_10997,N_7414,N_6394);
nand U10998 (N_10998,N_6267,N_7613);
xor U10999 (N_10999,N_7196,N_7541);
nor U11000 (N_11000,N_6623,N_7142);
xnor U11001 (N_11001,N_6135,N_8311);
nand U11002 (N_11002,N_8265,N_7394);
and U11003 (N_11003,N_7390,N_8154);
xor U11004 (N_11004,N_8016,N_7381);
nand U11005 (N_11005,N_7434,N_8554);
nor U11006 (N_11006,N_6298,N_7023);
or U11007 (N_11007,N_6849,N_7738);
and U11008 (N_11008,N_8004,N_8692);
nand U11009 (N_11009,N_7715,N_6025);
nand U11010 (N_11010,N_8769,N_7605);
or U11011 (N_11011,N_6939,N_8108);
nand U11012 (N_11012,N_7802,N_7815);
or U11013 (N_11013,N_7701,N_7986);
nand U11014 (N_11014,N_8118,N_8516);
and U11015 (N_11015,N_6387,N_8609);
and U11016 (N_11016,N_6881,N_6764);
xnor U11017 (N_11017,N_6337,N_6671);
nor U11018 (N_11018,N_8555,N_7572);
nor U11019 (N_11019,N_6794,N_6772);
or U11020 (N_11020,N_8397,N_7412);
and U11021 (N_11021,N_7999,N_8457);
and U11022 (N_11022,N_7125,N_6988);
xor U11023 (N_11023,N_6501,N_8559);
or U11024 (N_11024,N_8856,N_8703);
nand U11025 (N_11025,N_8975,N_8551);
nor U11026 (N_11026,N_7261,N_8996);
nor U11027 (N_11027,N_6641,N_8932);
nor U11028 (N_11028,N_6451,N_7867);
and U11029 (N_11029,N_7113,N_6468);
xnor U11030 (N_11030,N_6326,N_7989);
or U11031 (N_11031,N_7915,N_8329);
and U11032 (N_11032,N_6715,N_6878);
or U11033 (N_11033,N_6180,N_8076);
xor U11034 (N_11034,N_8398,N_6832);
or U11035 (N_11035,N_6678,N_6631);
or U11036 (N_11036,N_6502,N_6694);
nor U11037 (N_11037,N_8486,N_8974);
or U11038 (N_11038,N_8856,N_8380);
nor U11039 (N_11039,N_7672,N_7968);
xor U11040 (N_11040,N_7795,N_8155);
nor U11041 (N_11041,N_8002,N_8058);
and U11042 (N_11042,N_6149,N_6511);
nand U11043 (N_11043,N_8615,N_7035);
nor U11044 (N_11044,N_6123,N_8414);
and U11045 (N_11045,N_6248,N_6725);
nor U11046 (N_11046,N_6386,N_8919);
and U11047 (N_11047,N_7211,N_6129);
nor U11048 (N_11048,N_6522,N_6719);
nand U11049 (N_11049,N_8851,N_6507);
or U11050 (N_11050,N_6732,N_8332);
nor U11051 (N_11051,N_6890,N_8999);
xnor U11052 (N_11052,N_6862,N_8950);
xor U11053 (N_11053,N_6514,N_8236);
and U11054 (N_11054,N_7655,N_7366);
and U11055 (N_11055,N_7970,N_8793);
nand U11056 (N_11056,N_6509,N_6034);
or U11057 (N_11057,N_6417,N_8179);
xor U11058 (N_11058,N_6769,N_6088);
xor U11059 (N_11059,N_7562,N_6336);
or U11060 (N_11060,N_6408,N_6926);
or U11061 (N_11061,N_6543,N_7484);
nand U11062 (N_11062,N_8910,N_6867);
and U11063 (N_11063,N_7139,N_7642);
nor U11064 (N_11064,N_8671,N_6860);
or U11065 (N_11065,N_7647,N_7442);
xnor U11066 (N_11066,N_8840,N_6641);
nand U11067 (N_11067,N_7155,N_6801);
or U11068 (N_11068,N_7186,N_8385);
nor U11069 (N_11069,N_7792,N_7996);
or U11070 (N_11070,N_6814,N_7275);
nand U11071 (N_11071,N_8943,N_6225);
xnor U11072 (N_11072,N_8651,N_7032);
nor U11073 (N_11073,N_8538,N_8574);
nand U11074 (N_11074,N_8296,N_6798);
xnor U11075 (N_11075,N_7422,N_7160);
and U11076 (N_11076,N_6350,N_7822);
xnor U11077 (N_11077,N_6533,N_8521);
or U11078 (N_11078,N_8662,N_6153);
and U11079 (N_11079,N_7666,N_6213);
or U11080 (N_11080,N_8510,N_8340);
or U11081 (N_11081,N_8582,N_7562);
xor U11082 (N_11082,N_7516,N_8260);
or U11083 (N_11083,N_7329,N_8190);
and U11084 (N_11084,N_6017,N_8707);
and U11085 (N_11085,N_7375,N_7420);
or U11086 (N_11086,N_7720,N_8964);
or U11087 (N_11087,N_6694,N_7237);
xnor U11088 (N_11088,N_6778,N_7843);
xor U11089 (N_11089,N_8939,N_6004);
nor U11090 (N_11090,N_7905,N_6888);
xnor U11091 (N_11091,N_7261,N_7661);
nor U11092 (N_11092,N_7907,N_7411);
and U11093 (N_11093,N_7864,N_6421);
and U11094 (N_11094,N_6023,N_8133);
and U11095 (N_11095,N_8637,N_8278);
or U11096 (N_11096,N_8963,N_6434);
and U11097 (N_11097,N_7510,N_6302);
xnor U11098 (N_11098,N_6479,N_8196);
or U11099 (N_11099,N_7950,N_7524);
nor U11100 (N_11100,N_8767,N_6582);
nor U11101 (N_11101,N_7189,N_6867);
and U11102 (N_11102,N_7898,N_7717);
or U11103 (N_11103,N_8787,N_6934);
and U11104 (N_11104,N_6206,N_7489);
xnor U11105 (N_11105,N_6528,N_7144);
nand U11106 (N_11106,N_7138,N_6129);
and U11107 (N_11107,N_6843,N_7243);
nand U11108 (N_11108,N_6335,N_6938);
nor U11109 (N_11109,N_8293,N_6003);
xor U11110 (N_11110,N_6191,N_7549);
or U11111 (N_11111,N_7966,N_6401);
nor U11112 (N_11112,N_8921,N_6956);
and U11113 (N_11113,N_8861,N_6636);
and U11114 (N_11114,N_8114,N_7839);
nor U11115 (N_11115,N_6736,N_6647);
nor U11116 (N_11116,N_7837,N_8163);
or U11117 (N_11117,N_6077,N_8690);
nand U11118 (N_11118,N_6580,N_7266);
and U11119 (N_11119,N_7346,N_6319);
or U11120 (N_11120,N_6880,N_8238);
xnor U11121 (N_11121,N_8035,N_6991);
nor U11122 (N_11122,N_7242,N_8819);
nand U11123 (N_11123,N_8718,N_8901);
xor U11124 (N_11124,N_6681,N_6630);
xnor U11125 (N_11125,N_6923,N_8194);
and U11126 (N_11126,N_8365,N_6798);
and U11127 (N_11127,N_6868,N_8008);
nor U11128 (N_11128,N_7779,N_6079);
and U11129 (N_11129,N_8410,N_6405);
or U11130 (N_11130,N_6973,N_8146);
or U11131 (N_11131,N_8331,N_8453);
xnor U11132 (N_11132,N_6676,N_8028);
xnor U11133 (N_11133,N_8188,N_7525);
and U11134 (N_11134,N_8876,N_6006);
and U11135 (N_11135,N_7439,N_8989);
nand U11136 (N_11136,N_8384,N_7695);
nor U11137 (N_11137,N_7168,N_7251);
xnor U11138 (N_11138,N_6826,N_8591);
xnor U11139 (N_11139,N_8322,N_7608);
nand U11140 (N_11140,N_6028,N_7957);
nor U11141 (N_11141,N_8583,N_6544);
and U11142 (N_11142,N_6425,N_6039);
or U11143 (N_11143,N_6198,N_8924);
and U11144 (N_11144,N_6580,N_7471);
or U11145 (N_11145,N_8143,N_8321);
xnor U11146 (N_11146,N_6115,N_7369);
or U11147 (N_11147,N_6777,N_8148);
nor U11148 (N_11148,N_8544,N_8324);
and U11149 (N_11149,N_6129,N_6158);
nor U11150 (N_11150,N_7697,N_7637);
and U11151 (N_11151,N_7952,N_7383);
nand U11152 (N_11152,N_8490,N_7317);
nand U11153 (N_11153,N_6338,N_6716);
and U11154 (N_11154,N_6826,N_6066);
nand U11155 (N_11155,N_6264,N_8734);
nor U11156 (N_11156,N_6477,N_7140);
nor U11157 (N_11157,N_8453,N_8027);
or U11158 (N_11158,N_8541,N_6997);
and U11159 (N_11159,N_7267,N_7877);
and U11160 (N_11160,N_7071,N_8736);
nand U11161 (N_11161,N_6331,N_8800);
nor U11162 (N_11162,N_8549,N_8323);
nand U11163 (N_11163,N_6835,N_8564);
or U11164 (N_11164,N_8580,N_8842);
nor U11165 (N_11165,N_6434,N_8478);
nand U11166 (N_11166,N_8957,N_8346);
and U11167 (N_11167,N_7060,N_8266);
or U11168 (N_11168,N_8690,N_7472);
or U11169 (N_11169,N_8484,N_6547);
and U11170 (N_11170,N_8153,N_7325);
nand U11171 (N_11171,N_6278,N_8529);
nand U11172 (N_11172,N_7654,N_6131);
xnor U11173 (N_11173,N_7087,N_7004);
or U11174 (N_11174,N_8889,N_7272);
and U11175 (N_11175,N_6229,N_7329);
or U11176 (N_11176,N_6998,N_6457);
nand U11177 (N_11177,N_7416,N_7353);
xor U11178 (N_11178,N_7369,N_7338);
or U11179 (N_11179,N_7575,N_7057);
and U11180 (N_11180,N_6733,N_8534);
nand U11181 (N_11181,N_6179,N_6724);
xnor U11182 (N_11182,N_7354,N_6289);
xor U11183 (N_11183,N_6897,N_8917);
and U11184 (N_11184,N_7077,N_6804);
nand U11185 (N_11185,N_7897,N_7832);
xor U11186 (N_11186,N_8691,N_6128);
nor U11187 (N_11187,N_7679,N_8864);
nor U11188 (N_11188,N_8424,N_7774);
nor U11189 (N_11189,N_8180,N_6302);
nor U11190 (N_11190,N_8122,N_8945);
nand U11191 (N_11191,N_7134,N_8704);
xor U11192 (N_11192,N_8734,N_7259);
nor U11193 (N_11193,N_7034,N_7144);
xor U11194 (N_11194,N_8357,N_8646);
nor U11195 (N_11195,N_6329,N_7758);
xor U11196 (N_11196,N_6587,N_8650);
nor U11197 (N_11197,N_8336,N_8464);
or U11198 (N_11198,N_8722,N_7582);
or U11199 (N_11199,N_6278,N_8003);
and U11200 (N_11200,N_6779,N_7560);
and U11201 (N_11201,N_8426,N_7711);
or U11202 (N_11202,N_6403,N_8963);
nand U11203 (N_11203,N_6524,N_6640);
nor U11204 (N_11204,N_8239,N_7312);
or U11205 (N_11205,N_8366,N_8538);
nand U11206 (N_11206,N_7664,N_8210);
xor U11207 (N_11207,N_6943,N_7655);
nor U11208 (N_11208,N_6903,N_7714);
and U11209 (N_11209,N_6228,N_7475);
and U11210 (N_11210,N_7865,N_6303);
xor U11211 (N_11211,N_7465,N_7508);
or U11212 (N_11212,N_6586,N_7364);
and U11213 (N_11213,N_8081,N_6200);
nor U11214 (N_11214,N_8499,N_7546);
xor U11215 (N_11215,N_7538,N_8702);
xnor U11216 (N_11216,N_7147,N_6504);
xor U11217 (N_11217,N_7568,N_7113);
nor U11218 (N_11218,N_8592,N_8503);
nor U11219 (N_11219,N_7661,N_8471);
nand U11220 (N_11220,N_6105,N_7953);
and U11221 (N_11221,N_8922,N_8871);
or U11222 (N_11222,N_6315,N_6862);
or U11223 (N_11223,N_8851,N_7303);
nand U11224 (N_11224,N_8364,N_7134);
nor U11225 (N_11225,N_6475,N_7786);
or U11226 (N_11226,N_8258,N_6658);
nor U11227 (N_11227,N_7447,N_7979);
or U11228 (N_11228,N_7988,N_6175);
nor U11229 (N_11229,N_6339,N_6796);
xor U11230 (N_11230,N_7283,N_7138);
nand U11231 (N_11231,N_8302,N_8823);
xnor U11232 (N_11232,N_7797,N_8137);
or U11233 (N_11233,N_6581,N_7808);
xor U11234 (N_11234,N_8175,N_6242);
and U11235 (N_11235,N_7828,N_7727);
nand U11236 (N_11236,N_8478,N_8626);
and U11237 (N_11237,N_6077,N_7332);
and U11238 (N_11238,N_7099,N_7110);
nand U11239 (N_11239,N_8187,N_6618);
xnor U11240 (N_11240,N_7210,N_6610);
or U11241 (N_11241,N_6892,N_6634);
nor U11242 (N_11242,N_8795,N_7553);
xnor U11243 (N_11243,N_8324,N_7103);
or U11244 (N_11244,N_7729,N_6302);
and U11245 (N_11245,N_7147,N_6618);
nor U11246 (N_11246,N_8749,N_6357);
nand U11247 (N_11247,N_8925,N_8495);
nor U11248 (N_11248,N_6525,N_8060);
and U11249 (N_11249,N_8895,N_8790);
or U11250 (N_11250,N_7547,N_7849);
and U11251 (N_11251,N_8396,N_6551);
and U11252 (N_11252,N_7274,N_7957);
xnor U11253 (N_11253,N_8503,N_8004);
and U11254 (N_11254,N_7639,N_6747);
or U11255 (N_11255,N_7648,N_7244);
or U11256 (N_11256,N_7903,N_8810);
or U11257 (N_11257,N_7041,N_8328);
nand U11258 (N_11258,N_7314,N_6773);
xor U11259 (N_11259,N_7734,N_7669);
nor U11260 (N_11260,N_8525,N_8889);
or U11261 (N_11261,N_8988,N_7735);
xor U11262 (N_11262,N_6939,N_7372);
xnor U11263 (N_11263,N_6123,N_6182);
nand U11264 (N_11264,N_8592,N_6323);
nand U11265 (N_11265,N_6434,N_8967);
and U11266 (N_11266,N_8841,N_7970);
nor U11267 (N_11267,N_8665,N_6977);
and U11268 (N_11268,N_6116,N_7263);
nor U11269 (N_11269,N_8143,N_7326);
xnor U11270 (N_11270,N_7432,N_7092);
xor U11271 (N_11271,N_6461,N_7647);
nand U11272 (N_11272,N_7304,N_8152);
nand U11273 (N_11273,N_7344,N_6392);
xnor U11274 (N_11274,N_7978,N_8629);
or U11275 (N_11275,N_8224,N_6071);
nor U11276 (N_11276,N_7640,N_8993);
or U11277 (N_11277,N_7733,N_8091);
nor U11278 (N_11278,N_7860,N_6587);
or U11279 (N_11279,N_8428,N_7799);
xor U11280 (N_11280,N_7133,N_6940);
or U11281 (N_11281,N_6626,N_7015);
nand U11282 (N_11282,N_7103,N_8541);
and U11283 (N_11283,N_8593,N_6260);
or U11284 (N_11284,N_7093,N_6000);
nor U11285 (N_11285,N_7927,N_6342);
or U11286 (N_11286,N_6133,N_8655);
nor U11287 (N_11287,N_7157,N_6269);
nor U11288 (N_11288,N_6271,N_6661);
or U11289 (N_11289,N_6011,N_7534);
and U11290 (N_11290,N_8412,N_6182);
and U11291 (N_11291,N_6493,N_8490);
nand U11292 (N_11292,N_6079,N_8275);
and U11293 (N_11293,N_8564,N_8050);
and U11294 (N_11294,N_6166,N_8129);
and U11295 (N_11295,N_7759,N_7406);
nor U11296 (N_11296,N_8879,N_7892);
nand U11297 (N_11297,N_8476,N_7086);
or U11298 (N_11298,N_6113,N_8444);
nor U11299 (N_11299,N_6526,N_7089);
nand U11300 (N_11300,N_7783,N_7565);
xor U11301 (N_11301,N_7846,N_8008);
nor U11302 (N_11302,N_7374,N_7206);
nand U11303 (N_11303,N_8630,N_7758);
xor U11304 (N_11304,N_8173,N_6259);
nand U11305 (N_11305,N_6118,N_7450);
or U11306 (N_11306,N_8378,N_6732);
nand U11307 (N_11307,N_8192,N_7137);
nor U11308 (N_11308,N_6407,N_6724);
nor U11309 (N_11309,N_7693,N_8472);
xnor U11310 (N_11310,N_8987,N_7142);
or U11311 (N_11311,N_6074,N_6123);
and U11312 (N_11312,N_7745,N_7135);
nand U11313 (N_11313,N_8248,N_8822);
and U11314 (N_11314,N_7764,N_6884);
or U11315 (N_11315,N_6906,N_6741);
nand U11316 (N_11316,N_8784,N_8586);
xor U11317 (N_11317,N_6255,N_8582);
and U11318 (N_11318,N_6076,N_8466);
or U11319 (N_11319,N_6543,N_7224);
nor U11320 (N_11320,N_6484,N_7635);
and U11321 (N_11321,N_7945,N_6882);
xnor U11322 (N_11322,N_7590,N_6687);
nor U11323 (N_11323,N_8964,N_7592);
nor U11324 (N_11324,N_6582,N_8953);
nor U11325 (N_11325,N_7755,N_6611);
nand U11326 (N_11326,N_7855,N_8319);
and U11327 (N_11327,N_6442,N_7994);
xnor U11328 (N_11328,N_8618,N_6379);
xnor U11329 (N_11329,N_8193,N_7339);
nand U11330 (N_11330,N_6476,N_7218);
or U11331 (N_11331,N_7936,N_8522);
xor U11332 (N_11332,N_8357,N_7920);
and U11333 (N_11333,N_8156,N_7051);
xor U11334 (N_11334,N_6812,N_7602);
or U11335 (N_11335,N_7497,N_6734);
or U11336 (N_11336,N_8559,N_6526);
nand U11337 (N_11337,N_8410,N_7228);
xor U11338 (N_11338,N_6111,N_6806);
nand U11339 (N_11339,N_6029,N_8952);
or U11340 (N_11340,N_8897,N_8877);
nand U11341 (N_11341,N_8195,N_7305);
nand U11342 (N_11342,N_7615,N_7535);
or U11343 (N_11343,N_6907,N_8062);
and U11344 (N_11344,N_8662,N_6934);
xor U11345 (N_11345,N_8639,N_8174);
nand U11346 (N_11346,N_6500,N_8731);
and U11347 (N_11347,N_8153,N_6439);
or U11348 (N_11348,N_7984,N_6796);
or U11349 (N_11349,N_7617,N_7570);
nor U11350 (N_11350,N_6683,N_7952);
nand U11351 (N_11351,N_8246,N_8221);
nand U11352 (N_11352,N_7749,N_7775);
or U11353 (N_11353,N_6372,N_7445);
nor U11354 (N_11354,N_6949,N_8377);
nand U11355 (N_11355,N_8052,N_8474);
or U11356 (N_11356,N_6009,N_8784);
xnor U11357 (N_11357,N_8706,N_8251);
or U11358 (N_11358,N_8499,N_8479);
xor U11359 (N_11359,N_8923,N_6374);
xnor U11360 (N_11360,N_6090,N_6086);
nand U11361 (N_11361,N_6417,N_7546);
nand U11362 (N_11362,N_6253,N_6121);
nor U11363 (N_11363,N_8247,N_8198);
nor U11364 (N_11364,N_6285,N_8097);
nand U11365 (N_11365,N_6796,N_7278);
nand U11366 (N_11366,N_6901,N_6946);
xnor U11367 (N_11367,N_8136,N_8584);
xor U11368 (N_11368,N_7287,N_8708);
or U11369 (N_11369,N_8898,N_8961);
and U11370 (N_11370,N_6740,N_7995);
or U11371 (N_11371,N_7232,N_8105);
nor U11372 (N_11372,N_8205,N_8383);
and U11373 (N_11373,N_8333,N_8341);
nor U11374 (N_11374,N_6885,N_6147);
xor U11375 (N_11375,N_6000,N_7650);
or U11376 (N_11376,N_8611,N_8274);
xor U11377 (N_11377,N_7945,N_7949);
and U11378 (N_11378,N_7296,N_7658);
and U11379 (N_11379,N_7724,N_7670);
nand U11380 (N_11380,N_8723,N_8147);
nand U11381 (N_11381,N_8858,N_6613);
or U11382 (N_11382,N_7066,N_8594);
nand U11383 (N_11383,N_6830,N_6946);
and U11384 (N_11384,N_7168,N_7390);
or U11385 (N_11385,N_7569,N_7026);
or U11386 (N_11386,N_6961,N_6679);
and U11387 (N_11387,N_6698,N_8111);
nand U11388 (N_11388,N_8335,N_6933);
nor U11389 (N_11389,N_7116,N_6500);
and U11390 (N_11390,N_7743,N_7262);
nand U11391 (N_11391,N_8034,N_6062);
or U11392 (N_11392,N_8615,N_8359);
or U11393 (N_11393,N_7944,N_6183);
and U11394 (N_11394,N_7969,N_6909);
xor U11395 (N_11395,N_6692,N_8038);
or U11396 (N_11396,N_7238,N_7416);
or U11397 (N_11397,N_6752,N_6352);
or U11398 (N_11398,N_8892,N_7253);
nor U11399 (N_11399,N_8049,N_8286);
or U11400 (N_11400,N_6194,N_7108);
nor U11401 (N_11401,N_7630,N_8618);
nand U11402 (N_11402,N_7668,N_6495);
nor U11403 (N_11403,N_6929,N_7796);
nor U11404 (N_11404,N_8880,N_6967);
nand U11405 (N_11405,N_7600,N_7688);
nor U11406 (N_11406,N_8731,N_7087);
or U11407 (N_11407,N_6957,N_6522);
and U11408 (N_11408,N_8333,N_8161);
and U11409 (N_11409,N_7170,N_8173);
xnor U11410 (N_11410,N_8859,N_8720);
nor U11411 (N_11411,N_6566,N_8374);
and U11412 (N_11412,N_8679,N_7164);
xor U11413 (N_11413,N_8889,N_6107);
xnor U11414 (N_11414,N_7003,N_6322);
nand U11415 (N_11415,N_8939,N_7922);
xor U11416 (N_11416,N_7802,N_8293);
and U11417 (N_11417,N_7147,N_8814);
or U11418 (N_11418,N_6274,N_6224);
nand U11419 (N_11419,N_8990,N_8258);
nor U11420 (N_11420,N_8130,N_7275);
xor U11421 (N_11421,N_6511,N_7896);
xnor U11422 (N_11422,N_6881,N_7109);
and U11423 (N_11423,N_6141,N_6300);
and U11424 (N_11424,N_7488,N_7627);
nand U11425 (N_11425,N_7721,N_6592);
nand U11426 (N_11426,N_8774,N_6540);
nor U11427 (N_11427,N_8987,N_6499);
nand U11428 (N_11428,N_7642,N_6667);
or U11429 (N_11429,N_7495,N_8885);
and U11430 (N_11430,N_7712,N_6754);
xor U11431 (N_11431,N_6532,N_7064);
xnor U11432 (N_11432,N_7258,N_8970);
nand U11433 (N_11433,N_8096,N_6279);
nor U11434 (N_11434,N_6995,N_7801);
nor U11435 (N_11435,N_7677,N_8868);
nand U11436 (N_11436,N_7424,N_8593);
or U11437 (N_11437,N_7561,N_8820);
nor U11438 (N_11438,N_8351,N_8070);
nand U11439 (N_11439,N_8845,N_6530);
nor U11440 (N_11440,N_6019,N_6266);
or U11441 (N_11441,N_7154,N_7839);
nand U11442 (N_11442,N_8659,N_6018);
xnor U11443 (N_11443,N_7768,N_6889);
or U11444 (N_11444,N_8893,N_6592);
nor U11445 (N_11445,N_6338,N_8698);
and U11446 (N_11446,N_7156,N_6284);
xnor U11447 (N_11447,N_7559,N_8612);
xor U11448 (N_11448,N_6507,N_6894);
and U11449 (N_11449,N_7736,N_6770);
and U11450 (N_11450,N_7731,N_8304);
xnor U11451 (N_11451,N_6224,N_8780);
or U11452 (N_11452,N_8748,N_6309);
nand U11453 (N_11453,N_8942,N_6910);
nand U11454 (N_11454,N_7648,N_6181);
or U11455 (N_11455,N_8983,N_8236);
and U11456 (N_11456,N_7999,N_7876);
or U11457 (N_11457,N_8663,N_7542);
and U11458 (N_11458,N_6001,N_6599);
or U11459 (N_11459,N_8967,N_7882);
nor U11460 (N_11460,N_8807,N_8852);
and U11461 (N_11461,N_7023,N_7785);
and U11462 (N_11462,N_6332,N_8597);
xor U11463 (N_11463,N_6331,N_6155);
nand U11464 (N_11464,N_8657,N_6391);
xnor U11465 (N_11465,N_7581,N_6009);
xnor U11466 (N_11466,N_8994,N_8688);
nand U11467 (N_11467,N_7627,N_8466);
or U11468 (N_11468,N_7535,N_7552);
and U11469 (N_11469,N_8213,N_8913);
and U11470 (N_11470,N_7965,N_6886);
xnor U11471 (N_11471,N_8708,N_7503);
nand U11472 (N_11472,N_6708,N_7129);
and U11473 (N_11473,N_8439,N_7469);
and U11474 (N_11474,N_6105,N_8558);
or U11475 (N_11475,N_7282,N_7891);
nor U11476 (N_11476,N_8800,N_6348);
xnor U11477 (N_11477,N_6116,N_6616);
xor U11478 (N_11478,N_6842,N_8455);
xnor U11479 (N_11479,N_7842,N_8429);
nand U11480 (N_11480,N_8246,N_8203);
nor U11481 (N_11481,N_7320,N_7264);
nand U11482 (N_11482,N_8055,N_7154);
xor U11483 (N_11483,N_8876,N_6363);
and U11484 (N_11484,N_6960,N_7623);
or U11485 (N_11485,N_6699,N_7276);
nand U11486 (N_11486,N_7637,N_6925);
xnor U11487 (N_11487,N_8229,N_6164);
and U11488 (N_11488,N_6580,N_7143);
or U11489 (N_11489,N_6484,N_8714);
or U11490 (N_11490,N_6413,N_6685);
or U11491 (N_11491,N_8694,N_8753);
or U11492 (N_11492,N_6656,N_8385);
xnor U11493 (N_11493,N_7258,N_8833);
or U11494 (N_11494,N_7387,N_8787);
or U11495 (N_11495,N_7262,N_6197);
nand U11496 (N_11496,N_6577,N_8802);
and U11497 (N_11497,N_6187,N_6889);
or U11498 (N_11498,N_6880,N_7055);
xnor U11499 (N_11499,N_8076,N_8758);
xor U11500 (N_11500,N_7364,N_6782);
xnor U11501 (N_11501,N_6578,N_6779);
and U11502 (N_11502,N_8330,N_6247);
or U11503 (N_11503,N_6390,N_6135);
xor U11504 (N_11504,N_7069,N_7394);
xor U11505 (N_11505,N_8370,N_7952);
nand U11506 (N_11506,N_7351,N_6059);
or U11507 (N_11507,N_6709,N_8237);
or U11508 (N_11508,N_8789,N_7690);
or U11509 (N_11509,N_6743,N_7203);
nand U11510 (N_11510,N_7014,N_7828);
nand U11511 (N_11511,N_6055,N_6095);
or U11512 (N_11512,N_6373,N_8168);
xnor U11513 (N_11513,N_8777,N_8914);
nor U11514 (N_11514,N_6814,N_8159);
and U11515 (N_11515,N_8399,N_8429);
nand U11516 (N_11516,N_6032,N_7728);
and U11517 (N_11517,N_8533,N_6503);
xor U11518 (N_11518,N_7557,N_8563);
nor U11519 (N_11519,N_7891,N_6527);
or U11520 (N_11520,N_8204,N_6639);
xor U11521 (N_11521,N_6342,N_8464);
nand U11522 (N_11522,N_6675,N_8448);
and U11523 (N_11523,N_6018,N_8848);
xnor U11524 (N_11524,N_7998,N_8726);
and U11525 (N_11525,N_7401,N_7843);
xor U11526 (N_11526,N_8120,N_7178);
xnor U11527 (N_11527,N_7806,N_6430);
xor U11528 (N_11528,N_6278,N_6595);
and U11529 (N_11529,N_8489,N_6448);
xor U11530 (N_11530,N_8291,N_7185);
xor U11531 (N_11531,N_7924,N_6513);
xor U11532 (N_11532,N_6117,N_8603);
and U11533 (N_11533,N_7182,N_8504);
or U11534 (N_11534,N_6951,N_6816);
xnor U11535 (N_11535,N_7099,N_8298);
nand U11536 (N_11536,N_7833,N_7738);
or U11537 (N_11537,N_8859,N_6171);
xnor U11538 (N_11538,N_8552,N_8795);
or U11539 (N_11539,N_8879,N_7343);
or U11540 (N_11540,N_7187,N_7648);
xnor U11541 (N_11541,N_8110,N_7811);
and U11542 (N_11542,N_6105,N_8862);
and U11543 (N_11543,N_6406,N_8886);
nand U11544 (N_11544,N_8602,N_7583);
and U11545 (N_11545,N_8921,N_7909);
or U11546 (N_11546,N_7093,N_7386);
or U11547 (N_11547,N_8133,N_6349);
and U11548 (N_11548,N_6825,N_8073);
nor U11549 (N_11549,N_7332,N_6196);
nor U11550 (N_11550,N_8186,N_6258);
or U11551 (N_11551,N_7614,N_6437);
or U11552 (N_11552,N_8962,N_6424);
and U11553 (N_11553,N_8727,N_7769);
and U11554 (N_11554,N_7055,N_6296);
and U11555 (N_11555,N_8670,N_7248);
nor U11556 (N_11556,N_7505,N_6145);
nand U11557 (N_11557,N_7214,N_7516);
or U11558 (N_11558,N_6359,N_8531);
and U11559 (N_11559,N_6952,N_8995);
and U11560 (N_11560,N_7750,N_8452);
xnor U11561 (N_11561,N_8609,N_6350);
and U11562 (N_11562,N_8586,N_8150);
nand U11563 (N_11563,N_7517,N_8313);
nand U11564 (N_11564,N_8930,N_8488);
or U11565 (N_11565,N_7182,N_8467);
xor U11566 (N_11566,N_6798,N_6105);
nand U11567 (N_11567,N_6259,N_6300);
nand U11568 (N_11568,N_7492,N_7547);
nor U11569 (N_11569,N_6153,N_8362);
nand U11570 (N_11570,N_6543,N_8755);
nor U11571 (N_11571,N_7055,N_7940);
nor U11572 (N_11572,N_6432,N_8198);
and U11573 (N_11573,N_6864,N_8938);
or U11574 (N_11574,N_6297,N_6248);
nor U11575 (N_11575,N_6589,N_7437);
xnor U11576 (N_11576,N_6882,N_7927);
nand U11577 (N_11577,N_8970,N_6023);
nor U11578 (N_11578,N_6250,N_8773);
nor U11579 (N_11579,N_8371,N_6873);
xnor U11580 (N_11580,N_6736,N_7101);
xor U11581 (N_11581,N_8641,N_8103);
and U11582 (N_11582,N_7719,N_8583);
xnor U11583 (N_11583,N_8523,N_8480);
and U11584 (N_11584,N_8859,N_6533);
or U11585 (N_11585,N_8807,N_8539);
or U11586 (N_11586,N_8165,N_6996);
nor U11587 (N_11587,N_6067,N_7008);
and U11588 (N_11588,N_8754,N_8162);
and U11589 (N_11589,N_8325,N_8902);
nand U11590 (N_11590,N_8395,N_8697);
xnor U11591 (N_11591,N_7767,N_7464);
or U11592 (N_11592,N_8604,N_6782);
xnor U11593 (N_11593,N_8990,N_6468);
xnor U11594 (N_11594,N_7033,N_6338);
or U11595 (N_11595,N_8897,N_8428);
nor U11596 (N_11596,N_6843,N_6756);
or U11597 (N_11597,N_8243,N_8286);
xnor U11598 (N_11598,N_7663,N_7412);
nor U11599 (N_11599,N_7602,N_7586);
and U11600 (N_11600,N_7991,N_6871);
xor U11601 (N_11601,N_7909,N_8114);
and U11602 (N_11602,N_6189,N_7874);
xnor U11603 (N_11603,N_6756,N_7416);
nor U11604 (N_11604,N_8187,N_8576);
or U11605 (N_11605,N_8329,N_8587);
nand U11606 (N_11606,N_8653,N_6004);
xnor U11607 (N_11607,N_8735,N_7125);
and U11608 (N_11608,N_6931,N_6433);
nor U11609 (N_11609,N_8538,N_7461);
or U11610 (N_11610,N_7621,N_6477);
xnor U11611 (N_11611,N_7840,N_6763);
or U11612 (N_11612,N_6755,N_7059);
and U11613 (N_11613,N_6942,N_6268);
and U11614 (N_11614,N_7507,N_7076);
nand U11615 (N_11615,N_6262,N_6842);
or U11616 (N_11616,N_6830,N_6987);
or U11617 (N_11617,N_8326,N_7909);
nand U11618 (N_11618,N_7215,N_6573);
or U11619 (N_11619,N_6163,N_8913);
and U11620 (N_11620,N_7893,N_7833);
nand U11621 (N_11621,N_7497,N_8559);
and U11622 (N_11622,N_7919,N_8765);
nor U11623 (N_11623,N_6050,N_6662);
xnor U11624 (N_11624,N_8930,N_6009);
xor U11625 (N_11625,N_7978,N_8865);
nand U11626 (N_11626,N_8701,N_8159);
nor U11627 (N_11627,N_8596,N_7074);
nor U11628 (N_11628,N_8098,N_7532);
nand U11629 (N_11629,N_6146,N_7454);
xnor U11630 (N_11630,N_7595,N_8108);
nor U11631 (N_11631,N_8435,N_7181);
and U11632 (N_11632,N_7203,N_6151);
nand U11633 (N_11633,N_7483,N_8964);
xnor U11634 (N_11634,N_6277,N_7251);
or U11635 (N_11635,N_7241,N_7368);
nor U11636 (N_11636,N_7756,N_7686);
xnor U11637 (N_11637,N_6364,N_8113);
xor U11638 (N_11638,N_6962,N_7497);
xnor U11639 (N_11639,N_8700,N_6356);
nand U11640 (N_11640,N_8425,N_6700);
and U11641 (N_11641,N_7397,N_7722);
nor U11642 (N_11642,N_6205,N_8595);
nand U11643 (N_11643,N_7232,N_6523);
and U11644 (N_11644,N_6339,N_7264);
or U11645 (N_11645,N_8287,N_7834);
and U11646 (N_11646,N_8878,N_8942);
nand U11647 (N_11647,N_6996,N_8994);
xnor U11648 (N_11648,N_6239,N_8303);
or U11649 (N_11649,N_8168,N_6572);
nand U11650 (N_11650,N_8954,N_7821);
xor U11651 (N_11651,N_6882,N_8972);
and U11652 (N_11652,N_8318,N_8369);
nand U11653 (N_11653,N_6867,N_7854);
and U11654 (N_11654,N_7540,N_8830);
nand U11655 (N_11655,N_6091,N_8490);
and U11656 (N_11656,N_7167,N_8335);
xnor U11657 (N_11657,N_8143,N_6396);
and U11658 (N_11658,N_8797,N_7608);
xnor U11659 (N_11659,N_8585,N_8237);
nor U11660 (N_11660,N_8668,N_6832);
nand U11661 (N_11661,N_7872,N_7158);
nand U11662 (N_11662,N_7874,N_8778);
and U11663 (N_11663,N_8525,N_6029);
and U11664 (N_11664,N_6043,N_8829);
nand U11665 (N_11665,N_7060,N_6451);
or U11666 (N_11666,N_7580,N_8407);
or U11667 (N_11667,N_8050,N_8804);
nand U11668 (N_11668,N_8655,N_6867);
or U11669 (N_11669,N_8078,N_7121);
and U11670 (N_11670,N_6952,N_7725);
xnor U11671 (N_11671,N_8992,N_6297);
xnor U11672 (N_11672,N_8896,N_6697);
or U11673 (N_11673,N_8040,N_7390);
or U11674 (N_11674,N_7550,N_7181);
xnor U11675 (N_11675,N_7740,N_6548);
and U11676 (N_11676,N_7078,N_6701);
xnor U11677 (N_11677,N_6358,N_7698);
nor U11678 (N_11678,N_8420,N_7447);
nand U11679 (N_11679,N_6733,N_8852);
or U11680 (N_11680,N_8947,N_7140);
nor U11681 (N_11681,N_8330,N_8718);
or U11682 (N_11682,N_7744,N_8004);
xor U11683 (N_11683,N_6172,N_6026);
or U11684 (N_11684,N_8011,N_8967);
nand U11685 (N_11685,N_6356,N_6424);
or U11686 (N_11686,N_8146,N_7687);
nor U11687 (N_11687,N_7708,N_8739);
and U11688 (N_11688,N_8098,N_8944);
or U11689 (N_11689,N_8413,N_7560);
nor U11690 (N_11690,N_8574,N_7468);
nor U11691 (N_11691,N_6489,N_7198);
or U11692 (N_11692,N_7286,N_6221);
nand U11693 (N_11693,N_6158,N_7562);
nand U11694 (N_11694,N_8393,N_8694);
nor U11695 (N_11695,N_6222,N_6471);
or U11696 (N_11696,N_8872,N_8103);
or U11697 (N_11697,N_8107,N_6491);
or U11698 (N_11698,N_8663,N_8417);
nor U11699 (N_11699,N_8528,N_8030);
nor U11700 (N_11700,N_6813,N_8327);
nand U11701 (N_11701,N_8790,N_8824);
and U11702 (N_11702,N_8448,N_6540);
xnor U11703 (N_11703,N_7850,N_6929);
nand U11704 (N_11704,N_7483,N_6047);
or U11705 (N_11705,N_8953,N_7447);
xnor U11706 (N_11706,N_8920,N_6223);
or U11707 (N_11707,N_6745,N_6555);
or U11708 (N_11708,N_6685,N_6811);
nand U11709 (N_11709,N_7087,N_6503);
and U11710 (N_11710,N_7827,N_7377);
or U11711 (N_11711,N_8423,N_6032);
xor U11712 (N_11712,N_6205,N_7483);
and U11713 (N_11713,N_8680,N_6144);
or U11714 (N_11714,N_7568,N_7370);
or U11715 (N_11715,N_8288,N_8725);
nand U11716 (N_11716,N_6047,N_8487);
nor U11717 (N_11717,N_7870,N_6542);
xor U11718 (N_11718,N_7638,N_8090);
or U11719 (N_11719,N_7555,N_7303);
nor U11720 (N_11720,N_7374,N_6370);
or U11721 (N_11721,N_8417,N_7249);
and U11722 (N_11722,N_8386,N_6541);
and U11723 (N_11723,N_6895,N_8980);
xnor U11724 (N_11724,N_7732,N_8083);
or U11725 (N_11725,N_7879,N_8540);
nand U11726 (N_11726,N_7715,N_8687);
nand U11727 (N_11727,N_6920,N_6180);
nand U11728 (N_11728,N_7509,N_6741);
or U11729 (N_11729,N_6956,N_6654);
xor U11730 (N_11730,N_6098,N_6159);
and U11731 (N_11731,N_7673,N_6937);
nor U11732 (N_11732,N_6049,N_8010);
and U11733 (N_11733,N_6911,N_6469);
or U11734 (N_11734,N_6250,N_6987);
nand U11735 (N_11735,N_8161,N_7709);
or U11736 (N_11736,N_8997,N_8517);
or U11737 (N_11737,N_7714,N_7307);
and U11738 (N_11738,N_7136,N_6729);
nand U11739 (N_11739,N_7557,N_7285);
xor U11740 (N_11740,N_6779,N_8358);
xnor U11741 (N_11741,N_8019,N_6537);
xnor U11742 (N_11742,N_8906,N_8072);
nor U11743 (N_11743,N_8975,N_8188);
nand U11744 (N_11744,N_7588,N_8910);
nor U11745 (N_11745,N_7336,N_6038);
or U11746 (N_11746,N_8936,N_6291);
nand U11747 (N_11747,N_7448,N_8093);
nand U11748 (N_11748,N_8576,N_8838);
nor U11749 (N_11749,N_7487,N_7027);
nand U11750 (N_11750,N_8003,N_7234);
xor U11751 (N_11751,N_8162,N_7895);
or U11752 (N_11752,N_7146,N_6502);
and U11753 (N_11753,N_6148,N_8941);
and U11754 (N_11754,N_6061,N_7844);
nor U11755 (N_11755,N_8084,N_8247);
or U11756 (N_11756,N_7965,N_6464);
nor U11757 (N_11757,N_6842,N_8927);
or U11758 (N_11758,N_8263,N_7512);
nor U11759 (N_11759,N_7737,N_7944);
or U11760 (N_11760,N_6135,N_8003);
nor U11761 (N_11761,N_8534,N_6225);
or U11762 (N_11762,N_8762,N_7904);
nand U11763 (N_11763,N_6093,N_6443);
nand U11764 (N_11764,N_7479,N_7073);
nor U11765 (N_11765,N_6361,N_8655);
nand U11766 (N_11766,N_6453,N_8229);
nor U11767 (N_11767,N_7585,N_6945);
or U11768 (N_11768,N_7948,N_6385);
xor U11769 (N_11769,N_7562,N_7282);
xor U11770 (N_11770,N_8579,N_6317);
or U11771 (N_11771,N_7988,N_7576);
and U11772 (N_11772,N_6075,N_6101);
xnor U11773 (N_11773,N_6312,N_8552);
and U11774 (N_11774,N_8111,N_7809);
nand U11775 (N_11775,N_7180,N_6475);
and U11776 (N_11776,N_6968,N_8690);
nor U11777 (N_11777,N_8392,N_6765);
or U11778 (N_11778,N_7241,N_8011);
xnor U11779 (N_11779,N_7684,N_8175);
xor U11780 (N_11780,N_8651,N_8541);
or U11781 (N_11781,N_8917,N_8777);
xnor U11782 (N_11782,N_6069,N_7119);
nand U11783 (N_11783,N_6936,N_7966);
nand U11784 (N_11784,N_8520,N_7712);
nand U11785 (N_11785,N_7465,N_7281);
or U11786 (N_11786,N_8339,N_7533);
xnor U11787 (N_11787,N_6669,N_7856);
xor U11788 (N_11788,N_8041,N_6786);
xnor U11789 (N_11789,N_6581,N_7711);
and U11790 (N_11790,N_6683,N_8507);
or U11791 (N_11791,N_8027,N_6096);
xor U11792 (N_11792,N_8221,N_8916);
xnor U11793 (N_11793,N_7225,N_6453);
xnor U11794 (N_11794,N_7717,N_6718);
or U11795 (N_11795,N_6732,N_6498);
or U11796 (N_11796,N_8587,N_7378);
nand U11797 (N_11797,N_7395,N_6367);
nor U11798 (N_11798,N_7288,N_6495);
xnor U11799 (N_11799,N_7772,N_7079);
and U11800 (N_11800,N_8683,N_8834);
nand U11801 (N_11801,N_8426,N_8162);
nor U11802 (N_11802,N_8451,N_6413);
xnor U11803 (N_11803,N_8622,N_8018);
nor U11804 (N_11804,N_6573,N_7852);
nand U11805 (N_11805,N_8486,N_8993);
xor U11806 (N_11806,N_7217,N_7868);
or U11807 (N_11807,N_6746,N_6876);
or U11808 (N_11808,N_6289,N_8427);
nand U11809 (N_11809,N_6880,N_7301);
or U11810 (N_11810,N_7043,N_8212);
nor U11811 (N_11811,N_8242,N_8194);
and U11812 (N_11812,N_8925,N_6835);
xnor U11813 (N_11813,N_8600,N_7622);
or U11814 (N_11814,N_6651,N_6648);
or U11815 (N_11815,N_7013,N_8699);
nand U11816 (N_11816,N_6307,N_6551);
nand U11817 (N_11817,N_7122,N_8730);
nand U11818 (N_11818,N_8953,N_7687);
nand U11819 (N_11819,N_6114,N_6954);
and U11820 (N_11820,N_6043,N_7236);
xnor U11821 (N_11821,N_6794,N_6354);
nand U11822 (N_11822,N_7902,N_6565);
and U11823 (N_11823,N_6957,N_6412);
or U11824 (N_11824,N_6927,N_6169);
nand U11825 (N_11825,N_6740,N_7774);
nand U11826 (N_11826,N_8546,N_7092);
and U11827 (N_11827,N_6497,N_7202);
and U11828 (N_11828,N_6658,N_7683);
or U11829 (N_11829,N_7761,N_7034);
and U11830 (N_11830,N_7284,N_7766);
nor U11831 (N_11831,N_8610,N_7074);
xor U11832 (N_11832,N_8730,N_7702);
or U11833 (N_11833,N_6389,N_8548);
nand U11834 (N_11834,N_6955,N_6053);
and U11835 (N_11835,N_8641,N_6900);
xor U11836 (N_11836,N_6995,N_6288);
xnor U11837 (N_11837,N_7562,N_7778);
nand U11838 (N_11838,N_6752,N_8470);
nor U11839 (N_11839,N_7982,N_6618);
nor U11840 (N_11840,N_8676,N_8607);
nor U11841 (N_11841,N_7202,N_8468);
nand U11842 (N_11842,N_8554,N_8086);
xor U11843 (N_11843,N_6049,N_8312);
xor U11844 (N_11844,N_7008,N_6807);
nand U11845 (N_11845,N_7381,N_7161);
nand U11846 (N_11846,N_8610,N_6098);
or U11847 (N_11847,N_6001,N_8138);
xor U11848 (N_11848,N_6763,N_8690);
or U11849 (N_11849,N_8882,N_6184);
and U11850 (N_11850,N_6153,N_8344);
and U11851 (N_11851,N_8739,N_6088);
xnor U11852 (N_11852,N_7377,N_6725);
nor U11853 (N_11853,N_6912,N_7273);
or U11854 (N_11854,N_7544,N_8208);
xnor U11855 (N_11855,N_7358,N_6121);
and U11856 (N_11856,N_8616,N_6661);
xnor U11857 (N_11857,N_6184,N_6435);
and U11858 (N_11858,N_7806,N_8651);
nand U11859 (N_11859,N_7114,N_7942);
xnor U11860 (N_11860,N_7228,N_7733);
nor U11861 (N_11861,N_6753,N_6396);
or U11862 (N_11862,N_8462,N_6210);
and U11863 (N_11863,N_8405,N_7007);
nand U11864 (N_11864,N_8659,N_7744);
and U11865 (N_11865,N_6249,N_8443);
or U11866 (N_11866,N_7865,N_8753);
nor U11867 (N_11867,N_8420,N_6721);
nand U11868 (N_11868,N_7368,N_6061);
and U11869 (N_11869,N_8162,N_8763);
and U11870 (N_11870,N_6606,N_6922);
xnor U11871 (N_11871,N_6057,N_8018);
nand U11872 (N_11872,N_8439,N_8989);
nand U11873 (N_11873,N_7687,N_6805);
nand U11874 (N_11874,N_6080,N_6326);
nand U11875 (N_11875,N_8962,N_6711);
and U11876 (N_11876,N_6694,N_8577);
nand U11877 (N_11877,N_8104,N_7858);
xnor U11878 (N_11878,N_8685,N_8818);
nor U11879 (N_11879,N_8075,N_7265);
and U11880 (N_11880,N_7424,N_6995);
nor U11881 (N_11881,N_8645,N_7127);
and U11882 (N_11882,N_6368,N_7963);
xor U11883 (N_11883,N_8557,N_8556);
or U11884 (N_11884,N_7067,N_7783);
or U11885 (N_11885,N_6654,N_6905);
or U11886 (N_11886,N_6858,N_8995);
nand U11887 (N_11887,N_7639,N_6600);
and U11888 (N_11888,N_6324,N_7803);
or U11889 (N_11889,N_7969,N_7014);
nor U11890 (N_11890,N_6898,N_7441);
and U11891 (N_11891,N_8972,N_7625);
xnor U11892 (N_11892,N_7311,N_7149);
or U11893 (N_11893,N_7792,N_7334);
or U11894 (N_11894,N_7199,N_6079);
nand U11895 (N_11895,N_8292,N_8707);
or U11896 (N_11896,N_6632,N_8578);
nand U11897 (N_11897,N_6777,N_7538);
nand U11898 (N_11898,N_7799,N_6075);
or U11899 (N_11899,N_6022,N_7171);
and U11900 (N_11900,N_8263,N_7209);
nor U11901 (N_11901,N_7844,N_7687);
and U11902 (N_11902,N_8867,N_7959);
nand U11903 (N_11903,N_7300,N_6106);
nand U11904 (N_11904,N_7516,N_6699);
nand U11905 (N_11905,N_8358,N_6275);
nor U11906 (N_11906,N_8171,N_8616);
nor U11907 (N_11907,N_7265,N_7433);
nand U11908 (N_11908,N_6047,N_8801);
xnor U11909 (N_11909,N_8492,N_6350);
nand U11910 (N_11910,N_6613,N_8275);
and U11911 (N_11911,N_7364,N_7633);
and U11912 (N_11912,N_7073,N_7087);
or U11913 (N_11913,N_6547,N_6369);
or U11914 (N_11914,N_6335,N_6271);
nor U11915 (N_11915,N_6804,N_7054);
xnor U11916 (N_11916,N_7636,N_7041);
xor U11917 (N_11917,N_7387,N_8235);
nor U11918 (N_11918,N_6294,N_7323);
xnor U11919 (N_11919,N_8205,N_7085);
nand U11920 (N_11920,N_8544,N_6487);
nor U11921 (N_11921,N_7911,N_6310);
or U11922 (N_11922,N_8410,N_6920);
nor U11923 (N_11923,N_8446,N_7252);
or U11924 (N_11924,N_8958,N_6266);
nand U11925 (N_11925,N_6227,N_7165);
nor U11926 (N_11926,N_7575,N_8748);
or U11927 (N_11927,N_7707,N_7731);
and U11928 (N_11928,N_8748,N_6348);
or U11929 (N_11929,N_6850,N_7197);
or U11930 (N_11930,N_7285,N_6443);
nand U11931 (N_11931,N_7985,N_7514);
nand U11932 (N_11932,N_7306,N_6065);
or U11933 (N_11933,N_8468,N_8080);
nand U11934 (N_11934,N_6527,N_8498);
and U11935 (N_11935,N_8418,N_6566);
nand U11936 (N_11936,N_6578,N_8728);
and U11937 (N_11937,N_7115,N_7269);
and U11938 (N_11938,N_6967,N_6653);
or U11939 (N_11939,N_6329,N_6105);
nor U11940 (N_11940,N_7705,N_8459);
or U11941 (N_11941,N_7789,N_6362);
nand U11942 (N_11942,N_6503,N_8440);
nand U11943 (N_11943,N_7704,N_8178);
and U11944 (N_11944,N_8382,N_6255);
xor U11945 (N_11945,N_8985,N_8002);
and U11946 (N_11946,N_7404,N_7276);
and U11947 (N_11947,N_6122,N_7828);
and U11948 (N_11948,N_6411,N_7983);
xor U11949 (N_11949,N_6166,N_6726);
and U11950 (N_11950,N_6718,N_6576);
xor U11951 (N_11951,N_8177,N_8874);
nand U11952 (N_11952,N_8872,N_8854);
or U11953 (N_11953,N_8225,N_7290);
xor U11954 (N_11954,N_7468,N_6037);
or U11955 (N_11955,N_8938,N_8034);
and U11956 (N_11956,N_6149,N_8996);
nand U11957 (N_11957,N_8753,N_6878);
nor U11958 (N_11958,N_6854,N_7137);
nor U11959 (N_11959,N_7793,N_8198);
or U11960 (N_11960,N_8579,N_8774);
and U11961 (N_11961,N_7681,N_8707);
or U11962 (N_11962,N_7638,N_8419);
nand U11963 (N_11963,N_8170,N_8101);
nor U11964 (N_11964,N_8780,N_6348);
and U11965 (N_11965,N_8749,N_8521);
nor U11966 (N_11966,N_6779,N_7708);
nor U11967 (N_11967,N_7544,N_7368);
or U11968 (N_11968,N_6975,N_8257);
nor U11969 (N_11969,N_8272,N_7153);
nor U11970 (N_11970,N_7960,N_7586);
nor U11971 (N_11971,N_7701,N_7311);
or U11972 (N_11972,N_8316,N_8458);
nand U11973 (N_11973,N_8879,N_6356);
xor U11974 (N_11974,N_6213,N_6724);
and U11975 (N_11975,N_8443,N_6264);
and U11976 (N_11976,N_6278,N_6703);
nor U11977 (N_11977,N_8735,N_8279);
and U11978 (N_11978,N_8103,N_7397);
and U11979 (N_11979,N_8916,N_6363);
xnor U11980 (N_11980,N_8997,N_8555);
nor U11981 (N_11981,N_8305,N_6669);
xor U11982 (N_11982,N_8844,N_6234);
xnor U11983 (N_11983,N_6946,N_7826);
nor U11984 (N_11984,N_6936,N_8350);
or U11985 (N_11985,N_6569,N_7303);
nand U11986 (N_11986,N_8929,N_6105);
xnor U11987 (N_11987,N_6628,N_8091);
xnor U11988 (N_11988,N_6511,N_7084);
xnor U11989 (N_11989,N_6541,N_7444);
and U11990 (N_11990,N_6045,N_7968);
or U11991 (N_11991,N_7882,N_7519);
nor U11992 (N_11992,N_7100,N_6046);
xor U11993 (N_11993,N_7164,N_6010);
nand U11994 (N_11994,N_6358,N_8471);
nor U11995 (N_11995,N_7449,N_7388);
nor U11996 (N_11996,N_6301,N_6959);
nor U11997 (N_11997,N_7044,N_7264);
and U11998 (N_11998,N_7332,N_7510);
xnor U11999 (N_11999,N_6715,N_8893);
nor U12000 (N_12000,N_11756,N_9637);
nor U12001 (N_12001,N_10880,N_10247);
or U12002 (N_12002,N_9492,N_9003);
and U12003 (N_12003,N_11163,N_11052);
nor U12004 (N_12004,N_9377,N_11484);
xor U12005 (N_12005,N_11377,N_9677);
or U12006 (N_12006,N_10530,N_10606);
nand U12007 (N_12007,N_11728,N_10084);
nor U12008 (N_12008,N_9005,N_11942);
and U12009 (N_12009,N_10207,N_9487);
and U12010 (N_12010,N_10034,N_9110);
nand U12011 (N_12011,N_10169,N_9892);
or U12012 (N_12012,N_10386,N_11883);
or U12013 (N_12013,N_10324,N_11083);
or U12014 (N_12014,N_9545,N_9127);
and U12015 (N_12015,N_9548,N_11408);
nor U12016 (N_12016,N_10568,N_10409);
or U12017 (N_12017,N_10266,N_10866);
nand U12018 (N_12018,N_11050,N_11240);
nor U12019 (N_12019,N_10987,N_10039);
and U12020 (N_12020,N_9416,N_10674);
or U12021 (N_12021,N_11937,N_11281);
xnor U12022 (N_12022,N_11469,N_9042);
nand U12023 (N_12023,N_10273,N_9237);
nand U12024 (N_12024,N_9336,N_10467);
or U12025 (N_12025,N_10026,N_11591);
and U12026 (N_12026,N_11833,N_10691);
nand U12027 (N_12027,N_9284,N_9413);
or U12028 (N_12028,N_10572,N_9577);
nand U12029 (N_12029,N_11519,N_11238);
and U12030 (N_12030,N_11338,N_9804);
nand U12031 (N_12031,N_9306,N_11021);
nor U12032 (N_12032,N_10718,N_10204);
nand U12033 (N_12033,N_10206,N_11479);
nor U12034 (N_12034,N_9949,N_9040);
nand U12035 (N_12035,N_9950,N_9697);
xor U12036 (N_12036,N_11597,N_10818);
nand U12037 (N_12037,N_10624,N_11721);
and U12038 (N_12038,N_11701,N_11226);
and U12039 (N_12039,N_11569,N_9591);
nor U12040 (N_12040,N_9282,N_11199);
and U12041 (N_12041,N_10844,N_10633);
nor U12042 (N_12042,N_9676,N_9272);
and U12043 (N_12043,N_10146,N_9395);
and U12044 (N_12044,N_10407,N_9995);
nand U12045 (N_12045,N_10942,N_11537);
or U12046 (N_12046,N_11095,N_10177);
nand U12047 (N_12047,N_10198,N_11946);
or U12048 (N_12048,N_9461,N_9497);
and U12049 (N_12049,N_10233,N_9869);
and U12050 (N_12050,N_10044,N_10425);
or U12051 (N_12051,N_10265,N_9467);
xor U12052 (N_12052,N_10412,N_9004);
xnor U12053 (N_12053,N_10411,N_10185);
and U12054 (N_12054,N_11547,N_9787);
nor U12055 (N_12055,N_9552,N_10008);
nand U12056 (N_12056,N_9896,N_11960);
or U12057 (N_12057,N_10500,N_9133);
xor U12058 (N_12058,N_9354,N_10005);
and U12059 (N_12059,N_10330,N_10021);
xor U12060 (N_12060,N_11195,N_11253);
nor U12061 (N_12061,N_9459,N_10676);
xnor U12062 (N_12062,N_10363,N_11657);
or U12063 (N_12063,N_11441,N_9144);
or U12064 (N_12064,N_11840,N_11145);
or U12065 (N_12065,N_9060,N_9939);
and U12066 (N_12066,N_9396,N_9050);
or U12067 (N_12067,N_10344,N_10539);
nand U12068 (N_12068,N_10318,N_9843);
xor U12069 (N_12069,N_9798,N_10968);
nand U12070 (N_12070,N_11636,N_9313);
nand U12071 (N_12071,N_9394,N_10618);
and U12072 (N_12072,N_10751,N_11013);
nor U12073 (N_12073,N_9870,N_10667);
nand U12074 (N_12074,N_11324,N_11455);
nand U12075 (N_12075,N_10499,N_9222);
nand U12076 (N_12076,N_9528,N_11223);
or U12077 (N_12077,N_11466,N_11826);
or U12078 (N_12078,N_11473,N_10444);
and U12079 (N_12079,N_11369,N_9967);
and U12080 (N_12080,N_9737,N_9409);
or U12081 (N_12081,N_10703,N_11637);
and U12082 (N_12082,N_11108,N_9700);
or U12083 (N_12083,N_10393,N_9599);
and U12084 (N_12084,N_10155,N_11036);
and U12085 (N_12085,N_10243,N_9520);
nor U12086 (N_12086,N_9088,N_9605);
and U12087 (N_12087,N_11870,N_11925);
xor U12088 (N_12088,N_10013,N_11702);
and U12089 (N_12089,N_10228,N_11571);
nor U12090 (N_12090,N_10000,N_9542);
xnor U12091 (N_12091,N_9997,N_11898);
nand U12092 (N_12092,N_10404,N_11328);
and U12093 (N_12093,N_9472,N_11385);
nor U12094 (N_12094,N_9634,N_10215);
nand U12095 (N_12095,N_10768,N_10298);
xor U12096 (N_12096,N_11011,N_11995);
and U12097 (N_12097,N_10470,N_11334);
or U12098 (N_12098,N_11517,N_10195);
or U12099 (N_12099,N_11761,N_10834);
nand U12100 (N_12100,N_11081,N_9357);
or U12101 (N_12101,N_9479,N_9859);
nand U12102 (N_12102,N_9549,N_11462);
nand U12103 (N_12103,N_10263,N_11394);
nor U12104 (N_12104,N_9578,N_11184);
nand U12105 (N_12105,N_10682,N_9941);
nand U12106 (N_12106,N_9176,N_10194);
or U12107 (N_12107,N_9688,N_11889);
nand U12108 (N_12108,N_9242,N_11438);
nand U12109 (N_12109,N_9699,N_10496);
and U12110 (N_12110,N_9143,N_11296);
nor U12111 (N_12111,N_11291,N_11370);
xnor U12112 (N_12112,N_11332,N_9275);
or U12113 (N_12113,N_11178,N_9296);
or U12114 (N_12114,N_10153,N_11719);
xor U12115 (N_12115,N_11396,N_10382);
nor U12116 (N_12116,N_10351,N_9830);
nand U12117 (N_12117,N_11677,N_9371);
and U12118 (N_12118,N_11648,N_9048);
and U12119 (N_12119,N_10434,N_10437);
xor U12120 (N_12120,N_10851,N_9214);
or U12121 (N_12121,N_10604,N_9958);
and U12122 (N_12122,N_11235,N_10917);
and U12123 (N_12123,N_10927,N_10174);
and U12124 (N_12124,N_11953,N_10646);
and U12125 (N_12125,N_9126,N_9182);
nand U12126 (N_12126,N_11128,N_11956);
and U12127 (N_12127,N_11232,N_9861);
xor U12128 (N_12128,N_10523,N_9929);
nor U12129 (N_12129,N_9157,N_11373);
or U12130 (N_12130,N_10649,N_11666);
xnor U12131 (N_12131,N_9235,N_9172);
and U12132 (N_12132,N_11687,N_9732);
nor U12133 (N_12133,N_9819,N_10203);
and U12134 (N_12134,N_10037,N_10004);
nand U12135 (N_12135,N_11974,N_10240);
nor U12136 (N_12136,N_9831,N_10454);
or U12137 (N_12137,N_9992,N_10085);
and U12138 (N_12138,N_9072,N_9417);
nand U12139 (N_12139,N_11650,N_9146);
or U12140 (N_12140,N_9428,N_9298);
nand U12141 (N_12141,N_11678,N_9671);
nor U12142 (N_12142,N_10657,N_11839);
or U12143 (N_12143,N_11938,N_11550);
nand U12144 (N_12144,N_9116,N_10669);
nor U12145 (N_12145,N_9855,N_9132);
or U12146 (N_12146,N_11825,N_11808);
or U12147 (N_12147,N_10133,N_9419);
nor U12148 (N_12148,N_9691,N_9736);
and U12149 (N_12149,N_9293,N_10850);
and U12150 (N_12150,N_9962,N_11543);
and U12151 (N_12151,N_11325,N_10733);
and U12152 (N_12152,N_10424,N_10126);
or U12153 (N_12153,N_11776,N_9833);
or U12154 (N_12154,N_10287,N_9550);
nor U12155 (N_12155,N_10841,N_9277);
or U12156 (N_12156,N_11759,N_9233);
nand U12157 (N_12157,N_11186,N_11963);
and U12158 (N_12158,N_9669,N_10871);
and U12159 (N_12159,N_11002,N_9337);
nor U12160 (N_12160,N_9627,N_10800);
nand U12161 (N_12161,N_10257,N_10825);
nor U12162 (N_12162,N_10217,N_9572);
or U12163 (N_12163,N_9083,N_11010);
or U12164 (N_12164,N_10782,N_9231);
or U12165 (N_12165,N_10867,N_10612);
nor U12166 (N_12166,N_10309,N_10060);
or U12167 (N_12167,N_9759,N_10190);
xnor U12168 (N_12168,N_11765,N_11945);
and U12169 (N_12169,N_9940,N_11748);
xor U12170 (N_12170,N_9292,N_10744);
nor U12171 (N_12171,N_9478,N_10959);
nand U12172 (N_12172,N_11802,N_10459);
xnor U12173 (N_12173,N_9730,N_9103);
nor U12174 (N_12174,N_9886,N_11255);
nand U12175 (N_12175,N_9837,N_9925);
or U12176 (N_12176,N_10954,N_10801);
and U12177 (N_12177,N_9903,N_9529);
nor U12178 (N_12178,N_9376,N_9164);
xor U12179 (N_12179,N_9712,N_10750);
or U12180 (N_12180,N_10123,N_9809);
and U12181 (N_12181,N_11426,N_10130);
and U12182 (N_12182,N_11201,N_11400);
xnor U12183 (N_12183,N_11490,N_10541);
nand U12184 (N_12184,N_10717,N_11922);
and U12185 (N_12185,N_10684,N_10585);
and U12186 (N_12186,N_9476,N_9986);
nand U12187 (N_12187,N_11156,N_10946);
xor U12188 (N_12188,N_11869,N_11451);
nand U12189 (N_12189,N_11770,N_9425);
or U12190 (N_12190,N_9551,N_9918);
xnor U12191 (N_12191,N_11531,N_9738);
and U12192 (N_12192,N_9801,N_9555);
xor U12193 (N_12193,N_11985,N_11881);
xor U12194 (N_12194,N_9255,N_9288);
and U12195 (N_12195,N_11970,N_9025);
xnor U12196 (N_12196,N_11935,N_10574);
xor U12197 (N_12197,N_11848,N_11845);
nand U12198 (N_12198,N_10565,N_11135);
and U12199 (N_12199,N_9573,N_9885);
nand U12200 (N_12200,N_9215,N_9031);
nand U12201 (N_12201,N_11535,N_9734);
nor U12202 (N_12202,N_10975,N_11061);
nand U12203 (N_12203,N_9104,N_11605);
nand U12204 (N_12204,N_11056,N_11769);
or U12205 (N_12205,N_9266,N_10930);
and U12206 (N_12206,N_10161,N_11307);
xnor U12207 (N_12207,N_10697,N_10030);
nand U12208 (N_12208,N_10028,N_11518);
or U12209 (N_12209,N_11185,N_9561);
and U12210 (N_12210,N_11006,N_9657);
and U12211 (N_12211,N_11358,N_9991);
nand U12212 (N_12212,N_10753,N_11754);
or U12213 (N_12213,N_11936,N_11198);
nor U12214 (N_12214,N_10051,N_9366);
or U12215 (N_12215,N_9244,N_10367);
or U12216 (N_12216,N_11681,N_9335);
xnor U12217 (N_12217,N_11810,N_9068);
xor U12218 (N_12218,N_10116,N_9727);
nor U12219 (N_12219,N_9097,N_9444);
nor U12220 (N_12220,N_9808,N_10889);
or U12221 (N_12221,N_10197,N_10908);
nor U12222 (N_12222,N_9169,N_11387);
nor U12223 (N_12223,N_10708,N_9364);
xnor U12224 (N_12224,N_10741,N_11801);
nand U12225 (N_12225,N_11794,N_11117);
nand U12226 (N_12226,N_9204,N_11697);
nor U12227 (N_12227,N_10128,N_9447);
xnor U12228 (N_12228,N_10003,N_10352);
xor U12229 (N_12229,N_9020,N_10808);
or U12230 (N_12230,N_9027,N_11376);
xor U12231 (N_12231,N_10857,N_9350);
xnor U12232 (N_12232,N_9230,N_10507);
or U12233 (N_12233,N_10977,N_10230);
or U12234 (N_12234,N_10339,N_9443);
or U12235 (N_12235,N_9841,N_9483);
or U12236 (N_12236,N_10898,N_11587);
nor U12237 (N_12237,N_9674,N_11835);
or U12238 (N_12238,N_11532,N_11092);
nor U12239 (N_12239,N_11818,N_11094);
nand U12240 (N_12240,N_9516,N_9867);
nor U12241 (N_12241,N_10734,N_11347);
xnor U12242 (N_12242,N_10902,N_10370);
xor U12243 (N_12243,N_10780,N_11402);
and U12244 (N_12244,N_9239,N_9713);
or U12245 (N_12245,N_11897,N_11608);
nand U12246 (N_12246,N_11622,N_10790);
xor U12247 (N_12247,N_11330,N_9912);
nor U12248 (N_12248,N_9557,N_10487);
xnor U12249 (N_12249,N_10432,N_10192);
xor U12250 (N_12250,N_11667,N_9032);
or U12251 (N_12251,N_9465,N_11318);
or U12252 (N_12252,N_10599,N_11814);
and U12253 (N_12253,N_9408,N_9778);
and U12254 (N_12254,N_10639,N_9315);
nor U12255 (N_12255,N_11965,N_10609);
and U12256 (N_12256,N_10570,N_11724);
xor U12257 (N_12257,N_9217,N_10304);
xor U12258 (N_12258,N_11924,N_11523);
nor U12259 (N_12259,N_9802,N_9562);
or U12260 (N_12260,N_11862,N_10332);
xnor U12261 (N_12261,N_9576,N_11626);
or U12262 (N_12262,N_9094,N_10290);
and U12263 (N_12263,N_9565,N_10985);
xor U12264 (N_12264,N_11691,N_11866);
and U12265 (N_12265,N_9347,N_11422);
or U12266 (N_12266,N_10251,N_9763);
xor U12267 (N_12267,N_9630,N_10635);
nand U12268 (N_12268,N_10057,N_11110);
nor U12269 (N_12269,N_10219,N_11066);
xnor U12270 (N_12270,N_9165,N_11404);
or U12271 (N_12271,N_11350,N_11023);
or U12272 (N_12272,N_10100,N_11431);
and U12273 (N_12273,N_10664,N_11111);
or U12274 (N_12274,N_10286,N_11796);
and U12275 (N_12275,N_11046,N_10439);
or U12276 (N_12276,N_10474,N_11355);
nor U12277 (N_12277,N_10179,N_10678);
xnor U12278 (N_12278,N_9075,N_11189);
nor U12279 (N_12279,N_11661,N_10774);
nand U12280 (N_12280,N_11986,N_10157);
nand U12281 (N_12281,N_10885,N_10694);
nand U12282 (N_12282,N_10456,N_10278);
nor U12283 (N_12283,N_11710,N_11785);
or U12284 (N_12284,N_10865,N_10956);
or U12285 (N_12285,N_10242,N_10491);
xor U12286 (N_12286,N_11244,N_10214);
and U12287 (N_12287,N_11913,N_10299);
and U12288 (N_12288,N_11266,N_10595);
or U12289 (N_12289,N_9571,N_9036);
nor U12290 (N_12290,N_10879,N_10271);
or U12291 (N_12291,N_10868,N_11017);
nand U12292 (N_12292,N_10244,N_9829);
nor U12293 (N_12293,N_9754,N_9325);
and U12294 (N_12294,N_11811,N_11236);
or U12295 (N_12295,N_9302,N_9742);
or U12296 (N_12296,N_11300,N_9806);
or U12297 (N_12297,N_9744,N_11208);
nand U12298 (N_12298,N_10325,N_11509);
and U12299 (N_12299,N_11288,N_9570);
nor U12300 (N_12300,N_11638,N_11498);
nand U12301 (N_12301,N_10521,N_10756);
and U12302 (N_12302,N_11948,N_10275);
or U12303 (N_12303,N_9342,N_11653);
nand U12304 (N_12304,N_11912,N_9010);
and U12305 (N_12305,N_11161,N_10566);
or U12306 (N_12306,N_10118,N_10593);
xnor U12307 (N_12307,N_10001,N_9089);
nor U12308 (N_12308,N_10069,N_11842);
and U12309 (N_12309,N_10605,N_10952);
nand U12310 (N_12310,N_11162,N_10912);
nand U12311 (N_12311,N_9439,N_11193);
xor U12312 (N_12312,N_10261,N_11410);
nand U12313 (N_12313,N_11172,N_10073);
and U12314 (N_12314,N_10607,N_10732);
nor U12315 (N_12315,N_11939,N_10740);
nand U12316 (N_12316,N_9460,N_10969);
or U12317 (N_12317,N_10476,N_10279);
and U12318 (N_12318,N_11289,N_9748);
and U12319 (N_12319,N_9948,N_9910);
and U12320 (N_12320,N_10110,N_9877);
and U12321 (N_12321,N_11767,N_11560);
nand U12322 (N_12322,N_10571,N_10150);
and U12323 (N_12323,N_9085,N_11405);
nand U12324 (N_12324,N_10443,N_10302);
or U12325 (N_12325,N_10763,N_11690);
nor U12326 (N_12326,N_10726,N_11106);
nand U12327 (N_12327,N_11616,N_11252);
nand U12328 (N_12328,N_11173,N_10414);
nor U12329 (N_12329,N_9777,N_10364);
xor U12330 (N_12330,N_11465,N_11228);
nor U12331 (N_12331,N_10581,N_10514);
or U12332 (N_12332,N_9526,N_9253);
nor U12333 (N_12333,N_9052,N_10743);
nand U12334 (N_12334,N_9747,N_10453);
xnor U12335 (N_12335,N_9803,N_11642);
nand U12336 (N_12336,N_9294,N_9814);
or U12337 (N_12337,N_9194,N_10321);
nand U12338 (N_12338,N_10970,N_11070);
xor U12339 (N_12339,N_9705,N_10375);
xor U12340 (N_12340,N_10184,N_9056);
xor U12341 (N_12341,N_11641,N_10679);
nand U12342 (N_12342,N_11844,N_11467);
xor U12343 (N_12343,N_10512,N_11285);
or U12344 (N_12344,N_9767,N_11619);
nand U12345 (N_12345,N_10522,N_9595);
nor U12346 (N_12346,N_9218,N_9149);
nand U12347 (N_12347,N_10504,N_9639);
nor U12348 (N_12348,N_9345,N_9823);
xnor U12349 (N_12349,N_10140,N_11975);
xnor U12350 (N_12350,N_11249,N_11284);
nor U12351 (N_12351,N_10516,N_10209);
or U12352 (N_12352,N_9435,N_10596);
nand U12353 (N_12353,N_9195,N_10928);
nor U12354 (N_12354,N_10899,N_11651);
nand U12355 (N_12355,N_11420,N_10145);
nor U12356 (N_12356,N_11436,N_9380);
and U12357 (N_12357,N_11160,N_10087);
and U12358 (N_12358,N_11034,N_10757);
or U12359 (N_12359,N_10587,N_11314);
xnor U12360 (N_12360,N_10365,N_9265);
and U12361 (N_12361,N_10652,N_11596);
xnor U12362 (N_12362,N_9000,N_11472);
and U12363 (N_12363,N_9598,N_11363);
nand U12364 (N_12364,N_11918,N_11439);
nor U12365 (N_12365,N_11468,N_10922);
or U12366 (N_12366,N_9251,N_10445);
nor U12367 (N_12367,N_9168,N_9160);
and U12368 (N_12368,N_9611,N_9708);
or U12369 (N_12369,N_9091,N_9106);
nand U12370 (N_12370,N_11545,N_11962);
nor U12371 (N_12371,N_10925,N_9720);
nor U12372 (N_12372,N_11361,N_9874);
or U12373 (N_12373,N_11816,N_10955);
or U12374 (N_12374,N_11087,N_11432);
or U12375 (N_12375,N_11142,N_11039);
xor U12376 (N_12376,N_9422,N_9642);
nand U12377 (N_12377,N_9876,N_11584);
or U12378 (N_12378,N_11944,N_10199);
and U12379 (N_12379,N_11610,N_9984);
or U12380 (N_12380,N_10272,N_9619);
nor U12381 (N_12381,N_9844,N_10113);
or U12382 (N_12382,N_10096,N_9314);
nor U12383 (N_12383,N_11708,N_10584);
xor U12384 (N_12384,N_10359,N_9324);
nand U12385 (N_12385,N_10259,N_10097);
and U12386 (N_12386,N_9916,N_10471);
nor U12387 (N_12387,N_11071,N_10144);
nor U12388 (N_12388,N_10109,N_10877);
or U12389 (N_12389,N_9725,N_11647);
xnor U12390 (N_12390,N_9170,N_10075);
or U12391 (N_12391,N_10237,N_10253);
xor U12392 (N_12392,N_9062,N_9220);
and U12393 (N_12393,N_11099,N_10268);
nand U12394 (N_12394,N_11494,N_10510);
or U12395 (N_12395,N_9658,N_10211);
nor U12396 (N_12396,N_11231,N_10699);
and U12397 (N_12397,N_10495,N_9961);
nand U12398 (N_12398,N_9491,N_9729);
nor U12399 (N_12399,N_11475,N_11401);
nor U12400 (N_12400,N_10137,N_9782);
xor U12401 (N_12401,N_10115,N_9615);
and U12402 (N_12402,N_9928,N_10035);
nor U12403 (N_12403,N_10563,N_10068);
nor U12404 (N_12404,N_9596,N_11764);
xor U12405 (N_12405,N_11860,N_9457);
and U12406 (N_12406,N_10460,N_10569);
and U12407 (N_12407,N_9706,N_9970);
xnor U12408 (N_12408,N_11908,N_10660);
xor U12409 (N_12409,N_9769,N_10941);
nor U12410 (N_12410,N_9678,N_9946);
nor U12411 (N_12411,N_9659,N_11072);
nand U12412 (N_12412,N_11820,N_10559);
nor U12413 (N_12413,N_9064,N_10874);
nand U12414 (N_12414,N_11896,N_10226);
and U12415 (N_12415,N_9207,N_11220);
nand U12416 (N_12416,N_11245,N_9305);
nand U12417 (N_12417,N_11575,N_10630);
or U12418 (N_12418,N_10907,N_10032);
and U12419 (N_12419,N_9684,N_9383);
nand U12420 (N_12420,N_10971,N_9035);
and U12421 (N_12421,N_11480,N_11578);
nor U12422 (N_12422,N_9338,N_11695);
and U12423 (N_12423,N_10833,N_11564);
nand U12424 (N_12424,N_11206,N_10297);
nor U12425 (N_12425,N_11428,N_10427);
xor U12426 (N_12426,N_10189,N_10688);
or U12427 (N_12427,N_11621,N_10814);
or U12428 (N_12428,N_11372,N_10550);
xnor U12429 (N_12429,N_11976,N_9319);
nor U12430 (N_12430,N_11088,N_10043);
nor U12431 (N_12431,N_11459,N_9496);
or U12432 (N_12432,N_11298,N_10422);
or U12433 (N_12433,N_11850,N_10720);
nor U12434 (N_12434,N_10742,N_10435);
and U12435 (N_12435,N_9622,N_11313);
xnor U12436 (N_12436,N_10371,N_9848);
nand U12437 (N_12437,N_9386,N_11791);
nor U12438 (N_12438,N_9635,N_9556);
nor U12439 (N_12439,N_9190,N_9559);
nand U12440 (N_12440,N_9758,N_11541);
nor U12441 (N_12441,N_11980,N_9564);
nor U12442 (N_12442,N_9308,N_9860);
and U12443 (N_12443,N_11675,N_9994);
or U12444 (N_12444,N_11403,N_10173);
nand U12445 (N_12445,N_9602,N_11594);
and U12446 (N_12446,N_11452,N_9714);
and U12447 (N_12447,N_10093,N_10458);
or U12448 (N_12448,N_10081,N_10502);
and U12449 (N_12449,N_11655,N_10735);
xnor U12450 (N_12450,N_11557,N_10547);
nor U12451 (N_12451,N_11750,N_9438);
nor U12452 (N_12452,N_10493,N_10558);
xor U12453 (N_12453,N_9192,N_11316);
nand U12454 (N_12454,N_11194,N_10716);
nor U12455 (N_12455,N_9638,N_10863);
and U12456 (N_12456,N_9155,N_10457);
and U12457 (N_12457,N_11470,N_10934);
xor U12458 (N_12458,N_9074,N_9963);
and U12459 (N_12459,N_9101,N_11735);
or U12460 (N_12460,N_10246,N_10527);
nand U12461 (N_12461,N_10884,N_11684);
xnor U12462 (N_12462,N_9440,N_11994);
nand U12463 (N_12463,N_10088,N_10769);
xnor U12464 (N_12464,N_9073,N_11795);
xnor U12465 (N_12465,N_11640,N_10564);
or U12466 (N_12466,N_11778,N_11744);
nand U12467 (N_12467,N_9560,N_9931);
xor U12468 (N_12468,N_9718,N_11805);
nor U12469 (N_12469,N_11141,N_11280);
and U12470 (N_12470,N_9477,N_11340);
or U12471 (N_12471,N_11819,N_9490);
nand U12472 (N_12472,N_11736,N_11222);
or U12473 (N_12473,N_10838,N_10151);
or U12474 (N_12474,N_9077,N_9617);
or U12475 (N_12475,N_11580,N_10962);
nand U12476 (N_12476,N_9452,N_10136);
xnor U12477 (N_12477,N_10854,N_11649);
and U12478 (N_12478,N_9026,N_9623);
xnor U12479 (N_12479,N_11533,N_11342);
nor U12480 (N_12480,N_10931,N_10793);
xnor U12481 (N_12481,N_10965,N_10562);
or U12482 (N_12482,N_11474,N_9884);
or U12483 (N_12483,N_11694,N_10120);
nor U12484 (N_12484,N_9361,N_9716);
xnor U12485 (N_12485,N_11008,N_10816);
or U12486 (N_12486,N_10236,N_11614);
and U12487 (N_12487,N_9586,N_10260);
or U12488 (N_12488,N_11115,N_9102);
and U12489 (N_12489,N_9118,N_10142);
and U12490 (N_12490,N_10945,N_9188);
nand U12491 (N_12491,N_11093,N_9015);
nor U12492 (N_12492,N_10683,N_10705);
xnor U12493 (N_12493,N_11511,N_10138);
or U12494 (N_12494,N_10442,N_9406);
or U12495 (N_12495,N_11991,N_11923);
or U12496 (N_12496,N_9648,N_10022);
nor U12497 (N_12497,N_9202,N_10845);
xor U12498 (N_12498,N_11384,N_10231);
xor U12499 (N_12499,N_10187,N_11997);
and U12500 (N_12500,N_11672,N_10340);
and U12501 (N_12501,N_11295,N_11873);
and U12502 (N_12502,N_9989,N_11147);
nand U12503 (N_12503,N_10314,N_9261);
nand U12504 (N_12504,N_11456,N_10821);
nand U12505 (N_12505,N_10362,N_10208);
and U12506 (N_12506,N_11630,N_11048);
nand U12507 (N_12507,N_11855,N_10916);
nor U12508 (N_12508,N_9531,N_9140);
or U12509 (N_12509,N_10525,N_10640);
xnor U12510 (N_12510,N_9175,N_11287);
nor U12511 (N_12511,N_10811,N_9745);
and U12512 (N_12512,N_10989,N_9254);
xor U12513 (N_12513,N_10738,N_11894);
nor U12514 (N_12514,N_10376,N_9426);
xnor U12515 (N_12515,N_9661,N_10468);
nand U12516 (N_12516,N_9276,N_11134);
nor U12517 (N_12517,N_10799,N_11078);
xor U12518 (N_12518,N_10319,N_9612);
nor U12519 (N_12519,N_10603,N_9739);
and U12520 (N_12520,N_9248,N_10710);
xor U12521 (N_12521,N_10752,N_11977);
nor U12522 (N_12522,N_10310,N_9681);
and U12523 (N_12523,N_11731,N_10101);
nand U12524 (N_12524,N_10175,N_11514);
and U12525 (N_12525,N_11512,N_10575);
or U12526 (N_12526,N_11783,N_9935);
xnor U12527 (N_12527,N_9411,N_11504);
nor U12528 (N_12528,N_11229,N_10963);
xor U12529 (N_12529,N_9836,N_10728);
and U12530 (N_12530,N_10687,N_9245);
nor U12531 (N_12531,N_11001,N_10589);
and U12532 (N_12532,N_11158,N_9709);
xor U12533 (N_12533,N_11782,N_9174);
nand U12534 (N_12534,N_11282,N_10836);
and U12535 (N_12535,N_10131,N_11521);
nor U12536 (N_12536,N_11927,N_9330);
nor U12537 (N_12537,N_11283,N_9437);
or U12538 (N_12538,N_11804,N_9640);
nand U12539 (N_12539,N_9488,N_10357);
and U12540 (N_12540,N_9385,N_10341);
xor U12541 (N_12541,N_10706,N_9150);
nand U12542 (N_12542,N_10937,N_11746);
and U12543 (N_12543,N_10006,N_9498);
xnor U12544 (N_12544,N_11683,N_11685);
or U12545 (N_12545,N_9756,N_11020);
or U12546 (N_12546,N_11872,N_11957);
xnor U12547 (N_12547,N_10887,N_9504);
xor U12548 (N_12548,N_9232,N_10846);
or U12549 (N_12549,N_9733,N_10410);
nor U12550 (N_12550,N_11607,N_11563);
nand U12551 (N_12551,N_10615,N_10695);
nor U12552 (N_12552,N_10653,N_10897);
or U12553 (N_12553,N_9500,N_10245);
and U12554 (N_12554,N_10360,N_10295);
nor U12555 (N_12555,N_9346,N_9311);
xor U12556 (N_12556,N_11955,N_9981);
and U12557 (N_12557,N_9866,N_11030);
nor U12558 (N_12558,N_9554,N_11016);
nand U12559 (N_12559,N_9193,N_9594);
or U12560 (N_12560,N_9122,N_10225);
and U12561 (N_12561,N_9125,N_9014);
xnor U12562 (N_12562,N_11992,N_11018);
nor U12563 (N_12563,N_9061,N_9820);
or U12564 (N_12564,N_10837,N_9173);
and U12565 (N_12565,N_11191,N_11832);
xor U12566 (N_12566,N_11487,N_10167);
and U12567 (N_12567,N_9813,N_9793);
nand U12568 (N_12568,N_11983,N_10438);
nand U12569 (N_12569,N_11217,N_9179);
nor U12570 (N_12570,N_11067,N_10374);
and U12571 (N_12571,N_9965,N_10685);
nand U12572 (N_12572,N_11035,N_11251);
nand U12573 (N_12573,N_9295,N_11027);
and U12574 (N_12574,N_10932,N_11038);
nand U12575 (N_12575,N_11743,N_10778);
and U12576 (N_12576,N_9980,N_11843);
xor U12577 (N_12577,N_9973,N_11155);
xnor U12578 (N_12578,N_9585,N_11526);
or U12579 (N_12579,N_10578,N_10401);
or U12580 (N_12580,N_9002,N_9505);
nor U12581 (N_12581,N_10358,N_11720);
and U12582 (N_12582,N_11256,N_10737);
xor U12583 (N_12583,N_11751,N_11242);
nand U12584 (N_12584,N_9783,N_11887);
or U12585 (N_12585,N_11321,N_9303);
xor U12586 (N_12586,N_9864,N_9943);
nor U12587 (N_12587,N_9079,N_9373);
or U12588 (N_12588,N_10770,N_9887);
xnor U12589 (N_12589,N_9022,N_10518);
nor U12590 (N_12590,N_9795,N_10413);
nor U12591 (N_12591,N_9343,N_9321);
nor U12592 (N_12592,N_9041,N_9001);
or U12593 (N_12593,N_11262,N_9894);
xor U12594 (N_12594,N_11453,N_10385);
nand U12595 (N_12595,N_11349,N_10843);
nor U12596 (N_12596,N_10315,N_10979);
nand U12597 (N_12597,N_11190,N_11993);
and U12598 (N_12598,N_11871,N_9650);
nor U12599 (N_12599,N_10306,N_9226);
nand U12600 (N_12600,N_10526,N_10764);
or U12601 (N_12601,N_10625,N_10632);
or U12602 (N_12602,N_11259,N_9100);
nor U12603 (N_12603,N_10729,N_10634);
nor U12604 (N_12604,N_11540,N_10997);
and U12605 (N_12605,N_11566,N_11143);
or U12606 (N_12606,N_9045,N_9664);
xnor U12607 (N_12607,N_9663,N_10803);
nand U12608 (N_12608,N_9875,N_9049);
xnor U12609 (N_12609,N_11775,N_11076);
xor U12610 (N_12610,N_10895,N_9872);
nand U12611 (N_12611,N_10395,N_11577);
nand U12612 (N_12612,N_11230,N_11952);
or U12613 (N_12613,N_9423,N_11722);
or U12614 (N_12614,N_10111,N_11762);
and U12615 (N_12615,N_11668,N_11959);
nor U12616 (N_12616,N_11506,N_10249);
and U12617 (N_12617,N_11704,N_10397);
and U12618 (N_12618,N_9982,N_10842);
or U12619 (N_12619,N_11073,N_11322);
or U12620 (N_12620,N_9348,N_11628);
and U12621 (N_12621,N_9507,N_11265);
or U12622 (N_12622,N_10010,N_10610);
xor U12623 (N_12623,N_11773,N_10772);
xor U12624 (N_12624,N_9185,N_9656);
xnor U12625 (N_12625,N_11042,N_10668);
xnor U12626 (N_12626,N_10505,N_11771);
nand U12627 (N_12627,N_11268,N_9471);
and U12628 (N_12628,N_11861,N_9013);
xor U12629 (N_12629,N_11613,N_11154);
and U12630 (N_12630,N_11516,N_10806);
nand U12631 (N_12631,N_10862,N_11738);
xnor U12632 (N_12632,N_11045,N_9694);
xnor U12633 (N_12633,N_10680,N_9163);
nor U12634 (N_12634,N_10105,N_11781);
nor U12635 (N_12635,N_11429,N_11271);
and U12636 (N_12636,N_10222,N_10089);
xor U12637 (N_12637,N_9407,N_10629);
and U12638 (N_12638,N_11920,N_11634);
xor U12639 (N_12639,N_11170,N_10601);
nor U12640 (N_12640,N_9792,N_10285);
nand U12641 (N_12641,N_11264,N_11216);
nor U12642 (N_12642,N_9141,N_10662);
nand U12643 (N_12643,N_9880,N_9897);
xor U12644 (N_12644,N_9563,N_9030);
nand U12645 (N_12645,N_9271,N_9367);
nand U12646 (N_12646,N_11809,N_9124);
nand U12647 (N_12647,N_11457,N_11448);
nand U12648 (N_12648,N_11969,N_9054);
nand U12649 (N_12649,N_9743,N_9019);
xnor U12650 (N_12650,N_11928,N_11582);
xor U12651 (N_12651,N_10592,N_9198);
and U12652 (N_12652,N_10121,N_11546);
nor U12653 (N_12653,N_9234,N_11583);
nor U12654 (N_12654,N_11495,N_9956);
nand U12655 (N_12655,N_11343,N_11091);
and U12656 (N_12656,N_9012,N_11421);
nand U12657 (N_12657,N_10869,N_10802);
or U12658 (N_12658,N_10591,N_11180);
xnor U12659 (N_12659,N_9082,N_11454);
nand U12660 (N_12660,N_10213,N_10531);
or U12661 (N_12661,N_11435,N_10538);
nor U12662 (N_12662,N_10933,N_10430);
xor U12663 (N_12663,N_11799,N_9147);
nor U12664 (N_12664,N_11907,N_11567);
nor U12665 (N_12665,N_10156,N_11181);
or U12666 (N_12666,N_11169,N_9121);
xor U12667 (N_12667,N_10450,N_11753);
nor U12668 (N_12668,N_11824,N_9544);
nand U12669 (N_12669,N_10848,N_9112);
or U12670 (N_12670,N_9685,N_10515);
xor U12671 (N_12671,N_11290,N_11879);
nand U12672 (N_12672,N_10041,N_10451);
nand U12673 (N_12673,N_10642,N_10648);
or U12674 (N_12674,N_9468,N_9539);
or U12675 (N_12675,N_11164,N_10719);
or U12676 (N_12676,N_9590,N_11635);
or U12677 (N_12677,N_11633,N_10380);
or U12678 (N_12678,N_9365,N_9735);
nand U12679 (N_12679,N_11849,N_10333);
nand U12680 (N_12680,N_9575,N_10795);
xnor U12681 (N_12681,N_11885,N_9043);
and U12682 (N_12682,N_10712,N_11065);
xor U12683 (N_12683,N_9281,N_10761);
nand U12684 (N_12684,N_10588,N_10307);
and U12685 (N_12685,N_10433,N_9382);
nand U12686 (N_12686,N_11418,N_9095);
xor U12687 (N_12687,N_11659,N_10481);
and U12688 (N_12688,N_11758,N_10560);
nand U12689 (N_12689,N_9252,N_10947);
nor U12690 (N_12690,N_11930,N_11415);
or U12691 (N_12691,N_11507,N_9517);
xnor U12692 (N_12692,N_9906,N_11388);
or U12693 (N_12693,N_9243,N_11964);
nor U12694 (N_12694,N_9201,N_9811);
xor U12695 (N_12695,N_11241,N_10127);
xor U12696 (N_12696,N_9926,N_11627);
nand U12697 (N_12697,N_9652,N_9312);
or U12698 (N_12698,N_9518,N_11312);
and U12699 (N_12699,N_9320,N_10730);
and U12700 (N_12700,N_10338,N_11481);
nor U12701 (N_12701,N_9329,N_11916);
nand U12702 (N_12702,N_10882,N_11033);
nor U12703 (N_12703,N_10098,N_11876);
xnor U12704 (N_12704,N_11692,N_10497);
or U12705 (N_12705,N_11139,N_11698);
xor U12706 (N_12706,N_11227,N_10715);
xnor U12707 (N_12707,N_9693,N_10775);
nor U12708 (N_12708,N_10964,N_11768);
xor U12709 (N_12709,N_10112,N_9021);
and U12710 (N_12710,N_11797,N_11440);
and U12711 (N_12711,N_11788,N_10573);
and U12712 (N_12712,N_10637,N_11700);
xnor U12713 (N_12713,N_11337,N_10170);
and U12714 (N_12714,N_11806,N_9816);
xor U12715 (N_12715,N_10464,N_10440);
and U12716 (N_12716,N_10293,N_10168);
nor U12717 (N_12717,N_11437,N_10094);
nand U12718 (N_12718,N_9588,N_11341);
xor U12719 (N_12719,N_10294,N_11492);
and U12720 (N_12720,N_9463,N_9352);
and U12721 (N_12721,N_10789,N_11553);
xnor U12722 (N_12722,N_9318,N_9726);
nor U12723 (N_12723,N_11623,N_11570);
nand U12724 (N_12724,N_9057,N_9270);
nor U12725 (N_12725,N_11915,N_10337);
nor U12726 (N_12726,N_9953,N_10675);
or U12727 (N_12727,N_9624,N_9279);
and U12728 (N_12728,N_11319,N_9260);
or U12729 (N_12729,N_9278,N_10053);
or U12730 (N_12730,N_9987,N_10048);
xor U12731 (N_12731,N_10503,N_10149);
nand U12732 (N_12732,N_10066,N_10501);
xor U12733 (N_12733,N_11917,N_10714);
nor U12734 (N_12734,N_9291,N_11837);
nor U12735 (N_12735,N_9776,N_10544);
or U12736 (N_12736,N_9223,N_9978);
and U12737 (N_12737,N_11124,N_10815);
xnor U12738 (N_12738,N_10805,N_11888);
nand U12739 (N_12739,N_9985,N_9372);
xor U12740 (N_12740,N_11606,N_10777);
xor U12741 (N_12741,N_10810,N_10701);
nor U12742 (N_12742,N_9148,N_10239);
and U12743 (N_12743,N_9878,N_9606);
xnor U12744 (N_12744,N_10178,N_9341);
or U12745 (N_12745,N_11209,N_11458);
nand U12746 (N_12746,N_11971,N_10533);
nand U12747 (N_12747,N_11471,N_10534);
nand U12748 (N_12748,N_10797,N_9374);
nand U12749 (N_12749,N_11269,N_9707);
or U12750 (N_12750,N_9785,N_11182);
nand U12751 (N_12751,N_9134,N_9462);
or U12752 (N_12752,N_9404,N_10813);
and U12753 (N_12753,N_9715,N_11853);
nand U12754 (N_12754,N_9740,N_9667);
nand U12755 (N_12755,N_11609,N_9501);
xor U12756 (N_12756,N_9250,N_10067);
nor U12757 (N_12757,N_11053,N_11947);
nand U12758 (N_12758,N_11880,N_9832);
nor U12759 (N_12759,N_9369,N_10608);
or U12760 (N_12760,N_10661,N_11365);
xor U12761 (N_12761,N_10614,N_11430);
nor U12762 (N_12762,N_11586,N_11987);
xor U12763 (N_12763,N_9209,N_9822);
nor U12764 (N_12764,N_9821,N_9269);
or U12765 (N_12765,N_11581,N_11737);
nor U12766 (N_12766,N_10991,N_11715);
and U12767 (N_12767,N_9711,N_9882);
nor U12768 (N_12768,N_9410,N_10475);
nor U12769 (N_12769,N_10090,N_9511);
nand U12770 (N_12770,N_10063,N_10948);
nand U12771 (N_12771,N_11168,N_10528);
nand U12772 (N_12772,N_10990,N_10906);
nand U12773 (N_12773,N_11741,N_11411);
xnor U12774 (N_12774,N_10015,N_9537);
xor U12775 (N_12775,N_10817,N_10702);
xor U12776 (N_12776,N_10045,N_9883);
nand U12777 (N_12777,N_9654,N_11967);
nor U12778 (N_12778,N_10220,N_10760);
nor U12779 (N_12779,N_9362,N_11998);
or U12780 (N_12780,N_11089,N_11188);
and U12781 (N_12781,N_9589,N_11603);
nand U12782 (N_12782,N_9818,N_9332);
or U12783 (N_12783,N_10950,N_9418);
or U12784 (N_12784,N_11780,N_10347);
or U12785 (N_12785,N_10949,N_11882);
nand U12786 (N_12786,N_11103,N_11118);
and U12787 (N_12787,N_9166,N_11755);
nor U12788 (N_12788,N_10164,N_11112);
nand U12789 (N_12789,N_10159,N_11856);
xnor U12790 (N_12790,N_11443,N_9105);
or U12791 (N_12791,N_9241,N_11699);
xor U12792 (N_12792,N_11989,N_10872);
nand U12793 (N_12793,N_9683,N_10320);
xor U12794 (N_12794,N_9568,N_10080);
nand U12795 (N_12795,N_9249,N_9835);
xnor U12796 (N_12796,N_9211,N_10461);
nor U12797 (N_12797,N_10829,N_9922);
and U12798 (N_12798,N_11274,N_10666);
or U12799 (N_12799,N_9868,N_10202);
nand U12800 (N_12800,N_10196,N_9764);
nand U12801 (N_12801,N_11503,N_10548);
xor U12802 (N_12802,N_11276,N_10016);
nand U12803 (N_12803,N_9710,N_9933);
xnor U12804 (N_12804,N_9024,N_11793);
nand U12805 (N_12805,N_11836,N_11149);
and U12806 (N_12806,N_10262,N_11090);
and U12807 (N_12807,N_10366,N_10288);
xnor U12808 (N_12808,N_9391,N_10506);
or U12809 (N_12809,N_10586,N_9527);
xnor U12810 (N_12810,N_11177,N_9139);
xnor U12811 (N_12811,N_9203,N_9904);
xor U12812 (N_12812,N_10804,N_10890);
or U12813 (N_12813,N_9379,N_11727);
or U12814 (N_12814,N_10455,N_11555);
or U12815 (N_12815,N_11416,N_10007);
nand U12816 (N_12816,N_11352,N_11055);
and U12817 (N_12817,N_9702,N_10696);
nor U12818 (N_12818,N_11620,N_11542);
or U12819 (N_12819,N_9399,N_11278);
or U12820 (N_12820,N_11382,N_10739);
nor U12821 (N_12821,N_11859,N_9774);
and U12822 (N_12822,N_11019,N_10361);
or U12823 (N_12823,N_11572,N_11629);
nor U12824 (N_12824,N_10773,N_9256);
xnor U12825 (N_12825,N_10415,N_11929);
xor U12826 (N_12826,N_9120,N_9310);
nor U12827 (N_12827,N_10059,N_9197);
and U12828 (N_12828,N_9375,N_9996);
xnor U12829 (N_12829,N_9065,N_9228);
nand U12830 (N_12830,N_9824,N_11905);
or U12831 (N_12831,N_11137,N_11323);
and U12832 (N_12832,N_9187,N_11822);
and U12833 (N_12833,N_11176,N_11729);
or U12834 (N_12834,N_10114,N_9017);
nand U12835 (N_12835,N_9206,N_9543);
nor U12836 (N_12836,N_10312,N_11450);
nand U12837 (N_12837,N_11333,N_9273);
or U12838 (N_12838,N_11084,N_9464);
or U12839 (N_12839,N_11573,N_10296);
or U12840 (N_12840,N_10670,N_9344);
and U12841 (N_12841,N_9964,N_10072);
nand U12842 (N_12842,N_10553,N_9770);
and U12843 (N_12843,N_11243,N_11497);
xnor U12844 (N_12844,N_9990,N_9071);
nand U12845 (N_12845,N_10771,N_11579);
nand U12846 (N_12846,N_9535,N_9521);
xor U12847 (N_12847,N_10748,N_10343);
and U12848 (N_12848,N_11015,N_10235);
xnor U12849 (N_12849,N_9287,N_11664);
nand U12850 (N_12850,N_10038,N_11525);
nor U12851 (N_12851,N_10355,N_11463);
nand U12852 (N_12852,N_10663,N_9480);
or U12853 (N_12853,N_11874,N_11120);
nor U12854 (N_12854,N_11921,N_11389);
xor U12855 (N_12855,N_10524,N_10070);
nor U12856 (N_12856,N_10331,N_9761);
nor U12857 (N_12857,N_10232,N_9534);
nor U12858 (N_12858,N_9757,N_10106);
and U12859 (N_12859,N_10996,N_9392);
or U12860 (N_12860,N_11852,N_11098);
nand U12861 (N_12861,N_11260,N_11445);
and U12862 (N_12862,N_11250,N_9009);
or U12863 (N_12863,N_10555,N_11212);
and U12864 (N_12864,N_10535,N_9900);
nor U12865 (N_12865,N_11904,N_10256);
or U12866 (N_12866,N_11100,N_10252);
or U12867 (N_12867,N_11131,N_11834);
or U12868 (N_12868,N_9264,N_9216);
xor U12869 (N_12869,N_9494,N_10019);
or U12870 (N_12870,N_11914,N_10620);
and U12871 (N_12871,N_11549,N_11375);
or U12872 (N_12872,N_10172,N_10891);
and U12873 (N_12873,N_11884,N_10758);
or U12874 (N_12874,N_10372,N_9161);
nor U12875 (N_12875,N_10617,N_11339);
nor U12876 (N_12876,N_9117,N_9567);
nand U12877 (N_12877,N_11096,N_9316);
nand U12878 (N_12878,N_10224,N_11900);
nand U12879 (N_12879,N_10827,N_10776);
xnor U12880 (N_12880,N_10600,N_11032);
nand U12881 (N_12881,N_9053,N_11079);
xnor U12882 (N_12882,N_10638,N_11499);
nor U12883 (N_12883,N_11275,N_9796);
nor U12884 (N_12884,N_11211,N_9828);
nor U12885 (N_12885,N_9184,N_10576);
nor U12886 (N_12886,N_9229,N_11326);
nor U12887 (N_12887,N_11551,N_11179);
nor U12888 (N_12888,N_10873,N_9370);
nor U12889 (N_12889,N_10165,N_11831);
and U12890 (N_12890,N_11488,N_11515);
xnor U12891 (N_12891,N_10967,N_9760);
or U12892 (N_12892,N_9553,N_10229);
and U12893 (N_12893,N_9533,N_9208);
nor U12894 (N_12894,N_9574,N_10704);
xor U12895 (N_12895,N_10216,N_10420);
nor U12896 (N_12896,N_11447,N_10580);
nand U12897 (N_12897,N_10431,N_10180);
and U12898 (N_12898,N_10210,N_11059);
nand U12899 (N_12899,N_10783,N_11075);
or U12900 (N_12900,N_9387,N_10405);
nand U12901 (N_12901,N_9246,N_11040);
or U12902 (N_12902,N_10855,N_9525);
or U12903 (N_12903,N_9039,N_11807);
nand U12904 (N_12904,N_11505,N_10709);
or U12905 (N_12905,N_10201,N_10160);
xor U12906 (N_12906,N_10692,N_9752);
xnor U12907 (N_12907,N_9899,N_11357);
nor U12908 (N_12908,N_9719,N_10147);
xor U12909 (N_12909,N_11272,N_10058);
or U12910 (N_12910,N_9503,N_11442);
or U12911 (N_12911,N_10556,N_9301);
nor U12912 (N_12912,N_10529,N_9236);
or U12913 (N_12913,N_11368,N_9384);
nand U12914 (N_12914,N_11943,N_11787);
or U12915 (N_12915,N_9080,N_10020);
nor U12916 (N_12916,N_9183,N_11893);
xor U12917 (N_12917,N_10994,N_10711);
nor U12918 (N_12918,N_10047,N_10973);
xor U12919 (N_12919,N_11152,N_9613);
nor U12920 (N_12920,N_10373,N_10482);
xnor U12921 (N_12921,N_9280,N_10264);
and U12922 (N_12922,N_10492,N_11501);
and U12923 (N_12923,N_11617,N_11865);
or U12924 (N_12924,N_11239,N_9162);
xnor U12925 (N_12925,N_9334,N_11593);
or U12926 (N_12926,N_9081,N_11237);
nand U12927 (N_12927,N_10077,N_9368);
nor U12928 (N_12928,N_11125,N_11107);
nor U12929 (N_12929,N_10943,N_9186);
xor U12930 (N_12930,N_11058,N_10417);
and U12931 (N_12931,N_9620,N_10408);
nand U12932 (N_12932,N_11346,N_11144);
xnor U12933 (N_12933,N_10983,N_10377);
nor U12934 (N_12934,N_11528,N_9842);
nand U12935 (N_12935,N_9633,N_9858);
nor U12936 (N_12936,N_10346,N_9358);
or U12937 (N_12937,N_11461,N_10972);
xor U12938 (N_12938,N_9258,N_9673);
or U12939 (N_12939,N_11080,N_10554);
xnor U12940 (N_12940,N_10308,N_11367);
nand U12941 (N_12941,N_11949,N_9846);
or U12942 (N_12942,N_9854,N_10721);
or U12943 (N_12943,N_11966,N_11130);
or U12944 (N_12944,N_9114,N_11234);
and U12945 (N_12945,N_9285,N_11978);
nand U12946 (N_12946,N_9096,N_11419);
and U12947 (N_12947,N_11345,N_11941);
xnor U12948 (N_12948,N_11336,N_9717);
nor U12949 (N_12949,N_11127,N_10832);
nand U12950 (N_12950,N_11706,N_9579);
nor U12951 (N_12951,N_11119,N_10270);
or U12952 (N_12952,N_11460,N_11200);
or U12953 (N_12953,N_11446,N_10920);
and U12954 (N_12954,N_10809,N_11359);
xor U12955 (N_12955,N_9363,N_11486);
or U12956 (N_12956,N_11292,N_9834);
and U12957 (N_12957,N_9695,N_10282);
or U12958 (N_12958,N_11552,N_11906);
nand U12959 (N_12959,N_10335,N_10436);
and U12960 (N_12960,N_10012,N_11972);
nand U12961 (N_12961,N_10014,N_11602);
nor U12962 (N_12962,N_10490,N_10792);
nand U12963 (N_12963,N_10040,N_11847);
and U12964 (N_12964,N_11696,N_11476);
nor U12965 (N_12965,N_9547,N_10767);
nand U12966 (N_12966,N_10291,N_11380);
xnor U12967 (N_12967,N_10546,N_9976);
or U12968 (N_12968,N_10747,N_9129);
or U12969 (N_12969,N_10241,N_9448);
or U12970 (N_12970,N_10641,N_9889);
xor U12971 (N_12971,N_9789,N_9655);
xnor U12972 (N_12972,N_11565,N_10905);
nor U12973 (N_12973,N_10543,N_9458);
nand U12974 (N_12974,N_11689,N_9879);
and U12975 (N_12975,N_9008,N_9046);
or U12976 (N_12976,N_11643,N_10725);
and U12977 (N_12977,N_10472,N_11028);
xor U12978 (N_12978,N_10536,N_11652);
nand U12979 (N_12979,N_10200,N_11961);
nor U12980 (N_12980,N_9532,N_9355);
or U12981 (N_12981,N_10915,N_11254);
nor U12982 (N_12982,N_11562,N_9090);
or U12983 (N_12983,N_11717,N_10292);
nand U12984 (N_12984,N_10129,N_11247);
and U12985 (N_12985,N_10064,N_11395);
or U12986 (N_12986,N_10656,N_11482);
xor U12987 (N_12987,N_11077,N_9450);
nor U12988 (N_12988,N_11772,N_9219);
or U12989 (N_12989,N_11417,N_9069);
nor U12990 (N_12990,N_10532,N_10655);
xor U12991 (N_12991,N_11747,N_11665);
nand U12992 (N_12992,N_10909,N_10749);
nor U12993 (N_12993,N_11676,N_9495);
nand U12994 (N_12994,N_10992,N_11277);
nor U12995 (N_12995,N_9429,N_11968);
nand U12996 (N_12996,N_9093,N_11493);
and U12997 (N_12997,N_9432,N_11996);
xnor U12998 (N_12998,N_10327,N_9812);
or U12999 (N_12999,N_10108,N_9672);
and U13000 (N_13000,N_11187,N_11561);
nand U13001 (N_13001,N_9636,N_9538);
nand U13002 (N_13002,N_10429,N_10250);
nor U13003 (N_13003,N_10095,N_9768);
nor U13004 (N_13004,N_10602,N_10033);
nand U13005 (N_13005,N_9016,N_10421);
and U13006 (N_13006,N_9339,N_10621);
nor U13007 (N_13007,N_9690,N_11901);
or U13008 (N_13008,N_10423,N_9200);
and U13009 (N_13009,N_9628,N_11982);
xnor U13010 (N_13010,N_10938,N_11726);
nor U13011 (N_13011,N_11777,N_10835);
and U13012 (N_13012,N_9023,N_10388);
nand U13013 (N_13013,N_11301,N_11984);
nand U13014 (N_13014,N_10031,N_9066);
nor U13015 (N_13015,N_9643,N_11536);
xnor U13016 (N_13016,N_10995,N_11669);
or U13017 (N_13017,N_9932,N_11539);
nor U13018 (N_13018,N_11789,N_10929);
or U13019 (N_13019,N_11423,N_11354);
and U13020 (N_13020,N_9267,N_9728);
nor U13021 (N_13021,N_9587,N_11654);
and U13022 (N_13022,N_10509,N_9297);
xnor U13023 (N_13023,N_10416,N_11204);
and U13024 (N_13024,N_9670,N_11378);
nand U13025 (N_13025,N_10993,N_11827);
or U13026 (N_13026,N_10188,N_11892);
or U13027 (N_13027,N_10976,N_11309);
nand U13028 (N_13028,N_10911,N_10074);
and U13029 (N_13029,N_10284,N_9442);
or U13030 (N_13030,N_11146,N_11114);
xnor U13031 (N_13031,N_9651,N_9840);
nand U13032 (N_13032,N_11151,N_10134);
nand U13033 (N_13033,N_10883,N_9268);
nor U13034 (N_13034,N_9509,N_9898);
or U13035 (N_13035,N_11604,N_10009);
or U13036 (N_13036,N_10418,N_10957);
nand U13037 (N_13037,N_11165,N_9199);
or U13038 (N_13038,N_10354,N_10171);
nand U13039 (N_13039,N_10369,N_11857);
or U13040 (N_13040,N_9755,N_10921);
and U13041 (N_13041,N_11166,N_9455);
xnor U13042 (N_13042,N_11502,N_9152);
and U13043 (N_13043,N_9849,N_10860);
or U13044 (N_13044,N_9136,N_11829);
xnor U13045 (N_13045,N_11159,N_11060);
xnor U13046 (N_13046,N_10301,N_10079);
and U13047 (N_13047,N_11940,N_10221);
and U13048 (N_13048,N_10486,N_10322);
nand U13049 (N_13049,N_11051,N_9945);
nand U13050 (N_13050,N_11348,N_11444);
nand U13051 (N_13051,N_9847,N_9238);
nand U13052 (N_13052,N_11412,N_9327);
nor U13053 (N_13053,N_11703,N_11723);
or U13054 (N_13054,N_11713,N_11335);
and U13055 (N_13055,N_9626,N_9975);
xor U13056 (N_13056,N_11302,N_10083);
nand U13057 (N_13057,N_10387,N_11733);
nor U13058 (N_13058,N_10788,N_11197);
and U13059 (N_13059,N_10779,N_10984);
nor U13060 (N_13060,N_9167,N_9240);
nand U13061 (N_13061,N_10658,N_9299);
nand U13062 (N_13062,N_9512,N_10645);
xor U13063 (N_13063,N_10049,N_9067);
or U13064 (N_13064,N_10381,N_11757);
nand U13065 (N_13065,N_10647,N_11174);
nand U13066 (N_13066,N_9862,N_11004);
or U13067 (N_13067,N_9130,N_11413);
nor U13068 (N_13068,N_9430,N_10886);
or U13069 (N_13069,N_9420,N_11911);
or U13070 (N_13070,N_11344,N_10313);
or U13071 (N_13071,N_10807,N_11297);
xnor U13072 (N_13072,N_11383,N_11203);
or U13073 (N_13073,N_11138,N_11205);
nor U13074 (N_13074,N_9665,N_11740);
and U13075 (N_13075,N_9262,N_10091);
xnor U13076 (N_13076,N_9349,N_11686);
or U13077 (N_13077,N_9582,N_9481);
nor U13078 (N_13078,N_9955,N_11126);
and U13079 (N_13079,N_9333,N_10870);
nand U13080 (N_13080,N_9449,N_10162);
or U13081 (N_13081,N_11397,N_10998);
nor U13082 (N_13082,N_10856,N_10023);
and U13083 (N_13083,N_11121,N_10822);
or U13084 (N_13084,N_9286,N_9901);
or U13085 (N_13085,N_10830,N_10400);
and U13086 (N_13086,N_9514,N_9649);
or U13087 (N_13087,N_11823,N_10182);
or U13088 (N_13088,N_9608,N_10686);
nor U13089 (N_13089,N_9540,N_11646);
xnor U13090 (N_13090,N_10269,N_9873);
xor U13091 (N_13091,N_9666,N_11958);
or U13092 (N_13092,N_11101,N_10143);
or U13093 (N_13093,N_10152,N_11311);
nand U13094 (N_13094,N_9653,N_11714);
nor U13095 (N_13095,N_9703,N_11990);
or U13096 (N_13096,N_11598,N_9289);
nand U13097 (N_13097,N_10665,N_11303);
nand U13098 (N_13098,N_10654,N_9109);
or U13099 (N_13099,N_11595,N_10218);
or U13100 (N_13100,N_11132,N_10223);
and U13101 (N_13101,N_10693,N_11294);
and U13102 (N_13102,N_9797,N_11786);
xor U13103 (N_13103,N_10186,N_11148);
nor U13104 (N_13104,N_9810,N_9087);
nand U13105 (N_13105,N_11183,N_9988);
and U13106 (N_13106,N_11062,N_9826);
nor U13107 (N_13107,N_10823,N_9212);
nand U13108 (N_13108,N_10402,N_9888);
or U13109 (N_13109,N_11221,N_9632);
nor U13110 (N_13110,N_11116,N_9323);
or U13111 (N_13111,N_10392,N_10677);
nand U13112 (N_13112,N_11371,N_9692);
nor U13113 (N_13113,N_9603,N_9513);
or U13114 (N_13114,N_9519,N_11489);
and U13115 (N_13115,N_9128,N_11381);
and U13116 (N_13116,N_9920,N_9304);
or U13117 (N_13117,N_11263,N_11693);
and U13118 (N_13118,N_11658,N_11558);
nor U13119 (N_13119,N_10465,N_11841);
or U13120 (N_13120,N_11730,N_10903);
and U13121 (N_13121,N_10616,N_9999);
xnor U13122 (N_13122,N_11932,N_10940);
xor U13123 (N_13123,N_10025,N_11068);
or U13124 (N_13124,N_10623,N_10577);
nor U13125 (N_13125,N_10052,N_9393);
nor U13126 (N_13126,N_11207,N_10479);
or U13127 (N_13127,N_9581,N_11749);
xnor U13128 (N_13128,N_10281,N_9536);
nand U13129 (N_13129,N_9466,N_11745);
nand U13130 (N_13130,N_10999,N_9969);
or U13131 (N_13131,N_10276,N_11122);
nand U13132 (N_13132,N_9937,N_11508);
nor U13133 (N_13133,N_10511,N_11414);
nor U13134 (N_13134,N_10901,N_9751);
nor U13135 (N_13135,N_9038,N_9971);
and U13136 (N_13136,N_9415,N_9178);
or U13137 (N_13137,N_9601,N_9400);
and U13138 (N_13138,N_11592,N_11478);
nor U13139 (N_13139,N_9660,N_9746);
nor U13140 (N_13140,N_9722,N_10448);
nand U13141 (N_13141,N_9780,N_9322);
nor U13142 (N_13142,N_9781,N_10029);
and U13143 (N_13143,N_11425,N_10027);
nand U13144 (N_13144,N_10820,N_9431);
xor U13145 (N_13145,N_11934,N_10477);
nand U13146 (N_13146,N_9871,N_10349);
xor U13147 (N_13147,N_10488,N_9750);
nand U13148 (N_13148,N_11086,N_9851);
nand U13149 (N_13149,N_11688,N_9927);
xor U13150 (N_13150,N_11576,N_11104);
nor U13151 (N_13151,N_10698,N_9156);
or U13152 (N_13152,N_11656,N_9078);
nor U13153 (N_13153,N_11246,N_10988);
and U13154 (N_13154,N_9414,N_9131);
or U13155 (N_13155,N_11085,N_10316);
nand U13156 (N_13156,N_10011,N_10626);
or U13157 (N_13157,N_9790,N_9723);
nor U13158 (N_13158,N_9196,N_11682);
and U13159 (N_13159,N_11379,N_10517);
or U13160 (N_13160,N_11351,N_10050);
nand U13161 (N_13161,N_9180,N_11513);
nor U13162 (N_13162,N_10132,N_10166);
and U13163 (N_13163,N_9515,N_10759);
nand U13164 (N_13164,N_11393,N_10859);
nor U13165 (N_13165,N_11210,N_11304);
xnor U13166 (N_13166,N_11779,N_11530);
xnor U13167 (N_13167,N_9850,N_11406);
nor U13168 (N_13168,N_10107,N_10944);
or U13169 (N_13169,N_11153,N_10724);
nor U13170 (N_13170,N_9773,N_9597);
nand U13171 (N_13171,N_9724,N_9580);
xnor U13172 (N_13172,N_11202,N_9356);
nor U13173 (N_13173,N_9137,N_9135);
or U13174 (N_13174,N_9213,N_11625);
nand U13175 (N_13175,N_9037,N_11434);
or U13176 (N_13176,N_10311,N_11022);
nand U13177 (N_13177,N_9915,N_9506);
nor U13178 (N_13178,N_9473,N_9469);
nand U13179 (N_13179,N_11286,N_9523);
nor U13180 (N_13180,N_9454,N_10238);
or U13181 (N_13181,N_10746,N_9569);
nand U13182 (N_13182,N_9959,N_9424);
nor U13183 (N_13183,N_11590,N_9484);
and U13184 (N_13184,N_9954,N_9489);
xor U13185 (N_13185,N_10076,N_11293);
or U13186 (N_13186,N_11049,N_10248);
nor U13187 (N_13187,N_9353,N_10781);
or U13188 (N_13188,N_9210,N_10428);
nand U13189 (N_13189,N_10918,N_9610);
nand U13190 (N_13190,N_11026,N_10480);
nor U13191 (N_13191,N_11662,N_9607);
and U13192 (N_13192,N_11973,N_9791);
nand U13193 (N_13193,N_9629,N_10082);
nand U13194 (N_13194,N_10328,N_11171);
nor U13195 (N_13195,N_11097,N_11279);
and U13196 (N_13196,N_11868,N_9592);
nor U13197 (N_13197,N_10552,N_9938);
nor U13198 (N_13198,N_10342,N_10958);
nand U13199 (N_13199,N_9817,N_9086);
or U13200 (N_13200,N_10583,N_9412);
or U13201 (N_13201,N_9433,N_9441);
xor U13202 (N_13202,N_10597,N_11909);
or U13203 (N_13203,N_11981,N_10254);
nor U13204 (N_13204,N_10334,N_10537);
and U13205 (N_13205,N_10489,N_10277);
nor U13206 (N_13206,N_9766,N_11063);
and U13207 (N_13207,N_9111,N_10300);
xnor U13208 (N_13208,N_10056,N_10124);
or U13209 (N_13209,N_10234,N_10545);
xnor U13210 (N_13210,N_11175,N_10690);
xor U13211 (N_13211,N_10892,N_10736);
nor U13212 (N_13212,N_11331,N_10824);
nor U13213 (N_13213,N_11390,N_10148);
nand U13214 (N_13214,N_11954,N_11574);
nor U13215 (N_13215,N_9905,N_9340);
nor U13216 (N_13216,N_11306,N_10485);
xnor U13217 (N_13217,N_9486,N_10672);
nand U13218 (N_13218,N_9784,N_11800);
nand U13219 (N_13219,N_10092,N_10540);
and U13220 (N_13220,N_11261,N_11424);
nor U13221 (N_13221,N_9189,N_11589);
nor U13222 (N_13222,N_10317,N_11858);
and U13223 (N_13223,N_9687,N_11477);
and U13224 (N_13224,N_11890,N_9960);
and U13225 (N_13225,N_10119,N_11054);
or U13226 (N_13226,N_10163,N_10831);
xor U13227 (N_13227,N_11483,N_11315);
nand U13228 (N_13228,N_11554,N_11784);
nand U13229 (N_13229,N_9224,N_9788);
or U13230 (N_13230,N_10348,N_11398);
and U13231 (N_13231,N_10598,N_9890);
nand U13232 (N_13232,N_9668,N_10707);
xnor U13233 (N_13233,N_9427,N_10794);
or U13234 (N_13234,N_11718,N_11867);
and U13235 (N_13235,N_11310,N_10731);
and U13236 (N_13236,N_11299,N_10303);
or U13237 (N_13237,N_10643,N_9151);
or U13238 (N_13238,N_10888,N_9944);
or U13239 (N_13239,N_11320,N_9646);
and U13240 (N_13240,N_11496,N_9786);
or U13241 (N_13241,N_11005,N_11705);
and U13242 (N_13242,N_9942,N_10141);
and U13243 (N_13243,N_11041,N_9621);
and U13244 (N_13244,N_11864,N_11732);
nand U13245 (N_13245,N_11707,N_9604);
xor U13246 (N_13246,N_10762,N_9119);
and U13247 (N_13247,N_9731,N_10727);
and U13248 (N_13248,N_10158,N_10852);
nand U13249 (N_13249,N_10305,N_9401);
or U13250 (N_13250,N_9328,N_11069);
or U13251 (N_13251,N_10787,N_9359);
xor U13252 (N_13252,N_9721,N_10267);
or U13253 (N_13253,N_9274,N_9799);
or U13254 (N_13254,N_10378,N_10117);
xnor U13255 (N_13255,N_9979,N_10722);
and U13256 (N_13256,N_11218,N_9446);
and U13257 (N_13257,N_10644,N_9070);
xnor U13258 (N_13258,N_11449,N_9998);
or U13259 (N_13259,N_9403,N_10054);
or U13260 (N_13260,N_10447,N_11043);
or U13261 (N_13261,N_11386,N_11308);
nand U13262 (N_13262,N_9625,N_11950);
nand U13263 (N_13263,N_10078,N_11774);
and U13264 (N_13264,N_9390,N_9436);
nor U13265 (N_13265,N_9845,N_10754);
nand U13266 (N_13266,N_10935,N_11233);
nand U13267 (N_13267,N_10062,N_10812);
xor U13268 (N_13268,N_10700,N_10951);
nor U13269 (N_13269,N_9309,N_9779);
or U13270 (N_13270,N_10391,N_10659);
xor U13271 (N_13271,N_10452,N_10713);
and U13272 (N_13272,N_9326,N_10042);
or U13273 (N_13273,N_11817,N_10765);
and U13274 (N_13274,N_9076,N_10102);
or U13275 (N_13275,N_9524,N_9033);
and U13276 (N_13276,N_9307,N_11113);
and U13277 (N_13277,N_10061,N_10636);
or U13278 (N_13278,N_9893,N_11886);
xnor U13279 (N_13279,N_11109,N_11933);
or U13280 (N_13280,N_11813,N_10936);
nor U13281 (N_13281,N_10323,N_9451);
and U13282 (N_13282,N_9902,N_10923);
xor U13283 (N_13283,N_11196,N_11599);
and U13284 (N_13284,N_11524,N_9113);
xnor U13285 (N_13285,N_10446,N_11712);
nand U13286 (N_13286,N_10896,N_9142);
or U13287 (N_13287,N_9863,N_10441);
and U13288 (N_13288,N_11219,N_11979);
nor U13289 (N_13289,N_11895,N_11267);
or U13290 (N_13290,N_10394,N_10861);
or U13291 (N_13291,N_10071,N_11851);
xnor U13292 (N_13292,N_10611,N_11009);
nand U13293 (N_13293,N_10419,N_9675);
and U13294 (N_13294,N_9600,N_11353);
xnor U13295 (N_13295,N_11891,N_11123);
xnor U13296 (N_13296,N_9696,N_11875);
xor U13297 (N_13297,N_10176,N_9593);
nand U13298 (N_13298,N_10193,N_10924);
xnor U13299 (N_13299,N_11798,N_9063);
xnor U13300 (N_13300,N_9701,N_9807);
nor U13301 (N_13301,N_11631,N_9662);
nand U13302 (N_13302,N_9680,N_9453);
nand U13303 (N_13303,N_9951,N_10671);
or U13304 (N_13304,N_10513,N_10681);
nand U13305 (N_13305,N_10673,N_10135);
xnor U13306 (N_13306,N_10798,N_10910);
nor U13307 (N_13307,N_11902,N_11910);
xor U13308 (N_13308,N_9762,N_10689);
or U13309 (N_13309,N_11003,N_11670);
nor U13310 (N_13310,N_11674,N_10398);
nand U13311 (N_13311,N_10594,N_10520);
and U13312 (N_13312,N_11716,N_11632);
xor U13313 (N_13313,N_11538,N_11391);
nor U13314 (N_13314,N_11711,N_9044);
xnor U13315 (N_13315,N_9153,N_10878);
and U13316 (N_13316,N_10893,N_10960);
and U13317 (N_13317,N_9609,N_11709);
nor U13318 (N_13318,N_10473,N_9800);
nor U13319 (N_13319,N_9977,N_11790);
nand U13320 (N_13320,N_10613,N_9936);
nand U13321 (N_13321,N_11270,N_10326);
nand U13322 (N_13322,N_9911,N_11317);
and U13323 (N_13323,N_11136,N_10881);
and U13324 (N_13324,N_10389,N_10212);
nand U13325 (N_13325,N_10104,N_11105);
and U13326 (N_13326,N_10839,N_11660);
xor U13327 (N_13327,N_10926,N_10449);
or U13328 (N_13328,N_11585,N_11568);
nand U13329 (N_13329,N_11213,N_9123);
nor U13330 (N_13330,N_9510,N_11742);
nand U13331 (N_13331,N_9028,N_10966);
nand U13332 (N_13332,N_10336,N_11364);
nand U13333 (N_13333,N_11491,N_11329);
nand U13334 (N_13334,N_9058,N_10622);
or U13335 (N_13335,N_11663,N_9968);
nor U13336 (N_13336,N_11374,N_11057);
and U13337 (N_13337,N_9247,N_10631);
and U13338 (N_13338,N_9389,N_9099);
and U13339 (N_13339,N_10953,N_11102);
nand U13340 (N_13340,N_11812,N_9138);
nor U13341 (N_13341,N_9749,N_9159);
nor U13342 (N_13342,N_9541,N_11167);
and U13343 (N_13343,N_9558,N_10900);
xnor U13344 (N_13344,N_10819,N_11082);
and U13345 (N_13345,N_11671,N_11433);
nor U13346 (N_13346,N_11899,N_11360);
nor U13347 (N_13347,N_11129,N_11356);
xor U13348 (N_13348,N_9983,N_9171);
and U13349 (N_13349,N_9482,N_10651);
and U13350 (N_13350,N_9397,N_9290);
nand U13351 (N_13351,N_9853,N_9913);
xnor U13352 (N_13352,N_9741,N_10350);
nor U13353 (N_13353,N_10255,N_9644);
xor U13354 (N_13354,N_9221,N_9402);
xor U13355 (N_13355,N_10484,N_11680);
and U13356 (N_13356,N_11510,N_9618);
nor U13357 (N_13357,N_10103,N_10002);
or U13358 (N_13358,N_10036,N_11815);
nor U13359 (N_13359,N_11830,N_11014);
or U13360 (N_13360,N_10384,N_9225);
xor U13361 (N_13361,N_9947,N_9405);
nand U13362 (N_13362,N_11673,N_9047);
nor U13363 (N_13363,N_10542,N_9753);
or U13364 (N_13364,N_10875,N_10939);
xnor U13365 (N_13365,N_9181,N_10980);
nor U13366 (N_13366,N_9029,N_11639);
nor U13367 (N_13367,N_9805,N_9263);
nand U13368 (N_13368,N_11224,N_10904);
or U13369 (N_13369,N_9011,N_10368);
nor U13370 (N_13370,N_9378,N_9689);
and U13371 (N_13371,N_9919,N_11064);
nor U13372 (N_13372,N_9434,N_11157);
nand U13373 (N_13373,N_10961,N_9154);
xor U13374 (N_13374,N_9825,N_10274);
nand U13375 (N_13375,N_9794,N_10055);
and U13376 (N_13376,N_11522,N_11846);
and U13377 (N_13377,N_10549,N_9084);
nand U13378 (N_13378,N_11029,N_10864);
nor U13379 (N_13379,N_11534,N_11031);
nor U13380 (N_13380,N_9839,N_10469);
or U13381 (N_13381,N_11409,N_11215);
or U13382 (N_13382,N_10379,N_11615);
or U13383 (N_13383,N_9530,N_11427);
and U13384 (N_13384,N_10024,N_10463);
xor U13385 (N_13385,N_10390,N_11803);
xnor U13386 (N_13386,N_11828,N_11000);
or U13387 (N_13387,N_11007,N_10122);
xnor U13388 (N_13388,N_11618,N_9331);
xor U13389 (N_13389,N_9923,N_10913);
and U13390 (N_13390,N_9682,N_10498);
xnor U13391 (N_13391,N_11588,N_9924);
or U13392 (N_13392,N_11527,N_10986);
and U13393 (N_13393,N_11485,N_9158);
xnor U13394 (N_13394,N_11821,N_10086);
xor U13395 (N_13395,N_10154,N_11612);
nor U13396 (N_13396,N_11760,N_11362);
nor U13397 (N_13397,N_9421,N_9018);
nor U13398 (N_13398,N_10345,N_11399);
nor U13399 (N_13399,N_11679,N_9205);
or U13400 (N_13400,N_9059,N_11258);
and U13401 (N_13401,N_9259,N_9686);
nand U13402 (N_13402,N_9474,N_11037);
and U13403 (N_13403,N_11766,N_10356);
nor U13404 (N_13404,N_10462,N_11999);
nand U13405 (N_13405,N_10508,N_10283);
xnor U13406 (N_13406,N_9966,N_10628);
nor U13407 (N_13407,N_10494,N_11024);
xor U13408 (N_13408,N_10914,N_10786);
xor U13409 (N_13409,N_11520,N_9679);
or U13410 (N_13410,N_10191,N_11392);
nand U13411 (N_13411,N_10280,N_10981);
nand U13412 (N_13412,N_9857,N_9972);
nor U13413 (N_13413,N_9508,N_11624);
xnor U13414 (N_13414,N_9815,N_9838);
xnor U13415 (N_13415,N_9502,N_11150);
xnor U13416 (N_13416,N_10826,N_10982);
xnor U13417 (N_13417,N_10426,N_10399);
xor U13418 (N_13418,N_11877,N_10483);
and U13419 (N_13419,N_10858,N_9227);
nand U13420 (N_13420,N_9856,N_9566);
or U13421 (N_13421,N_11133,N_10876);
or U13422 (N_13422,N_11556,N_9974);
xor U13423 (N_13423,N_11192,N_10766);
nand U13424 (N_13424,N_10125,N_9092);
nor U13425 (N_13425,N_11464,N_10396);
nor U13426 (N_13426,N_11273,N_9360);
nand U13427 (N_13427,N_9930,N_9907);
or U13428 (N_13428,N_10478,N_11752);
nand U13429 (N_13429,N_11951,N_11214);
nand U13430 (N_13430,N_9257,N_11863);
nor U13431 (N_13431,N_11407,N_11248);
nand U13432 (N_13432,N_10551,N_11763);
and U13433 (N_13433,N_11926,N_9007);
and U13434 (N_13434,N_10828,N_9381);
and U13435 (N_13435,N_10650,N_10018);
nand U13436 (N_13436,N_11327,N_11919);
or U13437 (N_13437,N_9775,N_9616);
and U13438 (N_13438,N_11903,N_10919);
xor U13439 (N_13439,N_11792,N_10183);
or U13440 (N_13440,N_10840,N_10406);
nand U13441 (N_13441,N_10557,N_9283);
xnor U13442 (N_13442,N_9445,N_9614);
xor U13443 (N_13443,N_11225,N_9891);
nand U13444 (N_13444,N_9909,N_11559);
nor U13445 (N_13445,N_10582,N_9470);
xor U13446 (N_13446,N_9300,N_9917);
nand U13447 (N_13447,N_9351,N_10181);
xnor U13448 (N_13448,N_9914,N_9895);
nor U13449 (N_13449,N_10784,N_9934);
or U13450 (N_13450,N_11500,N_9107);
xnor U13451 (N_13451,N_11544,N_10046);
or U13452 (N_13452,N_9108,N_10847);
nor U13453 (N_13453,N_9098,N_9704);
nor U13454 (N_13454,N_11854,N_11044);
nand U13455 (N_13455,N_9145,N_9485);
nor U13456 (N_13456,N_11548,N_10403);
or U13457 (N_13457,N_9645,N_9398);
or U13458 (N_13458,N_11645,N_9055);
or U13459 (N_13459,N_9881,N_9993);
and U13460 (N_13460,N_9952,N_11074);
xnor U13461 (N_13461,N_11988,N_10065);
nand U13462 (N_13462,N_9921,N_10227);
nor U13463 (N_13463,N_10791,N_9631);
and U13464 (N_13464,N_10139,N_9475);
nor U13465 (N_13465,N_11838,N_10978);
nor U13466 (N_13466,N_9522,N_9765);
nor U13467 (N_13467,N_9317,N_10853);
and U13468 (N_13468,N_11529,N_10205);
and U13469 (N_13469,N_11644,N_11600);
or U13470 (N_13470,N_10017,N_10567);
nand U13471 (N_13471,N_10466,N_10796);
xnor U13472 (N_13472,N_11878,N_9584);
and U13473 (N_13473,N_9191,N_9051);
nand U13474 (N_13474,N_10099,N_9647);
or U13475 (N_13475,N_10561,N_11601);
xnor U13476 (N_13476,N_11931,N_9698);
or U13477 (N_13477,N_10974,N_9499);
nor U13478 (N_13478,N_9771,N_9115);
nor U13479 (N_13479,N_9827,N_10894);
nor U13480 (N_13480,N_9852,N_11012);
and U13481 (N_13481,N_10289,N_11025);
or U13482 (N_13482,N_11366,N_9546);
nand U13483 (N_13483,N_10590,N_11611);
and U13484 (N_13484,N_10745,N_10849);
xnor U13485 (N_13485,N_9006,N_10579);
nor U13486 (N_13486,N_9772,N_9493);
xnor U13487 (N_13487,N_11739,N_10383);
nor U13488 (N_13488,N_9957,N_9641);
xnor U13489 (N_13489,N_10627,N_9865);
nor U13490 (N_13490,N_11734,N_11257);
nand U13491 (N_13491,N_10353,N_10329);
and U13492 (N_13492,N_9177,N_9908);
xor U13493 (N_13493,N_9034,N_11140);
nor U13494 (N_13494,N_9388,N_10519);
xnor U13495 (N_13495,N_11305,N_11047);
nor U13496 (N_13496,N_10258,N_9583);
nor U13497 (N_13497,N_10619,N_9456);
or U13498 (N_13498,N_10755,N_10785);
or U13499 (N_13499,N_11725,N_10723);
and U13500 (N_13500,N_10199,N_9575);
nor U13501 (N_13501,N_9625,N_9660);
nor U13502 (N_13502,N_10202,N_9843);
nor U13503 (N_13503,N_11076,N_10627);
nand U13504 (N_13504,N_9954,N_10127);
xor U13505 (N_13505,N_9254,N_10690);
or U13506 (N_13506,N_11109,N_10253);
nand U13507 (N_13507,N_9458,N_11948);
or U13508 (N_13508,N_10721,N_9224);
nand U13509 (N_13509,N_10661,N_9133);
nand U13510 (N_13510,N_9313,N_11406);
or U13511 (N_13511,N_10222,N_10011);
nand U13512 (N_13512,N_9546,N_11255);
nand U13513 (N_13513,N_11853,N_9681);
and U13514 (N_13514,N_10395,N_9619);
nor U13515 (N_13515,N_10076,N_11124);
or U13516 (N_13516,N_11972,N_9721);
or U13517 (N_13517,N_10911,N_9524);
or U13518 (N_13518,N_9183,N_9631);
or U13519 (N_13519,N_11472,N_9682);
and U13520 (N_13520,N_10549,N_10785);
or U13521 (N_13521,N_9578,N_11522);
nand U13522 (N_13522,N_9803,N_9081);
and U13523 (N_13523,N_11600,N_10779);
and U13524 (N_13524,N_9998,N_9354);
nor U13525 (N_13525,N_10241,N_9609);
nand U13526 (N_13526,N_9072,N_9222);
xnor U13527 (N_13527,N_11855,N_10106);
nand U13528 (N_13528,N_9626,N_11154);
nor U13529 (N_13529,N_9056,N_10149);
and U13530 (N_13530,N_9644,N_10671);
nor U13531 (N_13531,N_11113,N_10305);
nand U13532 (N_13532,N_11584,N_9923);
or U13533 (N_13533,N_11565,N_11761);
xnor U13534 (N_13534,N_10100,N_9598);
nor U13535 (N_13535,N_11896,N_9125);
and U13536 (N_13536,N_11912,N_9627);
nand U13537 (N_13537,N_11966,N_9957);
xnor U13538 (N_13538,N_10034,N_11120);
or U13539 (N_13539,N_11538,N_10838);
nand U13540 (N_13540,N_11920,N_10186);
or U13541 (N_13541,N_11004,N_11384);
nor U13542 (N_13542,N_11360,N_9574);
and U13543 (N_13543,N_11565,N_9131);
or U13544 (N_13544,N_11410,N_11217);
nor U13545 (N_13545,N_9218,N_11230);
or U13546 (N_13546,N_11520,N_9251);
and U13547 (N_13547,N_11376,N_10997);
nand U13548 (N_13548,N_10180,N_11890);
or U13549 (N_13549,N_11023,N_9877);
and U13550 (N_13550,N_11026,N_10557);
nand U13551 (N_13551,N_10218,N_10254);
and U13552 (N_13552,N_9447,N_11785);
nand U13553 (N_13553,N_10107,N_10991);
or U13554 (N_13554,N_11855,N_9449);
and U13555 (N_13555,N_11037,N_10552);
xor U13556 (N_13556,N_10358,N_9807);
and U13557 (N_13557,N_9974,N_9949);
and U13558 (N_13558,N_10054,N_9078);
xor U13559 (N_13559,N_9060,N_9448);
and U13560 (N_13560,N_10726,N_9036);
xor U13561 (N_13561,N_11675,N_10792);
or U13562 (N_13562,N_11283,N_11710);
nor U13563 (N_13563,N_11521,N_10661);
or U13564 (N_13564,N_11633,N_10814);
nor U13565 (N_13565,N_10992,N_9880);
nor U13566 (N_13566,N_10321,N_10701);
nor U13567 (N_13567,N_10266,N_10180);
or U13568 (N_13568,N_9180,N_10702);
nor U13569 (N_13569,N_11006,N_10060);
nand U13570 (N_13570,N_10717,N_9657);
nand U13571 (N_13571,N_10103,N_11980);
nand U13572 (N_13572,N_10270,N_11677);
nand U13573 (N_13573,N_11761,N_10240);
xor U13574 (N_13574,N_9014,N_10179);
xnor U13575 (N_13575,N_11398,N_10402);
xnor U13576 (N_13576,N_11662,N_10043);
or U13577 (N_13577,N_10201,N_10354);
or U13578 (N_13578,N_10990,N_10721);
and U13579 (N_13579,N_11807,N_11071);
and U13580 (N_13580,N_9003,N_9421);
nor U13581 (N_13581,N_11689,N_11629);
and U13582 (N_13582,N_9123,N_11019);
xor U13583 (N_13583,N_11595,N_9776);
nand U13584 (N_13584,N_11718,N_10021);
xor U13585 (N_13585,N_9752,N_10407);
xor U13586 (N_13586,N_10020,N_10669);
and U13587 (N_13587,N_10016,N_10022);
and U13588 (N_13588,N_9275,N_9205);
xor U13589 (N_13589,N_10062,N_10597);
nor U13590 (N_13590,N_9039,N_10820);
or U13591 (N_13591,N_9801,N_11599);
xnor U13592 (N_13592,N_9984,N_11215);
nand U13593 (N_13593,N_10533,N_10923);
xor U13594 (N_13594,N_11012,N_11858);
xnor U13595 (N_13595,N_10489,N_11318);
and U13596 (N_13596,N_9069,N_10820);
or U13597 (N_13597,N_9623,N_11419);
or U13598 (N_13598,N_11652,N_10772);
and U13599 (N_13599,N_10491,N_9913);
or U13600 (N_13600,N_10295,N_10316);
nor U13601 (N_13601,N_9111,N_9127);
or U13602 (N_13602,N_9373,N_9180);
xor U13603 (N_13603,N_9422,N_9519);
or U13604 (N_13604,N_10825,N_10514);
nand U13605 (N_13605,N_11794,N_10246);
xnor U13606 (N_13606,N_11632,N_9410);
and U13607 (N_13607,N_10274,N_11432);
or U13608 (N_13608,N_10962,N_9550);
xnor U13609 (N_13609,N_10955,N_9559);
nor U13610 (N_13610,N_9198,N_11336);
nand U13611 (N_13611,N_10412,N_11720);
nand U13612 (N_13612,N_11044,N_11073);
xnor U13613 (N_13613,N_11626,N_9406);
xnor U13614 (N_13614,N_11578,N_11523);
or U13615 (N_13615,N_10655,N_10921);
nand U13616 (N_13616,N_11021,N_9638);
nand U13617 (N_13617,N_11530,N_10896);
nand U13618 (N_13618,N_11930,N_10308);
xor U13619 (N_13619,N_11802,N_9076);
xor U13620 (N_13620,N_11693,N_10897);
nor U13621 (N_13621,N_10900,N_10771);
nor U13622 (N_13622,N_10580,N_11960);
nand U13623 (N_13623,N_10634,N_10846);
or U13624 (N_13624,N_9709,N_9417);
and U13625 (N_13625,N_11986,N_9370);
and U13626 (N_13626,N_10087,N_11141);
and U13627 (N_13627,N_9037,N_11323);
and U13628 (N_13628,N_11560,N_10883);
xnor U13629 (N_13629,N_10987,N_10096);
xnor U13630 (N_13630,N_10488,N_9575);
nor U13631 (N_13631,N_11894,N_10326);
and U13632 (N_13632,N_11792,N_10271);
and U13633 (N_13633,N_9125,N_9366);
xor U13634 (N_13634,N_9251,N_11540);
nor U13635 (N_13635,N_9001,N_9089);
xor U13636 (N_13636,N_10234,N_10164);
xor U13637 (N_13637,N_9813,N_9755);
or U13638 (N_13638,N_10642,N_11061);
or U13639 (N_13639,N_10943,N_11897);
nor U13640 (N_13640,N_9135,N_11860);
xnor U13641 (N_13641,N_9053,N_9888);
xor U13642 (N_13642,N_11865,N_10631);
nand U13643 (N_13643,N_10687,N_11337);
nand U13644 (N_13644,N_10956,N_9597);
xnor U13645 (N_13645,N_9891,N_11579);
nor U13646 (N_13646,N_11223,N_9294);
and U13647 (N_13647,N_11637,N_10648);
nor U13648 (N_13648,N_10469,N_11633);
nand U13649 (N_13649,N_11084,N_10582);
and U13650 (N_13650,N_10141,N_11320);
xor U13651 (N_13651,N_9594,N_10554);
nand U13652 (N_13652,N_11690,N_9988);
and U13653 (N_13653,N_9952,N_9441);
xor U13654 (N_13654,N_11092,N_11802);
or U13655 (N_13655,N_11203,N_9093);
nand U13656 (N_13656,N_9404,N_11217);
nand U13657 (N_13657,N_10454,N_9963);
and U13658 (N_13658,N_10133,N_9481);
nor U13659 (N_13659,N_11123,N_11570);
or U13660 (N_13660,N_11892,N_11920);
nor U13661 (N_13661,N_10435,N_10297);
nor U13662 (N_13662,N_10092,N_11636);
or U13663 (N_13663,N_9675,N_9820);
and U13664 (N_13664,N_11578,N_11272);
xnor U13665 (N_13665,N_10308,N_9311);
xnor U13666 (N_13666,N_9025,N_11285);
or U13667 (N_13667,N_11276,N_11099);
nor U13668 (N_13668,N_11547,N_11637);
nand U13669 (N_13669,N_11797,N_9851);
and U13670 (N_13670,N_9579,N_10403);
and U13671 (N_13671,N_10053,N_10577);
or U13672 (N_13672,N_11650,N_9084);
nand U13673 (N_13673,N_10125,N_11645);
nor U13674 (N_13674,N_9997,N_9649);
xnor U13675 (N_13675,N_11981,N_11496);
nand U13676 (N_13676,N_10932,N_10098);
and U13677 (N_13677,N_9987,N_10091);
nand U13678 (N_13678,N_9733,N_10322);
xor U13679 (N_13679,N_10957,N_11041);
nor U13680 (N_13680,N_9729,N_10223);
or U13681 (N_13681,N_11902,N_9063);
xor U13682 (N_13682,N_11948,N_10707);
nand U13683 (N_13683,N_11970,N_10882);
xor U13684 (N_13684,N_9153,N_9603);
and U13685 (N_13685,N_9415,N_11914);
or U13686 (N_13686,N_11055,N_10418);
and U13687 (N_13687,N_9089,N_11923);
or U13688 (N_13688,N_11325,N_10609);
nor U13689 (N_13689,N_10026,N_9511);
nand U13690 (N_13690,N_10402,N_9847);
nand U13691 (N_13691,N_10098,N_11441);
xor U13692 (N_13692,N_10819,N_11561);
nor U13693 (N_13693,N_10257,N_11409);
nor U13694 (N_13694,N_9713,N_11824);
xor U13695 (N_13695,N_9814,N_11718);
xor U13696 (N_13696,N_11196,N_11843);
nand U13697 (N_13697,N_11066,N_10357);
nor U13698 (N_13698,N_11586,N_9408);
or U13699 (N_13699,N_9157,N_9330);
xor U13700 (N_13700,N_9674,N_9208);
nor U13701 (N_13701,N_10015,N_11318);
nor U13702 (N_13702,N_9986,N_10392);
xnor U13703 (N_13703,N_9944,N_10581);
xnor U13704 (N_13704,N_10984,N_11451);
and U13705 (N_13705,N_9413,N_10694);
and U13706 (N_13706,N_10168,N_11155);
and U13707 (N_13707,N_11454,N_9345);
nor U13708 (N_13708,N_11301,N_9868);
nand U13709 (N_13709,N_11711,N_9464);
and U13710 (N_13710,N_11311,N_9784);
nor U13711 (N_13711,N_9790,N_10977);
or U13712 (N_13712,N_10588,N_9435);
or U13713 (N_13713,N_11990,N_11250);
nand U13714 (N_13714,N_9716,N_11438);
and U13715 (N_13715,N_11457,N_9276);
or U13716 (N_13716,N_11064,N_10587);
nand U13717 (N_13717,N_9847,N_9488);
nor U13718 (N_13718,N_11995,N_11122);
nand U13719 (N_13719,N_10817,N_11777);
or U13720 (N_13720,N_10682,N_9919);
nand U13721 (N_13721,N_9285,N_9338);
or U13722 (N_13722,N_10497,N_11461);
and U13723 (N_13723,N_11234,N_11501);
or U13724 (N_13724,N_10937,N_10538);
xnor U13725 (N_13725,N_10200,N_11989);
nor U13726 (N_13726,N_9608,N_10578);
nor U13727 (N_13727,N_9048,N_11836);
and U13728 (N_13728,N_11239,N_11078);
xnor U13729 (N_13729,N_11180,N_9099);
nand U13730 (N_13730,N_11192,N_11158);
and U13731 (N_13731,N_11985,N_11585);
nand U13732 (N_13732,N_9756,N_11226);
nand U13733 (N_13733,N_11285,N_9478);
xnor U13734 (N_13734,N_10702,N_10846);
xnor U13735 (N_13735,N_11110,N_9051);
nor U13736 (N_13736,N_9054,N_11568);
nand U13737 (N_13737,N_9838,N_9850);
xor U13738 (N_13738,N_10891,N_9527);
xor U13739 (N_13739,N_9282,N_9437);
or U13740 (N_13740,N_10196,N_9116);
nand U13741 (N_13741,N_9056,N_11071);
nand U13742 (N_13742,N_9784,N_10580);
nand U13743 (N_13743,N_10301,N_11656);
nor U13744 (N_13744,N_11571,N_9156);
or U13745 (N_13745,N_10212,N_9659);
and U13746 (N_13746,N_11937,N_10547);
nand U13747 (N_13747,N_10182,N_11992);
or U13748 (N_13748,N_11548,N_9599);
nand U13749 (N_13749,N_10228,N_10779);
and U13750 (N_13750,N_10176,N_11378);
or U13751 (N_13751,N_9155,N_9824);
and U13752 (N_13752,N_9657,N_9640);
nor U13753 (N_13753,N_11504,N_10886);
nor U13754 (N_13754,N_10387,N_10311);
nand U13755 (N_13755,N_11305,N_11527);
nand U13756 (N_13756,N_9125,N_9793);
xnor U13757 (N_13757,N_10980,N_11957);
and U13758 (N_13758,N_9849,N_11491);
nor U13759 (N_13759,N_11614,N_10012);
xor U13760 (N_13760,N_11935,N_11074);
nand U13761 (N_13761,N_9558,N_9938);
xor U13762 (N_13762,N_10017,N_11268);
nand U13763 (N_13763,N_10033,N_9375);
nand U13764 (N_13764,N_10869,N_9460);
nand U13765 (N_13765,N_10141,N_10289);
and U13766 (N_13766,N_9285,N_9715);
or U13767 (N_13767,N_10056,N_11001);
and U13768 (N_13768,N_9307,N_11393);
xnor U13769 (N_13769,N_11303,N_10038);
nand U13770 (N_13770,N_11060,N_10212);
xor U13771 (N_13771,N_9552,N_11872);
and U13772 (N_13772,N_11794,N_9456);
and U13773 (N_13773,N_9109,N_10428);
or U13774 (N_13774,N_10167,N_10899);
nor U13775 (N_13775,N_9767,N_11437);
and U13776 (N_13776,N_9570,N_10807);
or U13777 (N_13777,N_9222,N_10122);
xor U13778 (N_13778,N_9977,N_9851);
nand U13779 (N_13779,N_10068,N_10982);
or U13780 (N_13780,N_10516,N_11884);
and U13781 (N_13781,N_11991,N_10831);
nor U13782 (N_13782,N_11248,N_9503);
nor U13783 (N_13783,N_10818,N_10597);
nor U13784 (N_13784,N_9326,N_11112);
xnor U13785 (N_13785,N_11060,N_9373);
xnor U13786 (N_13786,N_9714,N_11765);
xnor U13787 (N_13787,N_11576,N_10910);
nor U13788 (N_13788,N_11725,N_9110);
nor U13789 (N_13789,N_11486,N_9387);
nand U13790 (N_13790,N_11237,N_9417);
nor U13791 (N_13791,N_9075,N_11427);
xor U13792 (N_13792,N_11138,N_9797);
and U13793 (N_13793,N_10744,N_11050);
or U13794 (N_13794,N_11510,N_11109);
xnor U13795 (N_13795,N_11515,N_9549);
and U13796 (N_13796,N_11634,N_10787);
nor U13797 (N_13797,N_10891,N_9140);
and U13798 (N_13798,N_11217,N_10576);
xor U13799 (N_13799,N_9822,N_11150);
or U13800 (N_13800,N_10940,N_10995);
or U13801 (N_13801,N_10735,N_10962);
and U13802 (N_13802,N_10419,N_11242);
nor U13803 (N_13803,N_10535,N_10170);
nand U13804 (N_13804,N_10382,N_10942);
xnor U13805 (N_13805,N_10354,N_9706);
nor U13806 (N_13806,N_10742,N_10527);
xor U13807 (N_13807,N_11554,N_11534);
nor U13808 (N_13808,N_10219,N_11846);
nand U13809 (N_13809,N_10021,N_11797);
or U13810 (N_13810,N_9045,N_11091);
nor U13811 (N_13811,N_11692,N_11683);
nor U13812 (N_13812,N_11868,N_10490);
xnor U13813 (N_13813,N_11475,N_10121);
or U13814 (N_13814,N_10947,N_11627);
and U13815 (N_13815,N_9694,N_11590);
xor U13816 (N_13816,N_11139,N_9532);
xnor U13817 (N_13817,N_11057,N_9656);
or U13818 (N_13818,N_11234,N_11768);
or U13819 (N_13819,N_9797,N_10302);
nand U13820 (N_13820,N_9769,N_9575);
and U13821 (N_13821,N_9162,N_11128);
nand U13822 (N_13822,N_11932,N_9327);
and U13823 (N_13823,N_11644,N_11699);
nand U13824 (N_13824,N_11730,N_9006);
and U13825 (N_13825,N_11182,N_11869);
and U13826 (N_13826,N_10118,N_9704);
or U13827 (N_13827,N_9885,N_11108);
nor U13828 (N_13828,N_10582,N_9660);
or U13829 (N_13829,N_10996,N_10269);
xor U13830 (N_13830,N_9115,N_9046);
nor U13831 (N_13831,N_9191,N_11847);
nor U13832 (N_13832,N_10571,N_9824);
or U13833 (N_13833,N_10276,N_11967);
or U13834 (N_13834,N_11420,N_10147);
or U13835 (N_13835,N_9009,N_11843);
or U13836 (N_13836,N_9188,N_9732);
xor U13837 (N_13837,N_10968,N_9148);
xor U13838 (N_13838,N_9028,N_10049);
nor U13839 (N_13839,N_9206,N_11760);
nor U13840 (N_13840,N_9517,N_11708);
nor U13841 (N_13841,N_11106,N_11751);
nor U13842 (N_13842,N_9362,N_9003);
nand U13843 (N_13843,N_10846,N_9703);
nor U13844 (N_13844,N_11749,N_11648);
or U13845 (N_13845,N_10306,N_10855);
or U13846 (N_13846,N_11711,N_11714);
and U13847 (N_13847,N_10038,N_11129);
nand U13848 (N_13848,N_9401,N_10562);
xnor U13849 (N_13849,N_9169,N_9335);
or U13850 (N_13850,N_10139,N_10429);
nand U13851 (N_13851,N_10551,N_11421);
xnor U13852 (N_13852,N_11791,N_9066);
nand U13853 (N_13853,N_11172,N_10530);
and U13854 (N_13854,N_9340,N_9808);
nor U13855 (N_13855,N_10501,N_11663);
or U13856 (N_13856,N_9316,N_9823);
or U13857 (N_13857,N_10369,N_9350);
or U13858 (N_13858,N_11254,N_11125);
or U13859 (N_13859,N_10197,N_11549);
xnor U13860 (N_13860,N_9344,N_9364);
xnor U13861 (N_13861,N_10410,N_9618);
nand U13862 (N_13862,N_9715,N_10259);
or U13863 (N_13863,N_9699,N_10835);
and U13864 (N_13864,N_9724,N_10417);
nor U13865 (N_13865,N_9010,N_9925);
xnor U13866 (N_13866,N_11705,N_11653);
or U13867 (N_13867,N_9410,N_9576);
nor U13868 (N_13868,N_9878,N_9090);
nor U13869 (N_13869,N_11879,N_10512);
and U13870 (N_13870,N_10696,N_9800);
xor U13871 (N_13871,N_11859,N_11240);
or U13872 (N_13872,N_9083,N_9526);
nor U13873 (N_13873,N_9189,N_11639);
nor U13874 (N_13874,N_11383,N_11915);
and U13875 (N_13875,N_9246,N_11183);
nand U13876 (N_13876,N_9197,N_11267);
and U13877 (N_13877,N_10832,N_10397);
or U13878 (N_13878,N_10410,N_11885);
xnor U13879 (N_13879,N_10566,N_11605);
nor U13880 (N_13880,N_9722,N_11557);
nand U13881 (N_13881,N_10342,N_11330);
xnor U13882 (N_13882,N_9568,N_9187);
nor U13883 (N_13883,N_10269,N_11300);
or U13884 (N_13884,N_10888,N_11056);
and U13885 (N_13885,N_10987,N_10528);
or U13886 (N_13886,N_10532,N_10811);
or U13887 (N_13887,N_9929,N_10697);
or U13888 (N_13888,N_10320,N_9351);
xnor U13889 (N_13889,N_9143,N_11348);
and U13890 (N_13890,N_11420,N_9584);
nand U13891 (N_13891,N_10522,N_9058);
or U13892 (N_13892,N_10532,N_11325);
xor U13893 (N_13893,N_10557,N_11855);
and U13894 (N_13894,N_10235,N_10455);
and U13895 (N_13895,N_11830,N_9701);
or U13896 (N_13896,N_11093,N_10205);
nor U13897 (N_13897,N_9479,N_11111);
and U13898 (N_13898,N_9639,N_11397);
or U13899 (N_13899,N_9970,N_9238);
xor U13900 (N_13900,N_10257,N_11781);
nor U13901 (N_13901,N_10666,N_10554);
nor U13902 (N_13902,N_9942,N_10871);
xor U13903 (N_13903,N_10749,N_11331);
xor U13904 (N_13904,N_9904,N_9763);
or U13905 (N_13905,N_10374,N_11677);
xor U13906 (N_13906,N_9467,N_11766);
nor U13907 (N_13907,N_9482,N_10345);
and U13908 (N_13908,N_9699,N_10008);
and U13909 (N_13909,N_9297,N_9015);
or U13910 (N_13910,N_11063,N_11645);
and U13911 (N_13911,N_11515,N_11768);
xnor U13912 (N_13912,N_11245,N_10016);
nand U13913 (N_13913,N_11462,N_11273);
or U13914 (N_13914,N_10436,N_9047);
nor U13915 (N_13915,N_9813,N_10331);
nor U13916 (N_13916,N_11953,N_9940);
xnor U13917 (N_13917,N_11635,N_9467);
nand U13918 (N_13918,N_11954,N_11336);
and U13919 (N_13919,N_9349,N_11862);
nand U13920 (N_13920,N_10523,N_11117);
nand U13921 (N_13921,N_11657,N_11587);
or U13922 (N_13922,N_9369,N_9609);
and U13923 (N_13923,N_11598,N_11834);
nor U13924 (N_13924,N_9411,N_9809);
xnor U13925 (N_13925,N_9502,N_11898);
or U13926 (N_13926,N_11704,N_10290);
nor U13927 (N_13927,N_10389,N_9797);
nor U13928 (N_13928,N_11695,N_9051);
and U13929 (N_13929,N_11018,N_11632);
nand U13930 (N_13930,N_11026,N_11300);
xnor U13931 (N_13931,N_10854,N_11993);
nand U13932 (N_13932,N_9881,N_9039);
xnor U13933 (N_13933,N_11202,N_11323);
nand U13934 (N_13934,N_11308,N_11945);
xnor U13935 (N_13935,N_10902,N_10648);
nor U13936 (N_13936,N_10953,N_9476);
xnor U13937 (N_13937,N_9263,N_11244);
xnor U13938 (N_13938,N_9111,N_10454);
nor U13939 (N_13939,N_10357,N_9929);
nand U13940 (N_13940,N_11283,N_11905);
and U13941 (N_13941,N_11960,N_9059);
nor U13942 (N_13942,N_9632,N_9444);
or U13943 (N_13943,N_10705,N_11922);
nor U13944 (N_13944,N_11090,N_11678);
xor U13945 (N_13945,N_10808,N_10843);
nor U13946 (N_13946,N_11693,N_11537);
nor U13947 (N_13947,N_9166,N_11117);
nor U13948 (N_13948,N_10584,N_9453);
or U13949 (N_13949,N_10330,N_10053);
nand U13950 (N_13950,N_10192,N_10430);
and U13951 (N_13951,N_9638,N_9337);
and U13952 (N_13952,N_11127,N_10627);
nand U13953 (N_13953,N_10882,N_9980);
or U13954 (N_13954,N_11687,N_9637);
xor U13955 (N_13955,N_11652,N_11265);
xor U13956 (N_13956,N_10958,N_11986);
or U13957 (N_13957,N_10474,N_11680);
nand U13958 (N_13958,N_11380,N_10085);
or U13959 (N_13959,N_11798,N_9265);
or U13960 (N_13960,N_11121,N_11029);
xnor U13961 (N_13961,N_9365,N_10158);
or U13962 (N_13962,N_10335,N_11553);
nand U13963 (N_13963,N_9782,N_10295);
nor U13964 (N_13964,N_9748,N_11548);
nor U13965 (N_13965,N_11385,N_11299);
and U13966 (N_13966,N_9826,N_9961);
and U13967 (N_13967,N_11332,N_11978);
nor U13968 (N_13968,N_11894,N_11909);
nor U13969 (N_13969,N_11901,N_9088);
xnor U13970 (N_13970,N_9852,N_11262);
or U13971 (N_13971,N_10327,N_10660);
nor U13972 (N_13972,N_9258,N_9557);
xnor U13973 (N_13973,N_11815,N_9935);
and U13974 (N_13974,N_10052,N_9054);
nor U13975 (N_13975,N_9636,N_11371);
xnor U13976 (N_13976,N_9556,N_9845);
nor U13977 (N_13977,N_11731,N_10914);
xnor U13978 (N_13978,N_11306,N_11038);
and U13979 (N_13979,N_11810,N_10555);
nand U13980 (N_13980,N_11206,N_9759);
nor U13981 (N_13981,N_9564,N_10974);
nor U13982 (N_13982,N_11140,N_11396);
or U13983 (N_13983,N_9952,N_10412);
nand U13984 (N_13984,N_10944,N_11822);
and U13985 (N_13985,N_11563,N_10589);
xnor U13986 (N_13986,N_11284,N_9364);
and U13987 (N_13987,N_9662,N_9888);
nand U13988 (N_13988,N_9239,N_9326);
and U13989 (N_13989,N_9762,N_9410);
nor U13990 (N_13990,N_11247,N_9664);
xnor U13991 (N_13991,N_10226,N_9397);
xor U13992 (N_13992,N_9783,N_9611);
or U13993 (N_13993,N_10790,N_9712);
nor U13994 (N_13994,N_9263,N_11681);
or U13995 (N_13995,N_10907,N_9505);
nand U13996 (N_13996,N_10959,N_11269);
and U13997 (N_13997,N_10413,N_9730);
nor U13998 (N_13998,N_11810,N_9422);
xnor U13999 (N_13999,N_11259,N_10367);
and U14000 (N_14000,N_10841,N_11456);
nand U14001 (N_14001,N_9345,N_11830);
or U14002 (N_14002,N_9880,N_11662);
and U14003 (N_14003,N_10010,N_11567);
and U14004 (N_14004,N_9496,N_10296);
or U14005 (N_14005,N_10305,N_9028);
xor U14006 (N_14006,N_10557,N_10941);
xnor U14007 (N_14007,N_9374,N_11038);
nand U14008 (N_14008,N_9538,N_11884);
and U14009 (N_14009,N_10548,N_9364);
xor U14010 (N_14010,N_10327,N_9448);
and U14011 (N_14011,N_10035,N_9268);
nand U14012 (N_14012,N_10036,N_11359);
nand U14013 (N_14013,N_10988,N_10883);
and U14014 (N_14014,N_9684,N_11754);
or U14015 (N_14015,N_11953,N_10685);
xnor U14016 (N_14016,N_11839,N_11597);
or U14017 (N_14017,N_11709,N_11310);
and U14018 (N_14018,N_10877,N_9043);
and U14019 (N_14019,N_9204,N_10855);
and U14020 (N_14020,N_11573,N_10250);
and U14021 (N_14021,N_10836,N_10229);
nor U14022 (N_14022,N_9411,N_11916);
and U14023 (N_14023,N_11530,N_10683);
or U14024 (N_14024,N_9461,N_10144);
nor U14025 (N_14025,N_9654,N_11499);
nand U14026 (N_14026,N_11237,N_11408);
xnor U14027 (N_14027,N_11433,N_9359);
nor U14028 (N_14028,N_11851,N_11064);
xor U14029 (N_14029,N_9929,N_11820);
and U14030 (N_14030,N_10444,N_10770);
nand U14031 (N_14031,N_10546,N_11734);
nor U14032 (N_14032,N_9693,N_11408);
xnor U14033 (N_14033,N_9351,N_10763);
or U14034 (N_14034,N_11243,N_9015);
nand U14035 (N_14035,N_9810,N_11303);
nand U14036 (N_14036,N_9815,N_10604);
nand U14037 (N_14037,N_9944,N_11326);
or U14038 (N_14038,N_11645,N_9200);
xnor U14039 (N_14039,N_11096,N_9283);
xnor U14040 (N_14040,N_11081,N_10779);
or U14041 (N_14041,N_9585,N_10584);
nor U14042 (N_14042,N_9589,N_10385);
xnor U14043 (N_14043,N_11266,N_10192);
or U14044 (N_14044,N_9679,N_10703);
or U14045 (N_14045,N_11517,N_11458);
xnor U14046 (N_14046,N_9802,N_9457);
nor U14047 (N_14047,N_10260,N_9271);
xnor U14048 (N_14048,N_9484,N_11448);
nor U14049 (N_14049,N_10658,N_10827);
nand U14050 (N_14050,N_11454,N_9034);
and U14051 (N_14051,N_10767,N_11467);
nand U14052 (N_14052,N_9660,N_10265);
or U14053 (N_14053,N_9012,N_10974);
nor U14054 (N_14054,N_11713,N_10410);
xor U14055 (N_14055,N_10327,N_11058);
and U14056 (N_14056,N_9852,N_9054);
nand U14057 (N_14057,N_9997,N_9912);
and U14058 (N_14058,N_10840,N_11014);
xnor U14059 (N_14059,N_10255,N_10102);
nor U14060 (N_14060,N_9654,N_11905);
and U14061 (N_14061,N_11022,N_10681);
xnor U14062 (N_14062,N_9048,N_9801);
xnor U14063 (N_14063,N_9812,N_9666);
xor U14064 (N_14064,N_10528,N_10791);
nand U14065 (N_14065,N_11752,N_9779);
xnor U14066 (N_14066,N_10082,N_11254);
nor U14067 (N_14067,N_9289,N_11049);
nand U14068 (N_14068,N_11739,N_10451);
or U14069 (N_14069,N_9235,N_11264);
nand U14070 (N_14070,N_11192,N_9166);
and U14071 (N_14071,N_10124,N_11474);
nor U14072 (N_14072,N_9811,N_11469);
or U14073 (N_14073,N_11885,N_11610);
nand U14074 (N_14074,N_11166,N_11275);
xnor U14075 (N_14075,N_10021,N_9976);
or U14076 (N_14076,N_11779,N_9908);
nand U14077 (N_14077,N_11782,N_11599);
or U14078 (N_14078,N_10867,N_9977);
xnor U14079 (N_14079,N_10161,N_10992);
and U14080 (N_14080,N_9255,N_10722);
and U14081 (N_14081,N_11195,N_11878);
or U14082 (N_14082,N_10176,N_11001);
nor U14083 (N_14083,N_11757,N_10164);
or U14084 (N_14084,N_11050,N_11292);
xnor U14085 (N_14085,N_9054,N_9537);
nor U14086 (N_14086,N_11323,N_11777);
xnor U14087 (N_14087,N_10218,N_10041);
nand U14088 (N_14088,N_9016,N_11151);
or U14089 (N_14089,N_9926,N_11749);
or U14090 (N_14090,N_9126,N_9888);
xor U14091 (N_14091,N_9019,N_10040);
or U14092 (N_14092,N_10186,N_10200);
nor U14093 (N_14093,N_9929,N_10174);
xor U14094 (N_14094,N_11799,N_9756);
or U14095 (N_14095,N_9540,N_10350);
or U14096 (N_14096,N_10455,N_10083);
xor U14097 (N_14097,N_9090,N_11167);
xor U14098 (N_14098,N_11398,N_11652);
nand U14099 (N_14099,N_10560,N_11329);
and U14100 (N_14100,N_11678,N_9641);
xor U14101 (N_14101,N_11512,N_10102);
nor U14102 (N_14102,N_10774,N_9243);
nor U14103 (N_14103,N_11638,N_11332);
or U14104 (N_14104,N_9058,N_9355);
nand U14105 (N_14105,N_11860,N_9349);
and U14106 (N_14106,N_10518,N_9102);
and U14107 (N_14107,N_10530,N_10426);
nand U14108 (N_14108,N_11972,N_10312);
nor U14109 (N_14109,N_11613,N_10399);
xor U14110 (N_14110,N_11887,N_9960);
nand U14111 (N_14111,N_10321,N_11807);
or U14112 (N_14112,N_11137,N_11643);
and U14113 (N_14113,N_9617,N_9681);
xnor U14114 (N_14114,N_11232,N_9925);
and U14115 (N_14115,N_10094,N_11627);
xnor U14116 (N_14116,N_10482,N_11902);
or U14117 (N_14117,N_11204,N_10880);
or U14118 (N_14118,N_10374,N_9530);
or U14119 (N_14119,N_11020,N_11458);
nor U14120 (N_14120,N_10912,N_9542);
or U14121 (N_14121,N_9309,N_9494);
and U14122 (N_14122,N_10091,N_9257);
xor U14123 (N_14123,N_11015,N_9455);
xor U14124 (N_14124,N_11745,N_10528);
and U14125 (N_14125,N_11137,N_9585);
nand U14126 (N_14126,N_10459,N_11730);
nor U14127 (N_14127,N_9916,N_9187);
and U14128 (N_14128,N_10634,N_9889);
nor U14129 (N_14129,N_10626,N_10106);
nor U14130 (N_14130,N_9200,N_11566);
nor U14131 (N_14131,N_9752,N_11365);
nand U14132 (N_14132,N_10014,N_11215);
nor U14133 (N_14133,N_10670,N_11980);
nor U14134 (N_14134,N_9836,N_10270);
or U14135 (N_14135,N_10572,N_10374);
nand U14136 (N_14136,N_9997,N_11402);
or U14137 (N_14137,N_10838,N_11701);
nand U14138 (N_14138,N_9577,N_10604);
nand U14139 (N_14139,N_9153,N_9296);
xor U14140 (N_14140,N_11877,N_9720);
nor U14141 (N_14141,N_10340,N_10439);
and U14142 (N_14142,N_11496,N_9124);
and U14143 (N_14143,N_11629,N_9122);
nand U14144 (N_14144,N_10260,N_10221);
and U14145 (N_14145,N_9270,N_9482);
nand U14146 (N_14146,N_11178,N_9834);
nor U14147 (N_14147,N_10450,N_11011);
and U14148 (N_14148,N_10705,N_10812);
nand U14149 (N_14149,N_9297,N_10908);
and U14150 (N_14150,N_9906,N_10716);
xnor U14151 (N_14151,N_9570,N_9747);
nand U14152 (N_14152,N_11621,N_11702);
xor U14153 (N_14153,N_9757,N_10844);
nand U14154 (N_14154,N_10461,N_10273);
or U14155 (N_14155,N_9624,N_11160);
nand U14156 (N_14156,N_10750,N_10957);
or U14157 (N_14157,N_10683,N_10882);
or U14158 (N_14158,N_11483,N_10651);
nor U14159 (N_14159,N_10303,N_10238);
and U14160 (N_14160,N_9067,N_11153);
and U14161 (N_14161,N_10551,N_10924);
nor U14162 (N_14162,N_10280,N_11200);
or U14163 (N_14163,N_9646,N_9195);
nor U14164 (N_14164,N_9279,N_10333);
nand U14165 (N_14165,N_11007,N_9711);
or U14166 (N_14166,N_11420,N_10743);
nor U14167 (N_14167,N_10147,N_10639);
or U14168 (N_14168,N_9474,N_10245);
or U14169 (N_14169,N_9052,N_9967);
nand U14170 (N_14170,N_11441,N_11148);
xor U14171 (N_14171,N_11746,N_9798);
xnor U14172 (N_14172,N_9486,N_9102);
nor U14173 (N_14173,N_10981,N_11793);
or U14174 (N_14174,N_11640,N_9890);
nand U14175 (N_14175,N_10866,N_10494);
xor U14176 (N_14176,N_10475,N_11568);
and U14177 (N_14177,N_11098,N_9407);
xnor U14178 (N_14178,N_11572,N_10849);
nand U14179 (N_14179,N_11907,N_11251);
or U14180 (N_14180,N_9912,N_9024);
nor U14181 (N_14181,N_10001,N_11875);
and U14182 (N_14182,N_9191,N_9836);
and U14183 (N_14183,N_11408,N_9246);
nor U14184 (N_14184,N_10226,N_11422);
or U14185 (N_14185,N_11287,N_11063);
and U14186 (N_14186,N_9175,N_11261);
nand U14187 (N_14187,N_9352,N_11491);
and U14188 (N_14188,N_11587,N_9936);
or U14189 (N_14189,N_11935,N_9204);
nand U14190 (N_14190,N_9763,N_9678);
xor U14191 (N_14191,N_11251,N_10589);
or U14192 (N_14192,N_10629,N_9811);
and U14193 (N_14193,N_11239,N_9111);
xnor U14194 (N_14194,N_11597,N_9644);
nand U14195 (N_14195,N_9699,N_10950);
nand U14196 (N_14196,N_11117,N_9806);
and U14197 (N_14197,N_10708,N_11346);
nor U14198 (N_14198,N_9014,N_11573);
or U14199 (N_14199,N_11589,N_11060);
and U14200 (N_14200,N_11825,N_11837);
nand U14201 (N_14201,N_10843,N_9686);
nor U14202 (N_14202,N_11824,N_11278);
and U14203 (N_14203,N_11214,N_10849);
or U14204 (N_14204,N_11730,N_11011);
nand U14205 (N_14205,N_10734,N_10354);
or U14206 (N_14206,N_9580,N_11294);
or U14207 (N_14207,N_11699,N_10621);
nand U14208 (N_14208,N_10046,N_9206);
xor U14209 (N_14209,N_10168,N_10562);
or U14210 (N_14210,N_11071,N_10379);
and U14211 (N_14211,N_10632,N_10451);
nor U14212 (N_14212,N_11983,N_11100);
nand U14213 (N_14213,N_11029,N_9152);
or U14214 (N_14214,N_11815,N_9694);
xor U14215 (N_14215,N_9478,N_10136);
or U14216 (N_14216,N_9673,N_10873);
nor U14217 (N_14217,N_11671,N_11461);
and U14218 (N_14218,N_11286,N_10119);
nor U14219 (N_14219,N_9638,N_11074);
nand U14220 (N_14220,N_9969,N_10441);
or U14221 (N_14221,N_10647,N_11912);
and U14222 (N_14222,N_9067,N_9888);
or U14223 (N_14223,N_10834,N_10711);
or U14224 (N_14224,N_11928,N_11175);
nand U14225 (N_14225,N_9421,N_10048);
or U14226 (N_14226,N_10980,N_10035);
xnor U14227 (N_14227,N_10909,N_11074);
xnor U14228 (N_14228,N_9910,N_9214);
xor U14229 (N_14229,N_9509,N_11943);
nor U14230 (N_14230,N_11157,N_10967);
nor U14231 (N_14231,N_11995,N_11354);
nand U14232 (N_14232,N_9354,N_10596);
or U14233 (N_14233,N_11560,N_10583);
or U14234 (N_14234,N_9729,N_10975);
or U14235 (N_14235,N_11726,N_10670);
xnor U14236 (N_14236,N_10985,N_9084);
or U14237 (N_14237,N_11520,N_9928);
nor U14238 (N_14238,N_11287,N_11612);
nor U14239 (N_14239,N_10965,N_10870);
nand U14240 (N_14240,N_11296,N_9014);
nand U14241 (N_14241,N_11395,N_9544);
nor U14242 (N_14242,N_11882,N_10667);
nor U14243 (N_14243,N_10853,N_11550);
and U14244 (N_14244,N_9729,N_9525);
nand U14245 (N_14245,N_10537,N_10871);
and U14246 (N_14246,N_9214,N_9777);
nor U14247 (N_14247,N_9178,N_9350);
nor U14248 (N_14248,N_11576,N_10755);
and U14249 (N_14249,N_9442,N_9257);
or U14250 (N_14250,N_11877,N_10311);
nor U14251 (N_14251,N_9506,N_11765);
nand U14252 (N_14252,N_10028,N_10734);
and U14253 (N_14253,N_10400,N_11708);
nor U14254 (N_14254,N_11354,N_9711);
xnor U14255 (N_14255,N_9246,N_11427);
nand U14256 (N_14256,N_9940,N_10260);
or U14257 (N_14257,N_9964,N_11554);
or U14258 (N_14258,N_10498,N_9383);
and U14259 (N_14259,N_10685,N_10495);
nor U14260 (N_14260,N_11022,N_11598);
or U14261 (N_14261,N_9948,N_10096);
nor U14262 (N_14262,N_11607,N_11657);
or U14263 (N_14263,N_10006,N_9017);
nand U14264 (N_14264,N_10248,N_11222);
and U14265 (N_14265,N_11100,N_11321);
nand U14266 (N_14266,N_9296,N_9477);
and U14267 (N_14267,N_9568,N_10697);
nor U14268 (N_14268,N_11136,N_11091);
nor U14269 (N_14269,N_9018,N_10613);
xnor U14270 (N_14270,N_9537,N_9421);
or U14271 (N_14271,N_11984,N_9744);
or U14272 (N_14272,N_11368,N_10194);
or U14273 (N_14273,N_11619,N_11793);
and U14274 (N_14274,N_10069,N_11102);
nand U14275 (N_14275,N_10223,N_10011);
or U14276 (N_14276,N_11020,N_11100);
xor U14277 (N_14277,N_9020,N_10875);
or U14278 (N_14278,N_10590,N_11332);
nor U14279 (N_14279,N_9812,N_9506);
xnor U14280 (N_14280,N_10319,N_11293);
or U14281 (N_14281,N_11678,N_9194);
nor U14282 (N_14282,N_11900,N_11716);
and U14283 (N_14283,N_11272,N_10603);
nor U14284 (N_14284,N_9860,N_11751);
nor U14285 (N_14285,N_9387,N_11040);
nand U14286 (N_14286,N_11819,N_9728);
nor U14287 (N_14287,N_9976,N_9991);
nor U14288 (N_14288,N_10754,N_9303);
xor U14289 (N_14289,N_9072,N_11578);
nor U14290 (N_14290,N_10720,N_11453);
and U14291 (N_14291,N_10413,N_10580);
nand U14292 (N_14292,N_10527,N_11951);
nor U14293 (N_14293,N_10981,N_9126);
or U14294 (N_14294,N_9185,N_10126);
nor U14295 (N_14295,N_11985,N_10787);
nor U14296 (N_14296,N_9482,N_10352);
nand U14297 (N_14297,N_10066,N_10532);
xor U14298 (N_14298,N_11855,N_10481);
nor U14299 (N_14299,N_9154,N_10166);
and U14300 (N_14300,N_10368,N_9974);
nor U14301 (N_14301,N_11842,N_11030);
and U14302 (N_14302,N_11463,N_11242);
and U14303 (N_14303,N_9112,N_10664);
nor U14304 (N_14304,N_9416,N_9542);
and U14305 (N_14305,N_9436,N_9608);
nor U14306 (N_14306,N_11952,N_10572);
nand U14307 (N_14307,N_9394,N_11393);
xnor U14308 (N_14308,N_10720,N_10507);
xor U14309 (N_14309,N_10347,N_9409);
xor U14310 (N_14310,N_11570,N_9013);
or U14311 (N_14311,N_11306,N_9198);
nor U14312 (N_14312,N_9025,N_10403);
nand U14313 (N_14313,N_11182,N_9566);
nand U14314 (N_14314,N_10417,N_9892);
and U14315 (N_14315,N_10569,N_11168);
and U14316 (N_14316,N_9456,N_10908);
or U14317 (N_14317,N_10140,N_9536);
and U14318 (N_14318,N_9863,N_11703);
and U14319 (N_14319,N_10883,N_11613);
nand U14320 (N_14320,N_11177,N_11124);
nand U14321 (N_14321,N_10943,N_9870);
nor U14322 (N_14322,N_10683,N_10688);
nor U14323 (N_14323,N_10068,N_9003);
and U14324 (N_14324,N_10771,N_11845);
xor U14325 (N_14325,N_11221,N_11257);
or U14326 (N_14326,N_11665,N_9125);
xnor U14327 (N_14327,N_11254,N_11922);
or U14328 (N_14328,N_10906,N_9707);
nor U14329 (N_14329,N_9753,N_11759);
nor U14330 (N_14330,N_11633,N_10142);
nand U14331 (N_14331,N_10785,N_11301);
and U14332 (N_14332,N_10013,N_9531);
nand U14333 (N_14333,N_11115,N_11526);
or U14334 (N_14334,N_11135,N_10655);
or U14335 (N_14335,N_9191,N_11809);
or U14336 (N_14336,N_9333,N_11141);
nor U14337 (N_14337,N_10485,N_11981);
nor U14338 (N_14338,N_11874,N_10538);
and U14339 (N_14339,N_11338,N_10812);
and U14340 (N_14340,N_11069,N_9602);
and U14341 (N_14341,N_10213,N_9286);
or U14342 (N_14342,N_10008,N_10637);
or U14343 (N_14343,N_10217,N_11268);
xnor U14344 (N_14344,N_11640,N_10315);
nor U14345 (N_14345,N_9175,N_11307);
nand U14346 (N_14346,N_10689,N_9635);
nor U14347 (N_14347,N_10465,N_9280);
or U14348 (N_14348,N_11114,N_10861);
nor U14349 (N_14349,N_10798,N_9990);
nor U14350 (N_14350,N_10122,N_10993);
or U14351 (N_14351,N_11538,N_10587);
and U14352 (N_14352,N_11503,N_10428);
and U14353 (N_14353,N_11944,N_9563);
or U14354 (N_14354,N_9383,N_10169);
and U14355 (N_14355,N_11672,N_11829);
nor U14356 (N_14356,N_10686,N_9331);
nor U14357 (N_14357,N_10630,N_11667);
nand U14358 (N_14358,N_10839,N_9829);
nand U14359 (N_14359,N_9613,N_9734);
or U14360 (N_14360,N_9088,N_9326);
and U14361 (N_14361,N_11862,N_9159);
nand U14362 (N_14362,N_9246,N_9913);
nand U14363 (N_14363,N_9480,N_10295);
nor U14364 (N_14364,N_11840,N_9164);
nand U14365 (N_14365,N_9416,N_11497);
nor U14366 (N_14366,N_9535,N_9815);
nor U14367 (N_14367,N_9021,N_10646);
xnor U14368 (N_14368,N_9236,N_11470);
or U14369 (N_14369,N_11583,N_9704);
or U14370 (N_14370,N_9020,N_11338);
xor U14371 (N_14371,N_9530,N_11846);
or U14372 (N_14372,N_9084,N_9323);
xnor U14373 (N_14373,N_11964,N_10648);
nand U14374 (N_14374,N_11485,N_10025);
and U14375 (N_14375,N_11322,N_9771);
nand U14376 (N_14376,N_11329,N_10166);
xor U14377 (N_14377,N_11233,N_10161);
and U14378 (N_14378,N_10066,N_11434);
nand U14379 (N_14379,N_9643,N_9167);
and U14380 (N_14380,N_9877,N_10478);
or U14381 (N_14381,N_10163,N_10727);
and U14382 (N_14382,N_11024,N_10317);
nor U14383 (N_14383,N_9236,N_11417);
nor U14384 (N_14384,N_10611,N_9127);
and U14385 (N_14385,N_10046,N_9535);
nor U14386 (N_14386,N_10344,N_9778);
and U14387 (N_14387,N_10693,N_9104);
and U14388 (N_14388,N_11305,N_9713);
xnor U14389 (N_14389,N_11429,N_10217);
and U14390 (N_14390,N_9539,N_9234);
xnor U14391 (N_14391,N_10713,N_10321);
nor U14392 (N_14392,N_11367,N_11902);
and U14393 (N_14393,N_10680,N_9087);
xor U14394 (N_14394,N_10672,N_11655);
nand U14395 (N_14395,N_9854,N_10920);
xor U14396 (N_14396,N_11905,N_9727);
xor U14397 (N_14397,N_10048,N_10919);
or U14398 (N_14398,N_10156,N_11260);
and U14399 (N_14399,N_10658,N_10943);
nand U14400 (N_14400,N_11555,N_9661);
or U14401 (N_14401,N_9500,N_9963);
or U14402 (N_14402,N_11167,N_9177);
nand U14403 (N_14403,N_9321,N_9039);
nor U14404 (N_14404,N_11414,N_10024);
or U14405 (N_14405,N_10152,N_9064);
nor U14406 (N_14406,N_11560,N_9610);
nor U14407 (N_14407,N_10520,N_11849);
nand U14408 (N_14408,N_11301,N_11223);
nor U14409 (N_14409,N_9090,N_10736);
and U14410 (N_14410,N_10314,N_11971);
and U14411 (N_14411,N_9724,N_9529);
and U14412 (N_14412,N_11938,N_11669);
and U14413 (N_14413,N_9013,N_9330);
xor U14414 (N_14414,N_11439,N_10439);
nand U14415 (N_14415,N_11793,N_9961);
or U14416 (N_14416,N_10663,N_10173);
and U14417 (N_14417,N_11903,N_11051);
and U14418 (N_14418,N_11567,N_9189);
and U14419 (N_14419,N_10969,N_9098);
nand U14420 (N_14420,N_11939,N_10866);
nand U14421 (N_14421,N_11683,N_9768);
xnor U14422 (N_14422,N_10209,N_11444);
nor U14423 (N_14423,N_11219,N_10497);
and U14424 (N_14424,N_9619,N_9375);
and U14425 (N_14425,N_11336,N_11864);
xnor U14426 (N_14426,N_9190,N_10964);
or U14427 (N_14427,N_11985,N_9352);
nand U14428 (N_14428,N_9957,N_9418);
nand U14429 (N_14429,N_10969,N_11170);
and U14430 (N_14430,N_10306,N_10210);
xor U14431 (N_14431,N_9572,N_9762);
nand U14432 (N_14432,N_11880,N_10184);
or U14433 (N_14433,N_9053,N_10281);
nand U14434 (N_14434,N_9654,N_9685);
or U14435 (N_14435,N_9038,N_11970);
and U14436 (N_14436,N_10191,N_9474);
nor U14437 (N_14437,N_9635,N_11907);
and U14438 (N_14438,N_10109,N_10903);
xor U14439 (N_14439,N_9829,N_10288);
nor U14440 (N_14440,N_11820,N_10259);
nand U14441 (N_14441,N_11645,N_9377);
and U14442 (N_14442,N_10638,N_9532);
and U14443 (N_14443,N_10898,N_9565);
or U14444 (N_14444,N_11614,N_11727);
or U14445 (N_14445,N_9809,N_11285);
xor U14446 (N_14446,N_10854,N_9448);
nor U14447 (N_14447,N_9219,N_9045);
and U14448 (N_14448,N_11997,N_9028);
xnor U14449 (N_14449,N_10151,N_10939);
nand U14450 (N_14450,N_10721,N_9689);
nor U14451 (N_14451,N_10593,N_10099);
nand U14452 (N_14452,N_9624,N_10566);
nor U14453 (N_14453,N_10193,N_11094);
and U14454 (N_14454,N_11758,N_9474);
and U14455 (N_14455,N_10082,N_9221);
nand U14456 (N_14456,N_11006,N_9159);
nor U14457 (N_14457,N_11814,N_10040);
nand U14458 (N_14458,N_11516,N_9274);
or U14459 (N_14459,N_10301,N_10664);
nand U14460 (N_14460,N_9826,N_11693);
or U14461 (N_14461,N_9072,N_10672);
xor U14462 (N_14462,N_11123,N_9140);
nand U14463 (N_14463,N_9915,N_11133);
nand U14464 (N_14464,N_10556,N_10698);
nand U14465 (N_14465,N_9115,N_10757);
nor U14466 (N_14466,N_11416,N_10104);
nand U14467 (N_14467,N_10452,N_9840);
or U14468 (N_14468,N_10299,N_11370);
and U14469 (N_14469,N_11567,N_11968);
and U14470 (N_14470,N_10199,N_10303);
or U14471 (N_14471,N_10493,N_10658);
nor U14472 (N_14472,N_9116,N_10122);
and U14473 (N_14473,N_11407,N_9982);
xnor U14474 (N_14474,N_10984,N_10738);
nor U14475 (N_14475,N_9753,N_11118);
and U14476 (N_14476,N_11372,N_11711);
nor U14477 (N_14477,N_11168,N_11290);
xor U14478 (N_14478,N_10333,N_11424);
nand U14479 (N_14479,N_11049,N_11347);
and U14480 (N_14480,N_10423,N_10755);
nand U14481 (N_14481,N_9960,N_10534);
and U14482 (N_14482,N_11616,N_10186);
nor U14483 (N_14483,N_11137,N_11633);
and U14484 (N_14484,N_9107,N_10630);
nor U14485 (N_14485,N_9043,N_9338);
nor U14486 (N_14486,N_9302,N_9338);
or U14487 (N_14487,N_10625,N_11656);
and U14488 (N_14488,N_9638,N_10978);
nor U14489 (N_14489,N_10652,N_11523);
nand U14490 (N_14490,N_11757,N_10724);
xnor U14491 (N_14491,N_9367,N_9677);
nand U14492 (N_14492,N_10747,N_9895);
nand U14493 (N_14493,N_10350,N_10170);
nand U14494 (N_14494,N_10797,N_10285);
xnor U14495 (N_14495,N_11311,N_11733);
nor U14496 (N_14496,N_11196,N_9641);
nor U14497 (N_14497,N_11274,N_9206);
nor U14498 (N_14498,N_9703,N_9159);
or U14499 (N_14499,N_11271,N_10077);
xor U14500 (N_14500,N_10679,N_11721);
and U14501 (N_14501,N_10868,N_10842);
xor U14502 (N_14502,N_10032,N_10210);
nand U14503 (N_14503,N_9820,N_11175);
nand U14504 (N_14504,N_9959,N_9916);
and U14505 (N_14505,N_11411,N_9251);
xor U14506 (N_14506,N_9817,N_11066);
nand U14507 (N_14507,N_11064,N_10383);
nor U14508 (N_14508,N_9097,N_9629);
xnor U14509 (N_14509,N_10657,N_11608);
or U14510 (N_14510,N_10950,N_11486);
nor U14511 (N_14511,N_10716,N_10041);
or U14512 (N_14512,N_10258,N_11474);
and U14513 (N_14513,N_10540,N_10623);
or U14514 (N_14514,N_10018,N_10549);
nor U14515 (N_14515,N_9029,N_10336);
and U14516 (N_14516,N_10423,N_10797);
and U14517 (N_14517,N_11031,N_10052);
nand U14518 (N_14518,N_10119,N_10767);
nor U14519 (N_14519,N_10898,N_9010);
nor U14520 (N_14520,N_9356,N_9986);
or U14521 (N_14521,N_9102,N_10741);
and U14522 (N_14522,N_10904,N_11468);
nor U14523 (N_14523,N_11514,N_10059);
nor U14524 (N_14524,N_11026,N_10171);
or U14525 (N_14525,N_9098,N_9226);
or U14526 (N_14526,N_9229,N_9811);
nor U14527 (N_14527,N_10403,N_11595);
xnor U14528 (N_14528,N_9785,N_9325);
nor U14529 (N_14529,N_10970,N_9034);
and U14530 (N_14530,N_11079,N_11646);
nand U14531 (N_14531,N_9640,N_11561);
nand U14532 (N_14532,N_9145,N_10750);
or U14533 (N_14533,N_11672,N_10053);
xor U14534 (N_14534,N_11543,N_9648);
nand U14535 (N_14535,N_10352,N_11207);
nand U14536 (N_14536,N_9256,N_11392);
or U14537 (N_14537,N_10859,N_9941);
xnor U14538 (N_14538,N_9257,N_9771);
nand U14539 (N_14539,N_11015,N_9108);
xor U14540 (N_14540,N_9976,N_9016);
xor U14541 (N_14541,N_11054,N_11196);
and U14542 (N_14542,N_9236,N_11636);
nand U14543 (N_14543,N_10473,N_10330);
nor U14544 (N_14544,N_11762,N_10710);
nor U14545 (N_14545,N_11884,N_11849);
nand U14546 (N_14546,N_10614,N_9150);
nor U14547 (N_14547,N_11197,N_9876);
and U14548 (N_14548,N_11277,N_10448);
and U14549 (N_14549,N_11637,N_9613);
and U14550 (N_14550,N_9794,N_10677);
nand U14551 (N_14551,N_11740,N_11689);
nand U14552 (N_14552,N_10498,N_9978);
and U14553 (N_14553,N_11088,N_10980);
xor U14554 (N_14554,N_11383,N_9719);
nor U14555 (N_14555,N_11430,N_9466);
and U14556 (N_14556,N_10564,N_11495);
xnor U14557 (N_14557,N_9985,N_11274);
nand U14558 (N_14558,N_9437,N_10762);
nor U14559 (N_14559,N_11561,N_10116);
nand U14560 (N_14560,N_11042,N_9545);
nor U14561 (N_14561,N_10326,N_9326);
xor U14562 (N_14562,N_11171,N_11402);
nand U14563 (N_14563,N_10085,N_9096);
and U14564 (N_14564,N_10203,N_10224);
and U14565 (N_14565,N_10100,N_9020);
nand U14566 (N_14566,N_9866,N_11052);
xor U14567 (N_14567,N_9701,N_11783);
nand U14568 (N_14568,N_10697,N_11824);
nor U14569 (N_14569,N_10720,N_9416);
nand U14570 (N_14570,N_9400,N_11844);
and U14571 (N_14571,N_11717,N_10144);
nand U14572 (N_14572,N_11725,N_11498);
or U14573 (N_14573,N_11476,N_9246);
nor U14574 (N_14574,N_10275,N_9859);
and U14575 (N_14575,N_10257,N_11702);
and U14576 (N_14576,N_11001,N_11966);
nor U14577 (N_14577,N_9623,N_11031);
and U14578 (N_14578,N_9621,N_10715);
nor U14579 (N_14579,N_9652,N_11601);
xnor U14580 (N_14580,N_11827,N_9679);
nor U14581 (N_14581,N_11066,N_11139);
xnor U14582 (N_14582,N_9717,N_10500);
xor U14583 (N_14583,N_10845,N_11433);
nand U14584 (N_14584,N_11233,N_10270);
nand U14585 (N_14585,N_10128,N_11506);
nand U14586 (N_14586,N_9953,N_10017);
or U14587 (N_14587,N_11026,N_11518);
and U14588 (N_14588,N_11672,N_11352);
and U14589 (N_14589,N_11321,N_11012);
nor U14590 (N_14590,N_11579,N_11272);
xnor U14591 (N_14591,N_9533,N_10126);
nor U14592 (N_14592,N_11983,N_11040);
or U14593 (N_14593,N_11285,N_9994);
or U14594 (N_14594,N_9394,N_9423);
nor U14595 (N_14595,N_10731,N_9460);
nor U14596 (N_14596,N_10101,N_10219);
nand U14597 (N_14597,N_9821,N_11654);
and U14598 (N_14598,N_9421,N_11243);
xnor U14599 (N_14599,N_11099,N_10805);
nor U14600 (N_14600,N_11085,N_9018);
nor U14601 (N_14601,N_9198,N_11952);
xor U14602 (N_14602,N_11473,N_11724);
nor U14603 (N_14603,N_10195,N_10405);
and U14604 (N_14604,N_11312,N_11649);
xnor U14605 (N_14605,N_10216,N_9798);
nor U14606 (N_14606,N_10234,N_9557);
nand U14607 (N_14607,N_9433,N_9507);
nor U14608 (N_14608,N_9107,N_11359);
nor U14609 (N_14609,N_10047,N_11900);
and U14610 (N_14610,N_9860,N_11375);
nand U14611 (N_14611,N_9580,N_10670);
and U14612 (N_14612,N_10781,N_11082);
and U14613 (N_14613,N_9913,N_11111);
nor U14614 (N_14614,N_9394,N_10720);
xnor U14615 (N_14615,N_10902,N_11970);
and U14616 (N_14616,N_9537,N_9041);
nor U14617 (N_14617,N_11040,N_11854);
nand U14618 (N_14618,N_9412,N_10675);
nand U14619 (N_14619,N_11963,N_10666);
xor U14620 (N_14620,N_11287,N_11759);
nor U14621 (N_14621,N_9487,N_11967);
nand U14622 (N_14622,N_11308,N_9823);
nand U14623 (N_14623,N_9017,N_11699);
nor U14624 (N_14624,N_11370,N_10807);
and U14625 (N_14625,N_11675,N_11712);
xnor U14626 (N_14626,N_9709,N_11060);
and U14627 (N_14627,N_9124,N_9021);
nor U14628 (N_14628,N_9762,N_9443);
nand U14629 (N_14629,N_10410,N_11211);
nand U14630 (N_14630,N_9559,N_9096);
and U14631 (N_14631,N_10991,N_9161);
nor U14632 (N_14632,N_11468,N_11180);
or U14633 (N_14633,N_10991,N_11475);
xor U14634 (N_14634,N_11439,N_9835);
nor U14635 (N_14635,N_10669,N_11580);
nor U14636 (N_14636,N_11998,N_10382);
nor U14637 (N_14637,N_9573,N_9831);
nand U14638 (N_14638,N_9848,N_9661);
and U14639 (N_14639,N_10181,N_10894);
or U14640 (N_14640,N_11939,N_11653);
or U14641 (N_14641,N_10506,N_9250);
xor U14642 (N_14642,N_11098,N_10956);
or U14643 (N_14643,N_9606,N_9208);
or U14644 (N_14644,N_9554,N_9270);
and U14645 (N_14645,N_9661,N_11784);
or U14646 (N_14646,N_9856,N_9451);
or U14647 (N_14647,N_11631,N_10324);
xor U14648 (N_14648,N_9471,N_11502);
nand U14649 (N_14649,N_9411,N_9410);
nand U14650 (N_14650,N_9070,N_11423);
and U14651 (N_14651,N_9099,N_9629);
nor U14652 (N_14652,N_9848,N_9215);
xor U14653 (N_14653,N_9745,N_9876);
or U14654 (N_14654,N_11776,N_11878);
nor U14655 (N_14655,N_10931,N_10126);
xnor U14656 (N_14656,N_11325,N_11544);
nand U14657 (N_14657,N_10006,N_9464);
nand U14658 (N_14658,N_10696,N_10228);
or U14659 (N_14659,N_10705,N_9618);
nand U14660 (N_14660,N_11192,N_10994);
xor U14661 (N_14661,N_10816,N_9411);
and U14662 (N_14662,N_9448,N_10718);
nor U14663 (N_14663,N_9969,N_9786);
and U14664 (N_14664,N_9257,N_9464);
and U14665 (N_14665,N_10992,N_10163);
nor U14666 (N_14666,N_10494,N_10851);
or U14667 (N_14667,N_11148,N_9002);
and U14668 (N_14668,N_10684,N_9331);
and U14669 (N_14669,N_9575,N_10453);
xnor U14670 (N_14670,N_11863,N_10941);
or U14671 (N_14671,N_10821,N_11561);
xnor U14672 (N_14672,N_9364,N_11710);
xnor U14673 (N_14673,N_9784,N_9369);
nor U14674 (N_14674,N_9218,N_11833);
xor U14675 (N_14675,N_11631,N_11203);
nor U14676 (N_14676,N_11989,N_9814);
xor U14677 (N_14677,N_9549,N_11097);
or U14678 (N_14678,N_10581,N_10190);
and U14679 (N_14679,N_10378,N_11488);
nand U14680 (N_14680,N_11940,N_11541);
nor U14681 (N_14681,N_11349,N_10568);
nand U14682 (N_14682,N_10713,N_11774);
xnor U14683 (N_14683,N_9660,N_9332);
nand U14684 (N_14684,N_10863,N_9768);
xor U14685 (N_14685,N_11192,N_10545);
and U14686 (N_14686,N_10853,N_10133);
nor U14687 (N_14687,N_11496,N_10638);
or U14688 (N_14688,N_10168,N_9818);
and U14689 (N_14689,N_9256,N_10729);
nand U14690 (N_14690,N_11427,N_10056);
nand U14691 (N_14691,N_9273,N_10375);
or U14692 (N_14692,N_9765,N_9237);
or U14693 (N_14693,N_11770,N_9430);
or U14694 (N_14694,N_9257,N_11807);
nand U14695 (N_14695,N_11750,N_10687);
and U14696 (N_14696,N_10682,N_9646);
or U14697 (N_14697,N_9066,N_9115);
or U14698 (N_14698,N_11884,N_11780);
nand U14699 (N_14699,N_9714,N_11473);
nor U14700 (N_14700,N_11453,N_9293);
or U14701 (N_14701,N_9689,N_10166);
xor U14702 (N_14702,N_9732,N_11832);
nor U14703 (N_14703,N_10139,N_11310);
or U14704 (N_14704,N_10373,N_9152);
nor U14705 (N_14705,N_11651,N_9708);
or U14706 (N_14706,N_11043,N_11801);
nand U14707 (N_14707,N_10724,N_11914);
and U14708 (N_14708,N_10865,N_10036);
nand U14709 (N_14709,N_10590,N_9266);
or U14710 (N_14710,N_9022,N_10809);
or U14711 (N_14711,N_10036,N_10543);
nor U14712 (N_14712,N_11551,N_10464);
xor U14713 (N_14713,N_11435,N_11394);
xor U14714 (N_14714,N_9863,N_10316);
nor U14715 (N_14715,N_11810,N_11757);
nand U14716 (N_14716,N_9996,N_10411);
nand U14717 (N_14717,N_10433,N_10273);
nand U14718 (N_14718,N_9734,N_10097);
or U14719 (N_14719,N_9183,N_9695);
nand U14720 (N_14720,N_11348,N_10447);
nor U14721 (N_14721,N_9200,N_9862);
nor U14722 (N_14722,N_9680,N_10462);
nor U14723 (N_14723,N_10339,N_10482);
nor U14724 (N_14724,N_9704,N_9697);
or U14725 (N_14725,N_11531,N_10226);
nor U14726 (N_14726,N_11724,N_9113);
nand U14727 (N_14727,N_9332,N_10742);
and U14728 (N_14728,N_10575,N_10839);
xor U14729 (N_14729,N_9234,N_11055);
and U14730 (N_14730,N_10275,N_10248);
xnor U14731 (N_14731,N_9848,N_11997);
xnor U14732 (N_14732,N_10818,N_9836);
nor U14733 (N_14733,N_11318,N_9627);
and U14734 (N_14734,N_11072,N_11445);
or U14735 (N_14735,N_11842,N_11337);
or U14736 (N_14736,N_9228,N_10008);
and U14737 (N_14737,N_10863,N_9975);
and U14738 (N_14738,N_11180,N_11709);
and U14739 (N_14739,N_9501,N_11360);
and U14740 (N_14740,N_9530,N_10312);
nor U14741 (N_14741,N_11925,N_9302);
nor U14742 (N_14742,N_11331,N_9276);
or U14743 (N_14743,N_9809,N_11699);
nor U14744 (N_14744,N_11743,N_11605);
and U14745 (N_14745,N_9498,N_11520);
xnor U14746 (N_14746,N_9877,N_9160);
and U14747 (N_14747,N_9674,N_9700);
nor U14748 (N_14748,N_10607,N_9610);
nand U14749 (N_14749,N_10177,N_9937);
nor U14750 (N_14750,N_11307,N_10669);
and U14751 (N_14751,N_9690,N_11824);
and U14752 (N_14752,N_10028,N_10774);
and U14753 (N_14753,N_10707,N_11552);
nor U14754 (N_14754,N_9385,N_10035);
or U14755 (N_14755,N_9517,N_10864);
nand U14756 (N_14756,N_10684,N_9301);
nor U14757 (N_14757,N_10962,N_9577);
or U14758 (N_14758,N_9172,N_11542);
and U14759 (N_14759,N_10997,N_11086);
nor U14760 (N_14760,N_9094,N_9837);
and U14761 (N_14761,N_9291,N_9407);
xnor U14762 (N_14762,N_9492,N_10704);
nand U14763 (N_14763,N_9409,N_11119);
nor U14764 (N_14764,N_10956,N_11865);
or U14765 (N_14765,N_11504,N_9544);
xnor U14766 (N_14766,N_10638,N_10802);
and U14767 (N_14767,N_9053,N_11140);
nor U14768 (N_14768,N_10696,N_10900);
xor U14769 (N_14769,N_11869,N_10268);
or U14770 (N_14770,N_10070,N_10001);
and U14771 (N_14771,N_9906,N_10228);
nand U14772 (N_14772,N_9154,N_10768);
nand U14773 (N_14773,N_11623,N_10235);
xnor U14774 (N_14774,N_10619,N_9701);
nor U14775 (N_14775,N_11834,N_10287);
or U14776 (N_14776,N_9937,N_9914);
or U14777 (N_14777,N_9888,N_10811);
nor U14778 (N_14778,N_11716,N_11583);
nand U14779 (N_14779,N_9957,N_9736);
nand U14780 (N_14780,N_9404,N_11265);
or U14781 (N_14781,N_9909,N_10055);
xnor U14782 (N_14782,N_9361,N_11127);
or U14783 (N_14783,N_9608,N_10946);
nand U14784 (N_14784,N_10186,N_11751);
xnor U14785 (N_14785,N_9893,N_9377);
xnor U14786 (N_14786,N_9777,N_9363);
nor U14787 (N_14787,N_10073,N_11462);
nor U14788 (N_14788,N_9549,N_9655);
nand U14789 (N_14789,N_11658,N_11607);
and U14790 (N_14790,N_10297,N_11746);
nor U14791 (N_14791,N_9626,N_9016);
or U14792 (N_14792,N_11196,N_9789);
and U14793 (N_14793,N_9399,N_10269);
xnor U14794 (N_14794,N_10085,N_11530);
xor U14795 (N_14795,N_9310,N_11809);
nand U14796 (N_14796,N_11191,N_9352);
and U14797 (N_14797,N_11737,N_11829);
or U14798 (N_14798,N_11001,N_10120);
and U14799 (N_14799,N_9889,N_11207);
and U14800 (N_14800,N_9853,N_9665);
and U14801 (N_14801,N_10192,N_11785);
and U14802 (N_14802,N_9412,N_10771);
or U14803 (N_14803,N_11146,N_11423);
xnor U14804 (N_14804,N_10373,N_10385);
nand U14805 (N_14805,N_11830,N_11389);
xor U14806 (N_14806,N_10644,N_11121);
or U14807 (N_14807,N_10966,N_10281);
nand U14808 (N_14808,N_10884,N_9841);
nor U14809 (N_14809,N_9246,N_10630);
xor U14810 (N_14810,N_11890,N_10871);
nand U14811 (N_14811,N_9835,N_11751);
or U14812 (N_14812,N_10364,N_9960);
and U14813 (N_14813,N_10242,N_11203);
xnor U14814 (N_14814,N_11948,N_11138);
and U14815 (N_14815,N_10996,N_9349);
xnor U14816 (N_14816,N_11312,N_10342);
or U14817 (N_14817,N_10247,N_10676);
and U14818 (N_14818,N_9825,N_9487);
nor U14819 (N_14819,N_9217,N_10795);
and U14820 (N_14820,N_10165,N_10202);
nor U14821 (N_14821,N_11717,N_10538);
nor U14822 (N_14822,N_11021,N_10377);
nand U14823 (N_14823,N_9159,N_10314);
xnor U14824 (N_14824,N_9270,N_11186);
and U14825 (N_14825,N_10934,N_10809);
xnor U14826 (N_14826,N_9496,N_11388);
xnor U14827 (N_14827,N_10524,N_11833);
or U14828 (N_14828,N_10551,N_9177);
or U14829 (N_14829,N_10149,N_10941);
or U14830 (N_14830,N_11125,N_10202);
nor U14831 (N_14831,N_10295,N_11918);
nor U14832 (N_14832,N_10390,N_9250);
or U14833 (N_14833,N_10720,N_9278);
xnor U14834 (N_14834,N_9550,N_9317);
nand U14835 (N_14835,N_9365,N_9128);
nor U14836 (N_14836,N_11951,N_10937);
or U14837 (N_14837,N_10909,N_10302);
xor U14838 (N_14838,N_10785,N_9447);
xor U14839 (N_14839,N_9310,N_11611);
or U14840 (N_14840,N_10152,N_11926);
nor U14841 (N_14841,N_11578,N_10133);
or U14842 (N_14842,N_11095,N_10213);
and U14843 (N_14843,N_11235,N_9382);
or U14844 (N_14844,N_9567,N_9394);
or U14845 (N_14845,N_10999,N_10986);
or U14846 (N_14846,N_10176,N_10799);
and U14847 (N_14847,N_9647,N_9602);
nor U14848 (N_14848,N_10786,N_9473);
nand U14849 (N_14849,N_11934,N_9117);
nand U14850 (N_14850,N_11032,N_9296);
or U14851 (N_14851,N_11844,N_10266);
and U14852 (N_14852,N_10094,N_10698);
and U14853 (N_14853,N_10493,N_9487);
xor U14854 (N_14854,N_9511,N_10609);
or U14855 (N_14855,N_11772,N_11493);
and U14856 (N_14856,N_11004,N_11921);
and U14857 (N_14857,N_9408,N_9221);
nor U14858 (N_14858,N_11632,N_9894);
or U14859 (N_14859,N_10579,N_10478);
nand U14860 (N_14860,N_10282,N_9471);
nand U14861 (N_14861,N_9484,N_10913);
nor U14862 (N_14862,N_11931,N_10390);
xor U14863 (N_14863,N_10447,N_10550);
or U14864 (N_14864,N_9571,N_11810);
nand U14865 (N_14865,N_10836,N_10727);
nand U14866 (N_14866,N_9624,N_10010);
nor U14867 (N_14867,N_10728,N_11115);
nand U14868 (N_14868,N_11946,N_10502);
nand U14869 (N_14869,N_11313,N_11671);
or U14870 (N_14870,N_9018,N_11275);
and U14871 (N_14871,N_9323,N_9529);
xnor U14872 (N_14872,N_11498,N_11399);
and U14873 (N_14873,N_9951,N_9770);
or U14874 (N_14874,N_10287,N_11454);
or U14875 (N_14875,N_9149,N_10152);
and U14876 (N_14876,N_9146,N_11444);
nor U14877 (N_14877,N_11966,N_9362);
and U14878 (N_14878,N_9086,N_11834);
or U14879 (N_14879,N_9096,N_10474);
nor U14880 (N_14880,N_11368,N_10908);
xor U14881 (N_14881,N_9150,N_9142);
and U14882 (N_14882,N_11110,N_9225);
nor U14883 (N_14883,N_11918,N_10796);
and U14884 (N_14884,N_11937,N_11762);
nand U14885 (N_14885,N_9355,N_10254);
nand U14886 (N_14886,N_9428,N_10873);
and U14887 (N_14887,N_9650,N_10805);
or U14888 (N_14888,N_11152,N_9593);
and U14889 (N_14889,N_9220,N_10608);
or U14890 (N_14890,N_9459,N_11724);
and U14891 (N_14891,N_11170,N_11480);
or U14892 (N_14892,N_11975,N_9843);
or U14893 (N_14893,N_9830,N_11992);
and U14894 (N_14894,N_9421,N_11310);
or U14895 (N_14895,N_11315,N_9767);
nor U14896 (N_14896,N_9243,N_10770);
nand U14897 (N_14897,N_10261,N_10903);
nor U14898 (N_14898,N_10853,N_10939);
or U14899 (N_14899,N_11501,N_9025);
nand U14900 (N_14900,N_10524,N_10538);
and U14901 (N_14901,N_11619,N_11404);
or U14902 (N_14902,N_9240,N_10278);
nand U14903 (N_14903,N_11931,N_11860);
xor U14904 (N_14904,N_10060,N_11406);
or U14905 (N_14905,N_11589,N_11101);
and U14906 (N_14906,N_9017,N_10721);
and U14907 (N_14907,N_11397,N_10631);
and U14908 (N_14908,N_9060,N_11894);
nand U14909 (N_14909,N_10888,N_10322);
nand U14910 (N_14910,N_11900,N_10174);
or U14911 (N_14911,N_11238,N_11241);
or U14912 (N_14912,N_11573,N_11187);
xnor U14913 (N_14913,N_10518,N_9397);
and U14914 (N_14914,N_9987,N_11450);
xnor U14915 (N_14915,N_9099,N_11712);
xnor U14916 (N_14916,N_11830,N_10757);
or U14917 (N_14917,N_10768,N_10791);
nor U14918 (N_14918,N_9627,N_9677);
xnor U14919 (N_14919,N_10393,N_9676);
nor U14920 (N_14920,N_11748,N_11769);
and U14921 (N_14921,N_10233,N_11078);
and U14922 (N_14922,N_9220,N_10358);
nor U14923 (N_14923,N_11244,N_10179);
nand U14924 (N_14924,N_10598,N_9460);
or U14925 (N_14925,N_11133,N_11798);
and U14926 (N_14926,N_10590,N_11703);
or U14927 (N_14927,N_11060,N_9953);
nor U14928 (N_14928,N_10850,N_10840);
nand U14929 (N_14929,N_10525,N_9150);
and U14930 (N_14930,N_11096,N_9337);
and U14931 (N_14931,N_11316,N_11396);
or U14932 (N_14932,N_11871,N_11893);
or U14933 (N_14933,N_9707,N_9667);
and U14934 (N_14934,N_11144,N_10963);
nand U14935 (N_14935,N_9834,N_10996);
nor U14936 (N_14936,N_10395,N_11598);
nand U14937 (N_14937,N_10456,N_9236);
nand U14938 (N_14938,N_11711,N_11810);
or U14939 (N_14939,N_10225,N_10431);
nor U14940 (N_14940,N_9402,N_10036);
nand U14941 (N_14941,N_9715,N_11306);
xor U14942 (N_14942,N_9768,N_10082);
xnor U14943 (N_14943,N_9577,N_11812);
or U14944 (N_14944,N_10298,N_11445);
nand U14945 (N_14945,N_9720,N_9476);
and U14946 (N_14946,N_9365,N_10795);
nand U14947 (N_14947,N_10478,N_9956);
and U14948 (N_14948,N_9457,N_10122);
xor U14949 (N_14949,N_11964,N_10502);
and U14950 (N_14950,N_9699,N_10949);
or U14951 (N_14951,N_11279,N_10132);
nand U14952 (N_14952,N_10513,N_9944);
and U14953 (N_14953,N_10868,N_10377);
and U14954 (N_14954,N_11866,N_10808);
nand U14955 (N_14955,N_10762,N_10111);
or U14956 (N_14956,N_10196,N_9673);
nor U14957 (N_14957,N_10789,N_9526);
xor U14958 (N_14958,N_10935,N_10829);
xor U14959 (N_14959,N_11217,N_9513);
xor U14960 (N_14960,N_9468,N_11537);
nand U14961 (N_14961,N_9508,N_10095);
and U14962 (N_14962,N_10123,N_11636);
and U14963 (N_14963,N_10667,N_11243);
nor U14964 (N_14964,N_9025,N_9255);
nand U14965 (N_14965,N_11209,N_11440);
xnor U14966 (N_14966,N_10744,N_10351);
and U14967 (N_14967,N_10263,N_11621);
and U14968 (N_14968,N_9382,N_11632);
nand U14969 (N_14969,N_11535,N_10126);
nand U14970 (N_14970,N_11099,N_9100);
nand U14971 (N_14971,N_10957,N_10290);
xor U14972 (N_14972,N_10245,N_9041);
xnor U14973 (N_14973,N_11189,N_11677);
nand U14974 (N_14974,N_10171,N_11963);
and U14975 (N_14975,N_10761,N_9597);
nand U14976 (N_14976,N_9921,N_9587);
xnor U14977 (N_14977,N_10160,N_10882);
xnor U14978 (N_14978,N_9147,N_10645);
nand U14979 (N_14979,N_10177,N_10575);
and U14980 (N_14980,N_10945,N_9007);
nor U14981 (N_14981,N_10547,N_9819);
and U14982 (N_14982,N_11326,N_11304);
or U14983 (N_14983,N_9738,N_10987);
nand U14984 (N_14984,N_11343,N_9971);
or U14985 (N_14985,N_11415,N_9719);
or U14986 (N_14986,N_10131,N_9169);
nand U14987 (N_14987,N_9640,N_11189);
nor U14988 (N_14988,N_9548,N_11249);
xnor U14989 (N_14989,N_10582,N_11313);
nor U14990 (N_14990,N_10440,N_9136);
nand U14991 (N_14991,N_11708,N_11837);
and U14992 (N_14992,N_10953,N_11677);
or U14993 (N_14993,N_10730,N_10227);
and U14994 (N_14994,N_9238,N_10501);
and U14995 (N_14995,N_9565,N_9356);
nor U14996 (N_14996,N_11373,N_11287);
or U14997 (N_14997,N_11776,N_10942);
xnor U14998 (N_14998,N_10757,N_9382);
nand U14999 (N_14999,N_9224,N_9533);
or U15000 (N_15000,N_13673,N_14239);
nor U15001 (N_15001,N_13114,N_14937);
or U15002 (N_15002,N_13829,N_13421);
nor U15003 (N_15003,N_12763,N_12936);
and U15004 (N_15004,N_14297,N_14316);
xor U15005 (N_15005,N_12105,N_13739);
or U15006 (N_15006,N_13084,N_13012);
and U15007 (N_15007,N_14412,N_14836);
nor U15008 (N_15008,N_12403,N_12682);
nor U15009 (N_15009,N_14182,N_14685);
or U15010 (N_15010,N_14413,N_14011);
and U15011 (N_15011,N_13688,N_13862);
nand U15012 (N_15012,N_13659,N_13431);
and U15013 (N_15013,N_14112,N_14126);
nand U15014 (N_15014,N_12008,N_13605);
nand U15015 (N_15015,N_13637,N_12916);
or U15016 (N_15016,N_14600,N_12494);
and U15017 (N_15017,N_12171,N_12317);
and U15018 (N_15018,N_14722,N_13093);
nand U15019 (N_15019,N_14441,N_12999);
xnor U15020 (N_15020,N_13604,N_13334);
and U15021 (N_15021,N_12113,N_12125);
or U15022 (N_15022,N_14783,N_13641);
or U15023 (N_15023,N_13456,N_13546);
xnor U15024 (N_15024,N_14569,N_14073);
or U15025 (N_15025,N_13824,N_13667);
nor U15026 (N_15026,N_12577,N_12284);
nand U15027 (N_15027,N_13757,N_13043);
or U15028 (N_15028,N_12003,N_13141);
or U15029 (N_15029,N_14451,N_12543);
xor U15030 (N_15030,N_14625,N_13991);
nor U15031 (N_15031,N_12186,N_14709);
or U15032 (N_15032,N_12115,N_14482);
and U15033 (N_15033,N_14474,N_14640);
nand U15034 (N_15034,N_12055,N_14276);
nand U15035 (N_15035,N_12587,N_12597);
xor U15036 (N_15036,N_14853,N_12191);
and U15037 (N_15037,N_14531,N_13969);
or U15038 (N_15038,N_13398,N_12004);
or U15039 (N_15039,N_13860,N_14325);
nor U15040 (N_15040,N_13483,N_13965);
or U15041 (N_15041,N_13014,N_13317);
nor U15042 (N_15042,N_12283,N_13285);
and U15043 (N_15043,N_12194,N_13802);
xor U15044 (N_15044,N_13407,N_14875);
xor U15045 (N_15045,N_12993,N_14938);
and U15046 (N_15046,N_14442,N_13235);
nor U15047 (N_15047,N_12820,N_13409);
nor U15048 (N_15048,N_12533,N_12301);
xor U15049 (N_15049,N_12904,N_12336);
xor U15050 (N_15050,N_12885,N_13689);
nor U15051 (N_15051,N_13946,N_12552);
nand U15052 (N_15052,N_12431,N_14496);
nand U15053 (N_15053,N_13226,N_14332);
nor U15054 (N_15054,N_12232,N_13386);
nand U15055 (N_15055,N_13397,N_13363);
or U15056 (N_15056,N_12260,N_13265);
and U15057 (N_15057,N_14661,N_14019);
xnor U15058 (N_15058,N_14494,N_14289);
nand U15059 (N_15059,N_13022,N_12505);
nor U15060 (N_15060,N_13584,N_12347);
xor U15061 (N_15061,N_13760,N_14885);
nor U15062 (N_15062,N_13052,N_12281);
nor U15063 (N_15063,N_13685,N_12429);
or U15064 (N_15064,N_13183,N_14717);
xor U15065 (N_15065,N_14448,N_13212);
xor U15066 (N_15066,N_13968,N_14894);
xor U15067 (N_15067,N_12894,N_12743);
nor U15068 (N_15068,N_14232,N_12493);
or U15069 (N_15069,N_13635,N_13440);
and U15070 (N_15070,N_14207,N_12244);
nor U15071 (N_15071,N_14897,N_12868);
xor U15072 (N_15072,N_12783,N_13989);
nor U15073 (N_15073,N_13799,N_12927);
or U15074 (N_15074,N_14830,N_14698);
nor U15075 (N_15075,N_13316,N_12741);
nand U15076 (N_15076,N_13875,N_13289);
nor U15077 (N_15077,N_14994,N_14725);
and U15078 (N_15078,N_13237,N_14505);
nand U15079 (N_15079,N_12684,N_12188);
nand U15080 (N_15080,N_12935,N_14014);
xnor U15081 (N_15081,N_12831,N_12507);
nand U15082 (N_15082,N_13777,N_13649);
nand U15083 (N_15083,N_14389,N_14761);
or U15084 (N_15084,N_12753,N_14032);
or U15085 (N_15085,N_12242,N_13896);
and U15086 (N_15086,N_14330,N_14561);
xnor U15087 (N_15087,N_14731,N_14815);
and U15088 (N_15088,N_14406,N_12071);
or U15089 (N_15089,N_13894,N_13331);
nor U15090 (N_15090,N_12848,N_12189);
or U15091 (N_15091,N_13501,N_12560);
and U15092 (N_15092,N_13510,N_13458);
nand U15093 (N_15093,N_12442,N_13203);
nand U15094 (N_15094,N_12694,N_12160);
and U15095 (N_15095,N_14873,N_14341);
or U15096 (N_15096,N_13074,N_13932);
or U15097 (N_15097,N_14596,N_13197);
and U15098 (N_15098,N_13952,N_13847);
or U15099 (N_15099,N_12031,N_14870);
xor U15100 (N_15100,N_13511,N_12340);
nor U15101 (N_15101,N_12022,N_13157);
nor U15102 (N_15102,N_13962,N_14492);
nand U15103 (N_15103,N_14410,N_12561);
or U15104 (N_15104,N_12940,N_14762);
xor U15105 (N_15105,N_12933,N_12314);
nor U15106 (N_15106,N_13481,N_12046);
and U15107 (N_15107,N_12737,N_14270);
and U15108 (N_15108,N_13999,N_12406);
and U15109 (N_15109,N_13547,N_14540);
nand U15110 (N_15110,N_13545,N_14524);
or U15111 (N_15111,N_12359,N_13292);
nand U15112 (N_15112,N_12615,N_12106);
xnor U15113 (N_15113,N_14757,N_12161);
nor U15114 (N_15114,N_12149,N_12591);
nor U15115 (N_15115,N_14529,N_13206);
or U15116 (N_15116,N_13949,N_12256);
xor U15117 (N_15117,N_14384,N_13240);
and U15118 (N_15118,N_13929,N_12837);
nand U15119 (N_15119,N_14321,N_13256);
nor U15120 (N_15120,N_13615,N_12129);
xor U15121 (N_15121,N_12768,N_12382);
xor U15122 (N_15122,N_14576,N_14436);
nand U15123 (N_15123,N_12104,N_12832);
and U15124 (N_15124,N_12423,N_12265);
xor U15125 (N_15125,N_13709,N_12328);
nor U15126 (N_15126,N_14613,N_12872);
nand U15127 (N_15127,N_14103,N_12599);
and U15128 (N_15128,N_13057,N_12653);
nor U15129 (N_15129,N_13764,N_13478);
nor U15130 (N_15130,N_14479,N_12729);
nor U15131 (N_15131,N_12208,N_13262);
nand U15132 (N_15132,N_14047,N_14707);
and U15133 (N_15133,N_14714,N_14984);
nand U15134 (N_15134,N_14301,N_13128);
nor U15135 (N_15135,N_12042,N_12020);
nor U15136 (N_15136,N_14280,N_13063);
xor U15137 (N_15137,N_12452,N_12138);
xnor U15138 (N_15138,N_14752,N_13914);
nand U15139 (N_15139,N_13002,N_12723);
or U15140 (N_15140,N_12642,N_14932);
xor U15141 (N_15141,N_14858,N_14295);
and U15142 (N_15142,N_14951,N_12175);
nand U15143 (N_15143,N_12229,N_13352);
nand U15144 (N_15144,N_13681,N_12294);
or U15145 (N_15145,N_13745,N_14357);
nor U15146 (N_15146,N_12972,N_12035);
nand U15147 (N_15147,N_13536,N_13754);
nand U15148 (N_15148,N_13789,N_13936);
and U15149 (N_15149,N_13840,N_14493);
nand U15150 (N_15150,N_13109,N_14857);
or U15151 (N_15151,N_13761,N_14883);
nand U15152 (N_15152,N_14835,N_14310);
nand U15153 (N_15153,N_14303,N_14539);
xor U15154 (N_15154,N_12366,N_13294);
or U15155 (N_15155,N_12291,N_12482);
nand U15156 (N_15156,N_12805,N_14005);
xor U15157 (N_15157,N_12226,N_12475);
nor U15158 (N_15158,N_12293,N_14841);
or U15159 (N_15159,N_12784,N_13140);
xor U15160 (N_15160,N_13696,N_12953);
or U15161 (N_15161,N_14801,N_13987);
xnor U15162 (N_15162,N_13198,N_12914);
or U15163 (N_15163,N_14425,N_14433);
nor U15164 (N_15164,N_14086,N_13476);
nor U15165 (N_15165,N_14485,N_13768);
nor U15166 (N_15166,N_12401,N_12801);
and U15167 (N_15167,N_13550,N_14864);
and U15168 (N_15168,N_13746,N_12398);
and U15169 (N_15169,N_12414,N_12666);
xor U15170 (N_15170,N_12376,N_12140);
nor U15171 (N_15171,N_14254,N_12379);
xnor U15172 (N_15172,N_14924,N_14810);
nor U15173 (N_15173,N_13591,N_13272);
and U15174 (N_15174,N_12739,N_13678);
or U15175 (N_15175,N_14617,N_12154);
nand U15176 (N_15176,N_14142,N_14712);
nand U15177 (N_15177,N_12459,N_12799);
nor U15178 (N_15178,N_13357,N_12973);
nand U15179 (N_15179,N_14128,N_14151);
nand U15180 (N_15180,N_13158,N_13100);
nor U15181 (N_15181,N_12588,N_13007);
xor U15182 (N_15182,N_14072,N_14519);
nor U15183 (N_15183,N_13451,N_13921);
and U15184 (N_15184,N_12852,N_12633);
xnor U15185 (N_15185,N_14087,N_13454);
nand U15186 (N_15186,N_12077,N_14631);
or U15187 (N_15187,N_13137,N_12460);
nand U15188 (N_15188,N_13135,N_14085);
nor U15189 (N_15189,N_13617,N_12703);
or U15190 (N_15190,N_13477,N_14383);
nor U15191 (N_15191,N_13561,N_13793);
xor U15192 (N_15192,N_13504,N_12818);
xnor U15193 (N_15193,N_12108,N_12043);
nand U15194 (N_15194,N_12133,N_12664);
nor U15195 (N_15195,N_14510,N_14823);
and U15196 (N_15196,N_14998,N_13601);
nand U15197 (N_15197,N_13134,N_13060);
and U15198 (N_15198,N_12255,N_14216);
nand U15199 (N_15199,N_12963,N_13775);
nand U15200 (N_15200,N_12209,N_13411);
or U15201 (N_15201,N_13147,N_14096);
nor U15202 (N_15202,N_14525,N_13049);
and U15203 (N_15203,N_12767,N_13073);
xor U15204 (N_15204,N_12858,N_14738);
nand U15205 (N_15205,N_13525,N_14246);
nor U15206 (N_15206,N_13078,N_13691);
nor U15207 (N_15207,N_13161,N_14397);
and U15208 (N_15208,N_13654,N_13018);
nor U15209 (N_15209,N_14804,N_13836);
or U15210 (N_15210,N_12902,N_12861);
xnor U15211 (N_15211,N_12248,N_12326);
xor U15212 (N_15212,N_13827,N_12481);
nor U15213 (N_15213,N_13027,N_12227);
nor U15214 (N_15214,N_13121,N_12596);
nand U15215 (N_15215,N_13001,N_13770);
xor U15216 (N_15216,N_13807,N_14826);
and U15217 (N_15217,N_13033,N_13371);
nor U15218 (N_15218,N_12734,N_13152);
or U15219 (N_15219,N_14748,N_13111);
and U15220 (N_15220,N_12532,N_14775);
or U15221 (N_15221,N_14939,N_12345);
nor U15222 (N_15222,N_12199,N_14820);
nand U15223 (N_15223,N_14809,N_14274);
xnor U15224 (N_15224,N_14922,N_14620);
xor U15225 (N_15225,N_14318,N_13488);
nor U15226 (N_15226,N_12950,N_14509);
and U15227 (N_15227,N_14997,N_13179);
and U15228 (N_15228,N_14372,N_14555);
or U15229 (N_15229,N_12254,N_12637);
or U15230 (N_15230,N_12766,N_14037);
nor U15231 (N_15231,N_12023,N_13077);
and U15232 (N_15232,N_14674,N_12860);
and U15233 (N_15233,N_14257,N_13716);
nand U15234 (N_15234,N_13951,N_12887);
and U15235 (N_15235,N_13577,N_12444);
nor U15236 (N_15236,N_13148,N_14486);
nand U15237 (N_15237,N_13647,N_12378);
and U15238 (N_15238,N_14568,N_14976);
or U15239 (N_15239,N_12526,N_13192);
nor U15240 (N_15240,N_13805,N_14075);
nand U15241 (N_15241,N_14850,N_13722);
nor U15242 (N_15242,N_13436,N_13580);
and U15243 (N_15243,N_12795,N_14470);
and U15244 (N_15244,N_13338,N_14007);
or U15245 (N_15245,N_13959,N_14822);
and U15246 (N_15246,N_13642,N_12117);
xnor U15247 (N_15247,N_14376,N_12467);
nor U15248 (N_15248,N_14958,N_12177);
nand U15249 (N_15249,N_14169,N_13420);
and U15250 (N_15250,N_14109,N_12236);
and U15251 (N_15251,N_14584,N_14347);
xnor U15252 (N_15252,N_12478,N_12280);
xor U15253 (N_15253,N_13964,N_13005);
or U15254 (N_15254,N_12400,N_12508);
nand U15255 (N_15255,N_14727,N_12640);
nor U15256 (N_15256,N_12439,N_13699);
xnor U15257 (N_15257,N_14803,N_14528);
nand U15258 (N_15258,N_12365,N_14351);
nand U15259 (N_15259,N_14691,N_14814);
nor U15260 (N_15260,N_14445,N_13231);
nand U15261 (N_15261,N_13487,N_12924);
nor U15262 (N_15262,N_12941,N_14025);
xor U15263 (N_15263,N_13070,N_14137);
and U15264 (N_15264,N_14668,N_14118);
xor U15265 (N_15265,N_14354,N_13657);
nand U15266 (N_15266,N_14192,N_12926);
and U15267 (N_15267,N_13622,N_12093);
and U15268 (N_15268,N_12908,N_13903);
xnor U15269 (N_15269,N_12221,N_14656);
or U15270 (N_15270,N_14946,N_14154);
and U15271 (N_15271,N_14364,N_12779);
nand U15272 (N_15272,N_12152,N_14959);
or U15273 (N_15273,N_12752,N_12083);
or U15274 (N_15274,N_12390,N_14972);
nor U15275 (N_15275,N_12794,N_14834);
xor U15276 (N_15276,N_13835,N_12495);
nand U15277 (N_15277,N_12239,N_14664);
or U15278 (N_15278,N_12688,N_12346);
or U15279 (N_15279,N_14807,N_13261);
and U15280 (N_15280,N_12305,N_13865);
or U15281 (N_15281,N_12590,N_13132);
or U15282 (N_15282,N_14653,N_14601);
xnor U15283 (N_15283,N_14292,N_12012);
and U15284 (N_15284,N_12971,N_13613);
or U15285 (N_15285,N_12869,N_12367);
nor U15286 (N_15286,N_12215,N_13742);
nor U15287 (N_15287,N_14267,N_14964);
nor U15288 (N_15288,N_12958,N_13496);
and U15289 (N_15289,N_14871,N_14700);
xnor U15290 (N_15290,N_14056,N_13733);
xor U15291 (N_15291,N_13195,N_13297);
or U15292 (N_15292,N_13505,N_14993);
xor U15293 (N_15293,N_14657,N_14012);
and U15294 (N_15294,N_14751,N_14468);
xor U15295 (N_15295,N_13718,N_14061);
nor U15296 (N_15296,N_13643,N_13349);
nor U15297 (N_15297,N_14624,N_12811);
and U15298 (N_15298,N_13234,N_14305);
and U15299 (N_15299,N_12079,N_12812);
nand U15300 (N_15300,N_13176,N_13337);
nor U15301 (N_15301,N_14405,N_13028);
nand U15302 (N_15302,N_14840,N_12519);
nand U15303 (N_15303,N_14888,N_14264);
or U15304 (N_15304,N_13223,N_12807);
or U15305 (N_15305,N_14309,N_12939);
nand U15306 (N_15306,N_14400,N_14298);
and U15307 (N_15307,N_12344,N_13000);
xnor U15308 (N_15308,N_12484,N_12730);
nand U15309 (N_15309,N_12318,N_12517);
and U15310 (N_15310,N_13821,N_12037);
nand U15311 (N_15311,N_13211,N_12700);
xor U15312 (N_15312,N_13646,N_12893);
nand U15313 (N_15313,N_12604,N_13246);
xnor U15314 (N_15314,N_14222,N_12196);
or U15315 (N_15315,N_12462,N_14575);
nand U15316 (N_15316,N_13486,N_13774);
or U15317 (N_15317,N_13834,N_14003);
nand U15318 (N_15318,N_13600,N_13755);
xnor U15319 (N_15319,N_13912,N_12915);
and U15320 (N_15320,N_14419,N_13815);
nand U15321 (N_15321,N_12369,N_14963);
or U15322 (N_15322,N_12976,N_13849);
or U15323 (N_15323,N_12551,N_13380);
nor U15324 (N_15324,N_13396,N_14114);
nor U15325 (N_15325,N_12165,N_12128);
nor U15326 (N_15326,N_13323,N_12479);
nand U15327 (N_15327,N_12372,N_12488);
nand U15328 (N_15328,N_12896,N_12120);
nor U15329 (N_15329,N_13618,N_14370);
nor U15330 (N_15330,N_14824,N_13167);
and U15331 (N_15331,N_14350,N_12297);
or U15332 (N_15332,N_13009,N_13326);
nor U15333 (N_15333,N_13971,N_12824);
nor U15334 (N_15334,N_14877,N_14346);
xnor U15335 (N_15335,N_14477,N_13820);
or U15336 (N_15336,N_14326,N_14024);
nor U15337 (N_15337,N_14084,N_13187);
nor U15338 (N_15338,N_13258,N_12449);
nor U15339 (N_15339,N_13166,N_12947);
nand U15340 (N_15340,N_12357,N_13529);
or U15341 (N_15341,N_12485,N_13332);
nor U15342 (N_15342,N_14193,N_14224);
xnor U15343 (N_15343,N_12780,N_12450);
nor U15344 (N_15344,N_13651,N_13494);
nor U15345 (N_15345,N_12015,N_12881);
and U15346 (N_15346,N_12573,N_12930);
nand U15347 (N_15347,N_14452,N_14812);
nand U15348 (N_15348,N_12471,N_14818);
nand U15349 (N_15349,N_14892,N_12850);
nand U15350 (N_15350,N_13705,N_12056);
or U15351 (N_15351,N_14360,N_12074);
xnor U15352 (N_15352,N_13645,N_12182);
nand U15353 (N_15353,N_14627,N_14049);
nor U15354 (N_15354,N_14184,N_13471);
xnor U15355 (N_15355,N_14427,N_14793);
nor U15356 (N_15356,N_14837,N_12644);
xnor U15357 (N_15357,N_12970,N_13679);
xor U15358 (N_15358,N_12570,N_14827);
nor U15359 (N_15359,N_12143,N_14337);
nand U15360 (N_15360,N_14764,N_12135);
nor U15361 (N_15361,N_12103,N_13650);
nand U15362 (N_15362,N_12262,N_12412);
xnor U15363 (N_15363,N_12327,N_13627);
nor U15364 (N_15364,N_14382,N_12628);
xor U15365 (N_15365,N_13828,N_12081);
nand U15366 (N_15366,N_14031,N_14038);
xor U15367 (N_15367,N_14729,N_12067);
xnor U15368 (N_15368,N_12536,N_12612);
nand U15369 (N_15369,N_14265,N_12371);
and U15370 (N_15370,N_12525,N_12000);
or U15371 (N_15371,N_12068,N_12058);
and U15372 (N_15372,N_14407,N_13098);
xor U15373 (N_15373,N_12960,N_14516);
nor U15374 (N_15374,N_12629,N_12237);
xor U15375 (N_15375,N_12986,N_14683);
xor U15376 (N_15376,N_13762,N_14272);
nand U15377 (N_15377,N_14900,N_12178);
nand U15378 (N_15378,N_12121,N_14366);
nand U15379 (N_15379,N_14753,N_12697);
and U15380 (N_15380,N_14015,N_13153);
nor U15381 (N_15381,N_14632,N_14317);
and U15382 (N_15382,N_13184,N_13703);
and U15383 (N_15383,N_12205,N_13720);
or U15384 (N_15384,N_13120,N_14832);
xnor U15385 (N_15385,N_13741,N_12251);
nand U15386 (N_15386,N_13302,N_12553);
xnor U15387 (N_15387,N_12009,N_13418);
xnor U15388 (N_15388,N_13706,N_12578);
and U15389 (N_15389,N_12010,N_12034);
xor U15390 (N_15390,N_12631,N_13123);
and U15391 (N_15391,N_14570,N_13978);
xnor U15392 (N_15392,N_14985,N_13267);
nand U15393 (N_15393,N_12634,N_12252);
and U15394 (N_15394,N_12951,N_12912);
nor U15395 (N_15395,N_14846,N_13259);
nand U15396 (N_15396,N_12102,N_14538);
and U15397 (N_15397,N_13264,N_14898);
nand U15398 (N_15398,N_13410,N_14769);
or U15399 (N_15399,N_13424,N_14797);
or U15400 (N_15400,N_13698,N_13562);
or U15401 (N_15401,N_14173,N_14484);
nand U15402 (N_15402,N_13489,N_13899);
or U15403 (N_15403,N_14549,N_13778);
and U15404 (N_15404,N_14336,N_14062);
nor U15405 (N_15405,N_12892,N_12621);
nand U15406 (N_15406,N_13151,N_13570);
or U15407 (N_15407,N_13794,N_14237);
and U15408 (N_15408,N_12446,N_12945);
xnor U15409 (N_15409,N_12396,N_14881);
and U15410 (N_15410,N_12061,N_14721);
nor U15411 (N_15411,N_14308,N_12504);
and U15412 (N_15412,N_12421,N_13887);
nand U15413 (N_15413,N_12555,N_14426);
and U15414 (N_15414,N_14618,N_12172);
nand U15415 (N_15415,N_14473,N_12410);
xor U15416 (N_15416,N_13110,N_13099);
nand U15417 (N_15417,N_14682,N_13516);
nand U15418 (N_15418,N_14578,N_14566);
nand U15419 (N_15419,N_13990,N_12044);
or U15420 (N_15420,N_13146,N_12674);
and U15421 (N_15421,N_12139,N_12325);
nand U15422 (N_15422,N_13886,N_13950);
and U15423 (N_15423,N_12045,N_13353);
nand U15424 (N_15424,N_12298,N_12802);
or U15425 (N_15425,N_12557,N_12777);
xnor U15426 (N_15426,N_13734,N_13801);
and U15427 (N_15427,N_14890,N_14490);
or U15428 (N_15428,N_13631,N_12238);
nor U15429 (N_15429,N_12920,N_13305);
nor U15430 (N_15430,N_14307,N_14511);
or U15431 (N_15431,N_12047,N_12875);
xor U15432 (N_15432,N_13871,N_12091);
nand U15433 (N_15433,N_14608,N_13020);
nand U15434 (N_15434,N_14811,N_12127);
nand U15435 (N_15435,N_13541,N_13927);
xnor U15436 (N_15436,N_14928,N_13872);
or U15437 (N_15437,N_14284,N_14115);
or U15438 (N_15438,N_14587,N_13714);
xnor U15439 (N_15439,N_12392,N_14686);
or U15440 (N_15440,N_12381,N_14536);
and U15441 (N_15441,N_13596,N_12635);
nand U15442 (N_15442,N_14716,N_14230);
nor U15443 (N_15443,N_12871,N_12051);
and U15444 (N_15444,N_12545,N_14915);
and U15445 (N_15445,N_13830,N_13245);
nor U15446 (N_15446,N_12322,N_14472);
and U15447 (N_15447,N_14718,N_12863);
nor U15448 (N_15448,N_13817,N_13026);
and U15449 (N_15449,N_13974,N_13031);
or U15450 (N_15450,N_14375,N_14863);
or U15451 (N_15451,N_12918,N_14217);
and U15452 (N_15452,N_14340,N_12413);
or U15453 (N_15453,N_14008,N_12619);
or U15454 (N_15454,N_12388,N_13016);
nand U15455 (N_15455,N_13064,N_14211);
xor U15456 (N_15456,N_13254,N_14663);
xor U15457 (N_15457,N_13606,N_13837);
nand U15458 (N_15458,N_14423,N_14331);
and U15459 (N_15459,N_14696,N_13611);
nor U15460 (N_15460,N_14323,N_13960);
and U15461 (N_15461,N_13599,N_14550);
nor U15462 (N_15462,N_12416,N_14101);
nand U15463 (N_15463,N_13908,N_13520);
xor U15464 (N_15464,N_13780,N_14659);
nor U15465 (N_15465,N_14560,N_13091);
xor U15466 (N_15466,N_13178,N_12220);
or U15467 (N_15467,N_13663,N_13958);
nor U15468 (N_15468,N_14638,N_14223);
nor U15469 (N_15469,N_13055,N_14278);
nor U15470 (N_15470,N_14458,N_13988);
nand U15471 (N_15471,N_13573,N_13416);
nor U15472 (N_15472,N_13973,N_12393);
nor U15473 (N_15473,N_12758,N_12897);
and U15474 (N_15474,N_13181,N_12564);
nor U15475 (N_15475,N_14076,N_13842);
and U15476 (N_15476,N_14228,N_14693);
and U15477 (N_15477,N_13839,N_14141);
nand U15478 (N_15478,N_12876,N_12692);
nor U15479 (N_15479,N_12002,N_12668);
nand U15480 (N_15480,N_12306,N_12955);
xor U15481 (N_15481,N_12595,N_14943);
xor U15482 (N_15482,N_14121,N_13552);
xor U15483 (N_15483,N_12681,N_14028);
nor U15484 (N_15484,N_14291,N_13271);
xor U15485 (N_15485,N_13163,N_14678);
nor U15486 (N_15486,N_14842,N_13373);
xnor U15487 (N_15487,N_13751,N_13788);
xor U15488 (N_15488,N_13662,N_14615);
nand U15489 (N_15489,N_12962,N_13207);
nand U15490 (N_15490,N_12276,N_13926);
and U15491 (N_15491,N_14602,N_12593);
xnor U15492 (N_15492,N_12632,N_13438);
or U15493 (N_15493,N_12320,N_14833);
xor U15494 (N_15494,N_14934,N_12840);
and U15495 (N_15495,N_14843,N_13406);
or U15496 (N_15496,N_14750,N_14929);
or U15497 (N_15497,N_13518,N_12053);
nor U15498 (N_15498,N_12898,N_13215);
nor U15499 (N_15499,N_14009,N_12202);
or U15500 (N_15500,N_13869,N_13726);
nand U15501 (N_15501,N_13076,N_13355);
nor U15502 (N_15502,N_13779,N_12755);
xor U15503 (N_15503,N_14160,N_12639);
nor U15504 (N_15504,N_13066,N_13776);
nand U15505 (N_15505,N_14467,N_14981);
xnor U15506 (N_15506,N_13360,N_12538);
and U15507 (N_15507,N_13329,N_14447);
nand U15508 (N_15508,N_12007,N_13602);
nand U15509 (N_15509,N_14099,N_12486);
nor U15510 (N_15510,N_12770,N_12522);
nor U15511 (N_15511,N_12200,N_14925);
and U15512 (N_15512,N_14065,N_12052);
nand U15513 (N_15513,N_12050,N_12706);
xnor U15514 (N_15514,N_13164,N_14562);
and U15515 (N_15515,N_14438,N_12606);
or U15516 (N_15516,N_14785,N_12821);
or U15517 (N_15517,N_13150,N_14595);
or U15518 (N_15518,N_14146,N_12563);
nor U15519 (N_15519,N_13484,N_14935);
and U15520 (N_15520,N_14196,N_13819);
nand U15521 (N_15521,N_12339,N_12195);
and U15522 (N_15522,N_14860,N_12019);
and U15523 (N_15523,N_13790,N_12788);
and U15524 (N_15524,N_13797,N_12649);
nand U15525 (N_15525,N_14916,N_13970);
xnor U15526 (N_15526,N_12663,N_14912);
nand U15527 (N_15527,N_14208,N_14831);
and U15528 (N_15528,N_13089,N_13177);
nor U15529 (N_15529,N_14692,N_14961);
xnor U15530 (N_15530,N_13686,N_12319);
or U15531 (N_15531,N_12515,N_12222);
or U15532 (N_15532,N_14446,N_14393);
nand U15533 (N_15533,N_13675,N_13040);
and U15534 (N_15534,N_12213,N_14746);
nand U15535 (N_15535,N_13058,N_14138);
and U15536 (N_15536,N_12480,N_14161);
nor U15537 (N_15537,N_12667,N_12643);
nor U15538 (N_15538,N_14449,N_14293);
and U15539 (N_15539,N_13890,N_12919);
nor U15540 (N_15540,N_13155,N_13115);
nand U15541 (N_15541,N_12982,N_12977);
nor U15542 (N_15542,N_12775,N_13037);
and U15543 (N_15543,N_14017,N_12271);
or U15544 (N_15544,N_13015,N_12264);
or U15545 (N_15545,N_12289,N_13430);
xor U15546 (N_15546,N_12647,N_14968);
xor U15547 (N_15547,N_12749,N_13088);
xnor U15548 (N_15548,N_12826,N_13916);
and U15549 (N_15549,N_13976,N_12620);
nor U15550 (N_15550,N_14920,N_13544);
nor U15551 (N_15551,N_13404,N_13222);
nor U15552 (N_15552,N_12218,N_14098);
or U15553 (N_15553,N_13661,N_13441);
nand U15554 (N_15554,N_14786,N_13102);
and U15555 (N_15555,N_14590,N_13273);
nor U15556 (N_15556,N_13560,N_14251);
nor U15557 (N_15557,N_13639,N_14794);
and U15558 (N_15558,N_12101,N_12499);
nor U15559 (N_15559,N_12333,N_14127);
or U15560 (N_15560,N_14475,N_14588);
xnor U15561 (N_15561,N_13086,N_12645);
and U15562 (N_15562,N_13224,N_12735);
xnor U15563 (N_15563,N_14865,N_12943);
nor U15564 (N_15564,N_14418,N_12437);
nor U15565 (N_15565,N_12025,N_13493);
and U15566 (N_15566,N_13185,N_13712);
nor U15567 (N_15567,N_13906,N_12888);
xnor U15568 (N_15568,N_13188,N_13979);
nand U15569 (N_15569,N_12744,N_13808);
and U15570 (N_15570,N_13280,N_14299);
nor U15571 (N_15571,N_14335,N_14165);
and U15572 (N_15572,N_14052,N_13480);
and U15573 (N_15573,N_13850,N_13193);
nand U15574 (N_15574,N_12395,N_12358);
nor U15575 (N_15575,N_14522,N_14002);
or U15576 (N_15576,N_14022,N_12114);
nor U15577 (N_15577,N_14805,N_12883);
xnor U15578 (N_15578,N_13414,N_13897);
xor U15579 (N_15579,N_14444,N_12554);
nor U15580 (N_15580,N_14779,N_13204);
nor U15581 (N_15581,N_12835,N_14166);
and U15582 (N_15582,N_13855,N_14113);
nor U15583 (N_15583,N_13995,N_13039);
nand U15584 (N_15584,N_13061,N_13106);
and U15585 (N_15585,N_14743,N_13888);
nor U15586 (N_15586,N_13374,N_12895);
or U15587 (N_15587,N_12033,N_12650);
and U15588 (N_15588,N_12440,N_12286);
nor U15589 (N_15589,N_14001,N_14344);
xnor U15590 (N_15590,N_13597,N_14036);
nand U15591 (N_15591,N_14244,N_13046);
or U15592 (N_15592,N_13225,N_12774);
nor U15593 (N_15593,N_12013,N_14240);
and U15594 (N_15594,N_12503,N_13130);
nand U15595 (N_15595,N_13883,N_13526);
xor U15596 (N_15596,N_12028,N_12889);
and U15597 (N_15597,N_14772,N_14591);
nor U15598 (N_15598,N_12384,N_12605);
nor U15599 (N_15599,N_14489,N_12792);
nor U15600 (N_15600,N_14004,N_14057);
and U15601 (N_15601,N_12514,N_12321);
and U15602 (N_15602,N_14592,N_14093);
nor U15603 (N_15603,N_12761,N_12405);
and U15604 (N_15604,N_12026,N_14186);
nand U15605 (N_15605,N_14260,N_12404);
and U15606 (N_15606,N_14965,N_14175);
nand U15607 (N_15607,N_14609,N_14271);
and U15608 (N_15608,N_12419,N_12862);
and U15609 (N_15609,N_14349,N_14749);
nor U15610 (N_15610,N_14081,N_14909);
or U15611 (N_15611,N_12166,N_14198);
nor U15612 (N_15612,N_14255,N_12849);
xor U15613 (N_15613,N_14839,N_12701);
nor U15614 (N_15614,N_13555,N_14921);
nand U15615 (N_15615,N_13295,N_13354);
or U15616 (N_15616,N_14952,N_12434);
and U15617 (N_15617,N_14654,N_14582);
xnor U15618 (N_15618,N_13136,N_14636);
and U15619 (N_15619,N_14789,N_14060);
and U15620 (N_15620,N_13165,N_14163);
or U15621 (N_15621,N_12428,N_12698);
nand U15622 (N_15622,N_13450,N_14579);
nor U15623 (N_15623,N_12678,N_12934);
and U15624 (N_15624,N_13378,N_14042);
nor U15625 (N_15625,N_13462,N_12448);
or U15626 (N_15626,N_13876,N_14428);
or U15627 (N_15627,N_14432,N_12441);
xnor U15628 (N_15628,N_12424,N_14719);
nand U15629 (N_15629,N_12348,N_14675);
nand U15630 (N_15630,N_13882,N_12387);
nor U15631 (N_15631,N_12558,N_14917);
and U15632 (N_15632,N_13540,N_14203);
xnor U15633 (N_15633,N_12689,N_13809);
and U15634 (N_15634,N_12738,N_14124);
nand U15635 (N_15635,N_12447,N_14051);
xor U15636 (N_15636,N_13011,N_12827);
or U15637 (N_15637,N_12842,N_14107);
nor U15638 (N_15638,N_12594,N_14954);
xor U15639 (N_15639,N_12817,N_14497);
nor U15640 (N_15640,N_13448,N_14744);
or U15641 (N_15641,N_13619,N_14899);
or U15642 (N_15642,N_14443,N_13963);
or U15643 (N_15643,N_13290,N_13664);
xnor U15644 (N_15644,N_13648,N_12151);
nor U15645 (N_15645,N_12278,N_13117);
nor U15646 (N_15646,N_12268,N_14955);
nor U15647 (N_15647,N_12064,N_14673);
and U15648 (N_15648,N_13693,N_13400);
or U15649 (N_15649,N_14420,N_12655);
nor U15650 (N_15650,N_12296,N_14261);
nor U15651 (N_15651,N_13343,N_12959);
xnor U15652 (N_15652,N_14726,N_13528);
and U15653 (N_15653,N_13507,N_12652);
or U15654 (N_15654,N_12589,N_12386);
xor U15655 (N_15655,N_14471,N_12833);
and U15656 (N_15656,N_13377,N_13913);
nand U15657 (N_15657,N_14742,N_12310);
nand U15658 (N_15658,N_13732,N_14950);
xor U15659 (N_15659,N_14766,N_13364);
nor U15660 (N_15660,N_14206,N_13595);
nand U15661 (N_15661,N_12435,N_13350);
and U15662 (N_15662,N_14134,N_13571);
xor U15663 (N_15663,N_13335,N_12828);
nand U15664 (N_15664,N_14745,N_12956);
xnor U15665 (N_15665,N_14120,N_12803);
nand U15666 (N_15666,N_14799,N_13426);
xor U15667 (N_15667,N_12746,N_13472);
and U15668 (N_15668,N_12080,N_12981);
xor U15669 (N_15669,N_14253,N_12214);
nand U15670 (N_15670,N_12714,N_13253);
nand U15671 (N_15671,N_13748,N_13918);
xnor U15672 (N_15672,N_14641,N_14701);
nor U15673 (N_15673,N_13993,N_14190);
nor U15674 (N_15674,N_14880,N_14737);
nor U15675 (N_15675,N_14333,N_14463);
nand U15676 (N_15676,N_14637,N_13866);
xor U15677 (N_15677,N_14914,N_14978);
or U15678 (N_15678,N_12535,N_12676);
nor U15679 (N_15679,N_14802,N_13180);
xnor U15680 (N_15680,N_12231,N_13923);
nor U15681 (N_15681,N_14844,N_14907);
nand U15682 (N_15682,N_14247,N_12230);
or U15683 (N_15683,N_14537,N_12461);
nand U15684 (N_15684,N_12806,N_12075);
nor U15685 (N_15685,N_12665,N_13900);
nand U15686 (N_15686,N_12201,N_13213);
nand U15687 (N_15687,N_13509,N_13854);
and U15688 (N_15688,N_13791,N_13523);
nor U15689 (N_15689,N_14110,N_14355);
or U15690 (N_15690,N_14982,N_13403);
or U15691 (N_15691,N_14374,N_14594);
nor U15692 (N_15692,N_13513,N_14936);
xor U15693 (N_15693,N_13144,N_13202);
and U15694 (N_15694,N_12901,N_13947);
or U15695 (N_15695,N_12131,N_13942);
xnor U15696 (N_15696,N_12742,N_14642);
xor U15697 (N_15697,N_13574,N_12469);
or U15698 (N_15698,N_13864,N_13607);
nor U15699 (N_15699,N_12983,N_12072);
xor U15700 (N_15700,N_14687,N_14715);
nor U15701 (N_15701,N_13998,N_13500);
or U15702 (N_15702,N_13495,N_13515);
xnor U15703 (N_15703,N_12696,N_13719);
nand U15704 (N_15704,N_14235,N_12859);
nor U15705 (N_15705,N_13948,N_14248);
nor U15706 (N_15706,N_13934,N_13831);
xnor U15707 (N_15707,N_13563,N_13314);
nor U15708 (N_15708,N_12176,N_14523);
xor U15709 (N_15709,N_12917,N_12078);
nand U15710 (N_15710,N_13687,N_12713);
nand U15711 (N_15711,N_14913,N_14868);
xor U15712 (N_15712,N_14045,N_12740);
xor U15713 (N_15713,N_12122,N_13274);
or U15714 (N_15714,N_12630,N_13931);
nand U15715 (N_15715,N_13895,N_13743);
xor U15716 (N_15716,N_12913,N_14953);
nand U15717 (N_15717,N_13787,N_12097);
and U15718 (N_15718,N_14847,N_12477);
or U15719 (N_15719,N_13557,N_12245);
or U15720 (N_15720,N_13497,N_13533);
or U15721 (N_15721,N_12672,N_12069);
or U15722 (N_15722,N_13189,N_14966);
xnor U15723 (N_15723,N_14895,N_14515);
xor U15724 (N_15724,N_12954,N_14290);
and U15725 (N_15725,N_13937,N_12747);
nand U15726 (N_15726,N_14283,N_13892);
and U15727 (N_15727,N_12731,N_12693);
and U15728 (N_15728,N_12636,N_14225);
nand U15729 (N_15729,N_13035,N_12890);
or U15730 (N_15730,N_14461,N_14116);
and U15731 (N_15731,N_14586,N_14940);
nand U15732 (N_15732,N_12190,N_14989);
xnor U15733 (N_15733,N_12617,N_14504);
xnor U15734 (N_15734,N_14800,N_13346);
and U15735 (N_15735,N_13125,N_14153);
and U15736 (N_15736,N_12377,N_13381);
nand U15737 (N_15737,N_12292,N_12352);
nor U15738 (N_15738,N_14302,N_14218);
nand U15739 (N_15739,N_12453,N_13214);
xor U15740 (N_15740,N_12964,N_13858);
nand U15741 (N_15741,N_13677,N_14356);
nor U15742 (N_15742,N_13917,N_14174);
nor U15743 (N_15743,N_12925,N_13437);
or U15744 (N_15744,N_12759,N_12343);
or U15745 (N_15745,N_12211,N_14630);
or U15746 (N_15746,N_12524,N_14720);
xnor U15747 (N_15747,N_14429,N_13008);
xnor U15748 (N_15748,N_13752,N_14245);
or U15749 (N_15749,N_13833,N_14557);
nor U15750 (N_15750,N_12946,N_14699);
and U15751 (N_15751,N_12839,N_12228);
xnor U15752 (N_15752,N_13771,N_13798);
nor U15753 (N_15753,N_14534,N_12162);
xor U15754 (N_15754,N_14105,N_12415);
xor U15755 (N_15755,N_13356,N_14250);
nand U15756 (N_15756,N_14133,N_14266);
nand U15757 (N_15757,N_14327,N_14209);
nor U15758 (N_15758,N_12279,N_14996);
or U15759 (N_15759,N_13149,N_12882);
and U15760 (N_15760,N_13107,N_14611);
nor U15761 (N_15761,N_13499,N_13473);
or U15762 (N_15762,N_13636,N_13530);
and U15763 (N_15763,N_13464,N_13263);
nor U15764 (N_15764,N_14435,N_13048);
nor U15765 (N_15765,N_12845,N_12879);
xor U15766 (N_15766,N_14829,N_13823);
xnor U15767 (N_15767,N_12341,N_13630);
nand U15768 (N_15768,N_14059,N_14168);
nor U15769 (N_15769,N_12287,N_13405);
nand U15770 (N_15770,N_14083,N_14886);
nor U15771 (N_15771,N_13924,N_14359);
xor U15772 (N_15772,N_12662,N_14589);
nand U15773 (N_15773,N_14454,N_12234);
nor U15774 (N_15774,N_14697,N_13460);
nor U15775 (N_15775,N_12705,N_13731);
nand U15776 (N_15776,N_14102,N_12408);
nand U15777 (N_15777,N_12511,N_13154);
nor U15778 (N_15778,N_13825,N_14041);
nor U15779 (N_15779,N_12586,N_13461);
and U15780 (N_15780,N_14852,N_14183);
or U15781 (N_15781,N_13928,N_12880);
nor U15782 (N_15782,N_13867,N_12364);
nor U15783 (N_15783,N_12335,N_13390);
nor U15784 (N_15784,N_14622,N_14437);
nor U15785 (N_15785,N_14033,N_12411);
and U15786 (N_15786,N_14100,N_14358);
and U15787 (N_15787,N_14279,N_12324);
nor U15788 (N_15788,N_13594,N_13402);
nand U15789 (N_15789,N_13408,N_13233);
nand U15790 (N_15790,N_12994,N_12598);
nand U15791 (N_15791,N_12119,N_12311);
nand U15792 (N_15792,N_13318,N_12562);
nor U15793 (N_15793,N_12062,N_14381);
xor U15794 (N_15794,N_13104,N_14188);
and U15795 (N_15795,N_14987,N_12995);
nand U15796 (N_15796,N_14385,N_13992);
or U15797 (N_15797,N_13395,N_14520);
and U15798 (N_15798,N_13583,N_14439);
nand U15799 (N_15799,N_12516,N_14453);
xnor U15800 (N_15800,N_14770,N_13549);
or U15801 (N_15801,N_13051,N_14214);
and U15802 (N_15802,N_13812,N_14197);
and U15803 (N_15803,N_12259,N_12312);
nand U15804 (N_15804,N_12764,N_13491);
and U15805 (N_15805,N_13575,N_12204);
or U15806 (N_15806,N_12070,N_12006);
or U15807 (N_15807,N_13683,N_13512);
nand U15808 (N_15808,N_13766,N_14106);
or U15809 (N_15809,N_14066,N_14199);
nand U15810 (N_15810,N_13313,N_13653);
or U15811 (N_15811,N_14821,N_14242);
xor U15812 (N_15812,N_12702,N_13502);
nor U15813 (N_15813,N_13843,N_13090);
and U15814 (N_15814,N_12719,N_13803);
or U15815 (N_15815,N_13019,N_12675);
xnor U15816 (N_15816,N_14910,N_13845);
or U15817 (N_15817,N_14205,N_13392);
nand U15818 (N_15818,N_12373,N_14585);
nor U15819 (N_15819,N_14512,N_13168);
xnor U15820 (N_15820,N_14367,N_12657);
nor U15821 (N_15821,N_13248,N_12838);
xnor U15822 (N_15822,N_12542,N_14296);
xor U15823 (N_15823,N_14949,N_12397);
or U15824 (N_15824,N_14896,N_12991);
nor U15825 (N_15825,N_14619,N_12241);
or U15826 (N_15826,N_12017,N_12155);
or U15827 (N_15827,N_14689,N_13977);
xnor U15828 (N_15828,N_14572,N_12530);
nand U15829 (N_15829,N_12687,N_12704);
or U15830 (N_15830,N_12233,N_14050);
nand U15831 (N_15831,N_12353,N_13909);
xnor U15832 (N_15832,N_14417,N_14158);
xor U15833 (N_15833,N_13517,N_14991);
nor U15834 (N_15834,N_13094,N_13393);
xnor U15835 (N_15835,N_14088,N_13443);
nor U15836 (N_15836,N_14930,N_12539);
xnor U15837 (N_15837,N_12771,N_14828);
nor U15838 (N_15838,N_12054,N_13981);
nor U15839 (N_15839,N_12618,N_13620);
nand U15840 (N_15840,N_12502,N_12906);
xor U15841 (N_15841,N_12616,N_12432);
xnor U15842 (N_15842,N_12458,N_14070);
or U15843 (N_15843,N_12822,N_13730);
xor U15844 (N_15844,N_13537,N_14387);
and U15845 (N_15845,N_13453,N_14855);
nand U15846 (N_15846,N_12699,N_13945);
or U15847 (N_15847,N_12957,N_13208);
nor U15848 (N_15848,N_14483,N_14189);
and U15849 (N_15849,N_13365,N_14043);
nor U15850 (N_15850,N_13470,N_14533);
xnor U15851 (N_15851,N_13721,N_14013);
nand U15852 (N_15852,N_12173,N_13920);
and U15853 (N_15853,N_14662,N_12948);
xnor U15854 (N_15854,N_12607,N_13479);
nor U15855 (N_15855,N_13423,N_13826);
and U15856 (N_15856,N_13417,N_13439);
nand U15857 (N_15857,N_14287,N_13852);
and U15858 (N_15858,N_13362,N_12253);
or U15859 (N_15859,N_12250,N_12420);
xor U15860 (N_15860,N_13038,N_13103);
xor U15861 (N_15861,N_12534,N_13737);
xor U15862 (N_15862,N_14396,N_13284);
nor U15863 (N_15863,N_13535,N_14710);
nor U15864 (N_15864,N_13832,N_12965);
and U15865 (N_15865,N_12559,N_14227);
nor U15866 (N_15866,N_12585,N_12212);
nand U15867 (N_15867,N_14401,N_13032);
and U15868 (N_15868,N_14648,N_14460);
and U15869 (N_15869,N_14546,N_14304);
or U15870 (N_15870,N_13201,N_12059);
xor U15871 (N_15871,N_13465,N_14825);
and U15872 (N_15872,N_13065,N_12576);
xnor U15873 (N_15873,N_14532,N_14409);
or U15874 (N_15874,N_12087,N_13325);
nand U15875 (N_15875,N_13935,N_12571);
or U15876 (N_15876,N_12582,N_14094);
nand U15877 (N_15877,N_14259,N_14652);
xnor U15878 (N_15878,N_13626,N_12096);
and U15879 (N_15879,N_13708,N_14796);
nand U15880 (N_15880,N_14212,N_12041);
nor U15881 (N_15881,N_13644,N_13322);
and U15882 (N_15882,N_12350,N_12153);
nor U15883 (N_15883,N_13446,N_14459);
nand U15884 (N_15884,N_13182,N_14411);
and U15885 (N_15885,N_13041,N_12979);
and U15886 (N_15886,N_13986,N_13701);
nand U15887 (N_15887,N_12111,N_12095);
xor U15888 (N_15888,N_13425,N_13749);
xnor U15889 (N_15889,N_14681,N_14739);
xnor U15890 (N_15890,N_12791,N_14973);
nor U15891 (N_15891,N_13759,N_14029);
nand U15892 (N_15892,N_14879,N_13455);
xnor U15893 (N_15893,N_13822,N_12581);
xor U15894 (N_15894,N_12819,N_13818);
or U15895 (N_15895,N_13656,N_14455);
or U15896 (N_15896,N_13800,N_13283);
xnor U15897 (N_15897,N_14252,N_14565);
xor U15898 (N_15898,N_12216,N_14119);
nand U15899 (N_15899,N_12463,N_14501);
and U15900 (N_15900,N_14918,N_14684);
nand U15901 (N_15901,N_14500,N_13330);
and U15902 (N_15902,N_14313,N_13873);
nor U15903 (N_15903,N_13475,N_13053);
or U15904 (N_15904,N_13358,N_14213);
and U15905 (N_15905,N_14905,N_13796);
and U15906 (N_15906,N_14020,N_14792);
xor U15907 (N_15907,N_13707,N_13680);
and U15908 (N_15908,N_13050,N_13572);
and U15909 (N_15909,N_12032,N_13598);
xor U15910 (N_15910,N_14650,N_14893);
xor U15911 (N_15911,N_12658,N_12825);
xnor U15912 (N_15912,N_13848,N_12263);
or U15913 (N_15913,N_13127,N_12810);
or U15914 (N_15914,N_13288,N_13521);
or U15915 (N_15915,N_12611,N_14760);
nand U15916 (N_15916,N_14191,N_12600);
nor U15917 (N_15917,N_14498,N_12725);
nor U15918 (N_15918,N_12018,N_14777);
or U15919 (N_15919,N_12886,N_12464);
nor U15920 (N_15920,N_13804,N_14231);
nand U15921 (N_15921,N_14039,N_14063);
and U15922 (N_15922,N_12506,N_14424);
nand U15923 (N_15923,N_13442,N_12677);
or U15924 (N_15924,N_12720,N_14728);
and U15925 (N_15925,N_14933,N_12483);
nand U15926 (N_15926,N_13277,N_14948);
nand U15927 (N_15927,N_12996,N_14164);
and U15928 (N_15928,N_14962,N_12969);
nand U15929 (N_15929,N_12574,N_14567);
nor U15930 (N_15930,N_13059,N_12247);
xnor U15931 (N_15931,N_14754,N_14884);
nand U15932 (N_15932,N_14499,N_14776);
xnor U15933 (N_15933,N_12997,N_13108);
xor U15934 (N_15934,N_12267,N_12438);
and U15935 (N_15935,N_14564,N_12966);
or U15936 (N_15936,N_12800,N_13614);
or U15937 (N_15937,N_12769,N_13565);
or U15938 (N_15938,N_13668,N_12011);
nor U15939 (N_15939,N_13870,N_13608);
nor U15940 (N_15940,N_13341,N_12724);
or U15941 (N_15941,N_13503,N_13079);
and U15942 (N_15942,N_14132,N_14854);
or U15943 (N_15943,N_14027,N_12049);
nor U15944 (N_15944,N_14730,N_12246);
or U15945 (N_15945,N_13004,N_12624);
and U15946 (N_15946,N_13367,N_13838);
nand U15947 (N_15947,N_13907,N_12112);
and U15948 (N_15948,N_12001,N_13388);
xnor U15949 (N_15949,N_13697,N_14552);
or U15950 (N_15950,N_14635,N_12661);
or U15951 (N_15951,N_14677,N_13175);
xnor U15952 (N_15952,N_12005,N_12465);
nor U15953 (N_15953,N_12757,N_14348);
nand U15954 (N_15954,N_12454,N_12185);
xnor U15955 (N_15955,N_12866,N_14859);
nor U15956 (N_15956,N_14130,N_12527);
and U15957 (N_15957,N_14649,N_13634);
xor U15958 (N_15958,N_13713,N_14403);
xor U15959 (N_15959,N_14040,N_14711);
nand U15960 (N_15960,N_14944,N_12159);
and U15961 (N_15961,N_12544,N_13025);
and U15962 (N_15962,N_13846,N_13085);
xnor U15963 (N_15963,N_12710,N_13278);
xnor U15964 (N_15964,N_13943,N_14378);
nand U15965 (N_15965,N_14219,N_12929);
and U15966 (N_15966,N_14604,N_13676);
nor U15967 (N_15967,N_13539,N_13670);
nand U15968 (N_15968,N_13054,N_12938);
xor U15969 (N_15969,N_14607,N_12548);
or U15970 (N_15970,N_12985,N_12608);
and U15971 (N_15971,N_14535,N_13145);
xor U15972 (N_15972,N_13590,N_12110);
or U15973 (N_15973,N_14872,N_14583);
nor U15974 (N_15974,N_12726,N_12203);
nand U15975 (N_15975,N_14136,N_13216);
and U15976 (N_15976,N_12867,N_12443);
or U15977 (N_15977,N_12150,N_13324);
and U15978 (N_15978,N_14759,N_13853);
xor U15979 (N_15979,N_12865,N_12057);
nor U15980 (N_15980,N_12249,N_13782);
and U15981 (N_15981,N_13143,N_14365);
nor U15982 (N_15982,N_12931,N_14665);
nand U15983 (N_15983,N_13219,N_13017);
nor U15984 (N_15984,N_12385,N_12391);
nand U15985 (N_15985,N_12518,N_12354);
and U15986 (N_15986,N_13379,N_13361);
nor U15987 (N_15987,N_14530,N_12181);
xor U15988 (N_15988,N_12733,N_12030);
and U15989 (N_15989,N_13506,N_13047);
or U15990 (N_15990,N_14286,N_12659);
xnor U15991 (N_15991,N_13727,N_13399);
and U15992 (N_15992,N_13660,N_14975);
nand U15993 (N_15993,N_13044,N_14352);
nor U15994 (N_15994,N_12118,N_12466);
nor U15995 (N_15995,N_12445,N_13287);
nor U15996 (N_15996,N_13671,N_14646);
nand U15997 (N_15997,N_13092,N_14233);
or U15998 (N_15998,N_14767,N_12225);
nor U15999 (N_15999,N_13738,N_14551);
or U16000 (N_16000,N_12715,N_12844);
or U16001 (N_16001,N_12910,N_12789);
nand U16002 (N_16002,N_12891,N_12601);
and U16003 (N_16003,N_13893,N_12847);
nand U16004 (N_16004,N_13674,N_14518);
nor U16005 (N_16005,N_12451,N_14058);
nand U16006 (N_16006,N_12134,N_13369);
or U16007 (N_16007,N_12474,N_14992);
and U16008 (N_16008,N_12157,N_14018);
or U16009 (N_16009,N_13781,N_12669);
nand U16010 (N_16010,N_13301,N_12909);
xor U16011 (N_16011,N_13101,N_13160);
or U16012 (N_16012,N_14526,N_13228);
nor U16013 (N_16013,N_13919,N_13162);
nor U16014 (N_16014,N_12613,N_13159);
xor U16015 (N_16015,N_14135,N_12016);
and U16016 (N_16016,N_13879,N_13080);
xnor U16017 (N_16017,N_13312,N_12146);
nand U16018 (N_16018,N_13209,N_13482);
nor U16019 (N_16019,N_12967,N_13247);
nor U16020 (N_16020,N_12147,N_13375);
nor U16021 (N_16021,N_14734,N_12712);
xor U16022 (N_16022,N_13725,N_12174);
and U16023 (N_16023,N_13672,N_14694);
or U16024 (N_16024,N_13982,N_13953);
or U16025 (N_16025,N_12307,N_14314);
and U16026 (N_16026,N_13321,N_14732);
nor U16027 (N_16027,N_13444,N_13880);
and U16028 (N_16028,N_12473,N_13566);
nor U16029 (N_16029,N_13711,N_14139);
nor U16030 (N_16030,N_13030,N_12907);
xor U16031 (N_16031,N_12088,N_14178);
nor U16032 (N_16032,N_12797,N_12164);
nor U16033 (N_16033,N_13795,N_14140);
or U16034 (N_16034,N_14371,N_13105);
xor U16035 (N_16035,N_14942,N_14392);
or U16036 (N_16036,N_12277,N_12426);
and U16037 (N_16037,N_13538,N_13975);
nand U16038 (N_16038,N_13210,N_13633);
nor U16039 (N_16039,N_12680,N_14971);
or U16040 (N_16040,N_13172,N_13980);
nor U16041 (N_16041,N_13710,N_12132);
or U16042 (N_16042,N_14055,N_14404);
xnor U16043 (N_16043,N_13422,N_13199);
nand U16044 (N_16044,N_14181,N_12313);
xnor U16045 (N_16045,N_12836,N_14090);
nor U16046 (N_16046,N_13238,N_12834);
and U16047 (N_16047,N_14156,N_12987);
or U16048 (N_16048,N_12338,N_14238);
or U16049 (N_16049,N_13581,N_14778);
nand U16050 (N_16050,N_12099,N_12843);
or U16051 (N_16051,N_12040,N_14399);
nor U16052 (N_16052,N_12816,N_14695);
nand U16053 (N_16053,N_12855,N_12210);
and U16054 (N_16054,N_13071,N_12623);
or U16055 (N_16055,N_14414,N_12857);
and U16056 (N_16056,N_13728,N_12497);
nand U16057 (N_16057,N_12418,N_13753);
and U16058 (N_16058,N_13767,N_13632);
nor U16059 (N_16059,N_13972,N_14078);
and U16060 (N_16060,N_12148,N_14149);
xnor U16061 (N_16061,N_14666,N_13508);
xor U16062 (N_16062,N_12531,N_13531);
nor U16063 (N_16063,N_14503,N_14294);
or U16064 (N_16064,N_12796,N_14559);
and U16065 (N_16065,N_13474,N_12422);
and U16066 (N_16066,N_14275,N_12609);
xor U16067 (N_16067,N_14391,N_12565);
nor U16068 (N_16068,N_14957,N_14605);
or U16069 (N_16069,N_12425,N_12063);
and U16070 (N_16070,N_12417,N_12060);
and U16071 (N_16071,N_14945,N_14362);
nor U16072 (N_16072,N_12066,N_12206);
nand U16073 (N_16073,N_14788,N_12772);
xnor U16074 (N_16074,N_14319,N_14544);
and U16075 (N_16075,N_14513,N_12167);
nor U16076 (N_16076,N_13186,N_13655);
xnor U16077 (N_16077,N_12076,N_13119);
or U16078 (N_16078,N_14322,N_14969);
or U16079 (N_16079,N_13391,N_13112);
nor U16080 (N_16080,N_13382,N_13891);
nand U16081 (N_16081,N_13251,N_14263);
nand U16082 (N_16082,N_12989,N_14672);
nor U16083 (N_16083,N_12583,N_12765);
nor U16084 (N_16084,N_13621,N_12360);
and U16085 (N_16085,N_14282,N_13816);
nand U16086 (N_16086,N_14876,N_13967);
nand U16087 (N_16087,N_14603,N_14386);
nor U16088 (N_16088,N_14122,N_13003);
nor U16089 (N_16089,N_12911,N_13006);
nor U16090 (N_16090,N_14947,N_12540);
or U16091 (N_16091,N_13013,N_12456);
nand U16092 (N_16092,N_13029,N_14170);
or U16093 (N_16093,N_13551,N_12528);
or U16094 (N_16094,N_14074,N_13519);
xor U16095 (N_16095,N_12092,N_13616);
nor U16096 (N_16096,N_13554,N_14478);
nor U16097 (N_16097,N_14866,N_12361);
or U16098 (N_16098,N_14315,N_12782);
nor U16099 (N_16099,N_14514,N_14713);
or U16100 (N_16100,N_13559,N_14889);
nor U16101 (N_16101,N_13938,N_13652);
nor U16102 (N_16102,N_14874,N_13220);
and U16103 (N_16103,N_14806,N_13275);
nand U16104 (N_16104,N_13567,N_13682);
or U16105 (N_16105,N_12809,N_12529);
xor U16106 (N_16106,N_12673,N_12180);
xor U16107 (N_16107,N_13368,N_14988);
xnor U16108 (N_16108,N_13345,N_14089);
nand U16109 (N_16109,N_12878,N_12098);
or U16110 (N_16110,N_12240,N_12500);
nor U16111 (N_16111,N_12100,N_13695);
xor U16112 (N_16112,N_13056,N_14724);
nand U16113 (N_16113,N_13902,N_14626);
xnor U16114 (N_16114,N_14176,N_14144);
or U16115 (N_16115,N_14034,N_12375);
or U16116 (N_16116,N_13359,N_12036);
nor U16117 (N_16117,N_14481,N_12170);
or U16118 (N_16118,N_12928,N_12978);
nor U16119 (N_16119,N_14277,N_12711);
nor U16120 (N_16120,N_14621,N_13957);
xnor U16121 (N_16121,N_13469,N_12351);
and U16122 (N_16122,N_14995,N_13704);
nand U16123 (N_16123,N_13376,N_13230);
xor U16124 (N_16124,N_14269,N_12334);
and U16125 (N_16125,N_13578,N_14215);
nor U16126 (N_16126,N_14394,N_13534);
and U16127 (N_16127,N_14256,N_13384);
nor U16128 (N_16128,N_12922,N_13640);
and U16129 (N_16129,N_13785,N_14369);
nand U16130 (N_16130,N_12569,N_14345);
or U16131 (N_16131,N_13300,N_12038);
and U16132 (N_16132,N_14431,N_13700);
xnor U16133 (N_16133,N_13173,N_13985);
or U16134 (N_16134,N_12998,N_14740);
and U16135 (N_16135,N_12670,N_13279);
nor U16136 (N_16136,N_14092,N_12541);
and U16137 (N_16137,N_12512,N_14236);
and U16138 (N_16138,N_12580,N_14669);
nor U16139 (N_16139,N_13966,N_12039);
xor U16140 (N_16140,N_13142,N_13174);
nand U16141 (N_16141,N_13769,N_13097);
or U16142 (N_16142,N_13543,N_12109);
and U16143 (N_16143,N_12932,N_14495);
and U16144 (N_16144,N_14612,N_12523);
xor U16145 (N_16145,N_14064,N_12409);
xnor U16146 (N_16146,N_13638,N_14226);
nor U16147 (N_16147,N_13096,N_13492);
or U16148 (N_16148,N_14633,N_13348);
or U16149 (N_16149,N_14556,N_12829);
xor U16150 (N_16150,N_14152,N_12124);
nand U16151 (N_16151,N_12745,N_13266);
nand U16152 (N_16152,N_12223,N_12048);
xnor U16153 (N_16153,N_12065,N_12854);
xnor U16154 (N_16154,N_12086,N_14044);
xor U16155 (N_16155,N_14679,N_14507);
nor U16156 (N_16156,N_13592,N_13925);
xnor U16157 (N_16157,N_13311,N_13568);
and U16158 (N_16158,N_14035,N_12331);
and U16159 (N_16159,N_14960,N_13260);
or U16160 (N_16160,N_13196,N_14670);
or U16161 (N_16161,N_12270,N_13124);
or U16162 (N_16162,N_14660,N_13072);
and U16163 (N_16163,N_14143,N_13784);
nand U16164 (N_16164,N_12717,N_12492);
nor U16165 (N_16165,N_14311,N_13129);
xnor U16166 (N_16166,N_13729,N_14258);
or U16167 (N_16167,N_13589,N_13758);
or U16168 (N_16168,N_14220,N_13383);
and U16169 (N_16169,N_14787,N_14574);
xor U16170 (N_16170,N_13310,N_12566);
nand U16171 (N_16171,N_13612,N_14395);
nand U16172 (N_16172,N_14597,N_12905);
nor U16173 (N_16173,N_13684,N_13983);
or U16174 (N_16174,N_13466,N_12961);
nor U16175 (N_16175,N_12622,N_13861);
nor U16176 (N_16176,N_13252,N_12021);
nand U16177 (N_16177,N_12300,N_14361);
or U16178 (N_16178,N_13844,N_14201);
and U16179 (N_16179,N_13236,N_13715);
nand U16180 (N_16180,N_13281,N_12732);
or U16181 (N_16181,N_13315,N_13239);
xnor U16182 (N_16182,N_14545,N_13939);
xnor U16183 (N_16183,N_13610,N_13625);
xnor U16184 (N_16184,N_14388,N_14798);
nor U16185 (N_16185,N_14547,N_13585);
nand U16186 (N_16186,N_14791,N_12332);
nor U16187 (N_16187,N_14300,N_12760);
or U16188 (N_16188,N_14402,N_14457);
xor U16189 (N_16189,N_12776,N_14755);
xor U16190 (N_16190,N_13232,N_13954);
or U16191 (N_16191,N_12315,N_14148);
xor U16192 (N_16192,N_13270,N_13690);
xnor U16193 (N_16193,N_14908,N_13564);
and U16194 (N_16194,N_12798,N_13200);
and U16195 (N_16195,N_14104,N_12073);
xnor U16196 (N_16196,N_12785,N_14703);
xnor U16197 (N_16197,N_12853,N_12549);
and U16198 (N_16198,N_12877,N_12163);
xnor U16199 (N_16199,N_12374,N_13269);
xnor U16200 (N_16200,N_13692,N_12815);
and U16201 (N_16201,N_14628,N_14647);
nor U16202 (N_16202,N_13268,N_12094);
nor U16203 (N_16203,N_13490,N_12864);
nand U16204 (N_16204,N_13221,N_13432);
or U16205 (N_16205,N_12402,N_14655);
or U16206 (N_16206,N_13955,N_12754);
nand U16207 (N_16207,N_13944,N_14580);
xnor U16208 (N_16208,N_13190,N_12550);
or U16209 (N_16209,N_13898,N_13286);
nor U16210 (N_16210,N_12762,N_12363);
and U16211 (N_16211,N_12470,N_14867);
xnor U16212 (N_16212,N_12243,N_14465);
nor U16213 (N_16213,N_13841,N_14773);
or U16214 (N_16214,N_13131,N_14053);
nand U16215 (N_16215,N_14185,N_14558);
nor U16216 (N_16216,N_12496,N_14926);
nor U16217 (N_16217,N_12468,N_13122);
xnor U16218 (N_16218,N_13666,N_12407);
nor U16219 (N_16219,N_13394,N_14180);
and U16220 (N_16220,N_12394,N_13170);
or U16221 (N_16221,N_13878,N_12727);
and U16222 (N_16222,N_12567,N_12521);
xnor U16223 (N_16223,N_12123,N_13586);
nand U16224 (N_16224,N_12510,N_13773);
and U16225 (N_16225,N_12383,N_13930);
nor U16226 (N_16226,N_14464,N_13548);
and U16227 (N_16227,N_14645,N_13319);
nand U16228 (N_16228,N_12685,N_12579);
nand U16229 (N_16229,N_13553,N_13308);
xnor U16230 (N_16230,N_12851,N_12187);
nor U16231 (N_16231,N_13205,N_14923);
or U16232 (N_16232,N_13156,N_13658);
or U16233 (N_16233,N_14571,N_14733);
or U16234 (N_16234,N_14243,N_12169);
xor U16235 (N_16235,N_12903,N_14706);
or U16236 (N_16236,N_13250,N_12309);
nor U16237 (N_16237,N_13217,N_12654);
nand U16238 (N_16238,N_14329,N_13463);
and U16239 (N_16239,N_12126,N_12841);
and U16240 (N_16240,N_14903,N_13387);
or U16241 (N_16241,N_14202,N_13884);
nor U16242 (N_16242,N_12158,N_13524);
nand U16243 (N_16243,N_13296,N_13081);
or U16244 (N_16244,N_12592,N_14919);
nor U16245 (N_16245,N_13588,N_13603);
or U16246 (N_16246,N_12846,N_12130);
nor U16247 (N_16247,N_14542,N_14167);
and U16248 (N_16248,N_12141,N_13569);
nor U16249 (N_16249,N_14456,N_14048);
or U16250 (N_16250,N_13868,N_14644);
and U16251 (N_16251,N_13857,N_13255);
xnor U16252 (N_16252,N_12137,N_14200);
or U16253 (N_16253,N_14373,N_14342);
nand U16254 (N_16254,N_12304,N_12430);
or U16255 (N_16255,N_14488,N_12179);
xor U16256 (N_16256,N_13010,N_14097);
or U16257 (N_16257,N_13062,N_14904);
nor U16258 (N_16258,N_12856,N_12193);
or U16259 (N_16259,N_12329,N_14845);
nand U16260 (N_16260,N_12980,N_12787);
and U16261 (N_16261,N_14862,N_14006);
or U16262 (N_16262,N_12457,N_12156);
or U16263 (N_16263,N_13435,N_14819);
and U16264 (N_16264,N_12433,N_12316);
nand U16265 (N_16265,N_14838,N_13814);
nor U16266 (N_16266,N_13082,N_13904);
nor U16267 (N_16267,N_13922,N_12356);
and U16268 (N_16268,N_14756,N_12873);
xor U16269 (N_16269,N_12626,N_12547);
nand U16270 (N_16270,N_14434,N_12288);
and U16271 (N_16271,N_12489,N_13389);
or U16272 (N_16272,N_13307,N_14861);
nand U16273 (N_16273,N_12184,N_14368);
nor U16274 (N_16274,N_14765,N_14521);
and U16275 (N_16275,N_14780,N_13045);
and U16276 (N_16276,N_12874,N_12736);
and U16277 (N_16277,N_14131,N_13447);
xor U16278 (N_16278,N_12968,N_12952);
nor U16279 (N_16279,N_14977,N_13940);
xor U16280 (N_16280,N_13881,N_12556);
or U16281 (N_16281,N_14856,N_13527);
nor U16282 (N_16282,N_14517,N_12513);
xor U16283 (N_16283,N_12537,N_14927);
xnor U16284 (N_16284,N_14068,N_14069);
and U16285 (N_16285,N_14125,N_14416);
and U16286 (N_16286,N_14581,N_13427);
nor U16287 (N_16287,N_14979,N_12584);
nand U16288 (N_16288,N_13339,N_14848);
and U16289 (N_16289,N_12362,N_13665);
or U16290 (N_16290,N_14508,N_13717);
xor U16291 (N_16291,N_14390,N_12988);
nand U16292 (N_16292,N_12804,N_14285);
xnor U16293 (N_16293,N_12602,N_12641);
nor U16294 (N_16294,N_14983,N_12990);
nand U16295 (N_16295,N_13532,N_14817);
nand U16296 (N_16296,N_13587,N_13763);
or U16297 (N_16297,N_13340,N_12690);
nor U16298 (N_16298,N_12399,N_13428);
nor U16299 (N_16299,N_13306,N_12638);
nor U16300 (N_16300,N_14554,N_13792);
nor U16301 (N_16301,N_13735,N_14593);
or U16302 (N_16302,N_14150,N_13333);
xor U16303 (N_16303,N_13293,N_13522);
xor U16304 (N_16304,N_13218,N_14111);
xnor U16305 (N_16305,N_13291,N_13116);
nand U16306 (N_16306,N_13813,N_12224);
xnor U16307 (N_16307,N_12183,N_14306);
xor U16308 (N_16308,N_12472,N_13457);
or U16309 (N_16309,N_12786,N_13241);
nor U16310 (N_16310,N_12683,N_12721);
xnor U16311 (N_16311,N_13036,N_13118);
and U16312 (N_16312,N_13413,N_14651);
xor U16313 (N_16313,N_13514,N_13811);
or U16314 (N_16314,N_13901,N_12490);
nor U16315 (N_16315,N_12207,N_13810);
xnor U16316 (N_16316,N_13961,N_13401);
and U16317 (N_16317,N_14450,N_12082);
nand U16318 (N_16318,N_14281,N_13747);
or U16319 (N_16319,N_12921,N_12695);
nand U16320 (N_16320,N_13851,N_14723);
xor U16321 (N_16321,N_14195,N_13021);
nand U16322 (N_16322,N_13328,N_12648);
xnor U16323 (N_16323,N_12974,N_14221);
nand U16324 (N_16324,N_13372,N_14155);
and U16325 (N_16325,N_13126,N_12370);
or U16326 (N_16326,N_13783,N_14363);
or U16327 (N_16327,N_14187,N_12323);
nor U16328 (N_16328,N_14643,N_12546);
and U16329 (N_16329,N_12389,N_12823);
and U16330 (N_16330,N_14091,N_12024);
xnor U16331 (N_16331,N_14268,N_14082);
nor U16332 (N_16332,N_14598,N_14974);
xnor U16333 (N_16333,N_12707,N_14784);
and U16334 (N_16334,N_14813,N_12708);
nand U16335 (N_16335,N_14067,N_13244);
nand U16336 (N_16336,N_13191,N_12014);
xor U16337 (N_16337,N_12773,N_13412);
and U16338 (N_16338,N_13877,N_13485);
nor U16339 (N_16339,N_13138,N_13113);
xor U16340 (N_16340,N_14931,N_14380);
nand U16341 (N_16341,N_14320,N_14080);
nor U16342 (N_16342,N_13723,N_13750);
nor U16343 (N_16343,N_12501,N_12625);
nor U16344 (N_16344,N_12884,N_12029);
nand U16345 (N_16345,N_13786,N_14249);
xor U16346 (N_16346,N_12380,N_12299);
or U16347 (N_16347,N_12614,N_14676);
nor U16348 (N_16348,N_13298,N_13806);
nand U16349 (N_16349,N_12498,N_13905);
and U16350 (N_16350,N_13874,N_14851);
nand U16351 (N_16351,N_13756,N_13859);
xnor U16352 (N_16352,N_12168,N_13628);
and U16353 (N_16353,N_14108,N_14911);
or U16354 (N_16354,N_13467,N_14771);
and U16355 (N_16355,N_13429,N_13087);
nand U16356 (N_16356,N_14986,N_13694);
and U16357 (N_16357,N_14171,N_14000);
nor U16358 (N_16358,N_14629,N_14229);
xnor U16359 (N_16359,N_14768,N_14157);
nand U16360 (N_16360,N_14577,N_12830);
nand U16361 (N_16361,N_13299,N_13452);
or U16362 (N_16362,N_12269,N_14610);
and U16363 (N_16363,N_14147,N_12944);
and U16364 (N_16364,N_13933,N_14639);
xor U16365 (N_16365,N_13083,N_12295);
nor U16366 (N_16366,N_12142,N_14680);
nand U16367 (N_16367,N_13069,N_14781);
xor U16368 (N_16368,N_14599,N_12728);
xor U16369 (N_16369,N_13558,N_13623);
or U16370 (N_16370,N_14970,N_14177);
and U16371 (N_16371,N_12349,N_13956);
xor U16372 (N_16372,N_13075,N_13624);
xnor U16373 (N_16373,N_14849,N_14878);
and U16374 (N_16374,N_14541,N_14021);
nand U16375 (N_16375,N_12282,N_13556);
xor U16376 (N_16376,N_12487,N_14234);
nand U16377 (N_16377,N_14123,N_12709);
nor U16378 (N_16378,N_14430,N_12090);
or U16379 (N_16379,N_14324,N_13366);
and U16380 (N_16380,N_13941,N_14377);
xor U16381 (N_16381,N_13994,N_13910);
nand U16382 (N_16382,N_14353,N_12258);
nand U16383 (N_16383,N_13579,N_12793);
and U16384 (N_16384,N_12342,N_12778);
or U16385 (N_16385,N_12273,N_13740);
xnor U16386 (N_16386,N_14882,N_14408);
xor U16387 (N_16387,N_12900,N_14262);
or U16388 (N_16388,N_14634,N_14527);
nor U16389 (N_16389,N_14179,N_14763);
or U16390 (N_16390,N_14502,N_13576);
or U16391 (N_16391,N_14623,N_13282);
nor U16392 (N_16392,N_14690,N_13582);
and U16393 (N_16393,N_12870,N_14422);
nor U16394 (N_16394,N_12679,N_12455);
xnor U16395 (N_16395,N_14462,N_12603);
nand U16396 (N_16396,N_14476,N_13169);
xor U16397 (N_16397,N_13133,N_12813);
and U16398 (N_16398,N_14967,N_14343);
and U16399 (N_16399,N_12197,N_12716);
nand U16400 (N_16400,N_12691,N_13327);
and U16401 (N_16401,N_12509,N_14795);
nor U16402 (N_16402,N_14758,N_14658);
and U16403 (N_16403,N_12266,N_13445);
nand U16404 (N_16404,N_12217,N_13765);
xnor U16405 (N_16405,N_12751,N_12808);
nand U16406 (N_16406,N_14741,N_12671);
or U16407 (N_16407,N_13415,N_12303);
nand U16408 (N_16408,N_13351,N_14747);
and U16409 (N_16409,N_13772,N_12089);
and U16410 (N_16410,N_12790,N_13629);
xnor U16411 (N_16411,N_14736,N_12337);
nand U16412 (N_16412,N_14782,N_12756);
and U16413 (N_16413,N_12651,N_12923);
and U16414 (N_16414,N_13257,N_12814);
nand U16415 (N_16415,N_14688,N_14667);
xor U16416 (N_16416,N_12285,N_14506);
and U16417 (N_16417,N_12899,N_13997);
nor U16418 (N_16418,N_13459,N_13347);
nand U16419 (N_16419,N_12686,N_14421);
xnor U16420 (N_16420,N_14702,N_14079);
or U16421 (N_16421,N_13885,N_14162);
nand U16422 (N_16422,N_14906,N_13227);
nor U16423 (N_16423,N_14023,N_12198);
nand U16424 (N_16424,N_13024,N_13229);
nor U16425 (N_16425,N_13856,N_12355);
nor U16426 (N_16426,N_14705,N_12718);
xnor U16427 (N_16427,N_14030,N_14172);
or U16428 (N_16428,N_12610,N_12290);
nand U16429 (N_16429,N_14869,N_12656);
or U16430 (N_16430,N_14054,N_14339);
and U16431 (N_16431,N_14671,N_14334);
or U16432 (N_16432,N_14379,N_13342);
and U16433 (N_16433,N_14194,N_12330);
xor U16434 (N_16434,N_14704,N_13309);
nand U16435 (N_16435,N_14210,N_12136);
and U16436 (N_16436,N_12427,N_13702);
nor U16437 (N_16437,N_13863,N_12949);
or U16438 (N_16438,N_12145,N_14273);
xor U16439 (N_16439,N_12275,N_13736);
or U16440 (N_16440,N_14398,N_12274);
nand U16441 (N_16441,N_14415,N_14616);
nor U16442 (N_16442,N_12984,N_12085);
xnor U16443 (N_16443,N_12491,N_14328);
or U16444 (N_16444,N_13194,N_14466);
and U16445 (N_16445,N_12568,N_14548);
nor U16446 (N_16446,N_12107,N_14440);
nand U16447 (N_16447,N_12084,N_13915);
nor U16448 (N_16448,N_13385,N_12272);
xor U16449 (N_16449,N_13242,N_13304);
and U16450 (N_16450,N_14614,N_12302);
xnor U16451 (N_16451,N_12192,N_13498);
nor U16452 (N_16452,N_14956,N_12235);
nand U16453 (N_16453,N_14941,N_12748);
nand U16454 (N_16454,N_13434,N_12572);
and U16455 (N_16455,N_14563,N_12476);
xor U16456 (N_16456,N_14095,N_12520);
nand U16457 (N_16457,N_12144,N_12937);
nor U16458 (N_16458,N_14990,N_12436);
or U16459 (N_16459,N_14241,N_13034);
and U16460 (N_16460,N_13593,N_14480);
xor U16461 (N_16461,N_12722,N_13744);
nor U16462 (N_16462,N_13139,N_13243);
xnor U16463 (N_16463,N_12750,N_12992);
nor U16464 (N_16464,N_14010,N_12660);
or U16465 (N_16465,N_14312,N_14808);
nor U16466 (N_16466,N_14016,N_13724);
nor U16467 (N_16467,N_14487,N_14338);
nor U16468 (N_16468,N_12942,N_12261);
nand U16469 (N_16469,N_12219,N_13449);
and U16470 (N_16470,N_12627,N_13249);
xnor U16471 (N_16471,N_13419,N_13370);
xor U16472 (N_16472,N_14708,N_12027);
or U16473 (N_16473,N_13433,N_13468);
or U16474 (N_16474,N_13889,N_14891);
or U16475 (N_16475,N_14204,N_13911);
and U16476 (N_16476,N_12975,N_14077);
nand U16477 (N_16477,N_13067,N_14816);
nor U16478 (N_16478,N_14491,N_14774);
and U16479 (N_16479,N_14469,N_12575);
xor U16480 (N_16480,N_14071,N_13320);
and U16481 (N_16481,N_13068,N_13336);
nand U16482 (N_16482,N_13344,N_14980);
or U16483 (N_16483,N_12646,N_14145);
and U16484 (N_16484,N_14288,N_14999);
nor U16485 (N_16485,N_14129,N_14887);
nor U16486 (N_16486,N_14735,N_14159);
xnor U16487 (N_16487,N_13042,N_14117);
nor U16488 (N_16488,N_14790,N_13095);
and U16489 (N_16489,N_14553,N_13542);
and U16490 (N_16490,N_12116,N_13669);
xor U16491 (N_16491,N_14606,N_13171);
nand U16492 (N_16492,N_14046,N_14902);
nand U16493 (N_16493,N_13984,N_14901);
nor U16494 (N_16494,N_12257,N_13276);
nand U16495 (N_16495,N_12781,N_13303);
or U16496 (N_16496,N_13023,N_12368);
xor U16497 (N_16497,N_14573,N_12308);
and U16498 (N_16498,N_14026,N_14543);
xor U16499 (N_16499,N_13609,N_13996);
nand U16500 (N_16500,N_12281,N_14631);
and U16501 (N_16501,N_14228,N_14554);
nand U16502 (N_16502,N_12492,N_12977);
or U16503 (N_16503,N_14191,N_12388);
and U16504 (N_16504,N_12363,N_12904);
xor U16505 (N_16505,N_13644,N_14087);
and U16506 (N_16506,N_13007,N_14467);
xor U16507 (N_16507,N_13241,N_14842);
or U16508 (N_16508,N_12579,N_12573);
nand U16509 (N_16509,N_12418,N_14198);
xor U16510 (N_16510,N_12619,N_13977);
nand U16511 (N_16511,N_14564,N_14589);
xnor U16512 (N_16512,N_14810,N_14580);
nand U16513 (N_16513,N_12909,N_12592);
or U16514 (N_16514,N_12102,N_14677);
or U16515 (N_16515,N_12919,N_14007);
nand U16516 (N_16516,N_12751,N_14128);
nand U16517 (N_16517,N_14621,N_13578);
or U16518 (N_16518,N_13141,N_14944);
xnor U16519 (N_16519,N_13798,N_13581);
xor U16520 (N_16520,N_12595,N_14451);
or U16521 (N_16521,N_14979,N_13782);
nor U16522 (N_16522,N_12259,N_14469);
and U16523 (N_16523,N_14538,N_12559);
nor U16524 (N_16524,N_13789,N_13929);
or U16525 (N_16525,N_14081,N_14174);
nor U16526 (N_16526,N_12516,N_14734);
xnor U16527 (N_16527,N_13594,N_14277);
or U16528 (N_16528,N_13159,N_14786);
and U16529 (N_16529,N_14437,N_13935);
nand U16530 (N_16530,N_14583,N_14256);
or U16531 (N_16531,N_12762,N_12613);
nor U16532 (N_16532,N_14397,N_14971);
or U16533 (N_16533,N_14913,N_13244);
or U16534 (N_16534,N_14706,N_12676);
and U16535 (N_16535,N_14296,N_12312);
nand U16536 (N_16536,N_13975,N_13049);
and U16537 (N_16537,N_13398,N_14705);
or U16538 (N_16538,N_13167,N_12043);
xor U16539 (N_16539,N_13024,N_12072);
and U16540 (N_16540,N_14320,N_13105);
nor U16541 (N_16541,N_12645,N_14206);
xnor U16542 (N_16542,N_14708,N_13151);
or U16543 (N_16543,N_13343,N_14504);
nand U16544 (N_16544,N_13812,N_12622);
or U16545 (N_16545,N_13036,N_14203);
nand U16546 (N_16546,N_12740,N_14644);
or U16547 (N_16547,N_12274,N_13286);
or U16548 (N_16548,N_13211,N_12875);
nor U16549 (N_16549,N_14386,N_14200);
nor U16550 (N_16550,N_13634,N_12875);
nor U16551 (N_16551,N_12037,N_12714);
nand U16552 (N_16552,N_14910,N_13130);
xor U16553 (N_16553,N_12104,N_13505);
xnor U16554 (N_16554,N_12436,N_14475);
nand U16555 (N_16555,N_12421,N_12000);
and U16556 (N_16556,N_12001,N_12548);
or U16557 (N_16557,N_13185,N_14932);
or U16558 (N_16558,N_14264,N_13301);
and U16559 (N_16559,N_13374,N_14822);
nand U16560 (N_16560,N_12831,N_12532);
xnor U16561 (N_16561,N_12419,N_13697);
nand U16562 (N_16562,N_14919,N_14050);
or U16563 (N_16563,N_14432,N_14235);
nand U16564 (N_16564,N_14556,N_12906);
nor U16565 (N_16565,N_12714,N_13460);
nor U16566 (N_16566,N_12226,N_14612);
or U16567 (N_16567,N_14718,N_14167);
xor U16568 (N_16568,N_14851,N_12631);
or U16569 (N_16569,N_13764,N_14897);
nor U16570 (N_16570,N_14679,N_12334);
xnor U16571 (N_16571,N_13577,N_12368);
xor U16572 (N_16572,N_12861,N_13245);
nand U16573 (N_16573,N_14726,N_13854);
nand U16574 (N_16574,N_14572,N_13996);
or U16575 (N_16575,N_13181,N_13297);
nor U16576 (N_16576,N_12991,N_14077);
nor U16577 (N_16577,N_13868,N_12841);
nor U16578 (N_16578,N_12021,N_13026);
nor U16579 (N_16579,N_14535,N_12441);
nor U16580 (N_16580,N_13004,N_12342);
nand U16581 (N_16581,N_13963,N_12610);
or U16582 (N_16582,N_14122,N_12035);
nand U16583 (N_16583,N_13086,N_14873);
nor U16584 (N_16584,N_12597,N_14312);
or U16585 (N_16585,N_13093,N_13662);
nand U16586 (N_16586,N_12669,N_12336);
nand U16587 (N_16587,N_13086,N_14699);
or U16588 (N_16588,N_13364,N_13499);
and U16589 (N_16589,N_14749,N_12735);
xor U16590 (N_16590,N_13473,N_14283);
or U16591 (N_16591,N_12500,N_12218);
and U16592 (N_16592,N_13405,N_12215);
or U16593 (N_16593,N_13569,N_12761);
and U16594 (N_16594,N_12538,N_12104);
and U16595 (N_16595,N_13067,N_12169);
nor U16596 (N_16596,N_13726,N_14441);
nand U16597 (N_16597,N_12519,N_13536);
and U16598 (N_16598,N_12290,N_13260);
nand U16599 (N_16599,N_12033,N_13183);
xor U16600 (N_16600,N_13188,N_12658);
and U16601 (N_16601,N_14912,N_14165);
and U16602 (N_16602,N_12383,N_13957);
xnor U16603 (N_16603,N_13683,N_12064);
nor U16604 (N_16604,N_14840,N_14678);
nor U16605 (N_16605,N_13158,N_12738);
nor U16606 (N_16606,N_13356,N_13825);
xnor U16607 (N_16607,N_13746,N_13642);
and U16608 (N_16608,N_14777,N_13116);
or U16609 (N_16609,N_14074,N_14202);
xor U16610 (N_16610,N_13370,N_13185);
and U16611 (N_16611,N_13412,N_12633);
or U16612 (N_16612,N_13039,N_13017);
and U16613 (N_16613,N_14910,N_13244);
or U16614 (N_16614,N_13892,N_12544);
or U16615 (N_16615,N_14227,N_13772);
or U16616 (N_16616,N_12421,N_13310);
or U16617 (N_16617,N_14329,N_12989);
xnor U16618 (N_16618,N_14301,N_13589);
and U16619 (N_16619,N_12311,N_14941);
nor U16620 (N_16620,N_14010,N_13397);
xor U16621 (N_16621,N_12079,N_14948);
nand U16622 (N_16622,N_12708,N_12493);
and U16623 (N_16623,N_13398,N_14316);
or U16624 (N_16624,N_13336,N_13779);
nor U16625 (N_16625,N_12751,N_14908);
nor U16626 (N_16626,N_12211,N_12126);
nand U16627 (N_16627,N_13832,N_12522);
nand U16628 (N_16628,N_13404,N_12373);
nand U16629 (N_16629,N_12805,N_14391);
or U16630 (N_16630,N_12374,N_13014);
nor U16631 (N_16631,N_13178,N_12419);
xor U16632 (N_16632,N_14016,N_14739);
xnor U16633 (N_16633,N_12502,N_13457);
xnor U16634 (N_16634,N_14734,N_14604);
or U16635 (N_16635,N_12965,N_12195);
xor U16636 (N_16636,N_12236,N_14432);
and U16637 (N_16637,N_14628,N_12221);
nor U16638 (N_16638,N_13328,N_13612);
xnor U16639 (N_16639,N_12194,N_12445);
or U16640 (N_16640,N_14897,N_12737);
xnor U16641 (N_16641,N_13109,N_14087);
xnor U16642 (N_16642,N_13890,N_14472);
nand U16643 (N_16643,N_14823,N_13430);
nor U16644 (N_16644,N_12397,N_14311);
nor U16645 (N_16645,N_12983,N_13937);
nand U16646 (N_16646,N_14158,N_13162);
and U16647 (N_16647,N_13531,N_14163);
and U16648 (N_16648,N_14763,N_14629);
nand U16649 (N_16649,N_13190,N_12366);
xnor U16650 (N_16650,N_14755,N_13877);
and U16651 (N_16651,N_12418,N_14580);
nor U16652 (N_16652,N_13497,N_12059);
nand U16653 (N_16653,N_12719,N_12263);
nor U16654 (N_16654,N_14404,N_14570);
xnor U16655 (N_16655,N_13881,N_14450);
xnor U16656 (N_16656,N_13713,N_13930);
xnor U16657 (N_16657,N_13532,N_13215);
nor U16658 (N_16658,N_13161,N_12816);
xnor U16659 (N_16659,N_12567,N_12973);
or U16660 (N_16660,N_13096,N_14349);
nor U16661 (N_16661,N_14344,N_13670);
or U16662 (N_16662,N_13821,N_14859);
and U16663 (N_16663,N_12802,N_13836);
nor U16664 (N_16664,N_12434,N_14679);
nand U16665 (N_16665,N_13235,N_14201);
nand U16666 (N_16666,N_14114,N_12062);
nor U16667 (N_16667,N_12791,N_12351);
nand U16668 (N_16668,N_13346,N_13191);
nand U16669 (N_16669,N_14104,N_13277);
or U16670 (N_16670,N_13222,N_12295);
and U16671 (N_16671,N_12480,N_13062);
or U16672 (N_16672,N_14307,N_12730);
xnor U16673 (N_16673,N_13569,N_12759);
xor U16674 (N_16674,N_14289,N_12373);
or U16675 (N_16675,N_12786,N_13035);
or U16676 (N_16676,N_12684,N_14419);
nor U16677 (N_16677,N_14145,N_14814);
nor U16678 (N_16678,N_13150,N_12512);
xnor U16679 (N_16679,N_14558,N_12039);
nor U16680 (N_16680,N_12894,N_14886);
xor U16681 (N_16681,N_12859,N_12148);
xor U16682 (N_16682,N_12273,N_14301);
xor U16683 (N_16683,N_13917,N_13235);
and U16684 (N_16684,N_12050,N_13224);
and U16685 (N_16685,N_13440,N_13033);
or U16686 (N_16686,N_12294,N_12488);
and U16687 (N_16687,N_14218,N_14060);
nand U16688 (N_16688,N_12504,N_14217);
or U16689 (N_16689,N_14118,N_13205);
nand U16690 (N_16690,N_13420,N_13698);
and U16691 (N_16691,N_12804,N_14266);
nor U16692 (N_16692,N_14518,N_14310);
and U16693 (N_16693,N_12612,N_13468);
xnor U16694 (N_16694,N_13883,N_12956);
and U16695 (N_16695,N_14416,N_12499);
nand U16696 (N_16696,N_13533,N_12064);
nand U16697 (N_16697,N_13538,N_14801);
or U16698 (N_16698,N_12027,N_12653);
or U16699 (N_16699,N_12944,N_12902);
and U16700 (N_16700,N_13079,N_13126);
and U16701 (N_16701,N_14639,N_13293);
or U16702 (N_16702,N_14534,N_12516);
or U16703 (N_16703,N_14881,N_13387);
and U16704 (N_16704,N_13171,N_13480);
nand U16705 (N_16705,N_12348,N_13920);
or U16706 (N_16706,N_13268,N_13332);
or U16707 (N_16707,N_12271,N_14660);
or U16708 (N_16708,N_14534,N_14536);
xor U16709 (N_16709,N_12220,N_13543);
and U16710 (N_16710,N_13139,N_14304);
xnor U16711 (N_16711,N_13537,N_13755);
and U16712 (N_16712,N_13070,N_12049);
xor U16713 (N_16713,N_14611,N_13727);
and U16714 (N_16714,N_13301,N_14339);
or U16715 (N_16715,N_13562,N_12595);
and U16716 (N_16716,N_14134,N_13982);
nor U16717 (N_16717,N_14738,N_12917);
or U16718 (N_16718,N_12102,N_14880);
or U16719 (N_16719,N_12456,N_13713);
or U16720 (N_16720,N_12586,N_12265);
nor U16721 (N_16721,N_13675,N_12428);
xor U16722 (N_16722,N_12432,N_12854);
or U16723 (N_16723,N_14170,N_13326);
and U16724 (N_16724,N_14157,N_12504);
nor U16725 (N_16725,N_14820,N_12456);
nand U16726 (N_16726,N_14206,N_14537);
nand U16727 (N_16727,N_14256,N_12612);
or U16728 (N_16728,N_14659,N_14156);
or U16729 (N_16729,N_14556,N_13786);
or U16730 (N_16730,N_13883,N_13658);
xnor U16731 (N_16731,N_12401,N_14294);
nor U16732 (N_16732,N_13548,N_14625);
and U16733 (N_16733,N_14075,N_13406);
nor U16734 (N_16734,N_12933,N_13744);
nand U16735 (N_16735,N_14961,N_14170);
xor U16736 (N_16736,N_13281,N_12244);
nor U16737 (N_16737,N_13714,N_14992);
nor U16738 (N_16738,N_12637,N_14791);
nor U16739 (N_16739,N_14233,N_13412);
xor U16740 (N_16740,N_12791,N_13457);
xor U16741 (N_16741,N_12419,N_12998);
nand U16742 (N_16742,N_12992,N_13299);
xnor U16743 (N_16743,N_13161,N_13419);
and U16744 (N_16744,N_12890,N_14946);
nand U16745 (N_16745,N_12894,N_13473);
xor U16746 (N_16746,N_14346,N_12395);
nand U16747 (N_16747,N_13305,N_13730);
nand U16748 (N_16748,N_13301,N_14806);
and U16749 (N_16749,N_13242,N_13768);
or U16750 (N_16750,N_12000,N_12664);
or U16751 (N_16751,N_14526,N_14881);
xor U16752 (N_16752,N_12405,N_14847);
nor U16753 (N_16753,N_14632,N_14239);
and U16754 (N_16754,N_12588,N_13263);
nor U16755 (N_16755,N_13426,N_12559);
nand U16756 (N_16756,N_12098,N_14776);
and U16757 (N_16757,N_12501,N_12633);
and U16758 (N_16758,N_13171,N_12100);
nor U16759 (N_16759,N_12102,N_12927);
nand U16760 (N_16760,N_12988,N_12798);
or U16761 (N_16761,N_14025,N_14923);
nand U16762 (N_16762,N_12856,N_14869);
nor U16763 (N_16763,N_13719,N_12559);
or U16764 (N_16764,N_13629,N_13217);
and U16765 (N_16765,N_12403,N_12130);
nor U16766 (N_16766,N_12966,N_13473);
nor U16767 (N_16767,N_13608,N_12556);
nand U16768 (N_16768,N_12401,N_12853);
xor U16769 (N_16769,N_13686,N_14042);
nand U16770 (N_16770,N_12654,N_12715);
nor U16771 (N_16771,N_13330,N_13733);
nor U16772 (N_16772,N_13180,N_12272);
or U16773 (N_16773,N_13371,N_13359);
and U16774 (N_16774,N_14425,N_14581);
nor U16775 (N_16775,N_12044,N_12987);
nand U16776 (N_16776,N_14007,N_12813);
and U16777 (N_16777,N_12843,N_14812);
and U16778 (N_16778,N_14377,N_13590);
nand U16779 (N_16779,N_14433,N_12295);
nand U16780 (N_16780,N_12324,N_13031);
nand U16781 (N_16781,N_13161,N_14784);
and U16782 (N_16782,N_13650,N_13305);
nand U16783 (N_16783,N_14731,N_13731);
nor U16784 (N_16784,N_12478,N_14768);
or U16785 (N_16785,N_14568,N_12070);
and U16786 (N_16786,N_12534,N_13910);
nor U16787 (N_16787,N_14595,N_12541);
nand U16788 (N_16788,N_13297,N_14808);
xor U16789 (N_16789,N_12312,N_13595);
nand U16790 (N_16790,N_14074,N_13277);
and U16791 (N_16791,N_12222,N_13940);
nand U16792 (N_16792,N_14415,N_14157);
nand U16793 (N_16793,N_13887,N_12164);
and U16794 (N_16794,N_14777,N_12339);
xnor U16795 (N_16795,N_12870,N_12526);
or U16796 (N_16796,N_12017,N_12690);
and U16797 (N_16797,N_13069,N_14799);
nand U16798 (N_16798,N_14784,N_14585);
and U16799 (N_16799,N_13070,N_13058);
and U16800 (N_16800,N_14209,N_12661);
and U16801 (N_16801,N_13181,N_12282);
nand U16802 (N_16802,N_13094,N_13078);
xor U16803 (N_16803,N_12875,N_14030);
xnor U16804 (N_16804,N_14316,N_13729);
xnor U16805 (N_16805,N_14333,N_12889);
nor U16806 (N_16806,N_13416,N_13391);
and U16807 (N_16807,N_14176,N_13456);
xnor U16808 (N_16808,N_12383,N_13287);
nor U16809 (N_16809,N_12447,N_14047);
and U16810 (N_16810,N_13185,N_14776);
or U16811 (N_16811,N_13967,N_12961);
and U16812 (N_16812,N_12826,N_12524);
xnor U16813 (N_16813,N_14900,N_12786);
and U16814 (N_16814,N_13821,N_13588);
nand U16815 (N_16815,N_14933,N_12797);
nor U16816 (N_16816,N_12265,N_13682);
nand U16817 (N_16817,N_13802,N_12942);
and U16818 (N_16818,N_12071,N_13604);
nor U16819 (N_16819,N_13381,N_14754);
or U16820 (N_16820,N_13676,N_14706);
nand U16821 (N_16821,N_12811,N_14512);
nor U16822 (N_16822,N_14627,N_12974);
and U16823 (N_16823,N_12373,N_14592);
or U16824 (N_16824,N_13213,N_12857);
nand U16825 (N_16825,N_12661,N_14476);
or U16826 (N_16826,N_12386,N_14092);
nor U16827 (N_16827,N_14370,N_14175);
xor U16828 (N_16828,N_13156,N_14206);
nor U16829 (N_16829,N_13395,N_12597);
xnor U16830 (N_16830,N_12021,N_14913);
or U16831 (N_16831,N_14685,N_12870);
nor U16832 (N_16832,N_12523,N_14763);
xnor U16833 (N_16833,N_14920,N_12357);
or U16834 (N_16834,N_13667,N_14107);
and U16835 (N_16835,N_14883,N_12627);
nor U16836 (N_16836,N_13383,N_14651);
xnor U16837 (N_16837,N_12243,N_12641);
nor U16838 (N_16838,N_14265,N_12039);
nor U16839 (N_16839,N_12804,N_14730);
or U16840 (N_16840,N_14461,N_13595);
and U16841 (N_16841,N_14788,N_12369);
nor U16842 (N_16842,N_12408,N_14517);
nor U16843 (N_16843,N_12675,N_14453);
and U16844 (N_16844,N_14523,N_13765);
xor U16845 (N_16845,N_12157,N_12845);
nor U16846 (N_16846,N_12211,N_13911);
nor U16847 (N_16847,N_13886,N_12204);
nor U16848 (N_16848,N_13524,N_12499);
or U16849 (N_16849,N_13174,N_12656);
and U16850 (N_16850,N_13823,N_14477);
nor U16851 (N_16851,N_13677,N_12130);
and U16852 (N_16852,N_13647,N_13365);
xnor U16853 (N_16853,N_13990,N_12901);
or U16854 (N_16854,N_12298,N_13034);
nand U16855 (N_16855,N_12050,N_14732);
nand U16856 (N_16856,N_14004,N_13085);
and U16857 (N_16857,N_12062,N_14174);
xnor U16858 (N_16858,N_13477,N_13937);
xnor U16859 (N_16859,N_14175,N_14917);
nor U16860 (N_16860,N_13034,N_13220);
and U16861 (N_16861,N_14794,N_13774);
or U16862 (N_16862,N_14283,N_12823);
nor U16863 (N_16863,N_13896,N_13494);
nor U16864 (N_16864,N_13169,N_14308);
nor U16865 (N_16865,N_14797,N_13304);
and U16866 (N_16866,N_14811,N_14560);
nor U16867 (N_16867,N_14011,N_12725);
and U16868 (N_16868,N_12466,N_12059);
xnor U16869 (N_16869,N_13403,N_12627);
and U16870 (N_16870,N_14103,N_13558);
nor U16871 (N_16871,N_12326,N_12563);
nor U16872 (N_16872,N_14543,N_13305);
nor U16873 (N_16873,N_13128,N_14376);
nor U16874 (N_16874,N_12671,N_12270);
and U16875 (N_16875,N_14159,N_14420);
and U16876 (N_16876,N_14819,N_13301);
and U16877 (N_16877,N_14033,N_14100);
xor U16878 (N_16878,N_13883,N_13982);
nor U16879 (N_16879,N_14651,N_14866);
and U16880 (N_16880,N_14226,N_12451);
or U16881 (N_16881,N_12710,N_13776);
nor U16882 (N_16882,N_13895,N_12642);
or U16883 (N_16883,N_13816,N_13175);
or U16884 (N_16884,N_12768,N_13345);
or U16885 (N_16885,N_14133,N_13744);
nor U16886 (N_16886,N_12550,N_13488);
or U16887 (N_16887,N_14336,N_12814);
xnor U16888 (N_16888,N_13134,N_13069);
xnor U16889 (N_16889,N_14366,N_12947);
xor U16890 (N_16890,N_12438,N_14150);
and U16891 (N_16891,N_13844,N_12036);
xnor U16892 (N_16892,N_13005,N_13092);
xnor U16893 (N_16893,N_13523,N_12046);
nor U16894 (N_16894,N_12810,N_13353);
or U16895 (N_16895,N_13741,N_13178);
nor U16896 (N_16896,N_13144,N_13451);
and U16897 (N_16897,N_14871,N_13170);
or U16898 (N_16898,N_14297,N_14676);
or U16899 (N_16899,N_14935,N_14255);
or U16900 (N_16900,N_13410,N_12720);
xor U16901 (N_16901,N_12379,N_14970);
xnor U16902 (N_16902,N_12037,N_14677);
xor U16903 (N_16903,N_13440,N_14956);
and U16904 (N_16904,N_13367,N_12033);
and U16905 (N_16905,N_13314,N_14769);
xnor U16906 (N_16906,N_14505,N_13544);
and U16907 (N_16907,N_12909,N_12047);
xor U16908 (N_16908,N_14415,N_14939);
xnor U16909 (N_16909,N_12251,N_13446);
nor U16910 (N_16910,N_12079,N_13396);
xor U16911 (N_16911,N_12426,N_13056);
or U16912 (N_16912,N_13969,N_14200);
and U16913 (N_16913,N_14539,N_14691);
or U16914 (N_16914,N_14859,N_13588);
nand U16915 (N_16915,N_13506,N_14758);
or U16916 (N_16916,N_13510,N_13951);
and U16917 (N_16917,N_13088,N_12274);
and U16918 (N_16918,N_13544,N_14049);
and U16919 (N_16919,N_13376,N_14160);
nor U16920 (N_16920,N_13201,N_14993);
nor U16921 (N_16921,N_14256,N_14009);
nor U16922 (N_16922,N_12952,N_12705);
xnor U16923 (N_16923,N_13397,N_12019);
nand U16924 (N_16924,N_12073,N_14727);
and U16925 (N_16925,N_14075,N_13794);
and U16926 (N_16926,N_14268,N_13305);
nor U16927 (N_16927,N_14730,N_14762);
nor U16928 (N_16928,N_14710,N_12188);
xnor U16929 (N_16929,N_14681,N_13012);
or U16930 (N_16930,N_12431,N_12324);
nor U16931 (N_16931,N_13343,N_13553);
and U16932 (N_16932,N_14747,N_14083);
or U16933 (N_16933,N_12123,N_13271);
nor U16934 (N_16934,N_12069,N_13920);
or U16935 (N_16935,N_12652,N_13582);
nand U16936 (N_16936,N_14622,N_12235);
nand U16937 (N_16937,N_13627,N_14224);
xnor U16938 (N_16938,N_14681,N_12787);
and U16939 (N_16939,N_12213,N_12145);
and U16940 (N_16940,N_14556,N_14473);
xnor U16941 (N_16941,N_14782,N_12693);
nor U16942 (N_16942,N_14798,N_14626);
nand U16943 (N_16943,N_14409,N_13818);
nand U16944 (N_16944,N_12443,N_13386);
nand U16945 (N_16945,N_14906,N_14031);
xor U16946 (N_16946,N_13112,N_12605);
nor U16947 (N_16947,N_14995,N_13133);
nand U16948 (N_16948,N_13458,N_14321);
nand U16949 (N_16949,N_13312,N_12225);
nor U16950 (N_16950,N_13148,N_13359);
and U16951 (N_16951,N_14432,N_13435);
nand U16952 (N_16952,N_12148,N_12022);
or U16953 (N_16953,N_13415,N_13918);
nand U16954 (N_16954,N_13973,N_13710);
and U16955 (N_16955,N_14000,N_14990);
nor U16956 (N_16956,N_13100,N_13010);
xnor U16957 (N_16957,N_14145,N_12136);
or U16958 (N_16958,N_12687,N_12622);
and U16959 (N_16959,N_14923,N_14240);
or U16960 (N_16960,N_14714,N_13628);
or U16961 (N_16961,N_12049,N_14287);
nor U16962 (N_16962,N_14941,N_12546);
or U16963 (N_16963,N_13130,N_12759);
or U16964 (N_16964,N_12806,N_13981);
and U16965 (N_16965,N_12558,N_12799);
and U16966 (N_16966,N_14588,N_13242);
xnor U16967 (N_16967,N_12095,N_13172);
nor U16968 (N_16968,N_14778,N_13588);
xor U16969 (N_16969,N_12661,N_12165);
nor U16970 (N_16970,N_14830,N_14960);
nor U16971 (N_16971,N_14552,N_14784);
xnor U16972 (N_16972,N_13866,N_13995);
and U16973 (N_16973,N_14082,N_14490);
and U16974 (N_16974,N_13875,N_12583);
xor U16975 (N_16975,N_14182,N_14659);
nor U16976 (N_16976,N_13523,N_12345);
or U16977 (N_16977,N_14355,N_14605);
nor U16978 (N_16978,N_13119,N_14787);
nand U16979 (N_16979,N_13350,N_14436);
and U16980 (N_16980,N_13776,N_13543);
xor U16981 (N_16981,N_14595,N_13387);
nand U16982 (N_16982,N_14825,N_14056);
or U16983 (N_16983,N_13408,N_14371);
xnor U16984 (N_16984,N_13874,N_13753);
and U16985 (N_16985,N_13835,N_14370);
or U16986 (N_16986,N_12386,N_12028);
and U16987 (N_16987,N_12155,N_14005);
or U16988 (N_16988,N_12834,N_12069);
nand U16989 (N_16989,N_12846,N_12152);
nor U16990 (N_16990,N_13171,N_12630);
and U16991 (N_16991,N_12527,N_13887);
nand U16992 (N_16992,N_13054,N_12935);
nand U16993 (N_16993,N_14092,N_12561);
xnor U16994 (N_16994,N_13524,N_12454);
xor U16995 (N_16995,N_12903,N_13434);
and U16996 (N_16996,N_14344,N_12252);
nand U16997 (N_16997,N_13106,N_14806);
or U16998 (N_16998,N_14127,N_14873);
nor U16999 (N_16999,N_12232,N_14385);
xnor U17000 (N_17000,N_12785,N_13936);
nand U17001 (N_17001,N_14319,N_14351);
nand U17002 (N_17002,N_12220,N_13766);
and U17003 (N_17003,N_13292,N_12336);
and U17004 (N_17004,N_13658,N_13804);
nand U17005 (N_17005,N_12986,N_14440);
xnor U17006 (N_17006,N_14643,N_14928);
xor U17007 (N_17007,N_13830,N_12194);
nand U17008 (N_17008,N_12301,N_13078);
nand U17009 (N_17009,N_13395,N_14546);
xor U17010 (N_17010,N_12726,N_12420);
nor U17011 (N_17011,N_13666,N_12765);
or U17012 (N_17012,N_12828,N_14654);
and U17013 (N_17013,N_13611,N_13591);
nor U17014 (N_17014,N_14855,N_12278);
nor U17015 (N_17015,N_13615,N_12855);
nor U17016 (N_17016,N_12191,N_14959);
xor U17017 (N_17017,N_12081,N_13588);
nand U17018 (N_17018,N_13038,N_14380);
nand U17019 (N_17019,N_13545,N_13773);
nand U17020 (N_17020,N_14779,N_12437);
and U17021 (N_17021,N_13148,N_12824);
nand U17022 (N_17022,N_13496,N_13995);
or U17023 (N_17023,N_12322,N_13855);
nor U17024 (N_17024,N_13016,N_12564);
nor U17025 (N_17025,N_13608,N_14018);
nand U17026 (N_17026,N_14897,N_13403);
nor U17027 (N_17027,N_12052,N_12379);
nand U17028 (N_17028,N_12000,N_14369);
and U17029 (N_17029,N_12829,N_13309);
nor U17030 (N_17030,N_12844,N_14407);
nand U17031 (N_17031,N_12262,N_14834);
xnor U17032 (N_17032,N_14595,N_12947);
xnor U17033 (N_17033,N_14975,N_12352);
nor U17034 (N_17034,N_13673,N_12314);
xnor U17035 (N_17035,N_14612,N_13014);
nor U17036 (N_17036,N_13866,N_13731);
xnor U17037 (N_17037,N_14603,N_13433);
nand U17038 (N_17038,N_13662,N_12374);
xor U17039 (N_17039,N_14079,N_13439);
and U17040 (N_17040,N_13210,N_13553);
nor U17041 (N_17041,N_12827,N_14759);
nand U17042 (N_17042,N_14136,N_12135);
nand U17043 (N_17043,N_13764,N_14515);
and U17044 (N_17044,N_14905,N_12334);
and U17045 (N_17045,N_12892,N_13397);
nand U17046 (N_17046,N_12301,N_13229);
and U17047 (N_17047,N_14000,N_13709);
nor U17048 (N_17048,N_12453,N_13127);
xor U17049 (N_17049,N_13605,N_12855);
nor U17050 (N_17050,N_13831,N_14419);
or U17051 (N_17051,N_12264,N_14307);
and U17052 (N_17052,N_14107,N_12800);
or U17053 (N_17053,N_13140,N_12757);
and U17054 (N_17054,N_12592,N_14320);
or U17055 (N_17055,N_14817,N_13069);
or U17056 (N_17056,N_13693,N_13178);
xor U17057 (N_17057,N_14980,N_14199);
nand U17058 (N_17058,N_14970,N_12166);
xnor U17059 (N_17059,N_13576,N_12431);
nor U17060 (N_17060,N_13878,N_12477);
or U17061 (N_17061,N_14114,N_12680);
and U17062 (N_17062,N_12983,N_12161);
nor U17063 (N_17063,N_12957,N_12551);
nand U17064 (N_17064,N_12729,N_14143);
nor U17065 (N_17065,N_12525,N_12529);
and U17066 (N_17066,N_12927,N_14941);
and U17067 (N_17067,N_14809,N_13664);
nand U17068 (N_17068,N_12822,N_12356);
nand U17069 (N_17069,N_13108,N_14570);
nand U17070 (N_17070,N_14715,N_12903);
xnor U17071 (N_17071,N_14639,N_13611);
and U17072 (N_17072,N_13821,N_12365);
and U17073 (N_17073,N_12711,N_14407);
nor U17074 (N_17074,N_12503,N_12306);
or U17075 (N_17075,N_13977,N_12552);
nand U17076 (N_17076,N_13621,N_13214);
or U17077 (N_17077,N_12330,N_13846);
nor U17078 (N_17078,N_13645,N_13677);
or U17079 (N_17079,N_12836,N_12368);
nor U17080 (N_17080,N_14652,N_13725);
nand U17081 (N_17081,N_14632,N_13412);
nor U17082 (N_17082,N_14531,N_12868);
and U17083 (N_17083,N_13852,N_12730);
and U17084 (N_17084,N_14656,N_13138);
and U17085 (N_17085,N_14771,N_12852);
or U17086 (N_17086,N_14526,N_12110);
nand U17087 (N_17087,N_14118,N_12269);
and U17088 (N_17088,N_13638,N_14643);
or U17089 (N_17089,N_12593,N_12667);
or U17090 (N_17090,N_12946,N_14655);
or U17091 (N_17091,N_12876,N_14690);
or U17092 (N_17092,N_12193,N_12325);
and U17093 (N_17093,N_14872,N_13502);
nand U17094 (N_17094,N_14008,N_13378);
nand U17095 (N_17095,N_13949,N_14795);
or U17096 (N_17096,N_14586,N_12977);
xnor U17097 (N_17097,N_12074,N_12129);
xor U17098 (N_17098,N_14251,N_13394);
and U17099 (N_17099,N_12097,N_14260);
nand U17100 (N_17100,N_13012,N_14033);
and U17101 (N_17101,N_14690,N_12742);
or U17102 (N_17102,N_14151,N_13209);
nor U17103 (N_17103,N_13323,N_13911);
nor U17104 (N_17104,N_14038,N_12814);
and U17105 (N_17105,N_12376,N_13401);
and U17106 (N_17106,N_13205,N_14535);
xor U17107 (N_17107,N_12110,N_13750);
nor U17108 (N_17108,N_13308,N_14034);
or U17109 (N_17109,N_13282,N_14811);
xor U17110 (N_17110,N_13775,N_12215);
nor U17111 (N_17111,N_12711,N_12905);
nor U17112 (N_17112,N_14568,N_12386);
nand U17113 (N_17113,N_13523,N_14144);
or U17114 (N_17114,N_14281,N_13230);
or U17115 (N_17115,N_13929,N_13888);
nand U17116 (N_17116,N_14555,N_13527);
and U17117 (N_17117,N_12666,N_12246);
xnor U17118 (N_17118,N_14741,N_12403);
xnor U17119 (N_17119,N_14114,N_14955);
nand U17120 (N_17120,N_13420,N_12289);
xnor U17121 (N_17121,N_12237,N_13653);
xor U17122 (N_17122,N_12440,N_13242);
nor U17123 (N_17123,N_14468,N_13335);
xnor U17124 (N_17124,N_12582,N_12991);
xor U17125 (N_17125,N_13237,N_12103);
or U17126 (N_17126,N_13173,N_13729);
or U17127 (N_17127,N_12811,N_12798);
nand U17128 (N_17128,N_13857,N_13961);
nor U17129 (N_17129,N_14992,N_14816);
nor U17130 (N_17130,N_12640,N_12964);
nor U17131 (N_17131,N_13831,N_13342);
nor U17132 (N_17132,N_13804,N_12328);
and U17133 (N_17133,N_14250,N_14209);
xnor U17134 (N_17134,N_13875,N_12978);
or U17135 (N_17135,N_12392,N_13229);
nor U17136 (N_17136,N_13158,N_12407);
or U17137 (N_17137,N_13675,N_14828);
and U17138 (N_17138,N_14278,N_14069);
or U17139 (N_17139,N_13421,N_12039);
xor U17140 (N_17140,N_13016,N_13902);
and U17141 (N_17141,N_14882,N_12458);
and U17142 (N_17142,N_13742,N_12377);
and U17143 (N_17143,N_12109,N_13641);
nor U17144 (N_17144,N_13783,N_12929);
and U17145 (N_17145,N_12500,N_13575);
xor U17146 (N_17146,N_13620,N_14359);
nand U17147 (N_17147,N_13948,N_14280);
and U17148 (N_17148,N_14723,N_14727);
nor U17149 (N_17149,N_14522,N_12721);
and U17150 (N_17150,N_13517,N_12310);
and U17151 (N_17151,N_13935,N_13541);
nand U17152 (N_17152,N_13344,N_14734);
nand U17153 (N_17153,N_13813,N_14387);
and U17154 (N_17154,N_13738,N_13996);
or U17155 (N_17155,N_14216,N_14085);
or U17156 (N_17156,N_13863,N_12520);
and U17157 (N_17157,N_13493,N_14687);
or U17158 (N_17158,N_12195,N_12788);
xnor U17159 (N_17159,N_14588,N_14552);
xnor U17160 (N_17160,N_13634,N_13548);
nor U17161 (N_17161,N_13316,N_13487);
nor U17162 (N_17162,N_12909,N_14898);
xnor U17163 (N_17163,N_14050,N_12277);
xor U17164 (N_17164,N_12883,N_13792);
or U17165 (N_17165,N_13734,N_14412);
nor U17166 (N_17166,N_14775,N_13882);
or U17167 (N_17167,N_14589,N_14628);
nor U17168 (N_17168,N_14793,N_14403);
nor U17169 (N_17169,N_13420,N_12166);
nor U17170 (N_17170,N_12729,N_12330);
nand U17171 (N_17171,N_13864,N_13234);
xnor U17172 (N_17172,N_13295,N_12194);
or U17173 (N_17173,N_14821,N_14208);
or U17174 (N_17174,N_14360,N_13783);
nor U17175 (N_17175,N_12367,N_14982);
xor U17176 (N_17176,N_14528,N_12622);
nand U17177 (N_17177,N_14968,N_13050);
xor U17178 (N_17178,N_13184,N_13896);
xnor U17179 (N_17179,N_13702,N_12420);
or U17180 (N_17180,N_13941,N_13570);
and U17181 (N_17181,N_12010,N_13730);
nor U17182 (N_17182,N_12171,N_13115);
nand U17183 (N_17183,N_14436,N_14283);
nand U17184 (N_17184,N_13941,N_12195);
nand U17185 (N_17185,N_12796,N_12835);
xnor U17186 (N_17186,N_14631,N_13669);
nor U17187 (N_17187,N_13064,N_14364);
and U17188 (N_17188,N_14786,N_14557);
nor U17189 (N_17189,N_12294,N_12506);
and U17190 (N_17190,N_13967,N_14427);
nor U17191 (N_17191,N_14212,N_14293);
or U17192 (N_17192,N_13467,N_13822);
xnor U17193 (N_17193,N_14322,N_12351);
and U17194 (N_17194,N_12562,N_14713);
and U17195 (N_17195,N_14250,N_14594);
or U17196 (N_17196,N_12835,N_12244);
xnor U17197 (N_17197,N_14145,N_14368);
nor U17198 (N_17198,N_13686,N_14837);
nand U17199 (N_17199,N_12017,N_14378);
nor U17200 (N_17200,N_14229,N_12421);
and U17201 (N_17201,N_14304,N_14616);
and U17202 (N_17202,N_14775,N_14084);
xor U17203 (N_17203,N_12909,N_13608);
and U17204 (N_17204,N_13719,N_14478);
and U17205 (N_17205,N_14080,N_12841);
nor U17206 (N_17206,N_14542,N_13912);
and U17207 (N_17207,N_14484,N_12231);
nor U17208 (N_17208,N_13208,N_14643);
nand U17209 (N_17209,N_12062,N_13845);
or U17210 (N_17210,N_14489,N_13514);
xor U17211 (N_17211,N_13113,N_12038);
nor U17212 (N_17212,N_12999,N_14491);
xnor U17213 (N_17213,N_13697,N_12032);
nand U17214 (N_17214,N_14203,N_14160);
xnor U17215 (N_17215,N_12493,N_12593);
xor U17216 (N_17216,N_12873,N_12194);
nand U17217 (N_17217,N_14522,N_14521);
xnor U17218 (N_17218,N_12096,N_14788);
and U17219 (N_17219,N_12377,N_12517);
nand U17220 (N_17220,N_14544,N_12546);
xor U17221 (N_17221,N_12175,N_14696);
or U17222 (N_17222,N_13637,N_12435);
nor U17223 (N_17223,N_12807,N_12057);
nor U17224 (N_17224,N_13429,N_14306);
nand U17225 (N_17225,N_14688,N_13405);
xor U17226 (N_17226,N_14738,N_12561);
or U17227 (N_17227,N_12917,N_12244);
nor U17228 (N_17228,N_14199,N_14237);
and U17229 (N_17229,N_13175,N_13251);
and U17230 (N_17230,N_12102,N_12666);
nor U17231 (N_17231,N_14308,N_14697);
nor U17232 (N_17232,N_13651,N_13850);
or U17233 (N_17233,N_14126,N_12243);
or U17234 (N_17234,N_13300,N_13974);
or U17235 (N_17235,N_12493,N_14492);
nor U17236 (N_17236,N_13905,N_12625);
nand U17237 (N_17237,N_12878,N_12573);
xor U17238 (N_17238,N_14217,N_12960);
and U17239 (N_17239,N_13392,N_13257);
nor U17240 (N_17240,N_12541,N_14180);
nand U17241 (N_17241,N_14886,N_14116);
and U17242 (N_17242,N_13785,N_14868);
xnor U17243 (N_17243,N_13832,N_14087);
xor U17244 (N_17244,N_14913,N_12488);
and U17245 (N_17245,N_14814,N_13239);
and U17246 (N_17246,N_13056,N_12229);
xor U17247 (N_17247,N_14079,N_13721);
and U17248 (N_17248,N_13343,N_14712);
nor U17249 (N_17249,N_12953,N_12256);
and U17250 (N_17250,N_12172,N_13631);
xor U17251 (N_17251,N_12040,N_13206);
xnor U17252 (N_17252,N_12376,N_12923);
nor U17253 (N_17253,N_12781,N_12487);
xnor U17254 (N_17254,N_13982,N_12568);
nand U17255 (N_17255,N_12737,N_12885);
nand U17256 (N_17256,N_12971,N_13186);
xnor U17257 (N_17257,N_14884,N_13747);
or U17258 (N_17258,N_13588,N_14817);
xnor U17259 (N_17259,N_12346,N_14171);
nand U17260 (N_17260,N_13987,N_13382);
nand U17261 (N_17261,N_13433,N_13155);
or U17262 (N_17262,N_12862,N_14118);
and U17263 (N_17263,N_14827,N_13145);
nand U17264 (N_17264,N_13630,N_14713);
nor U17265 (N_17265,N_14464,N_12461);
xnor U17266 (N_17266,N_12827,N_14652);
nor U17267 (N_17267,N_14300,N_13023);
or U17268 (N_17268,N_12446,N_13517);
and U17269 (N_17269,N_14719,N_13381);
nand U17270 (N_17270,N_13419,N_13688);
nand U17271 (N_17271,N_12923,N_12419);
nor U17272 (N_17272,N_13812,N_12178);
nor U17273 (N_17273,N_12996,N_12944);
xor U17274 (N_17274,N_12057,N_12801);
xor U17275 (N_17275,N_14701,N_14167);
or U17276 (N_17276,N_14051,N_13857);
xor U17277 (N_17277,N_14761,N_13152);
nor U17278 (N_17278,N_12130,N_14676);
xnor U17279 (N_17279,N_12002,N_14268);
nand U17280 (N_17280,N_14245,N_12668);
and U17281 (N_17281,N_13339,N_14048);
and U17282 (N_17282,N_14968,N_13114);
nand U17283 (N_17283,N_13825,N_13223);
nand U17284 (N_17284,N_12384,N_14189);
or U17285 (N_17285,N_12150,N_13606);
nor U17286 (N_17286,N_13439,N_14095);
and U17287 (N_17287,N_14313,N_13726);
nor U17288 (N_17288,N_14552,N_13312);
nor U17289 (N_17289,N_12062,N_13587);
nand U17290 (N_17290,N_12488,N_12915);
and U17291 (N_17291,N_13672,N_14052);
nand U17292 (N_17292,N_13938,N_12501);
nor U17293 (N_17293,N_14959,N_14833);
xnor U17294 (N_17294,N_12412,N_13547);
xor U17295 (N_17295,N_13903,N_14641);
nor U17296 (N_17296,N_13015,N_14028);
and U17297 (N_17297,N_14485,N_13180);
and U17298 (N_17298,N_12137,N_14807);
xnor U17299 (N_17299,N_13758,N_14638);
nor U17300 (N_17300,N_12756,N_12562);
nand U17301 (N_17301,N_14095,N_12461);
nand U17302 (N_17302,N_12675,N_13029);
nor U17303 (N_17303,N_13618,N_14297);
nor U17304 (N_17304,N_13785,N_14347);
nor U17305 (N_17305,N_14887,N_13189);
xnor U17306 (N_17306,N_12606,N_13279);
nor U17307 (N_17307,N_14244,N_12655);
nand U17308 (N_17308,N_13872,N_13952);
nor U17309 (N_17309,N_12050,N_14466);
nor U17310 (N_17310,N_13783,N_12618);
nor U17311 (N_17311,N_13773,N_13889);
nor U17312 (N_17312,N_14162,N_13803);
or U17313 (N_17313,N_12822,N_14643);
and U17314 (N_17314,N_14596,N_12419);
nor U17315 (N_17315,N_13626,N_14888);
or U17316 (N_17316,N_12385,N_12135);
or U17317 (N_17317,N_13560,N_13769);
and U17318 (N_17318,N_14322,N_14470);
and U17319 (N_17319,N_12231,N_13232);
nor U17320 (N_17320,N_14784,N_14662);
nor U17321 (N_17321,N_13927,N_13251);
nor U17322 (N_17322,N_13823,N_12402);
nand U17323 (N_17323,N_12004,N_12353);
nand U17324 (N_17324,N_14521,N_12642);
or U17325 (N_17325,N_12280,N_12647);
and U17326 (N_17326,N_12959,N_13038);
nand U17327 (N_17327,N_13084,N_14650);
nor U17328 (N_17328,N_13522,N_12432);
or U17329 (N_17329,N_12663,N_12639);
nor U17330 (N_17330,N_14160,N_13798);
nor U17331 (N_17331,N_13396,N_12103);
nand U17332 (N_17332,N_12870,N_13732);
nand U17333 (N_17333,N_13632,N_12543);
nor U17334 (N_17334,N_14929,N_13878);
nand U17335 (N_17335,N_12309,N_12822);
or U17336 (N_17336,N_12315,N_12578);
or U17337 (N_17337,N_12172,N_14668);
nand U17338 (N_17338,N_13404,N_14776);
xnor U17339 (N_17339,N_13973,N_14055);
xor U17340 (N_17340,N_14676,N_13212);
nand U17341 (N_17341,N_13403,N_14336);
or U17342 (N_17342,N_12046,N_12073);
nand U17343 (N_17343,N_13793,N_12446);
or U17344 (N_17344,N_12270,N_12933);
and U17345 (N_17345,N_14814,N_12643);
nor U17346 (N_17346,N_12814,N_12420);
nor U17347 (N_17347,N_13279,N_14880);
nand U17348 (N_17348,N_14055,N_12996);
or U17349 (N_17349,N_14197,N_12849);
nor U17350 (N_17350,N_13147,N_12621);
nor U17351 (N_17351,N_13186,N_13577);
or U17352 (N_17352,N_13017,N_14019);
nor U17353 (N_17353,N_13131,N_13288);
nand U17354 (N_17354,N_14590,N_12433);
or U17355 (N_17355,N_14804,N_12058);
or U17356 (N_17356,N_12956,N_13933);
or U17357 (N_17357,N_12903,N_14381);
or U17358 (N_17358,N_14043,N_13547);
or U17359 (N_17359,N_12513,N_12690);
and U17360 (N_17360,N_14242,N_14523);
xor U17361 (N_17361,N_14490,N_14830);
nor U17362 (N_17362,N_12043,N_14698);
nand U17363 (N_17363,N_12961,N_13905);
nor U17364 (N_17364,N_13539,N_13894);
nor U17365 (N_17365,N_13866,N_13207);
nand U17366 (N_17366,N_12684,N_14910);
xnor U17367 (N_17367,N_13599,N_13795);
nor U17368 (N_17368,N_13060,N_12170);
nor U17369 (N_17369,N_14203,N_13777);
nand U17370 (N_17370,N_12284,N_12674);
xor U17371 (N_17371,N_14427,N_13143);
and U17372 (N_17372,N_13725,N_13200);
xnor U17373 (N_17373,N_12350,N_13994);
nand U17374 (N_17374,N_13264,N_14551);
nor U17375 (N_17375,N_12611,N_14828);
nand U17376 (N_17376,N_12857,N_12510);
and U17377 (N_17377,N_12946,N_13143);
xnor U17378 (N_17378,N_13796,N_12938);
xor U17379 (N_17379,N_12104,N_12059);
nor U17380 (N_17380,N_13969,N_14605);
xor U17381 (N_17381,N_13360,N_12081);
and U17382 (N_17382,N_14256,N_13439);
xor U17383 (N_17383,N_13864,N_12771);
xor U17384 (N_17384,N_13021,N_12702);
nor U17385 (N_17385,N_12976,N_13503);
nand U17386 (N_17386,N_12515,N_12027);
nor U17387 (N_17387,N_13882,N_14505);
nor U17388 (N_17388,N_12148,N_12417);
and U17389 (N_17389,N_12640,N_12017);
or U17390 (N_17390,N_12972,N_14079);
nand U17391 (N_17391,N_12431,N_12147);
xor U17392 (N_17392,N_13655,N_14802);
or U17393 (N_17393,N_13632,N_12421);
nor U17394 (N_17394,N_12323,N_13530);
xor U17395 (N_17395,N_14026,N_14426);
xor U17396 (N_17396,N_13860,N_12086);
nand U17397 (N_17397,N_13796,N_13179);
and U17398 (N_17398,N_14538,N_14848);
nor U17399 (N_17399,N_14482,N_14180);
or U17400 (N_17400,N_12870,N_13231);
nor U17401 (N_17401,N_14451,N_14352);
or U17402 (N_17402,N_13846,N_12211);
and U17403 (N_17403,N_13440,N_13341);
nand U17404 (N_17404,N_13404,N_12811);
xnor U17405 (N_17405,N_13842,N_14319);
nand U17406 (N_17406,N_13419,N_13867);
nand U17407 (N_17407,N_13645,N_12696);
nand U17408 (N_17408,N_14697,N_13973);
nor U17409 (N_17409,N_13886,N_12957);
and U17410 (N_17410,N_13750,N_13607);
nor U17411 (N_17411,N_14576,N_14093);
and U17412 (N_17412,N_14412,N_12904);
and U17413 (N_17413,N_14534,N_14066);
and U17414 (N_17414,N_12199,N_13195);
and U17415 (N_17415,N_12858,N_13451);
xor U17416 (N_17416,N_12580,N_12991);
nor U17417 (N_17417,N_13898,N_14162);
or U17418 (N_17418,N_12123,N_12693);
or U17419 (N_17419,N_14557,N_14178);
or U17420 (N_17420,N_13716,N_12018);
and U17421 (N_17421,N_12826,N_12363);
or U17422 (N_17422,N_13902,N_13875);
or U17423 (N_17423,N_14209,N_13766);
xor U17424 (N_17424,N_13266,N_12826);
and U17425 (N_17425,N_12099,N_12541);
or U17426 (N_17426,N_13041,N_13831);
and U17427 (N_17427,N_13971,N_13189);
or U17428 (N_17428,N_13752,N_13242);
nor U17429 (N_17429,N_12405,N_13950);
xnor U17430 (N_17430,N_13571,N_14921);
xnor U17431 (N_17431,N_13344,N_12740);
nand U17432 (N_17432,N_13733,N_14219);
nand U17433 (N_17433,N_14592,N_12835);
nor U17434 (N_17434,N_14191,N_13439);
and U17435 (N_17435,N_13345,N_14922);
and U17436 (N_17436,N_12802,N_12898);
xor U17437 (N_17437,N_12738,N_12413);
nand U17438 (N_17438,N_14578,N_13038);
nor U17439 (N_17439,N_13839,N_14928);
nor U17440 (N_17440,N_12216,N_13618);
and U17441 (N_17441,N_13422,N_13295);
nand U17442 (N_17442,N_13520,N_12202);
xor U17443 (N_17443,N_14143,N_13145);
and U17444 (N_17444,N_14629,N_12157);
and U17445 (N_17445,N_13172,N_12872);
or U17446 (N_17446,N_14544,N_14389);
nand U17447 (N_17447,N_13291,N_12462);
xor U17448 (N_17448,N_13657,N_12582);
and U17449 (N_17449,N_14488,N_14555);
xnor U17450 (N_17450,N_13389,N_14916);
and U17451 (N_17451,N_14728,N_13437);
nor U17452 (N_17452,N_12522,N_13713);
xor U17453 (N_17453,N_14065,N_13558);
or U17454 (N_17454,N_14795,N_12490);
xnor U17455 (N_17455,N_14019,N_12183);
xnor U17456 (N_17456,N_14159,N_14516);
nor U17457 (N_17457,N_14458,N_12957);
nand U17458 (N_17458,N_12663,N_13430);
and U17459 (N_17459,N_12601,N_12739);
xor U17460 (N_17460,N_12387,N_12579);
nor U17461 (N_17461,N_12418,N_14019);
and U17462 (N_17462,N_14455,N_12599);
nand U17463 (N_17463,N_12914,N_13457);
nor U17464 (N_17464,N_12858,N_12297);
xor U17465 (N_17465,N_13883,N_13697);
nor U17466 (N_17466,N_13992,N_14520);
or U17467 (N_17467,N_14597,N_12125);
and U17468 (N_17468,N_13960,N_14800);
nand U17469 (N_17469,N_12180,N_14999);
nor U17470 (N_17470,N_14009,N_12512);
and U17471 (N_17471,N_13767,N_14386);
nor U17472 (N_17472,N_14479,N_14490);
or U17473 (N_17473,N_13056,N_14950);
or U17474 (N_17474,N_14627,N_13218);
xnor U17475 (N_17475,N_14429,N_14050);
and U17476 (N_17476,N_13289,N_12813);
nand U17477 (N_17477,N_13826,N_14502);
nor U17478 (N_17478,N_14095,N_14030);
nand U17479 (N_17479,N_14140,N_14023);
nand U17480 (N_17480,N_14174,N_14415);
nor U17481 (N_17481,N_14998,N_14350);
nor U17482 (N_17482,N_13942,N_14192);
nor U17483 (N_17483,N_13292,N_12815);
nor U17484 (N_17484,N_13956,N_13363);
and U17485 (N_17485,N_14939,N_14201);
and U17486 (N_17486,N_14261,N_12495);
nor U17487 (N_17487,N_12490,N_12603);
xor U17488 (N_17488,N_13667,N_13324);
xnor U17489 (N_17489,N_12640,N_12301);
and U17490 (N_17490,N_13673,N_14015);
nor U17491 (N_17491,N_13392,N_13178);
xor U17492 (N_17492,N_12396,N_12811);
xor U17493 (N_17493,N_13483,N_14774);
and U17494 (N_17494,N_14189,N_14040);
xor U17495 (N_17495,N_13475,N_13970);
nor U17496 (N_17496,N_12695,N_14509);
nand U17497 (N_17497,N_14809,N_13547);
xor U17498 (N_17498,N_12668,N_12433);
and U17499 (N_17499,N_14565,N_13956);
nor U17500 (N_17500,N_14367,N_14923);
and U17501 (N_17501,N_13330,N_13341);
nand U17502 (N_17502,N_14279,N_12564);
nand U17503 (N_17503,N_14808,N_14458);
nand U17504 (N_17504,N_14593,N_12120);
nor U17505 (N_17505,N_14633,N_13258);
xnor U17506 (N_17506,N_12942,N_13599);
xor U17507 (N_17507,N_12197,N_12111);
nor U17508 (N_17508,N_13319,N_12793);
and U17509 (N_17509,N_12012,N_13392);
xnor U17510 (N_17510,N_14294,N_13836);
or U17511 (N_17511,N_12888,N_14278);
or U17512 (N_17512,N_13653,N_14438);
nor U17513 (N_17513,N_13480,N_12351);
nand U17514 (N_17514,N_12284,N_14170);
or U17515 (N_17515,N_12585,N_12599);
or U17516 (N_17516,N_12832,N_13336);
or U17517 (N_17517,N_13614,N_14754);
nor U17518 (N_17518,N_12937,N_14455);
nand U17519 (N_17519,N_14331,N_13147);
nand U17520 (N_17520,N_14257,N_13283);
or U17521 (N_17521,N_12227,N_14869);
or U17522 (N_17522,N_12583,N_12004);
nor U17523 (N_17523,N_14302,N_13403);
and U17524 (N_17524,N_12256,N_12715);
or U17525 (N_17525,N_13931,N_13700);
or U17526 (N_17526,N_14505,N_14349);
nor U17527 (N_17527,N_13979,N_14645);
nor U17528 (N_17528,N_14484,N_12222);
or U17529 (N_17529,N_14318,N_12535);
and U17530 (N_17530,N_12111,N_12992);
or U17531 (N_17531,N_14493,N_14317);
and U17532 (N_17532,N_14058,N_14633);
and U17533 (N_17533,N_12112,N_13627);
and U17534 (N_17534,N_12866,N_13661);
xnor U17535 (N_17535,N_13755,N_14218);
xnor U17536 (N_17536,N_12600,N_14973);
xnor U17537 (N_17537,N_14546,N_12579);
nand U17538 (N_17538,N_12394,N_13406);
nor U17539 (N_17539,N_13817,N_14594);
nand U17540 (N_17540,N_12730,N_14812);
xor U17541 (N_17541,N_12823,N_14630);
and U17542 (N_17542,N_14486,N_12587);
nand U17543 (N_17543,N_14246,N_13580);
nor U17544 (N_17544,N_14641,N_12021);
or U17545 (N_17545,N_14773,N_14383);
nand U17546 (N_17546,N_14560,N_13116);
nand U17547 (N_17547,N_12785,N_12134);
and U17548 (N_17548,N_13055,N_13024);
nor U17549 (N_17549,N_12737,N_13888);
nor U17550 (N_17550,N_12596,N_14582);
nor U17551 (N_17551,N_12462,N_13600);
xnor U17552 (N_17552,N_14326,N_12195);
nand U17553 (N_17553,N_14713,N_12818);
nor U17554 (N_17554,N_13208,N_13166);
and U17555 (N_17555,N_14073,N_14845);
xnor U17556 (N_17556,N_12745,N_14621);
or U17557 (N_17557,N_13922,N_14287);
nor U17558 (N_17558,N_12962,N_12970);
or U17559 (N_17559,N_13971,N_12566);
and U17560 (N_17560,N_14889,N_12810);
xor U17561 (N_17561,N_13893,N_14041);
nand U17562 (N_17562,N_12192,N_12840);
xnor U17563 (N_17563,N_14644,N_13113);
nor U17564 (N_17564,N_14108,N_13679);
nand U17565 (N_17565,N_12388,N_13392);
xor U17566 (N_17566,N_13354,N_12829);
xnor U17567 (N_17567,N_12815,N_12834);
or U17568 (N_17568,N_13700,N_13270);
nor U17569 (N_17569,N_12808,N_12144);
nor U17570 (N_17570,N_14454,N_14584);
xor U17571 (N_17571,N_12745,N_13398);
and U17572 (N_17572,N_13186,N_14701);
xor U17573 (N_17573,N_14452,N_12430);
xor U17574 (N_17574,N_12606,N_14630);
or U17575 (N_17575,N_13871,N_13676);
or U17576 (N_17576,N_12685,N_13832);
nand U17577 (N_17577,N_13686,N_13735);
nor U17578 (N_17578,N_14844,N_14178);
nand U17579 (N_17579,N_12585,N_14335);
or U17580 (N_17580,N_13271,N_12492);
xnor U17581 (N_17581,N_12830,N_13693);
nand U17582 (N_17582,N_13062,N_13295);
nor U17583 (N_17583,N_13664,N_14487);
or U17584 (N_17584,N_12613,N_12089);
nand U17585 (N_17585,N_12795,N_13227);
and U17586 (N_17586,N_13997,N_12405);
nand U17587 (N_17587,N_14935,N_14821);
or U17588 (N_17588,N_13592,N_14891);
nor U17589 (N_17589,N_13559,N_12735);
xor U17590 (N_17590,N_13110,N_12571);
nor U17591 (N_17591,N_13984,N_14016);
and U17592 (N_17592,N_14766,N_14739);
nand U17593 (N_17593,N_12452,N_12105);
nor U17594 (N_17594,N_12066,N_14303);
or U17595 (N_17595,N_13625,N_13801);
xor U17596 (N_17596,N_12376,N_14154);
and U17597 (N_17597,N_14029,N_13204);
or U17598 (N_17598,N_14863,N_13348);
nor U17599 (N_17599,N_13448,N_14542);
or U17600 (N_17600,N_12985,N_13528);
xor U17601 (N_17601,N_12890,N_13830);
and U17602 (N_17602,N_14718,N_13434);
xnor U17603 (N_17603,N_13154,N_13315);
nor U17604 (N_17604,N_13366,N_13532);
nand U17605 (N_17605,N_12026,N_14680);
xor U17606 (N_17606,N_12053,N_13879);
or U17607 (N_17607,N_13960,N_13200);
nor U17608 (N_17608,N_12559,N_14706);
nand U17609 (N_17609,N_12958,N_13901);
nor U17610 (N_17610,N_14044,N_13193);
or U17611 (N_17611,N_13522,N_14385);
xnor U17612 (N_17612,N_12219,N_14115);
and U17613 (N_17613,N_13009,N_13088);
nor U17614 (N_17614,N_13197,N_13098);
nand U17615 (N_17615,N_14012,N_13435);
and U17616 (N_17616,N_12938,N_13572);
and U17617 (N_17617,N_12309,N_14411);
xnor U17618 (N_17618,N_12403,N_13036);
and U17619 (N_17619,N_14215,N_13885);
nand U17620 (N_17620,N_13894,N_14982);
nand U17621 (N_17621,N_12818,N_12698);
nand U17622 (N_17622,N_12897,N_14791);
nand U17623 (N_17623,N_14813,N_12992);
xor U17624 (N_17624,N_14092,N_14567);
xnor U17625 (N_17625,N_13266,N_14213);
and U17626 (N_17626,N_14019,N_13682);
xnor U17627 (N_17627,N_12822,N_14348);
xor U17628 (N_17628,N_12200,N_13986);
or U17629 (N_17629,N_13269,N_13461);
and U17630 (N_17630,N_14646,N_14556);
nand U17631 (N_17631,N_13279,N_13320);
nand U17632 (N_17632,N_14254,N_14108);
and U17633 (N_17633,N_12207,N_12202);
or U17634 (N_17634,N_14298,N_12479);
and U17635 (N_17635,N_14072,N_13860);
nor U17636 (N_17636,N_12006,N_12090);
xor U17637 (N_17637,N_13184,N_14470);
and U17638 (N_17638,N_13265,N_14620);
or U17639 (N_17639,N_13442,N_14409);
nand U17640 (N_17640,N_14115,N_14960);
and U17641 (N_17641,N_14725,N_14931);
nor U17642 (N_17642,N_13776,N_12501);
nand U17643 (N_17643,N_14578,N_14398);
and U17644 (N_17644,N_14686,N_12363);
and U17645 (N_17645,N_13633,N_13584);
xor U17646 (N_17646,N_12751,N_13802);
or U17647 (N_17647,N_14314,N_14061);
and U17648 (N_17648,N_14125,N_14508);
or U17649 (N_17649,N_14697,N_13945);
and U17650 (N_17650,N_12408,N_13152);
nor U17651 (N_17651,N_12030,N_14717);
or U17652 (N_17652,N_12023,N_13608);
or U17653 (N_17653,N_13640,N_12283);
nor U17654 (N_17654,N_13626,N_14589);
xnor U17655 (N_17655,N_12337,N_14466);
and U17656 (N_17656,N_12096,N_14239);
xor U17657 (N_17657,N_14452,N_12943);
nor U17658 (N_17658,N_13846,N_12276);
nor U17659 (N_17659,N_14972,N_12199);
and U17660 (N_17660,N_14471,N_14667);
nor U17661 (N_17661,N_13294,N_13726);
nor U17662 (N_17662,N_12147,N_14674);
or U17663 (N_17663,N_14008,N_12350);
nand U17664 (N_17664,N_14507,N_14017);
xor U17665 (N_17665,N_14019,N_13852);
nor U17666 (N_17666,N_12586,N_12522);
xor U17667 (N_17667,N_12589,N_12649);
nor U17668 (N_17668,N_12164,N_14066);
and U17669 (N_17669,N_13924,N_12395);
xor U17670 (N_17670,N_12077,N_12656);
or U17671 (N_17671,N_14503,N_14917);
or U17672 (N_17672,N_14369,N_13432);
nor U17673 (N_17673,N_13914,N_12342);
or U17674 (N_17674,N_12886,N_14027);
xnor U17675 (N_17675,N_13288,N_12808);
or U17676 (N_17676,N_12424,N_12659);
nor U17677 (N_17677,N_13699,N_14923);
or U17678 (N_17678,N_13433,N_12915);
nand U17679 (N_17679,N_14876,N_12826);
and U17680 (N_17680,N_12827,N_14531);
nand U17681 (N_17681,N_13143,N_13657);
nor U17682 (N_17682,N_12220,N_12782);
nand U17683 (N_17683,N_12052,N_13898);
or U17684 (N_17684,N_12611,N_12846);
nor U17685 (N_17685,N_12017,N_14523);
nand U17686 (N_17686,N_14309,N_13869);
nand U17687 (N_17687,N_13697,N_12979);
nor U17688 (N_17688,N_12911,N_13907);
nor U17689 (N_17689,N_12874,N_14367);
nand U17690 (N_17690,N_12888,N_12890);
or U17691 (N_17691,N_14726,N_14422);
nand U17692 (N_17692,N_12204,N_14569);
or U17693 (N_17693,N_12470,N_14743);
and U17694 (N_17694,N_14604,N_14912);
or U17695 (N_17695,N_14016,N_13950);
xnor U17696 (N_17696,N_14101,N_12211);
xnor U17697 (N_17697,N_13346,N_13648);
and U17698 (N_17698,N_12804,N_14935);
or U17699 (N_17699,N_12080,N_12444);
xor U17700 (N_17700,N_13158,N_13683);
or U17701 (N_17701,N_12393,N_12021);
nor U17702 (N_17702,N_14233,N_14059);
nand U17703 (N_17703,N_13582,N_13881);
or U17704 (N_17704,N_12008,N_14791);
and U17705 (N_17705,N_14273,N_13659);
or U17706 (N_17706,N_14847,N_13068);
xor U17707 (N_17707,N_14808,N_12971);
xor U17708 (N_17708,N_13777,N_12989);
nand U17709 (N_17709,N_14439,N_14143);
or U17710 (N_17710,N_12100,N_13992);
xor U17711 (N_17711,N_12925,N_12525);
nand U17712 (N_17712,N_13657,N_14141);
nand U17713 (N_17713,N_14456,N_14555);
xor U17714 (N_17714,N_12782,N_14339);
xor U17715 (N_17715,N_14872,N_13917);
and U17716 (N_17716,N_12948,N_14666);
nor U17717 (N_17717,N_14842,N_12830);
or U17718 (N_17718,N_13138,N_12240);
or U17719 (N_17719,N_13608,N_14568);
nor U17720 (N_17720,N_13474,N_13191);
nor U17721 (N_17721,N_14016,N_12963);
and U17722 (N_17722,N_13981,N_13378);
xnor U17723 (N_17723,N_14130,N_13642);
and U17724 (N_17724,N_12850,N_13032);
nor U17725 (N_17725,N_14055,N_13365);
nand U17726 (N_17726,N_12277,N_12512);
nand U17727 (N_17727,N_14047,N_14271);
nor U17728 (N_17728,N_14013,N_12493);
or U17729 (N_17729,N_13755,N_14769);
and U17730 (N_17730,N_13774,N_14819);
and U17731 (N_17731,N_14291,N_14677);
and U17732 (N_17732,N_12870,N_12104);
and U17733 (N_17733,N_12841,N_14053);
nand U17734 (N_17734,N_14279,N_13016);
or U17735 (N_17735,N_14669,N_13053);
xor U17736 (N_17736,N_13771,N_13866);
nand U17737 (N_17737,N_14873,N_12712);
or U17738 (N_17738,N_12218,N_14557);
nand U17739 (N_17739,N_13799,N_13631);
nor U17740 (N_17740,N_12788,N_12998);
xnor U17741 (N_17741,N_12235,N_12023);
nor U17742 (N_17742,N_13333,N_13563);
or U17743 (N_17743,N_13514,N_14708);
nor U17744 (N_17744,N_13099,N_13189);
or U17745 (N_17745,N_12098,N_14940);
and U17746 (N_17746,N_13397,N_14015);
and U17747 (N_17747,N_14240,N_12987);
xnor U17748 (N_17748,N_14224,N_12623);
xnor U17749 (N_17749,N_12074,N_14811);
nor U17750 (N_17750,N_14991,N_13629);
nand U17751 (N_17751,N_13227,N_13024);
nand U17752 (N_17752,N_13481,N_12357);
or U17753 (N_17753,N_12482,N_12214);
or U17754 (N_17754,N_14824,N_12156);
or U17755 (N_17755,N_12243,N_12395);
and U17756 (N_17756,N_12009,N_12909);
nand U17757 (N_17757,N_14806,N_13282);
nand U17758 (N_17758,N_12394,N_14410);
xnor U17759 (N_17759,N_13986,N_13289);
and U17760 (N_17760,N_14171,N_13497);
or U17761 (N_17761,N_13912,N_12864);
nor U17762 (N_17762,N_12679,N_13576);
and U17763 (N_17763,N_14533,N_14463);
nand U17764 (N_17764,N_13020,N_12203);
xnor U17765 (N_17765,N_13156,N_13667);
or U17766 (N_17766,N_12449,N_12034);
nand U17767 (N_17767,N_14233,N_14541);
and U17768 (N_17768,N_14352,N_13304);
nor U17769 (N_17769,N_14002,N_14283);
xnor U17770 (N_17770,N_13740,N_14816);
nor U17771 (N_17771,N_13289,N_13199);
or U17772 (N_17772,N_12734,N_12549);
nand U17773 (N_17773,N_12455,N_13226);
and U17774 (N_17774,N_14566,N_14043);
nand U17775 (N_17775,N_13554,N_12603);
xor U17776 (N_17776,N_14988,N_14175);
and U17777 (N_17777,N_12885,N_14605);
xor U17778 (N_17778,N_13034,N_14633);
nand U17779 (N_17779,N_14200,N_14312);
and U17780 (N_17780,N_12384,N_12983);
nor U17781 (N_17781,N_12932,N_13762);
xor U17782 (N_17782,N_13376,N_14459);
xnor U17783 (N_17783,N_14060,N_13631);
nor U17784 (N_17784,N_12396,N_12747);
or U17785 (N_17785,N_14732,N_13664);
and U17786 (N_17786,N_14751,N_13062);
and U17787 (N_17787,N_12816,N_14009);
or U17788 (N_17788,N_12206,N_12031);
or U17789 (N_17789,N_14014,N_12012);
nor U17790 (N_17790,N_12678,N_13152);
nor U17791 (N_17791,N_13986,N_12802);
xnor U17792 (N_17792,N_13543,N_13619);
and U17793 (N_17793,N_12451,N_14349);
nor U17794 (N_17794,N_12789,N_12856);
or U17795 (N_17795,N_14704,N_14770);
and U17796 (N_17796,N_12008,N_12493);
and U17797 (N_17797,N_12725,N_12605);
or U17798 (N_17798,N_12184,N_14270);
and U17799 (N_17799,N_12598,N_12952);
or U17800 (N_17800,N_13825,N_13721);
or U17801 (N_17801,N_12794,N_13641);
nand U17802 (N_17802,N_13767,N_12814);
xnor U17803 (N_17803,N_13369,N_13718);
or U17804 (N_17804,N_12940,N_13512);
or U17805 (N_17805,N_13315,N_14739);
and U17806 (N_17806,N_12166,N_13722);
nand U17807 (N_17807,N_14554,N_13518);
nor U17808 (N_17808,N_14710,N_14318);
nand U17809 (N_17809,N_12451,N_12970);
nor U17810 (N_17810,N_13749,N_12723);
and U17811 (N_17811,N_12518,N_12074);
or U17812 (N_17812,N_12900,N_12202);
xor U17813 (N_17813,N_14738,N_13659);
nor U17814 (N_17814,N_12314,N_12452);
xor U17815 (N_17815,N_14232,N_13388);
or U17816 (N_17816,N_13862,N_12669);
or U17817 (N_17817,N_13200,N_12639);
nand U17818 (N_17818,N_14623,N_12010);
or U17819 (N_17819,N_12036,N_14871);
and U17820 (N_17820,N_12922,N_13249);
and U17821 (N_17821,N_12021,N_13374);
nor U17822 (N_17822,N_12490,N_12422);
nor U17823 (N_17823,N_12255,N_14664);
and U17824 (N_17824,N_14348,N_12746);
nand U17825 (N_17825,N_13720,N_13884);
xnor U17826 (N_17826,N_14209,N_12127);
or U17827 (N_17827,N_13378,N_14521);
and U17828 (N_17828,N_14095,N_13374);
or U17829 (N_17829,N_13136,N_14093);
xor U17830 (N_17830,N_14926,N_14528);
nor U17831 (N_17831,N_13550,N_14793);
nand U17832 (N_17832,N_14978,N_13396);
xnor U17833 (N_17833,N_12209,N_13826);
nor U17834 (N_17834,N_13922,N_12544);
or U17835 (N_17835,N_14766,N_12277);
nor U17836 (N_17836,N_13572,N_13037);
xnor U17837 (N_17837,N_14955,N_12221);
and U17838 (N_17838,N_14899,N_12193);
xnor U17839 (N_17839,N_13559,N_13203);
and U17840 (N_17840,N_13435,N_13543);
nand U17841 (N_17841,N_13255,N_12467);
nand U17842 (N_17842,N_12807,N_13054);
or U17843 (N_17843,N_14898,N_13084);
nand U17844 (N_17844,N_14771,N_12330);
or U17845 (N_17845,N_13904,N_12158);
xor U17846 (N_17846,N_14156,N_13808);
xor U17847 (N_17847,N_13281,N_13645);
nor U17848 (N_17848,N_14489,N_14321);
or U17849 (N_17849,N_13423,N_14468);
nand U17850 (N_17850,N_14514,N_13427);
nor U17851 (N_17851,N_13678,N_13494);
nand U17852 (N_17852,N_14569,N_14793);
and U17853 (N_17853,N_13923,N_14051);
and U17854 (N_17854,N_13922,N_12351);
xor U17855 (N_17855,N_13506,N_14265);
nor U17856 (N_17856,N_12197,N_12615);
or U17857 (N_17857,N_13936,N_13045);
or U17858 (N_17858,N_14756,N_13778);
and U17859 (N_17859,N_14486,N_13822);
xor U17860 (N_17860,N_13759,N_14489);
xnor U17861 (N_17861,N_13437,N_13571);
xor U17862 (N_17862,N_13881,N_14532);
and U17863 (N_17863,N_12095,N_14741);
nand U17864 (N_17864,N_13695,N_13176);
nand U17865 (N_17865,N_14920,N_13186);
nand U17866 (N_17866,N_14763,N_12788);
xnor U17867 (N_17867,N_14645,N_13353);
xnor U17868 (N_17868,N_13162,N_13797);
nor U17869 (N_17869,N_13591,N_14559);
and U17870 (N_17870,N_14081,N_14827);
or U17871 (N_17871,N_12943,N_13339);
nand U17872 (N_17872,N_14265,N_12720);
nand U17873 (N_17873,N_13830,N_13091);
or U17874 (N_17874,N_13947,N_14785);
or U17875 (N_17875,N_12517,N_14740);
nand U17876 (N_17876,N_13140,N_12223);
nand U17877 (N_17877,N_14457,N_12458);
nand U17878 (N_17878,N_14212,N_12646);
nand U17879 (N_17879,N_13817,N_13787);
xnor U17880 (N_17880,N_12622,N_12170);
nor U17881 (N_17881,N_13325,N_14838);
nand U17882 (N_17882,N_14530,N_12221);
and U17883 (N_17883,N_12284,N_12413);
or U17884 (N_17884,N_13402,N_13805);
nor U17885 (N_17885,N_14151,N_12176);
nand U17886 (N_17886,N_13095,N_14067);
or U17887 (N_17887,N_13040,N_12325);
and U17888 (N_17888,N_14199,N_13058);
or U17889 (N_17889,N_13879,N_12472);
nand U17890 (N_17890,N_14116,N_13264);
and U17891 (N_17891,N_14068,N_13226);
nand U17892 (N_17892,N_13367,N_12593);
and U17893 (N_17893,N_12696,N_14328);
and U17894 (N_17894,N_13425,N_13174);
nor U17895 (N_17895,N_12563,N_13873);
xnor U17896 (N_17896,N_12558,N_12064);
and U17897 (N_17897,N_13761,N_14937);
and U17898 (N_17898,N_14166,N_13643);
xor U17899 (N_17899,N_14763,N_13085);
nor U17900 (N_17900,N_13742,N_12521);
nand U17901 (N_17901,N_13351,N_14998);
or U17902 (N_17902,N_12063,N_12453);
nor U17903 (N_17903,N_12588,N_13407);
or U17904 (N_17904,N_12762,N_13245);
xnor U17905 (N_17905,N_12125,N_12298);
or U17906 (N_17906,N_14796,N_13833);
or U17907 (N_17907,N_13984,N_13127);
nand U17908 (N_17908,N_14626,N_14984);
or U17909 (N_17909,N_12611,N_12130);
nand U17910 (N_17910,N_13035,N_14006);
and U17911 (N_17911,N_12928,N_13148);
or U17912 (N_17912,N_12153,N_12387);
or U17913 (N_17913,N_12286,N_13375);
nand U17914 (N_17914,N_14414,N_14036);
nor U17915 (N_17915,N_14670,N_12964);
and U17916 (N_17916,N_12384,N_12845);
nand U17917 (N_17917,N_12244,N_12192);
or U17918 (N_17918,N_13040,N_12395);
and U17919 (N_17919,N_13520,N_13110);
nor U17920 (N_17920,N_14168,N_13478);
xor U17921 (N_17921,N_13804,N_14172);
and U17922 (N_17922,N_12847,N_13680);
xnor U17923 (N_17923,N_14663,N_14521);
nor U17924 (N_17924,N_13955,N_13468);
nand U17925 (N_17925,N_14395,N_14141);
nor U17926 (N_17926,N_13427,N_12896);
and U17927 (N_17927,N_14255,N_12704);
nor U17928 (N_17928,N_12550,N_14496);
xor U17929 (N_17929,N_14381,N_14134);
or U17930 (N_17930,N_13584,N_14782);
xnor U17931 (N_17931,N_13606,N_12811);
nand U17932 (N_17932,N_12277,N_12907);
nand U17933 (N_17933,N_13686,N_12253);
nor U17934 (N_17934,N_12650,N_12726);
nand U17935 (N_17935,N_12775,N_14695);
and U17936 (N_17936,N_13293,N_14408);
nor U17937 (N_17937,N_13614,N_13230);
nand U17938 (N_17938,N_13538,N_14017);
nor U17939 (N_17939,N_13634,N_12444);
nand U17940 (N_17940,N_12414,N_14370);
nand U17941 (N_17941,N_12374,N_13274);
xor U17942 (N_17942,N_13231,N_14102);
nor U17943 (N_17943,N_12909,N_14066);
nor U17944 (N_17944,N_14291,N_13317);
or U17945 (N_17945,N_13981,N_13194);
nand U17946 (N_17946,N_13125,N_13992);
xnor U17947 (N_17947,N_13347,N_13293);
nand U17948 (N_17948,N_12769,N_14558);
nor U17949 (N_17949,N_12107,N_12878);
nor U17950 (N_17950,N_12840,N_13307);
or U17951 (N_17951,N_13516,N_14720);
and U17952 (N_17952,N_12117,N_13694);
xor U17953 (N_17953,N_13344,N_14505);
xnor U17954 (N_17954,N_12741,N_13761);
nor U17955 (N_17955,N_13420,N_14859);
xor U17956 (N_17956,N_13928,N_12408);
nand U17957 (N_17957,N_14133,N_13968);
xnor U17958 (N_17958,N_12370,N_13621);
nor U17959 (N_17959,N_13221,N_13279);
nor U17960 (N_17960,N_13705,N_14704);
nand U17961 (N_17961,N_13900,N_14135);
nand U17962 (N_17962,N_12341,N_13410);
nand U17963 (N_17963,N_14346,N_13399);
xnor U17964 (N_17964,N_13404,N_12801);
nor U17965 (N_17965,N_13123,N_12014);
or U17966 (N_17966,N_14809,N_14415);
nor U17967 (N_17967,N_13510,N_14319);
nand U17968 (N_17968,N_12162,N_12600);
or U17969 (N_17969,N_12533,N_13849);
and U17970 (N_17970,N_14673,N_12407);
or U17971 (N_17971,N_14666,N_13176);
xor U17972 (N_17972,N_14339,N_12164);
or U17973 (N_17973,N_13120,N_12585);
and U17974 (N_17974,N_14616,N_12344);
xnor U17975 (N_17975,N_12845,N_12967);
nand U17976 (N_17976,N_14917,N_12425);
or U17977 (N_17977,N_12787,N_14012);
xor U17978 (N_17978,N_12678,N_13792);
nand U17979 (N_17979,N_12499,N_14042);
and U17980 (N_17980,N_14504,N_13327);
xor U17981 (N_17981,N_12589,N_12111);
xnor U17982 (N_17982,N_12746,N_12105);
or U17983 (N_17983,N_14465,N_14939);
and U17984 (N_17984,N_13157,N_13785);
and U17985 (N_17985,N_14141,N_12585);
nor U17986 (N_17986,N_13235,N_13908);
nand U17987 (N_17987,N_12044,N_12796);
nand U17988 (N_17988,N_14796,N_14276);
nor U17989 (N_17989,N_13918,N_13444);
and U17990 (N_17990,N_13308,N_14470);
nor U17991 (N_17991,N_13816,N_14536);
and U17992 (N_17992,N_12455,N_12733);
nand U17993 (N_17993,N_14898,N_12986);
nor U17994 (N_17994,N_12570,N_13263);
or U17995 (N_17995,N_14727,N_13127);
or U17996 (N_17996,N_12971,N_13044);
nand U17997 (N_17997,N_12068,N_13737);
and U17998 (N_17998,N_14074,N_13626);
or U17999 (N_17999,N_12033,N_12599);
xor U18000 (N_18000,N_16356,N_16838);
and U18001 (N_18001,N_15090,N_16725);
and U18002 (N_18002,N_15013,N_16919);
or U18003 (N_18003,N_15132,N_15184);
xnor U18004 (N_18004,N_15243,N_15197);
xnor U18005 (N_18005,N_15215,N_16002);
nand U18006 (N_18006,N_15112,N_17960);
and U18007 (N_18007,N_17985,N_17795);
or U18008 (N_18008,N_16449,N_15155);
nand U18009 (N_18009,N_15600,N_16055);
xor U18010 (N_18010,N_15791,N_17360);
nand U18011 (N_18011,N_17606,N_15628);
or U18012 (N_18012,N_17406,N_16817);
or U18013 (N_18013,N_17095,N_17261);
nand U18014 (N_18014,N_17479,N_16293);
or U18015 (N_18015,N_15104,N_17299);
nor U18016 (N_18016,N_16447,N_15658);
or U18017 (N_18017,N_16237,N_15669);
and U18018 (N_18018,N_15303,N_15762);
xnor U18019 (N_18019,N_15252,N_16963);
or U18020 (N_18020,N_16831,N_15569);
nor U18021 (N_18021,N_15420,N_15729);
and U18022 (N_18022,N_16450,N_17212);
and U18023 (N_18023,N_16133,N_16668);
nor U18024 (N_18024,N_17419,N_16728);
xnor U18025 (N_18025,N_15676,N_16713);
or U18026 (N_18026,N_15083,N_15626);
nor U18027 (N_18027,N_16021,N_16349);
nand U18028 (N_18028,N_15036,N_17461);
nor U18029 (N_18029,N_17339,N_15589);
and U18030 (N_18030,N_17823,N_16538);
nor U18031 (N_18031,N_16882,N_16484);
nand U18032 (N_18032,N_16360,N_16542);
and U18033 (N_18033,N_16398,N_16408);
xor U18034 (N_18034,N_17966,N_16918);
nand U18035 (N_18035,N_16631,N_15525);
and U18036 (N_18036,N_17306,N_17735);
and U18037 (N_18037,N_15091,N_15292);
xor U18038 (N_18038,N_16690,N_17983);
xor U18039 (N_18039,N_16067,N_15161);
xor U18040 (N_18040,N_16229,N_16269);
or U18041 (N_18041,N_15088,N_16783);
nand U18042 (N_18042,N_16122,N_15208);
xor U18043 (N_18043,N_15516,N_17748);
nand U18044 (N_18044,N_17399,N_17445);
and U18045 (N_18045,N_17117,N_17340);
and U18046 (N_18046,N_16079,N_15368);
xnor U18047 (N_18047,N_17045,N_17351);
and U18048 (N_18048,N_15202,N_15898);
or U18049 (N_18049,N_15214,N_16096);
or U18050 (N_18050,N_15545,N_17012);
xnor U18051 (N_18051,N_16962,N_15320);
nor U18052 (N_18052,N_15367,N_15205);
and U18053 (N_18053,N_15951,N_16483);
and U18054 (N_18054,N_17425,N_17503);
nor U18055 (N_18055,N_15805,N_17542);
nor U18056 (N_18056,N_15552,N_15983);
xor U18057 (N_18057,N_15334,N_17763);
nand U18058 (N_18058,N_16344,N_15757);
nand U18059 (N_18059,N_15493,N_16321);
xnor U18060 (N_18060,N_17081,N_17053);
xnor U18061 (N_18061,N_15255,N_17154);
or U18062 (N_18062,N_15051,N_17186);
xnor U18063 (N_18063,N_17847,N_15821);
or U18064 (N_18064,N_15187,N_15321);
xor U18065 (N_18065,N_15152,N_17885);
and U18066 (N_18066,N_15802,N_15747);
nor U18067 (N_18067,N_16111,N_15964);
and U18068 (N_18068,N_17662,N_15692);
or U18069 (N_18069,N_15424,N_16390);
xor U18070 (N_18070,N_15748,N_15625);
and U18071 (N_18071,N_17125,N_15509);
or U18072 (N_18072,N_15022,N_17901);
nor U18073 (N_18073,N_17502,N_15918);
nor U18074 (N_18074,N_16240,N_16495);
and U18075 (N_18075,N_16524,N_17938);
nor U18076 (N_18076,N_16766,N_16709);
and U18077 (N_18077,N_16743,N_17519);
nand U18078 (N_18078,N_16706,N_17264);
nand U18079 (N_18079,N_15151,N_16197);
nor U18080 (N_18080,N_17812,N_15884);
nand U18081 (N_18081,N_16585,N_17380);
and U18082 (N_18082,N_17840,N_15854);
xnor U18083 (N_18083,N_15572,N_16411);
nand U18084 (N_18084,N_16035,N_16640);
and U18085 (N_18085,N_17621,N_16412);
and U18086 (N_18086,N_17065,N_16930);
and U18087 (N_18087,N_17976,N_16172);
nor U18088 (N_18088,N_15019,N_16537);
xnor U18089 (N_18089,N_15488,N_15494);
nand U18090 (N_18090,N_15858,N_16849);
and U18091 (N_18091,N_16970,N_15687);
xnor U18092 (N_18092,N_16314,N_15661);
and U18093 (N_18093,N_17565,N_17547);
nor U18094 (N_18094,N_15558,N_17742);
and U18095 (N_18095,N_16512,N_15062);
nor U18096 (N_18096,N_17288,N_15198);
xor U18097 (N_18097,N_16072,N_17237);
nor U18098 (N_18098,N_15594,N_15142);
or U18099 (N_18099,N_17193,N_16442);
nand U18100 (N_18100,N_17324,N_15105);
and U18101 (N_18101,N_16206,N_15551);
and U18102 (N_18102,N_17040,N_16660);
or U18103 (N_18103,N_17513,N_17307);
and U18104 (N_18104,N_16150,N_16881);
nand U18105 (N_18105,N_17485,N_15627);
xor U18106 (N_18106,N_16801,N_16937);
and U18107 (N_18107,N_16897,N_17522);
nand U18108 (N_18108,N_16749,N_15557);
nor U18109 (N_18109,N_17342,N_16541);
or U18110 (N_18110,N_15351,N_16163);
nand U18111 (N_18111,N_16145,N_17162);
and U18112 (N_18112,N_15060,N_15440);
and U18113 (N_18113,N_15392,N_16103);
nor U18114 (N_18114,N_17977,N_17179);
and U18115 (N_18115,N_17329,N_16517);
nand U18116 (N_18116,N_15568,N_16959);
and U18117 (N_18117,N_17284,N_16260);
nand U18118 (N_18118,N_17036,N_17225);
nand U18119 (N_18119,N_17495,N_16380);
xor U18120 (N_18120,N_15719,N_17376);
nor U18121 (N_18121,N_16800,N_16754);
xnor U18122 (N_18122,N_16065,N_15879);
xor U18123 (N_18123,N_17838,N_16518);
and U18124 (N_18124,N_17855,N_16996);
and U18125 (N_18125,N_16702,N_17775);
nand U18126 (N_18126,N_17308,N_15196);
nand U18127 (N_18127,N_17844,N_15499);
nand U18128 (N_18128,N_15000,N_17630);
and U18129 (N_18129,N_15796,N_15310);
xor U18130 (N_18130,N_16926,N_15792);
xor U18131 (N_18131,N_15758,N_17296);
or U18132 (N_18132,N_17119,N_17070);
xor U18133 (N_18133,N_15576,N_17285);
nor U18134 (N_18134,N_15337,N_17878);
and U18135 (N_18135,N_15737,N_16992);
nand U18136 (N_18136,N_15213,N_15386);
xor U18137 (N_18137,N_16890,N_16679);
nor U18138 (N_18138,N_16530,N_15766);
or U18139 (N_18139,N_15853,N_16355);
xnor U18140 (N_18140,N_15738,N_15479);
and U18141 (N_18141,N_16940,N_15540);
and U18142 (N_18142,N_15904,N_16833);
nor U18143 (N_18143,N_16845,N_15253);
nor U18144 (N_18144,N_17021,N_17286);
nor U18145 (N_18145,N_15366,N_16603);
xnor U18146 (N_18146,N_16502,N_16346);
and U18147 (N_18147,N_15598,N_16835);
xnor U18148 (N_18148,N_17774,N_16182);
nand U18149 (N_18149,N_17037,N_16755);
xor U18150 (N_18150,N_17933,N_17917);
nor U18151 (N_18151,N_17431,N_17968);
nand U18152 (N_18152,N_17895,N_15108);
or U18153 (N_18153,N_16257,N_17403);
or U18154 (N_18154,N_17149,N_17879);
nand U18155 (N_18155,N_17508,N_16282);
nor U18156 (N_18156,N_16492,N_16654);
nand U18157 (N_18157,N_17592,N_15129);
nand U18158 (N_18158,N_16858,N_17739);
and U18159 (N_18159,N_17854,N_16906);
nand U18160 (N_18160,N_17539,N_15260);
and U18161 (N_18161,N_15886,N_17616);
nand U18162 (N_18162,N_15293,N_17669);
nor U18163 (N_18163,N_15346,N_17247);
nor U18164 (N_18164,N_17738,N_15369);
nor U18165 (N_18165,N_17255,N_16493);
xnor U18166 (N_18166,N_16094,N_16477);
xor U18167 (N_18167,N_17642,N_17991);
nand U18168 (N_18168,N_17241,N_16764);
or U18169 (N_18169,N_17319,N_15244);
or U18170 (N_18170,N_16956,N_15047);
nor U18171 (N_18171,N_16802,N_17348);
nand U18172 (N_18172,N_17220,N_17373);
nor U18173 (N_18173,N_15457,N_17083);
nor U18174 (N_18174,N_16826,N_15709);
nor U18175 (N_18175,N_17428,N_16922);
nand U18176 (N_18176,N_16460,N_15903);
or U18177 (N_18177,N_16899,N_17259);
and U18178 (N_18178,N_16457,N_16954);
or U18179 (N_18179,N_15847,N_17874);
xnor U18180 (N_18180,N_16830,N_16030);
or U18181 (N_18181,N_15164,N_16436);
xnor U18182 (N_18182,N_15041,N_16888);
and U18183 (N_18183,N_17104,N_17378);
nor U18184 (N_18184,N_16769,N_17741);
and U18185 (N_18185,N_17345,N_15373);
and U18186 (N_18186,N_15772,N_16203);
nor U18187 (N_18187,N_17275,N_17355);
nor U18188 (N_18188,N_16433,N_17369);
xor U18189 (N_18189,N_16128,N_15145);
nand U18190 (N_18190,N_15482,N_16470);
nor U18191 (N_18191,N_15442,N_16225);
nand U18192 (N_18192,N_17391,N_17454);
nand U18193 (N_18193,N_17200,N_16009);
nand U18194 (N_18194,N_16080,N_17128);
xor U18195 (N_18195,N_17004,N_16671);
and U18196 (N_18196,N_16400,N_17506);
nor U18197 (N_18197,N_16622,N_16135);
nand U18198 (N_18198,N_16676,N_15431);
or U18199 (N_18199,N_16183,N_15714);
and U18200 (N_18200,N_16733,N_15695);
nor U18201 (N_18201,N_17435,N_15110);
nor U18202 (N_18202,N_16594,N_15465);
or U18203 (N_18203,N_17514,N_17447);
nor U18204 (N_18204,N_16735,N_15793);
xor U18205 (N_18205,N_15941,N_17709);
nand U18206 (N_18206,N_17211,N_17463);
nand U18207 (N_18207,N_16313,N_17886);
nor U18208 (N_18208,N_16939,N_15359);
and U18209 (N_18209,N_17999,N_15732);
and U18210 (N_18210,N_15943,N_15524);
nor U18211 (N_18211,N_15584,N_17471);
and U18212 (N_18212,N_16961,N_17682);
or U18213 (N_18213,N_16138,N_17395);
or U18214 (N_18214,N_16144,N_17733);
xor U18215 (N_18215,N_16291,N_16815);
xor U18216 (N_18216,N_16259,N_15741);
or U18217 (N_18217,N_15451,N_15410);
xor U18218 (N_18218,N_15072,N_15938);
xor U18219 (N_18219,N_17880,N_17684);
or U18220 (N_18220,N_15402,N_16965);
or U18221 (N_18221,N_16839,N_17453);
xor U18222 (N_18222,N_15483,N_16990);
xnor U18223 (N_18223,N_15667,N_15262);
or U18224 (N_18224,N_17687,N_15287);
nand U18225 (N_18225,N_15588,N_16738);
or U18226 (N_18226,N_17014,N_17531);
nand U18227 (N_18227,N_17473,N_17597);
nand U18228 (N_18228,N_16562,N_16246);
xnor U18229 (N_18229,N_17618,N_15819);
xnor U18230 (N_18230,N_16781,N_15394);
xnor U18231 (N_18231,N_17677,N_15968);
or U18232 (N_18232,N_17404,N_16152);
nor U18233 (N_18233,N_15464,N_17054);
nor U18234 (N_18234,N_17668,N_15102);
or U18235 (N_18235,N_15562,N_17664);
xor U18236 (N_18236,N_16915,N_15115);
nor U18237 (N_18237,N_17566,N_17955);
or U18238 (N_18238,N_15840,N_17928);
or U18239 (N_18239,N_16157,N_17906);
or U18240 (N_18240,N_17957,N_16422);
nor U18241 (N_18241,N_15691,N_15206);
nand U18242 (N_18242,N_17759,N_17333);
nand U18243 (N_18243,N_16185,N_17517);
nor U18244 (N_18244,N_16564,N_15979);
xnor U18245 (N_18245,N_17254,N_16308);
nand U18246 (N_18246,N_15486,N_17323);
nand U18247 (N_18247,N_16461,N_15326);
xnor U18248 (N_18248,N_17632,N_15079);
or U18249 (N_18249,N_17312,N_16290);
xnor U18250 (N_18250,N_15607,N_16636);
or U18251 (N_18251,N_15146,N_17167);
nor U18252 (N_18252,N_16155,N_16479);
nor U18253 (N_18253,N_16184,N_17033);
or U18254 (N_18254,N_16490,N_15005);
nor U18255 (N_18255,N_17135,N_15702);
and U18256 (N_18256,N_17090,N_16768);
nand U18257 (N_18257,N_16993,N_17940);
or U18258 (N_18258,N_17359,N_17530);
xor U18259 (N_18259,N_15783,N_16375);
nor U18260 (N_18260,N_15230,N_17836);
or U18261 (N_18261,N_17913,N_16404);
xor U18262 (N_18262,N_15109,N_15400);
and U18263 (N_18263,N_16902,N_15784);
nand U18264 (N_18264,N_15289,N_15852);
nor U18265 (N_18265,N_17967,N_16244);
xor U18266 (N_18266,N_15118,N_15054);
nor U18267 (N_18267,N_17890,N_15043);
and U18268 (N_18268,N_15585,N_17510);
xor U18269 (N_18269,N_15612,N_15596);
or U18270 (N_18270,N_17227,N_15093);
and U18271 (N_18271,N_16011,N_16335);
or U18272 (N_18272,N_15902,N_15298);
or U18273 (N_18273,N_16431,N_15265);
and U18274 (N_18274,N_17035,N_15827);
nor U18275 (N_18275,N_16704,N_15236);
xnor U18276 (N_18276,N_17919,N_16262);
nand U18277 (N_18277,N_17246,N_15615);
and U18278 (N_18278,N_16909,N_16256);
or U18279 (N_18279,N_16731,N_16181);
nor U18280 (N_18280,N_15891,N_15001);
nor U18281 (N_18281,N_17258,N_15419);
and U18282 (N_18282,N_17696,N_17725);
or U18283 (N_18283,N_15209,N_15593);
or U18284 (N_18284,N_17007,N_17971);
xor U18285 (N_18285,N_15948,N_16266);
and U18286 (N_18286,N_17444,N_16586);
and U18287 (N_18287,N_15859,N_16329);
nor U18288 (N_18288,N_15481,N_15824);
nand U18289 (N_18289,N_17068,N_16843);
nand U18290 (N_18290,N_15534,N_16819);
and U18291 (N_18291,N_17010,N_17577);
nand U18292 (N_18292,N_17328,N_16070);
or U18293 (N_18293,N_15458,N_17136);
or U18294 (N_18294,N_17982,N_17166);
or U18295 (N_18295,N_17375,N_16292);
xor U18296 (N_18296,N_15657,N_17484);
xnor U18297 (N_18297,N_15634,N_16545);
and U18298 (N_18298,N_15125,N_15565);
and U18299 (N_18299,N_16787,N_17929);
or U18300 (N_18300,N_16642,N_16752);
nand U18301 (N_18301,N_15158,N_17835);
and U18302 (N_18302,N_16664,N_16678);
nand U18303 (N_18303,N_16651,N_16159);
or U18304 (N_18304,N_17272,N_15620);
or U18305 (N_18305,N_17800,N_15770);
nand U18306 (N_18306,N_16916,N_17325);
and U18307 (N_18307,N_16860,N_15679);
xor U18308 (N_18308,N_17151,N_15867);
or U18309 (N_18309,N_17223,N_15517);
xor U18310 (N_18310,N_15520,N_17724);
nor U18311 (N_18311,N_16462,N_17392);
nand U18312 (N_18312,N_15760,N_15307);
and U18313 (N_18313,N_17487,N_15388);
and U18314 (N_18314,N_16062,N_17785);
or U18315 (N_18315,N_15188,N_15135);
or U18316 (N_18316,N_17843,N_17633);
or U18317 (N_18317,N_15496,N_17310);
nand U18318 (N_18318,N_17683,N_17363);
and U18319 (N_18319,N_17361,N_16473);
xnor U18320 (N_18320,N_16068,N_17238);
xor U18321 (N_18321,N_16635,N_16033);
nor U18322 (N_18322,N_16058,N_16363);
xor U18323 (N_18323,N_17611,N_17573);
or U18324 (N_18324,N_15773,N_16267);
nor U18325 (N_18325,N_16855,N_17610);
nand U18326 (N_18326,N_16804,N_16165);
xor U18327 (N_18327,N_16550,N_17707);
xnor U18328 (N_18328,N_17975,N_17504);
nor U18329 (N_18329,N_16123,N_15582);
or U18330 (N_18330,N_16864,N_16101);
nand U18331 (N_18331,N_17019,N_17704);
xnor U18332 (N_18332,N_16786,N_16368);
xnor U18333 (N_18333,N_15272,N_16513);
or U18334 (N_18334,N_16113,N_16480);
and U18335 (N_18335,N_17280,N_16814);
xor U18336 (N_18336,N_15381,N_16988);
or U18337 (N_18337,N_16057,N_15817);
and U18338 (N_18338,N_16606,N_16298);
nor U18339 (N_18339,N_17870,N_17335);
nor U18340 (N_18340,N_17424,N_15357);
nand U18341 (N_18341,N_17047,N_17016);
and U18342 (N_18342,N_15429,N_16720);
nand U18343 (N_18343,N_15924,N_15319);
nand U18344 (N_18344,N_17121,N_17477);
nor U18345 (N_18345,N_17115,N_15996);
or U18346 (N_18346,N_17069,N_17464);
nand U18347 (N_18347,N_17056,N_17978);
nor U18348 (N_18348,N_15833,N_15536);
and U18349 (N_18349,N_16191,N_15573);
nor U18350 (N_18350,N_17766,N_15895);
and U18351 (N_18351,N_17239,N_15192);
or U18352 (N_18352,N_17302,N_15099);
nor U18353 (N_18353,N_17617,N_15871);
nand U18354 (N_18354,N_16928,N_17469);
or U18355 (N_18355,N_17139,N_15985);
nand U18356 (N_18356,N_15328,N_15191);
nor U18357 (N_18357,N_15156,N_15096);
or U18358 (N_18358,N_16509,N_15531);
nand U18359 (N_18359,N_15003,N_16539);
nand U18360 (N_18360,N_17123,N_17020);
xnor U18361 (N_18361,N_17198,N_16692);
xnor U18362 (N_18362,N_15502,N_17370);
and U18363 (N_18363,N_15354,N_15492);
xor U18364 (N_18364,N_17270,N_15722);
and U18365 (N_18365,N_15171,N_17234);
and U18366 (N_18366,N_17298,N_17429);
xnor U18367 (N_18367,N_15984,N_15268);
and U18368 (N_18368,N_16440,N_17075);
and U18369 (N_18369,N_15689,N_17882);
xor U18370 (N_18370,N_15131,N_16367);
or U18371 (N_18371,N_15278,N_17426);
xnor U18372 (N_18372,N_15782,N_17575);
xor U18373 (N_18373,N_15530,N_16972);
or U18374 (N_18374,N_17729,N_16551);
nand U18375 (N_18375,N_15374,N_16142);
nor U18376 (N_18376,N_15383,N_16997);
or U18377 (N_18377,N_16131,N_15314);
nor U18378 (N_18378,N_15219,N_16892);
or U18379 (N_18379,N_16580,N_16914);
and U18380 (N_18380,N_17923,N_16571);
nor U18381 (N_18381,N_15332,N_15274);
and U18382 (N_18382,N_15474,N_16018);
nand U18383 (N_18383,N_16452,N_15637);
nor U18384 (N_18384,N_17764,N_15324);
nand U18385 (N_18385,N_17685,N_17099);
nand U18386 (N_18386,N_16644,N_15663);
nor U18387 (N_18387,N_15797,N_17561);
nor U18388 (N_18388,N_15207,N_15365);
xor U18389 (N_18389,N_15010,N_16873);
nor U18390 (N_18390,N_17672,N_16283);
nor U18391 (N_18391,N_16666,N_16199);
and U18392 (N_18392,N_17556,N_16932);
nor U18393 (N_18393,N_17060,N_16040);
nor U18394 (N_18394,N_16141,N_17679);
nand U18395 (N_18395,N_16143,N_16385);
nor U18396 (N_18396,N_15727,N_17024);
or U18397 (N_18397,N_16805,N_15845);
or U18398 (N_18398,N_17316,N_17912);
or U18399 (N_18399,N_16074,N_15395);
nor U18400 (N_18400,N_15119,N_17641);
or U18401 (N_18401,N_17107,N_15799);
xnor U18402 (N_18402,N_16985,N_15945);
or U18403 (N_18403,N_15249,N_17645);
and U18404 (N_18404,N_16276,N_16024);
nand U18405 (N_18405,N_17173,N_15635);
nand U18406 (N_18406,N_17914,N_17073);
nand U18407 (N_18407,N_17598,N_17674);
nor U18408 (N_18408,N_16556,N_16354);
nand U18409 (N_18409,N_17232,N_17420);
or U18410 (N_18410,N_17266,N_17224);
nor U18411 (N_18411,N_16087,N_17727);
nand U18412 (N_18412,N_16763,N_15940);
and U18413 (N_18413,N_15767,N_16482);
and U18414 (N_18414,N_17860,N_16649);
nor U18415 (N_18415,N_16837,N_17777);
or U18416 (N_18416,N_17989,N_17528);
xnor U18417 (N_18417,N_17915,N_15232);
and U18418 (N_18418,N_17086,N_15982);
or U18419 (N_18419,N_16039,N_17660);
or U18420 (N_18420,N_17172,N_15034);
and U18421 (N_18421,N_17900,N_17658);
nand U18422 (N_18422,N_17767,N_16441);
nor U18423 (N_18423,N_16633,N_15123);
xor U18424 (N_18424,N_15407,N_17209);
xnor U18425 (N_18425,N_17374,N_16775);
and U18426 (N_18426,N_17364,N_16345);
and U18427 (N_18427,N_17711,N_17160);
nand U18428 (N_18428,N_17170,N_15350);
xor U18429 (N_18429,N_17935,N_16674);
or U18430 (N_18430,N_15873,N_15807);
xor U18431 (N_18431,N_15175,N_15027);
or U18432 (N_18432,N_15498,N_17137);
nor U18433 (N_18433,N_15467,N_15622);
nor U18434 (N_18434,N_16535,N_17898);
nand U18435 (N_18435,N_17267,N_16081);
and U18436 (N_18436,N_15353,N_17809);
and U18437 (N_18437,N_17398,N_15340);
or U18438 (N_18438,N_16170,N_16341);
or U18439 (N_18439,N_15245,N_15301);
or U18440 (N_18440,N_16444,N_15070);
and U18441 (N_18441,N_17690,N_17026);
nand U18442 (N_18442,N_16469,N_15275);
and U18443 (N_18443,N_15148,N_17410);
and U18444 (N_18444,N_16907,N_16230);
nor U18445 (N_18445,N_16813,N_16139);
nor U18446 (N_18446,N_15015,N_15756);
nor U18447 (N_18447,N_16696,N_17770);
nand U18448 (N_18448,N_17371,N_17092);
xnor U18449 (N_18449,N_15358,N_15623);
xor U18450 (N_18450,N_17581,N_17548);
or U18451 (N_18451,N_15566,N_16872);
or U18452 (N_18452,N_17124,N_16722);
nor U18453 (N_18453,N_17436,N_15503);
or U18454 (N_18454,N_15283,N_16397);
xnor U18455 (N_18455,N_15823,N_15443);
xor U18456 (N_18456,N_16741,N_15216);
and U18457 (N_18457,N_15874,N_15809);
nand U18458 (N_18458,N_15094,N_17875);
and U18459 (N_18459,N_15378,N_17482);
or U18460 (N_18460,N_16883,N_15708);
or U18461 (N_18461,N_16379,N_17175);
or U18462 (N_18462,N_16515,N_16526);
nand U18463 (N_18463,N_17931,N_17206);
xor U18464 (N_18464,N_16547,N_17958);
or U18465 (N_18465,N_17257,N_15844);
nand U18466 (N_18466,N_16004,N_17365);
or U18467 (N_18467,N_16521,N_16784);
xor U18468 (N_18468,N_16593,N_16395);
xor U18469 (N_18469,N_16685,N_16019);
and U18470 (N_18470,N_15361,N_17634);
nor U18471 (N_18471,N_17277,N_17341);
nand U18472 (N_18472,N_15250,N_15452);
and U18473 (N_18473,N_16546,N_17501);
and U18474 (N_18474,N_16245,N_15820);
and U18475 (N_18475,N_15480,N_16052);
and U18476 (N_18476,N_17497,N_17962);
nand U18477 (N_18477,N_16894,N_17817);
or U18478 (N_18478,N_17796,N_15510);
xor U18479 (N_18479,N_15703,N_16732);
and U18480 (N_18480,N_17511,N_15512);
xnor U18481 (N_18481,N_15097,N_15396);
nand U18482 (N_18482,N_15955,N_17350);
xor U18483 (N_18483,N_16661,N_15935);
nor U18484 (N_18484,N_15662,N_17920);
or U18485 (N_18485,N_17570,N_16264);
and U18486 (N_18486,N_16770,N_15270);
and U18487 (N_18487,N_15578,N_16730);
nor U18488 (N_18488,N_17944,N_17467);
nand U18489 (N_18489,N_15273,N_17820);
or U18490 (N_18490,N_17222,N_17169);
and U18491 (N_18491,N_15078,N_15678);
xor U18492 (N_18492,N_16866,N_16099);
nor U18493 (N_18493,N_17338,N_16984);
nand U18494 (N_18494,N_16616,N_15271);
and U18495 (N_18495,N_17784,N_17719);
nor U18496 (N_18496,N_16977,N_16966);
and U18497 (N_18497,N_17829,N_15960);
xnor U18498 (N_18498,N_15024,N_17861);
nor U18499 (N_18499,N_17387,N_16445);
nand U18500 (N_18500,N_15730,N_17405);
nor U18501 (N_18501,N_15040,N_16465);
or U18502 (N_18502,N_16132,N_17680);
or U18503 (N_18503,N_17188,N_17732);
and U18504 (N_18504,N_15694,N_16862);
nor U18505 (N_18505,N_16119,N_16707);
nand U18506 (N_18506,N_16413,N_16658);
xor U18507 (N_18507,N_15261,N_16796);
or U18508 (N_18508,N_16167,N_17049);
xnor U18509 (N_18509,N_16595,N_17907);
and U18510 (N_18510,N_17052,N_17715);
and U18511 (N_18511,N_15632,N_16893);
and U18512 (N_18512,N_16126,N_16265);
nand U18513 (N_18513,N_15280,N_17295);
and U18514 (N_18514,N_17720,N_15575);
and U18515 (N_18515,N_17953,N_16406);
and U18516 (N_18516,N_17031,N_15413);
and U18517 (N_18517,N_17718,N_15659);
nor U18518 (N_18518,N_15026,N_15789);
nor U18519 (N_18519,N_15543,N_16034);
or U18520 (N_18520,N_15939,N_16127);
and U18521 (N_18521,N_15954,N_17659);
xnor U18522 (N_18522,N_15059,N_17631);
nand U18523 (N_18523,N_17480,N_15300);
xor U18524 (N_18524,N_17076,N_17509);
nor U18525 (N_18525,N_15609,N_15291);
nand U18526 (N_18526,N_16389,N_17113);
nor U18527 (N_18527,N_16374,N_16703);
and U18528 (N_18528,N_16038,N_16980);
nand U18529 (N_18529,N_16721,N_15862);
and U18530 (N_18530,N_17273,N_17526);
nor U18531 (N_18531,N_17448,N_16130);
nor U18532 (N_18532,N_16532,N_15647);
xor U18533 (N_18533,N_17697,N_15136);
or U18534 (N_18534,N_16841,N_17969);
nor U18535 (N_18535,N_15580,N_17806);
or U18536 (N_18536,N_17622,N_16896);
xor U18537 (N_18537,N_15344,N_15134);
or U18538 (N_18538,N_17465,N_16964);
or U18539 (N_18539,N_16318,N_15591);
nor U18540 (N_18540,N_17862,N_15656);
nand U18541 (N_18541,N_16792,N_16592);
nand U18542 (N_18542,N_15315,N_15610);
or U18543 (N_18543,N_17476,N_16558);
xor U18544 (N_18544,N_16579,N_17155);
nor U18545 (N_18545,N_17552,N_17926);
xnor U18546 (N_18546,N_17551,N_16249);
xor U18547 (N_18547,N_17580,N_15032);
nor U18548 (N_18548,N_16423,N_17109);
or U18549 (N_18549,N_17423,N_16186);
or U18550 (N_18550,N_16584,N_16332);
and U18551 (N_18551,N_15563,N_16723);
or U18552 (N_18552,N_17187,N_15693);
or U18553 (N_18553,N_17712,N_15929);
nor U18554 (N_18554,N_17446,N_16421);
and U18555 (N_18555,N_16958,N_15619);
or U18556 (N_18556,N_16942,N_16285);
nor U18557 (N_18557,N_17022,N_17873);
xnor U18558 (N_18558,N_17451,N_15856);
or U18559 (N_18559,N_15470,N_17562);
and U18560 (N_18560,N_15974,N_17646);
and U18561 (N_18561,N_15006,N_15190);
and U18562 (N_18562,N_16861,N_16953);
nor U18563 (N_18563,N_16875,N_15199);
and U18564 (N_18564,N_17693,N_16471);
nor U18565 (N_18565,N_15035,N_16322);
xnor U18566 (N_18566,N_17152,N_17533);
nor U18567 (N_18567,N_17226,N_16639);
xor U18568 (N_18568,N_17305,N_16740);
nor U18569 (N_18569,N_16601,N_17427);
nand U18570 (N_18570,N_15815,N_15869);
xor U18571 (N_18571,N_17623,N_15876);
nor U18572 (N_18572,N_15379,N_17214);
nor U18573 (N_18573,N_16540,N_17974);
nor U18574 (N_18574,N_17643,N_17221);
xnor U18575 (N_18575,N_17251,N_16270);
xnor U18576 (N_18576,N_17582,N_15744);
nor U18577 (N_18577,N_17195,N_17993);
nor U18578 (N_18578,N_16427,N_17368);
and U18579 (N_18579,N_15352,N_15877);
nand U18580 (N_18580,N_15114,N_17269);
or U18581 (N_18581,N_16851,N_15890);
nor U18582 (N_18582,N_15527,N_15544);
and U18583 (N_18583,N_16543,N_15086);
nor U18584 (N_18584,N_15362,N_17337);
and U18585 (N_18585,N_17527,N_17082);
nand U18586 (N_18586,N_15495,N_17700);
nand U18587 (N_18587,N_15174,N_17180);
nand U18588 (N_18588,N_15677,N_16047);
and U18589 (N_18589,N_15547,N_17625);
or U18590 (N_18590,N_17415,N_15910);
xor U18591 (N_18591,N_16384,N_15745);
or U18592 (N_18592,N_15841,N_15140);
or U18593 (N_18593,N_17105,N_16794);
and U18594 (N_18594,N_17028,N_17013);
xnor U18595 (N_18595,N_16105,N_16823);
nand U18596 (N_18596,N_17791,N_15848);
nand U18597 (N_18597,N_15554,N_17867);
nor U18598 (N_18598,N_17930,N_17372);
nand U18599 (N_18599,N_16284,N_15515);
nor U18600 (N_18600,N_15801,N_17722);
nor U18601 (N_18601,N_15417,N_17908);
nand U18602 (N_18602,N_15029,N_17743);
and U18603 (N_18603,N_17789,N_17412);
and U18604 (N_18604,N_17230,N_16549);
and U18605 (N_18605,N_16924,N_17400);
or U18606 (N_18606,N_17753,N_15325);
nor U18607 (N_18607,N_17591,N_17433);
xor U18608 (N_18608,N_15690,N_15896);
and U18609 (N_18609,N_16487,N_15126);
nor U18610 (N_18610,N_15098,N_17803);
or U18611 (N_18611,N_17987,N_15716);
or U18612 (N_18612,N_15816,N_17343);
and U18613 (N_18613,N_17046,N_15713);
nor U18614 (N_18614,N_15698,N_17571);
xor U18615 (N_18615,N_16686,N_17554);
nand U18616 (N_18616,N_17945,N_16273);
xnor U18617 (N_18617,N_17747,N_15641);
xor U18618 (N_18618,N_17218,N_16913);
or U18619 (N_18619,N_16054,N_17922);
nand U18620 (N_18620,N_15808,N_16957);
or U18621 (N_18621,N_17951,N_15749);
nand U18622 (N_18622,N_17924,N_15810);
nand U18623 (N_18623,N_15909,N_15439);
nand U18624 (N_18624,N_15590,N_17321);
and U18625 (N_18625,N_17734,N_16560);
or U18626 (N_18626,N_15514,N_17141);
xnor U18627 (N_18627,N_16010,N_15345);
nand U18628 (N_18628,N_17201,N_17334);
nand U18629 (N_18629,N_16430,N_16627);
nand U18630 (N_18630,N_17274,N_15990);
xnor U18631 (N_18631,N_17072,N_16221);
nor U18632 (N_18632,N_15644,N_15277);
nor U18633 (N_18633,N_15751,N_16737);
or U18634 (N_18634,N_16761,N_15355);
nand U18635 (N_18635,N_17948,N_16497);
nand U18636 (N_18636,N_15836,N_15194);
xnor U18637 (N_18637,N_16618,N_15613);
xor U18638 (N_18638,N_15611,N_15276);
or U18639 (N_18639,N_16415,N_17786);
and U18640 (N_18640,N_16553,N_17637);
or U18641 (N_18641,N_17132,N_15861);
xnor U18642 (N_18642,N_15390,N_15489);
and U18643 (N_18643,N_17244,N_16147);
nand U18644 (N_18644,N_16905,N_17543);
and U18645 (N_18645,N_15932,N_16925);
and U18646 (N_18646,N_17096,N_16655);
xor U18647 (N_18647,N_15057,N_16015);
nand U18648 (N_18648,N_16921,N_17228);
xnor U18649 (N_18649,N_16222,N_15173);
or U18650 (N_18650,N_17604,N_15944);
nand U18651 (N_18651,N_15700,N_17129);
nor U18652 (N_18652,N_16582,N_16555);
or U18653 (N_18653,N_17005,N_16402);
xnor U18654 (N_18654,N_17217,N_15065);
xnor U18655 (N_18655,N_17904,N_15497);
nor U18656 (N_18656,N_16357,N_16056);
or U18657 (N_18657,N_15317,N_15269);
nor U18658 (N_18658,N_17394,N_15212);
xnor U18659 (N_18659,N_15887,N_17194);
xnor U18660 (N_18660,N_15372,N_16771);
nand U18661 (N_18661,N_17236,N_17011);
nor U18662 (N_18662,N_17456,N_17730);
nand U18663 (N_18663,N_15734,N_17171);
xor U18664 (N_18664,N_17490,N_16968);
nand U18665 (N_18665,N_17185,N_15672);
or U18666 (N_18666,N_15012,N_15038);
or U18667 (N_18667,N_15246,N_16351);
nand U18668 (N_18668,N_17950,N_15670);
nand U18669 (N_18669,N_16859,N_15654);
nand U18670 (N_18670,N_16149,N_17790);
nor U18671 (N_18671,N_16148,N_16714);
xor U18672 (N_18672,N_16288,N_17366);
nand U18673 (N_18673,N_17458,N_17174);
or U18674 (N_18674,N_16350,N_16286);
xnor U18675 (N_18675,N_16912,N_17721);
or U18676 (N_18676,N_16971,N_15581);
nand U18677 (N_18677,N_15798,N_17529);
or U18678 (N_18678,N_15406,N_16178);
xnor U18679 (N_18679,N_17276,N_15302);
or U18680 (N_18680,N_16619,N_15864);
and U18681 (N_18681,N_15831,N_15356);
and U18682 (N_18682,N_15966,N_16614);
nand U18683 (N_18683,N_17988,N_15322);
and U18684 (N_18684,N_16568,N_15200);
and U18685 (N_18685,N_15154,N_16213);
or U18686 (N_18686,N_16362,N_15247);
nor U18687 (N_18687,N_17686,N_17771);
or U18688 (N_18688,N_15103,N_16846);
or U18689 (N_18689,N_15925,N_16933);
and U18690 (N_18690,N_15595,N_17354);
or U18691 (N_18691,N_15401,N_17231);
and U18692 (N_18692,N_16917,N_15437);
nor U18693 (N_18693,N_17832,N_16935);
xnor U18694 (N_18694,N_15204,N_17614);
nor U18695 (N_18695,N_16719,N_15418);
nor U18696 (N_18696,N_15124,N_16020);
xor U18697 (N_18697,N_16337,N_15541);
nand U18698 (N_18698,N_17058,N_17661);
nand U18699 (N_18699,N_15056,N_17110);
nor U18700 (N_18700,N_16850,N_16453);
nand U18701 (N_18701,N_17810,N_15518);
and U18702 (N_18702,N_16125,N_15282);
nor U18703 (N_18703,N_16981,N_16842);
and U18704 (N_18704,N_15504,N_16648);
or U18705 (N_18705,N_16196,N_15999);
and U18706 (N_18706,N_17176,N_17970);
xnor U18707 (N_18707,N_16811,N_15736);
and U18708 (N_18708,N_15728,N_15240);
nand U18709 (N_18709,N_15264,N_15435);
nand U18710 (N_18710,N_15750,N_17972);
xnor U18711 (N_18711,N_16347,N_16392);
nand U18712 (N_18712,N_17569,N_17080);
nand U18713 (N_18713,N_15608,N_15139);
or U18714 (N_18714,N_16751,N_16757);
nand U18715 (N_18715,N_17842,N_16478);
or U18716 (N_18716,N_15911,N_16588);
nor U18717 (N_18717,N_17466,N_16112);
nor U18718 (N_18718,N_16428,N_15872);
or U18719 (N_18719,N_17758,N_16424);
or U18720 (N_18720,N_16153,N_15652);
and U18721 (N_18721,N_16190,N_16865);
xnor U18722 (N_18722,N_15153,N_16204);
or U18723 (N_18723,N_15606,N_15347);
and U18724 (N_18724,N_16782,N_17749);
xor U18725 (N_18725,N_16669,N_16945);
nand U18726 (N_18726,N_16974,N_16646);
and U18727 (N_18727,N_15343,N_16877);
xor U18728 (N_18728,N_16116,N_16840);
nand U18729 (N_18729,N_16334,N_16641);
xnor U18730 (N_18730,N_15523,N_15529);
nand U18731 (N_18731,N_15144,N_16863);
nand U18732 (N_18732,N_17142,N_16573);
nor U18733 (N_18733,N_16026,N_16060);
nor U18734 (N_18734,N_16193,N_15229);
nand U18735 (N_18735,N_15731,N_16536);
nand U18736 (N_18736,N_16005,N_15533);
and U18737 (N_18737,N_16369,N_16336);
xor U18738 (N_18738,N_17397,N_15463);
and U18739 (N_18739,N_16607,N_16003);
xor U18740 (N_18740,N_15333,N_16508);
or U18741 (N_18741,N_16693,N_17532);
or U18742 (N_18742,N_16816,N_16565);
nand U18743 (N_18743,N_17250,N_15159);
nand U18744 (N_18744,N_15830,N_17357);
xnor U18745 (N_18745,N_16085,N_16328);
and U18746 (N_18746,N_15128,N_17202);
or U18747 (N_18747,N_17902,N_15387);
nand U18748 (N_18748,N_16699,N_17640);
or U18749 (N_18749,N_15863,N_17794);
nor U18750 (N_18750,N_15288,N_16386);
nand U18751 (N_18751,N_15087,N_16758);
and U18752 (N_18752,N_17655,N_15052);
or U18753 (N_18753,N_17030,N_16438);
and U18754 (N_18754,N_16803,N_17671);
nand U18755 (N_18755,N_16154,N_17936);
nor U18756 (N_18756,N_17245,N_15806);
and U18757 (N_18757,N_17825,N_17439);
or U18758 (N_18758,N_17990,N_17032);
nor U18759 (N_18759,N_15915,N_16012);
and U18760 (N_18760,N_15950,N_15715);
or U18761 (N_18761,N_15583,N_17853);
and U18762 (N_18762,N_15849,N_17265);
nand U18763 (N_18763,N_15927,N_17705);
xor U18764 (N_18764,N_16596,N_15329);
xnor U18765 (N_18765,N_15989,N_15312);
and U18766 (N_18766,N_15226,N_17303);
and U18767 (N_18767,N_15138,N_15009);
and U18768 (N_18768,N_15223,N_17377);
xor U18769 (N_18769,N_17383,N_15765);
and U18770 (N_18770,N_17579,N_15906);
nor U18771 (N_18771,N_16202,N_17601);
nand U18772 (N_18772,N_15621,N_15147);
nand U18773 (N_18773,N_16778,N_15919);
nor U18774 (N_18774,N_16563,N_15028);
or U18775 (N_18775,N_15163,N_16330);
xnor U18776 (N_18776,N_16604,N_15237);
nand U18777 (N_18777,N_16243,N_17834);
nor U18778 (N_18778,N_17253,N_15014);
and U18779 (N_18779,N_16653,N_17402);
nand U18780 (N_18780,N_17535,N_17002);
or U18781 (N_18781,N_16700,N_17038);
xor U18782 (N_18782,N_15447,N_16014);
or U18783 (N_18783,N_15956,N_15776);
or U18784 (N_18784,N_15649,N_17094);
nor U18785 (N_18785,N_15281,N_16694);
and U18786 (N_18786,N_15085,N_16489);
nor U18787 (N_18787,N_16097,N_16634);
xnor U18788 (N_18788,N_16591,N_17893);
and U18789 (N_18789,N_16305,N_16295);
and U18790 (N_18790,N_16682,N_16405);
or U18791 (N_18791,N_16659,N_15221);
nand U18792 (N_18792,N_17263,N_17837);
nand U18793 (N_18793,N_16300,N_17761);
nor U18794 (N_18794,N_16053,N_15888);
and U18795 (N_18795,N_17041,N_15803);
xnor U18796 (N_18796,N_16211,N_15754);
or U18797 (N_18797,N_16514,N_17182);
xor U18798 (N_18798,N_17421,N_17863);
nor U18799 (N_18799,N_17788,N_16115);
xor U18800 (N_18800,N_17793,N_15506);
xnor U18801 (N_18801,N_17883,N_16691);
xor U18802 (N_18802,N_15934,N_15710);
nor U18803 (N_18803,N_17483,N_15428);
or U18804 (N_18804,N_16516,N_15603);
and U18805 (N_18805,N_17093,N_17567);
xnor U18806 (N_18806,N_15976,N_16226);
nor U18807 (N_18807,N_16911,N_16201);
or U18808 (N_18808,N_17889,N_17470);
nor U18809 (N_18809,N_17615,N_17887);
nor U18810 (N_18810,N_17078,N_15377);
and U18811 (N_18811,N_17001,N_16736);
nor U18812 (N_18812,N_15592,N_15681);
nand U18813 (N_18813,N_15432,N_17821);
and U18814 (N_18814,N_16742,N_16006);
nor U18815 (N_18815,N_15995,N_16338);
nand U18816 (N_18816,N_15016,N_16566);
nor U18817 (N_18817,N_16195,N_16976);
xnor U18818 (N_18818,N_16137,N_15037);
nand U18819 (N_18819,N_17491,N_16506);
nor U18820 (N_18820,N_17765,N_16106);
nand U18821 (N_18821,N_17818,N_16806);
or U18822 (N_18822,N_17710,N_15889);
nand U18823 (N_18823,N_15468,N_15217);
nor U18824 (N_18824,N_15546,N_16324);
nor U18825 (N_18825,N_17498,N_17892);
xor U18826 (N_18826,N_15892,N_16889);
or U18827 (N_18827,N_16683,N_16476);
xor U18828 (N_18828,N_16871,N_16795);
nor U18829 (N_18829,N_15137,N_17781);
nor U18830 (N_18830,N_15339,N_16399);
xnor U18831 (N_18831,N_16605,N_17585);
nor U18832 (N_18832,N_15564,N_16342);
nor U18833 (N_18833,N_17362,N_17884);
or U18834 (N_18834,N_16991,N_17390);
nor U18835 (N_18835,N_16501,N_16652);
nand U18836 (N_18836,N_17133,N_16409);
xnor U18837 (N_18837,N_16248,N_17087);
and U18838 (N_18838,N_16510,N_17596);
and U18839 (N_18839,N_15235,N_17851);
and U18840 (N_18840,N_17934,N_16432);
or U18841 (N_18841,N_16748,N_16110);
or U18842 (N_18842,N_17097,N_17204);
nor U18843 (N_18843,N_17586,N_17416);
or U18844 (N_18844,N_17869,N_17624);
and U18845 (N_18845,N_15779,N_15117);
nand U18846 (N_18846,N_15666,N_16886);
or U18847 (N_18847,N_15077,N_15643);
and U18848 (N_18848,N_15476,N_17691);
and U18849 (N_18849,N_15993,N_15179);
xnor U18850 (N_18850,N_17418,N_17744);
nor U18851 (N_18851,N_15684,N_17807);
nor U18852 (N_18852,N_16297,N_15411);
nor U18853 (N_18853,N_17588,N_16168);
and U18854 (N_18854,N_15165,N_17746);
nand U18855 (N_18855,N_16118,N_15456);
and U18856 (N_18856,N_16612,N_17112);
nand U18857 (N_18857,N_15972,N_16241);
nand U18858 (N_18858,N_16695,N_16684);
nor U18859 (N_18859,N_17163,N_15838);
xor U18860 (N_18860,N_15233,N_17760);
or U18861 (N_18861,N_16789,N_17714);
nor U18862 (N_18862,N_17252,N_17602);
xor U18863 (N_18863,N_16396,N_16504);
or U18864 (N_18864,N_16999,N_15577);
nor U18865 (N_18865,N_16410,N_15597);
xnor U18866 (N_18866,N_15908,N_15846);
nand U18867 (N_18867,N_16667,N_17460);
or U18868 (N_18868,N_17356,N_17507);
or U18869 (N_18869,N_17831,N_17589);
or U18870 (N_18870,N_15063,N_17116);
nand U18871 (N_18871,N_15150,N_15696);
and U18872 (N_18872,N_17422,N_16359);
xor U18873 (N_18873,N_17816,N_16073);
xnor U18874 (N_18874,N_17039,N_17197);
nand U18875 (N_18875,N_17414,N_17262);
and U18876 (N_18876,N_17157,N_15961);
xnor U18877 (N_18877,N_15701,N_16505);
and U18878 (N_18878,N_17568,N_16767);
and U18879 (N_18879,N_15201,N_17563);
or U18880 (N_18880,N_16383,N_17260);
and U18881 (N_18881,N_17089,N_15485);
and U18882 (N_18882,N_16299,N_15166);
and U18883 (N_18883,N_16121,N_15860);
xnor U18884 (N_18884,N_17098,N_16901);
or U18885 (N_18885,N_17158,N_16507);
xnor U18886 (N_18886,N_16929,N_15473);
nor U18887 (N_18887,N_16151,N_16095);
nor U18888 (N_18888,N_16156,N_16274);
nor U18889 (N_18889,N_15318,N_16180);
nor U18890 (N_18890,N_15399,N_17525);
xnor U18891 (N_18891,N_17156,N_15998);
or U18892 (N_18892,N_16227,N_16414);
and U18893 (N_18893,N_16534,N_17043);
xor U18894 (N_18894,N_15172,N_17281);
or U18895 (N_18895,N_16820,N_15986);
and U18896 (N_18896,N_16983,N_17042);
nor U18897 (N_18897,N_16844,N_15787);
nand U18898 (N_18898,N_15046,N_15636);
and U18899 (N_18899,N_15712,N_16254);
and U18900 (N_18900,N_17995,N_16785);
nor U18901 (N_18901,N_15875,N_17824);
xor U18902 (N_18902,N_15885,N_17126);
and U18903 (N_18903,N_17808,N_16715);
xnor U18904 (N_18904,N_16857,N_16561);
nor U18905 (N_18905,N_15258,N_17434);
xnor U18906 (N_18906,N_16657,N_15567);
nand U18907 (N_18907,N_15997,N_16468);
or U18908 (N_18908,N_16760,N_17085);
and U18909 (N_18909,N_17449,N_15818);
or U18910 (N_18910,N_16429,N_16548);
nand U18911 (N_18911,N_17932,N_15309);
xnor U18912 (N_18912,N_16982,N_15905);
or U18913 (N_18913,N_17752,N_15008);
nor U18914 (N_18914,N_17297,N_16310);
xnor U18915 (N_18915,N_15067,N_15828);
and U18916 (N_18916,N_16936,N_15682);
nand U18917 (N_18917,N_15304,N_16028);
nand U18918 (N_18918,N_17462,N_17165);
nor U18919 (N_18919,N_16231,N_16602);
nand U18920 (N_18920,N_15769,N_17587);
and U18921 (N_18921,N_16750,N_16044);
or U18922 (N_18922,N_15066,N_17216);
and U18923 (N_18923,N_16599,N_17779);
nand U18924 (N_18924,N_15685,N_15186);
and U18925 (N_18925,N_17998,N_16403);
nor U18926 (N_18926,N_15865,N_16281);
or U18927 (N_18927,N_17143,N_15299);
and U18928 (N_18928,N_15835,N_17153);
or U18929 (N_18929,N_17184,N_17911);
and U18930 (N_18930,N_17583,N_16910);
and U18931 (N_18931,N_15642,N_16710);
nor U18932 (N_18932,N_15618,N_15338);
and U18933 (N_18933,N_16474,N_17550);
and U18934 (N_18934,N_16610,N_16494);
nand U18935 (N_18935,N_17852,N_16711);
nor U18936 (N_18936,N_15375,N_16689);
xor U18937 (N_18937,N_17603,N_17557);
nor U18938 (N_18938,N_17612,N_17122);
nand U18939 (N_18939,N_16745,N_16301);
nor U18940 (N_18940,N_16998,N_17196);
or U18941 (N_18941,N_16989,N_15241);
and U18942 (N_18942,N_17074,N_15080);
nand U18943 (N_18943,N_15638,N_15256);
and U18944 (N_18944,N_16581,N_16223);
nor U18945 (N_18945,N_15398,N_16621);
nand U18946 (N_18946,N_16531,N_16451);
xnor U18947 (N_18947,N_16158,N_15069);
nor U18948 (N_18948,N_17322,N_16289);
or U18949 (N_18949,N_17499,N_16372);
xnor U18950 (N_18950,N_17131,N_16834);
nor U18951 (N_18951,N_15752,N_16779);
and U18952 (N_18952,N_15721,N_17706);
or U18953 (N_18953,N_16632,N_17332);
and U18954 (N_18954,N_16032,N_16808);
or U18955 (N_18955,N_17868,N_15313);
nand U18956 (N_18956,N_15341,N_15705);
nor U18957 (N_18957,N_17846,N_16868);
nand U18958 (N_18958,N_16464,N_15254);
nor U18959 (N_18959,N_15242,N_16967);
nand U18960 (N_18960,N_15064,N_16114);
xnor U18961 (N_18961,N_15002,N_16701);
xor U18962 (N_18962,N_16364,N_16934);
nand U18963 (N_18963,N_15639,N_17694);
nand U18964 (N_18964,N_17009,N_16117);
nand U18965 (N_18965,N_15239,N_17663);
and U18966 (N_18966,N_16756,N_17897);
xnor U18967 (N_18967,N_16587,N_17318);
and U18968 (N_18968,N_16029,N_17025);
nand U18969 (N_18969,N_16340,N_17797);
and U18970 (N_18970,N_17111,N_17102);
nor U18971 (N_18971,N_16232,N_16287);
or U18972 (N_18972,N_16093,N_16164);
xor U18973 (N_18973,N_16885,N_16608);
xor U18974 (N_18974,N_16278,N_16898);
nor U18975 (N_18975,N_16576,N_17408);
or U18976 (N_18976,N_17916,N_17815);
xnor U18977 (N_18977,N_15422,N_16378);
or U18978 (N_18978,N_16675,N_15786);
and U18979 (N_18979,N_15228,N_16059);
nor U18980 (N_18980,N_17352,N_16134);
xnor U18981 (N_18981,N_16016,N_17164);
and U18982 (N_18982,N_16590,N_17314);
nor U18983 (N_18983,N_17538,N_15089);
nand U18984 (N_18984,N_16744,N_15225);
xnor U18985 (N_18985,N_17651,N_15363);
nor U18986 (N_18986,N_16306,N_16774);
xor U18987 (N_18987,N_17688,N_17210);
nor U18988 (N_18988,N_15680,N_16272);
and U18989 (N_18989,N_16578,N_15183);
or U18990 (N_18990,N_15176,N_15605);
xor U18991 (N_18991,N_17866,N_17822);
and U18992 (N_18992,N_16776,N_16734);
nand U18993 (N_18993,N_16466,N_15049);
and U18994 (N_18994,N_17478,N_17762);
xor U18995 (N_18995,N_15408,N_17287);
or U18996 (N_18996,N_16448,N_15331);
or U18997 (N_18997,N_17077,N_16381);
nor U18998 (N_18998,N_16948,N_15071);
xnor U18999 (N_18999,N_17118,N_16960);
nand U19000 (N_19000,N_17388,N_16951);
nand U19001 (N_19001,N_17051,N_17703);
nor U19002 (N_19002,N_17857,N_17336);
nor U19003 (N_19003,N_16923,N_15947);
nor U19004 (N_19004,N_17787,N_15975);
nor U19005 (N_19005,N_16809,N_16041);
and U19006 (N_19006,N_17505,N_17347);
nand U19007 (N_19007,N_17475,N_17023);
or U19008 (N_19008,N_16665,N_15633);
or U19009 (N_19009,N_15507,N_17103);
nand U19010 (N_19010,N_17946,N_15897);
or U19011 (N_19011,N_17813,N_15122);
nor U19012 (N_19012,N_17802,N_15601);
or U19013 (N_19013,N_15735,N_16304);
or U19014 (N_19014,N_16947,N_17219);
and U19015 (N_19015,N_16252,N_17590);
or U19016 (N_19016,N_15461,N_17540);
nor U19017 (N_19017,N_15133,N_16326);
xor U19018 (N_19018,N_16177,N_17782);
or U19019 (N_19019,N_16645,N_16557);
nand U19020 (N_19020,N_16454,N_15931);
xnor U19021 (N_19021,N_16780,N_15311);
and U19022 (N_19022,N_15795,N_17941);
nor U19023 (N_19023,N_15655,N_15697);
and U19024 (N_19024,N_15106,N_17437);
xnor U19025 (N_19025,N_15393,N_15426);
and U19026 (N_19026,N_16697,N_15774);
or U19027 (N_19027,N_17349,N_15629);
or U19028 (N_19028,N_17177,N_17108);
or U19029 (N_19029,N_17848,N_17903);
nor U19030 (N_19030,N_16161,N_15017);
nor U19031 (N_19031,N_16554,N_17546);
or U19032 (N_19032,N_17064,N_17311);
or U19033 (N_19033,N_15843,N_16215);
xor U19034 (N_19034,N_15484,N_17698);
and U19035 (N_19035,N_15814,N_17367);
nor U19036 (N_19036,N_15445,N_15965);
or U19037 (N_19037,N_17949,N_16952);
xnor U19038 (N_19038,N_17756,N_15579);
or U19039 (N_19039,N_15455,N_15826);
and U19040 (N_19040,N_16867,N_15586);
nor U19041 (N_19041,N_16333,N_17864);
or U19042 (N_19042,N_17291,N_15459);
and U19043 (N_19043,N_16046,N_16025);
nand U19044 (N_19044,N_17979,N_17644);
and U19045 (N_19045,N_17578,N_16174);
xor U19046 (N_19046,N_17675,N_15084);
and U19047 (N_19047,N_17670,N_15316);
and U19048 (N_19048,N_17199,N_15403);
nor U19049 (N_19049,N_16496,N_15901);
xnor U19050 (N_19050,N_15023,N_15462);
nor U19051 (N_19051,N_17555,N_16488);
or U19052 (N_19052,N_17055,N_15914);
nand U19053 (N_19053,N_17652,N_17050);
nor U19054 (N_19054,N_16187,N_15532);
nor U19055 (N_19055,N_17438,N_15490);
and U19056 (N_19056,N_16228,N_17379);
nand U19057 (N_19057,N_16008,N_15189);
xnor U19058 (N_19058,N_15248,N_17327);
or U19059 (N_19059,N_15912,N_16628);
or U19060 (N_19060,N_17804,N_15923);
xor U19061 (N_19061,N_17385,N_15851);
and U19062 (N_19062,N_16620,N_15811);
or U19063 (N_19063,N_16904,N_15921);
nor U19064 (N_19064,N_15548,N_16361);
or U19065 (N_19065,N_16643,N_15959);
or U19066 (N_19066,N_15785,N_17240);
xnor U19067 (N_19067,N_16277,N_15971);
nor U19068 (N_19068,N_17396,N_17716);
nor U19069 (N_19069,N_15231,N_16309);
or U19070 (N_19070,N_15178,N_17994);
nor U19071 (N_19071,N_15936,N_15733);
and U19072 (N_19072,N_16847,N_16559);
xor U19073 (N_19073,N_17899,N_16773);
or U19074 (N_19074,N_17515,N_15211);
nand U19075 (N_19075,N_15631,N_17845);
nand U19076 (N_19076,N_15556,N_15740);
nor U19077 (N_19077,N_16275,N_15234);
xor U19078 (N_19078,N_15376,N_16900);
and U19079 (N_19079,N_17008,N_17320);
xnor U19080 (N_19080,N_17595,N_16078);
nor U19081 (N_19081,N_17067,N_17888);
nor U19082 (N_19082,N_15389,N_17894);
xor U19083 (N_19083,N_15042,N_17455);
xnor U19084 (N_19084,N_16188,N_17871);
and U19085 (N_19085,N_16253,N_15448);
nor U19086 (N_19086,N_17178,N_16102);
xnor U19087 (N_19087,N_15327,N_17636);
and U19088 (N_19088,N_17015,N_15267);
nand U19089 (N_19089,N_15599,N_16194);
nand U19090 (N_19090,N_16146,N_16472);
nor U19091 (N_19091,N_16066,N_16339);
xnor U19092 (N_19092,N_16533,N_16876);
nand U19093 (N_19093,N_15553,N_17120);
nand U19094 (N_19094,N_15761,N_16343);
xnor U19095 (N_19095,N_17256,N_17401);
and U19096 (N_19096,N_15780,N_15330);
nand U19097 (N_19097,N_16626,N_17205);
nand U19098 (N_19098,N_17678,N_17190);
or U19099 (N_19099,N_15519,N_16071);
or U19100 (N_19100,N_17751,N_17279);
xnor U19101 (N_19101,N_17798,N_17106);
and U19102 (N_19102,N_16376,N_16348);
or U19103 (N_19103,N_16136,N_17249);
xor U19104 (N_19104,N_17283,N_15193);
or U19105 (N_19105,N_17127,N_16486);
xnor U19106 (N_19106,N_17432,N_16443);
and U19107 (N_19107,N_17442,N_15794);
nand U19108 (N_19108,N_16656,N_16975);
nor U19109 (N_19109,N_16698,N_17841);
and U19110 (N_19110,N_16358,N_16629);
or U19111 (N_19111,N_15980,N_16394);
and U19112 (N_19112,N_15444,N_15755);
and U19113 (N_19113,N_16043,N_16124);
or U19114 (N_19114,N_16818,N_17676);
nand U19115 (N_19115,N_15169,N_17496);
or U19116 (N_19116,N_17997,N_16064);
nand U19117 (N_19117,N_17799,N_15711);
or U19118 (N_19118,N_15227,N_15706);
nand U19119 (N_19119,N_16000,N_15121);
xnor U19120 (N_19120,N_16050,N_16527);
nor U19121 (N_19121,N_15370,N_15180);
nor U19122 (N_19122,N_15937,N_15294);
nand U19123 (N_19123,N_16023,N_16129);
xnor U19124 (N_19124,N_16426,N_17939);
nor U19125 (N_19125,N_17027,N_15257);
and U19126 (N_19126,N_15290,N_15958);
nand U19127 (N_19127,N_15449,N_17150);
and U19128 (N_19128,N_16498,N_16416);
or U19129 (N_19129,N_15928,N_17523);
nand U19130 (N_19130,N_15053,N_15177);
or U19131 (N_19131,N_16007,N_16673);
nand U19132 (N_19132,N_15055,N_15210);
and U19133 (N_19133,N_16088,N_17161);
and U19134 (N_19134,N_16220,N_16822);
xnor U19135 (N_19135,N_15699,N_16878);
nor U19136 (N_19136,N_16832,N_15380);
nor U19137 (N_19137,N_15286,N_16100);
nor U19138 (N_19138,N_15007,N_17776);
and U19139 (N_19139,N_15839,N_17560);
and U19140 (N_19140,N_17638,N_16219);
xor U19141 (N_19141,N_16171,N_16224);
and U19142 (N_19142,N_17925,N_15073);
and U19143 (N_19143,N_15511,N_16049);
or U19144 (N_19144,N_15916,N_15296);
nor U19145 (N_19145,N_16944,N_17524);
nor U19146 (N_19146,N_16455,N_16762);
or U19147 (N_19147,N_15279,N_15724);
xor U19148 (N_19148,N_17084,N_16615);
nand U19149 (N_19149,N_16233,N_15946);
and U19150 (N_19150,N_15218,N_17629);
nor U19151 (N_19151,N_17138,N_16688);
nor U19152 (N_19152,N_16903,N_15651);
nand U19153 (N_19153,N_17147,N_17443);
nand U19154 (N_19154,N_17330,N_16746);
or U19155 (N_19155,N_17344,N_15305);
or U19156 (N_19156,N_17723,N_15742);
nor U19157 (N_19157,N_16987,N_15364);
nand U19158 (N_19158,N_15942,N_17304);
nor U19159 (N_19159,N_16577,N_16108);
or U19160 (N_19160,N_17489,N_17769);
xnor U19161 (N_19161,N_16160,N_17353);
nand U19162 (N_19162,N_17692,N_17981);
or U19163 (N_19163,N_17114,N_17833);
nand U19164 (N_19164,N_16852,N_16572);
or U19165 (N_19165,N_16891,N_15170);
and U19166 (N_19166,N_15021,N_15764);
and U19167 (N_19167,N_16887,N_17017);
or U19168 (N_19168,N_17229,N_16986);
nand U19169 (N_19169,N_15185,N_17881);
or U19170 (N_19170,N_15686,N_16013);
xnor U19171 (N_19171,N_16708,N_15238);
or U19172 (N_19172,N_16198,N_16420);
xnor U19173 (N_19173,N_16263,N_17271);
or U19174 (N_19174,N_17441,N_16503);
and U19175 (N_19175,N_16437,N_16307);
nor U19176 (N_19176,N_15306,N_17609);
xor U19177 (N_19177,N_17750,N_15949);
and U19178 (N_19178,N_16739,N_16417);
and U19179 (N_19179,N_17207,N_17839);
or U19180 (N_19180,N_17731,N_16938);
or U19181 (N_19181,N_15349,N_15913);
nor U19182 (N_19182,N_16212,N_17029);
nand U19183 (N_19183,N_17830,N_15450);
and U19184 (N_19184,N_15412,N_17650);
and U19185 (N_19185,N_16042,N_15962);
nor U19186 (N_19186,N_15537,N_15674);
xor U19187 (N_19187,N_17653,N_17654);
nand U19188 (N_19188,N_16393,N_17605);
or U19189 (N_19189,N_15048,N_16895);
nand U19190 (N_19190,N_17828,N_16373);
xor U19191 (N_19191,N_17599,N_15058);
nor U19192 (N_19192,N_16091,N_16523);
nand U19193 (N_19193,N_15834,N_16812);
nor U19194 (N_19194,N_16574,N_15168);
and U19195 (N_19195,N_16567,N_15430);
xor U19196 (N_19196,N_15160,N_17006);
nor U19197 (N_19197,N_16522,N_15471);
xor U19198 (N_19198,N_16061,N_15127);
or U19199 (N_19199,N_17865,N_17100);
and U19200 (N_19200,N_17984,N_16017);
nand U19201 (N_19201,N_15182,N_16810);
nand U19202 (N_19202,N_15777,N_17959);
nor U19203 (N_19203,N_17736,N_16825);
or U19204 (N_19204,N_17858,N_15920);
and U19205 (N_19205,N_16950,N_17726);
xnor U19206 (N_19206,N_16104,N_16552);
xnor U19207 (N_19207,N_17018,N_16037);
and U19208 (N_19208,N_15832,N_17964);
xor U19209 (N_19209,N_17626,N_16255);
nand U19210 (N_19210,N_15866,N_17057);
nor U19211 (N_19211,N_17181,N_15561);
nand U19212 (N_19212,N_17826,N_16235);
and U19213 (N_19213,N_15505,N_16218);
xnor U19214 (N_19214,N_16391,N_17317);
and U19215 (N_19215,N_16242,N_16192);
nand U19216 (N_19216,N_17921,N_16765);
nor U19217 (N_19217,N_17278,N_15336);
and U19218 (N_19218,N_16036,N_17290);
nand U19219 (N_19219,N_16439,N_17947);
xnor U19220 (N_19220,N_15894,N_15295);
nor U19221 (N_19221,N_15837,N_16279);
and U19222 (N_19222,N_15116,N_16941);
xor U19223 (N_19223,N_16092,N_17574);
xnor U19224 (N_19224,N_17326,N_16836);
and U19225 (N_19225,N_16663,N_15141);
xnor U19226 (N_19226,N_15574,N_15020);
nor U19227 (N_19227,N_17819,N_16529);
or U19228 (N_19228,N_16747,N_15804);
and U19229 (N_19229,N_16681,N_15668);
nand U19230 (N_19230,N_15778,N_17918);
nand U19231 (N_19231,N_15107,N_16205);
xnor U19232 (N_19232,N_17191,N_17063);
xor U19233 (N_19233,N_17859,N_16258);
or U19234 (N_19234,N_16425,N_16370);
xnor U19235 (N_19235,N_16583,N_16520);
and U19236 (N_19236,N_17695,N_15436);
and U19237 (N_19237,N_16611,N_16525);
nor U19238 (N_19238,N_15100,N_15665);
nand U19239 (N_19239,N_16908,N_15542);
nor U19240 (N_19240,N_16316,N_15397);
and U19241 (N_19241,N_16407,N_15522);
nand U19242 (N_19242,N_15500,N_15195);
and U19243 (N_19243,N_15528,N_15900);
xor U19244 (N_19244,N_16302,N_16377);
nor U19245 (N_19245,N_15917,N_16609);
nand U19246 (N_19246,N_16051,N_17537);
nor U19247 (N_19247,N_17294,N_15800);
or U19248 (N_19248,N_17358,N_17576);
or U19249 (N_19249,N_16467,N_16208);
or U19250 (N_19250,N_15263,N_16791);
or U19251 (N_19251,N_16637,N_17293);
nor U19252 (N_19252,N_15624,N_17620);
and U19253 (N_19253,N_17192,N_17091);
nand U19254 (N_19254,N_16320,N_15409);
and U19255 (N_19255,N_15812,N_17961);
and U19256 (N_19256,N_15587,N_17740);
and U19257 (N_19257,N_15478,N_16821);
nor U19258 (N_19258,N_15075,N_16869);
nand U19259 (N_19259,N_15342,N_17639);
xnor U19260 (N_19260,N_16045,N_16870);
xnor U19261 (N_19261,N_17411,N_16234);
or U19262 (N_19262,N_17856,N_17593);
nor U19263 (N_19263,N_16793,N_16854);
nor U19264 (N_19264,N_16250,N_15284);
and U19265 (N_19265,N_17992,N_17282);
and U19266 (N_19266,N_16303,N_17648);
or U19267 (N_19267,N_15415,N_17145);
xnor U19268 (N_19268,N_15870,N_15095);
and U19269 (N_19269,N_17814,N_15469);
and U19270 (N_19270,N_15039,N_16788);
or U19271 (N_19271,N_15893,N_17755);
xnor U19272 (N_19272,N_17520,N_16943);
and U19273 (N_19273,N_16098,N_16759);
xnor U19274 (N_19274,N_17600,N_16175);
xnor U19275 (N_19275,N_15549,N_15074);
xor U19276 (N_19276,N_17452,N_15688);
or U19277 (N_19277,N_17963,N_16729);
xnor U19278 (N_19278,N_16323,N_17044);
and U19279 (N_19279,N_16829,N_16879);
xor U19280 (N_19280,N_16216,N_17048);
and U19281 (N_19281,N_17909,N_17417);
or U19282 (N_19282,N_15384,N_16949);
and U19283 (N_19283,N_15491,N_17952);
nor U19284 (N_19284,N_15653,N_16459);
and U19285 (N_19285,N_17635,N_15790);
or U19286 (N_19286,N_15994,N_15308);
and U19287 (N_19287,N_17628,N_15266);
nor U19288 (N_19288,N_17943,N_17757);
nand U19289 (N_19289,N_17702,N_16261);
or U19290 (N_19290,N_17545,N_16209);
or U19291 (N_19291,N_15061,N_17500);
nand U19292 (N_19292,N_16173,N_17488);
nor U19293 (N_19293,N_16446,N_16777);
nor U19294 (N_19294,N_16294,N_17146);
and U19295 (N_19295,N_15788,N_15404);
xor U19296 (N_19296,N_15438,N_17457);
nor U19297 (N_19297,N_17071,N_17472);
and U19298 (N_19298,N_15602,N_16401);
nor U19299 (N_19299,N_15425,N_15617);
nand U19300 (N_19300,N_15385,N_17805);
nor U19301 (N_19301,N_16927,N_15878);
or U19302 (N_19302,N_15763,N_15825);
xnor U19303 (N_19303,N_17673,N_17309);
nand U19304 (N_19304,N_17134,N_17233);
nand U19305 (N_19305,N_16434,N_16617);
or U19306 (N_19306,N_15433,N_17667);
or U19307 (N_19307,N_15297,N_16799);
xnor U19308 (N_19308,N_16687,N_17413);
or U19309 (N_19309,N_17665,N_15746);
nor U19310 (N_19310,N_15648,N_17965);
xnor U19311 (N_19311,N_16371,N_15822);
or U19312 (N_19312,N_17492,N_16382);
xor U19313 (N_19313,N_15604,N_15725);
and U19314 (N_19314,N_16120,N_15526);
nand U19315 (N_19315,N_17996,N_17607);
and U19316 (N_19316,N_16236,N_15922);
nand U19317 (N_19317,N_15768,N_17235);
and U19318 (N_19318,N_17000,N_17849);
nor U19319 (N_19319,N_16419,N_16296);
and U19320 (N_19320,N_15130,N_16570);
nor U19321 (N_19321,N_16705,N_16214);
nor U19322 (N_19322,N_17544,N_15030);
and U19323 (N_19323,N_15673,N_16724);
and U19324 (N_19324,N_17905,N_15068);
xor U19325 (N_19325,N_16848,N_15446);
nand U19326 (N_19326,N_17486,N_16162);
or U19327 (N_19327,N_15421,N_16481);
and U19328 (N_19328,N_15162,N_16677);
nor U19329 (N_19329,N_17407,N_15957);
or U19330 (N_19330,N_17737,N_15423);
or U19331 (N_19331,N_15664,N_15285);
and U19332 (N_19332,N_17584,N_15973);
xnor U19333 (N_19333,N_16880,N_17973);
and U19334 (N_19334,N_17130,N_15718);
nand U19335 (N_19335,N_15453,N_17242);
nand U19336 (N_19336,N_17381,N_15460);
or U19337 (N_19337,N_16790,N_15081);
or U19338 (N_19338,N_16485,N_17148);
nor U19339 (N_19339,N_17384,N_17608);
nor U19340 (N_19340,N_15720,N_16874);
xnor U19341 (N_19341,N_16598,N_16499);
nor U19342 (N_19342,N_15025,N_15683);
or U19343 (N_19343,N_16069,N_16140);
or U19344 (N_19344,N_17553,N_17783);
and U19345 (N_19345,N_17459,N_15538);
or U19346 (N_19346,N_16856,N_15535);
and U19347 (N_19347,N_16076,N_17521);
or U19348 (N_19348,N_16268,N_17954);
and U19349 (N_19349,N_15011,N_17468);
and U19350 (N_19350,N_16717,N_17613);
nor U19351 (N_19351,N_17594,N_17215);
xnor U19352 (N_19352,N_16716,N_15391);
and U19353 (N_19353,N_15466,N_15050);
or U19354 (N_19354,N_16217,N_16247);
nor U19355 (N_19355,N_16312,N_16623);
and U19356 (N_19356,N_15630,N_15992);
and U19357 (N_19357,N_15650,N_17494);
nand U19358 (N_19358,N_16638,N_16672);
or U19359 (N_19359,N_16727,N_17518);
xnor U19360 (N_19360,N_15675,N_16353);
nand U19361 (N_19361,N_17292,N_15759);
xnor U19362 (N_19362,N_16027,N_15739);
and U19363 (N_19363,N_15963,N_17745);
xnor U19364 (N_19364,N_16239,N_16176);
nor U19365 (N_19365,N_16978,N_15977);
or U19366 (N_19366,N_15477,N_16650);
nand U19367 (N_19367,N_17910,N_15781);
and U19368 (N_19368,N_16662,N_16569);
nor U19369 (N_19369,N_16613,N_17189);
and U19370 (N_19370,N_15704,N_15614);
nand U19371 (N_19371,N_16048,N_17896);
or U19372 (N_19372,N_16001,N_17389);
xnor U19373 (N_19373,N_16189,N_16475);
and U19374 (N_19374,N_15224,N_16435);
and U19375 (N_19375,N_17512,N_15501);
nor U19376 (N_19376,N_17516,N_16544);
and U19377 (N_19377,N_17140,N_17159);
nand U19378 (N_19378,N_17534,N_15120);
nor U19379 (N_19379,N_16772,N_17541);
or U19380 (N_19380,N_15640,N_16458);
nand U19381 (N_19381,N_15157,N_15082);
and U19382 (N_19382,N_15616,N_16519);
and U19383 (N_19383,N_16853,N_17778);
nand U19384 (N_19384,N_17850,N_16084);
xnor U19385 (N_19385,N_15475,N_15360);
xor U19386 (N_19386,N_16280,N_17066);
nand U19387 (N_19387,N_17474,N_17876);
xnor U19388 (N_19388,N_16798,N_16418);
or U19389 (N_19389,N_15004,N_16031);
xor U19390 (N_19390,N_15033,N_16107);
xnor U19391 (N_19391,N_17440,N_17572);
nand U19392 (N_19392,N_16463,N_15771);
or U19393 (N_19393,N_15427,N_15203);
and U19394 (N_19394,N_17331,N_17986);
or U19395 (N_19395,N_16920,N_16200);
or U19396 (N_19396,N_16647,N_15953);
xnor U19397 (N_19397,N_17558,N_17827);
or U19398 (N_19398,N_15933,N_16317);
nand U19399 (N_19399,N_17699,N_16251);
nor U19400 (N_19400,N_17772,N_15899);
and U19401 (N_19401,N_15323,N_16352);
xor U19402 (N_19402,N_16589,N_16207);
and U19403 (N_19403,N_16797,N_15076);
nand U19404 (N_19404,N_15987,N_17564);
or U19405 (N_19405,N_17248,N_16387);
nor U19406 (N_19406,N_15045,N_16325);
nor U19407 (N_19407,N_16946,N_16824);
nor U19408 (N_19408,N_15018,N_17079);
nor U19409 (N_19409,N_16271,N_15414);
and U19410 (N_19410,N_15472,N_15726);
xor U19411 (N_19411,N_17956,N_15111);
or U19412 (N_19412,N_16955,N_17937);
and U19413 (N_19413,N_17666,N_16082);
xor U19414 (N_19414,N_17872,N_17382);
nand U19415 (N_19415,N_16500,N_16169);
and U19416 (N_19416,N_15743,N_16969);
or U19417 (N_19417,N_15143,N_17549);
or U19418 (N_19418,N_15371,N_17208);
or U19419 (N_19419,N_16109,N_15508);
or U19420 (N_19420,N_17754,N_17780);
xor U19421 (N_19421,N_17536,N_15521);
nand U19422 (N_19422,N_17450,N_17243);
or U19423 (N_19423,N_16979,N_15382);
or U19424 (N_19424,N_17792,N_15707);
xnor U19425 (N_19425,N_15149,N_15454);
or U19426 (N_19426,N_17927,N_16365);
xnor U19427 (N_19427,N_15850,N_15222);
xor U19428 (N_19428,N_17300,N_17183);
or U19429 (N_19429,N_17811,N_17801);
and U19430 (N_19430,N_15646,N_16366);
or U19431 (N_19431,N_17768,N_17681);
xnor U19432 (N_19432,N_15970,N_15978);
nor U19433 (N_19433,N_16807,N_17289);
nor U19434 (N_19434,N_15031,N_15882);
xnor U19435 (N_19435,N_15092,N_16166);
nand U19436 (N_19436,N_15813,N_15753);
nand U19437 (N_19437,N_15981,N_15926);
nand U19438 (N_19438,N_16680,N_16238);
nor U19439 (N_19439,N_15044,N_15550);
nor U19440 (N_19440,N_17877,N_15660);
nor U19441 (N_19441,N_15167,N_15855);
or U19442 (N_19442,N_17717,N_17088);
nand U19443 (N_19443,N_16625,N_17346);
or U19444 (N_19444,N_15251,N_15113);
and U19445 (N_19445,N_15571,N_16090);
or U19446 (N_19446,N_15416,N_17213);
xor U19447 (N_19447,N_15967,N_16075);
nand U19448 (N_19448,N_17313,N_15441);
nand U19449 (N_19449,N_16179,N_17430);
and U19450 (N_19450,N_16491,N_15513);
or U19451 (N_19451,N_17773,N_17481);
nand U19452 (N_19452,N_16528,N_17649);
nand U19453 (N_19453,N_17062,N_17059);
and U19454 (N_19454,N_17034,N_17980);
nand U19455 (N_19455,N_15555,N_15775);
xor U19456 (N_19456,N_15434,N_16077);
and U19457 (N_19457,N_17101,N_16388);
and U19458 (N_19458,N_17713,N_17619);
or U19459 (N_19459,N_16931,N_16597);
or U19460 (N_19460,N_17656,N_16086);
nor U19461 (N_19461,N_15101,N_15487);
and U19462 (N_19462,N_15645,N_15671);
or U19463 (N_19463,N_17942,N_15559);
and U19464 (N_19464,N_16624,N_17144);
nand U19465 (N_19465,N_16083,N_17689);
or U19466 (N_19466,N_16726,N_16319);
or U19467 (N_19467,N_16311,N_17559);
or U19468 (N_19468,N_16827,N_16994);
or U19469 (N_19469,N_15405,N_15988);
nor U19470 (N_19470,N_16315,N_17708);
nor U19471 (N_19471,N_17168,N_17003);
nand U19472 (N_19472,N_15560,N_16712);
xnor U19473 (N_19473,N_15829,N_15570);
xor U19474 (N_19474,N_17268,N_16511);
xnor U19475 (N_19475,N_16973,N_17647);
nand U19476 (N_19476,N_16884,N_15539);
nor U19477 (N_19477,N_15723,N_15348);
and U19478 (N_19478,N_17061,N_15880);
or U19479 (N_19479,N_15930,N_17627);
nand U19480 (N_19480,N_15907,N_16630);
xor U19481 (N_19481,N_15857,N_16331);
nand U19482 (N_19482,N_16327,N_15969);
nand U19483 (N_19483,N_16456,N_17203);
or U19484 (N_19484,N_16022,N_16753);
or U19485 (N_19485,N_16210,N_15868);
and U19486 (N_19486,N_16089,N_16063);
xnor U19487 (N_19487,N_17315,N_17701);
xor U19488 (N_19488,N_15717,N_17657);
nor U19489 (N_19489,N_16670,N_15335);
xnor U19490 (N_19490,N_16575,N_15181);
nand U19491 (N_19491,N_17386,N_16828);
and U19492 (N_19492,N_17891,N_16600);
nand U19493 (N_19493,N_17493,N_17728);
nand U19494 (N_19494,N_15259,N_15883);
nand U19495 (N_19495,N_17393,N_16995);
nand U19496 (N_19496,N_15991,N_17301);
nor U19497 (N_19497,N_15220,N_16718);
or U19498 (N_19498,N_17409,N_15952);
and U19499 (N_19499,N_15881,N_15842);
or U19500 (N_19500,N_16757,N_16277);
nor U19501 (N_19501,N_16377,N_17682);
or U19502 (N_19502,N_15101,N_17164);
nand U19503 (N_19503,N_17124,N_15862);
and U19504 (N_19504,N_15800,N_15612);
nor U19505 (N_19505,N_15020,N_15498);
xor U19506 (N_19506,N_15420,N_17639);
nor U19507 (N_19507,N_16745,N_16765);
xnor U19508 (N_19508,N_16752,N_16973);
or U19509 (N_19509,N_16082,N_16658);
xnor U19510 (N_19510,N_16148,N_16710);
nand U19511 (N_19511,N_15760,N_16804);
or U19512 (N_19512,N_17313,N_15498);
nand U19513 (N_19513,N_15823,N_15177);
or U19514 (N_19514,N_16951,N_17443);
nand U19515 (N_19515,N_17180,N_16070);
or U19516 (N_19516,N_17438,N_16983);
xor U19517 (N_19517,N_17025,N_17575);
or U19518 (N_19518,N_16499,N_17810);
or U19519 (N_19519,N_16473,N_16001);
xor U19520 (N_19520,N_15234,N_16176);
xnor U19521 (N_19521,N_15886,N_16674);
xor U19522 (N_19522,N_16829,N_17822);
nand U19523 (N_19523,N_15718,N_17546);
and U19524 (N_19524,N_17803,N_15219);
nand U19525 (N_19525,N_16669,N_17788);
xor U19526 (N_19526,N_17348,N_16308);
nand U19527 (N_19527,N_17348,N_15517);
nand U19528 (N_19528,N_17969,N_15573);
and U19529 (N_19529,N_17277,N_17178);
and U19530 (N_19530,N_16639,N_15956);
nand U19531 (N_19531,N_15732,N_17789);
nor U19532 (N_19532,N_16926,N_17665);
xnor U19533 (N_19533,N_16595,N_17762);
nand U19534 (N_19534,N_16616,N_15703);
or U19535 (N_19535,N_15200,N_15488);
nor U19536 (N_19536,N_16095,N_16998);
or U19537 (N_19537,N_15424,N_17449);
nand U19538 (N_19538,N_16078,N_15043);
or U19539 (N_19539,N_17302,N_16028);
nor U19540 (N_19540,N_15432,N_17551);
nor U19541 (N_19541,N_16883,N_17006);
or U19542 (N_19542,N_16325,N_17959);
and U19543 (N_19543,N_17510,N_16071);
nand U19544 (N_19544,N_16348,N_17585);
and U19545 (N_19545,N_15594,N_17687);
xnor U19546 (N_19546,N_16589,N_16350);
or U19547 (N_19547,N_17002,N_17621);
nand U19548 (N_19548,N_16053,N_15890);
nand U19549 (N_19549,N_15239,N_15153);
nand U19550 (N_19550,N_17804,N_16032);
and U19551 (N_19551,N_15383,N_16893);
nor U19552 (N_19552,N_16970,N_17636);
xor U19553 (N_19553,N_15091,N_16001);
and U19554 (N_19554,N_15667,N_15881);
or U19555 (N_19555,N_15561,N_16013);
nor U19556 (N_19556,N_17094,N_16644);
xor U19557 (N_19557,N_17236,N_17145);
nor U19558 (N_19558,N_15381,N_16690);
and U19559 (N_19559,N_17081,N_16195);
nor U19560 (N_19560,N_15039,N_16949);
nand U19561 (N_19561,N_16981,N_17535);
nand U19562 (N_19562,N_16771,N_17754);
nand U19563 (N_19563,N_16149,N_16806);
and U19564 (N_19564,N_16271,N_17583);
xnor U19565 (N_19565,N_15452,N_15805);
and U19566 (N_19566,N_15123,N_15799);
xnor U19567 (N_19567,N_16898,N_15605);
xor U19568 (N_19568,N_17564,N_15680);
nor U19569 (N_19569,N_15100,N_16185);
or U19570 (N_19570,N_15053,N_15912);
and U19571 (N_19571,N_16094,N_17561);
or U19572 (N_19572,N_15073,N_16650);
nor U19573 (N_19573,N_15922,N_16804);
nand U19574 (N_19574,N_15165,N_16688);
and U19575 (N_19575,N_15382,N_17230);
nor U19576 (N_19576,N_15842,N_17415);
or U19577 (N_19577,N_16258,N_15725);
or U19578 (N_19578,N_16221,N_15255);
xnor U19579 (N_19579,N_15429,N_17654);
nand U19580 (N_19580,N_17691,N_17029);
or U19581 (N_19581,N_17653,N_15424);
nor U19582 (N_19582,N_15712,N_17735);
xnor U19583 (N_19583,N_15517,N_15960);
and U19584 (N_19584,N_17623,N_17122);
and U19585 (N_19585,N_16758,N_16756);
nor U19586 (N_19586,N_15565,N_15824);
and U19587 (N_19587,N_17621,N_16623);
xor U19588 (N_19588,N_15019,N_16925);
or U19589 (N_19589,N_16727,N_16601);
nand U19590 (N_19590,N_16156,N_16460);
and U19591 (N_19591,N_16041,N_16057);
and U19592 (N_19592,N_17889,N_16034);
or U19593 (N_19593,N_15877,N_15021);
nand U19594 (N_19594,N_17713,N_17572);
and U19595 (N_19595,N_17606,N_16066);
or U19596 (N_19596,N_15785,N_17920);
and U19597 (N_19597,N_17874,N_16285);
and U19598 (N_19598,N_17732,N_16812);
nand U19599 (N_19599,N_17399,N_17010);
and U19600 (N_19600,N_17328,N_15180);
xor U19601 (N_19601,N_16623,N_16858);
xor U19602 (N_19602,N_16383,N_17777);
and U19603 (N_19603,N_17844,N_16980);
xor U19604 (N_19604,N_15982,N_15230);
and U19605 (N_19605,N_15549,N_15525);
and U19606 (N_19606,N_16753,N_16477);
xnor U19607 (N_19607,N_15040,N_15664);
nand U19608 (N_19608,N_15815,N_15919);
or U19609 (N_19609,N_17168,N_15259);
nor U19610 (N_19610,N_15301,N_17786);
nand U19611 (N_19611,N_15402,N_17868);
and U19612 (N_19612,N_15712,N_15055);
nand U19613 (N_19613,N_16460,N_16107);
and U19614 (N_19614,N_17212,N_16667);
nand U19615 (N_19615,N_17010,N_16829);
or U19616 (N_19616,N_17168,N_17621);
nand U19617 (N_19617,N_15493,N_15976);
xnor U19618 (N_19618,N_15003,N_15575);
xor U19619 (N_19619,N_17403,N_15867);
nor U19620 (N_19620,N_17964,N_16736);
or U19621 (N_19621,N_16743,N_17584);
and U19622 (N_19622,N_15719,N_17430);
xnor U19623 (N_19623,N_16401,N_15386);
or U19624 (N_19624,N_15046,N_17432);
nand U19625 (N_19625,N_15936,N_17185);
and U19626 (N_19626,N_15281,N_17276);
and U19627 (N_19627,N_15615,N_15698);
or U19628 (N_19628,N_16703,N_16510);
nand U19629 (N_19629,N_16205,N_17179);
nor U19630 (N_19630,N_17641,N_15057);
and U19631 (N_19631,N_16542,N_17490);
nand U19632 (N_19632,N_15309,N_17452);
and U19633 (N_19633,N_16472,N_17912);
or U19634 (N_19634,N_16465,N_17633);
nand U19635 (N_19635,N_16356,N_16113);
or U19636 (N_19636,N_17820,N_16899);
nand U19637 (N_19637,N_16097,N_16322);
nand U19638 (N_19638,N_15117,N_15965);
xor U19639 (N_19639,N_17397,N_15553);
xor U19640 (N_19640,N_17815,N_17041);
or U19641 (N_19641,N_17683,N_17657);
xnor U19642 (N_19642,N_17753,N_16057);
nand U19643 (N_19643,N_17258,N_15159);
xnor U19644 (N_19644,N_16176,N_17983);
and U19645 (N_19645,N_17001,N_16627);
and U19646 (N_19646,N_15565,N_16163);
nand U19647 (N_19647,N_17093,N_15297);
and U19648 (N_19648,N_17966,N_16180);
or U19649 (N_19649,N_16806,N_15711);
xnor U19650 (N_19650,N_17634,N_15929);
nor U19651 (N_19651,N_15915,N_17727);
nor U19652 (N_19652,N_16736,N_15423);
and U19653 (N_19653,N_17890,N_15096);
nand U19654 (N_19654,N_16616,N_17261);
nor U19655 (N_19655,N_15934,N_16321);
and U19656 (N_19656,N_16027,N_16722);
and U19657 (N_19657,N_16562,N_17253);
and U19658 (N_19658,N_16171,N_16579);
nand U19659 (N_19659,N_15350,N_17371);
xor U19660 (N_19660,N_16312,N_16648);
and U19661 (N_19661,N_15709,N_15872);
nand U19662 (N_19662,N_17178,N_15810);
and U19663 (N_19663,N_17371,N_16779);
nor U19664 (N_19664,N_16871,N_16834);
nand U19665 (N_19665,N_16657,N_16961);
xnor U19666 (N_19666,N_17354,N_17814);
nand U19667 (N_19667,N_16682,N_15055);
nor U19668 (N_19668,N_17005,N_16469);
or U19669 (N_19669,N_17688,N_17743);
nor U19670 (N_19670,N_16894,N_16923);
and U19671 (N_19671,N_17285,N_16086);
nand U19672 (N_19672,N_17675,N_16080);
nand U19673 (N_19673,N_15260,N_16844);
and U19674 (N_19674,N_16391,N_16075);
nor U19675 (N_19675,N_15356,N_17943);
and U19676 (N_19676,N_16007,N_15731);
or U19677 (N_19677,N_17988,N_15235);
nor U19678 (N_19678,N_16370,N_17286);
and U19679 (N_19679,N_16993,N_15456);
xnor U19680 (N_19680,N_17278,N_15311);
xnor U19681 (N_19681,N_17952,N_17836);
nand U19682 (N_19682,N_16389,N_15373);
xnor U19683 (N_19683,N_16658,N_15282);
and U19684 (N_19684,N_17765,N_16771);
or U19685 (N_19685,N_16339,N_16717);
or U19686 (N_19686,N_15894,N_15436);
and U19687 (N_19687,N_16331,N_16298);
xnor U19688 (N_19688,N_17575,N_16595);
nor U19689 (N_19689,N_16033,N_15256);
nand U19690 (N_19690,N_17141,N_17975);
nor U19691 (N_19691,N_16770,N_17121);
nand U19692 (N_19692,N_15287,N_15004);
xor U19693 (N_19693,N_15842,N_17045);
and U19694 (N_19694,N_15184,N_15573);
xor U19695 (N_19695,N_17165,N_15914);
or U19696 (N_19696,N_17601,N_16880);
xor U19697 (N_19697,N_16051,N_15619);
xnor U19698 (N_19698,N_17893,N_16023);
or U19699 (N_19699,N_17072,N_15625);
xor U19700 (N_19700,N_16352,N_17049);
and U19701 (N_19701,N_16530,N_17016);
and U19702 (N_19702,N_17290,N_17779);
xor U19703 (N_19703,N_17284,N_16890);
nand U19704 (N_19704,N_17486,N_16887);
nand U19705 (N_19705,N_15337,N_16119);
xor U19706 (N_19706,N_15382,N_15367);
or U19707 (N_19707,N_15961,N_17258);
nor U19708 (N_19708,N_16251,N_16778);
nand U19709 (N_19709,N_15554,N_15900);
xor U19710 (N_19710,N_16602,N_17005);
and U19711 (N_19711,N_16266,N_17688);
nand U19712 (N_19712,N_17650,N_17921);
and U19713 (N_19713,N_15056,N_16529);
or U19714 (N_19714,N_16441,N_15677);
xnor U19715 (N_19715,N_15650,N_17140);
nand U19716 (N_19716,N_17541,N_16386);
xnor U19717 (N_19717,N_17216,N_15124);
nor U19718 (N_19718,N_17875,N_16054);
or U19719 (N_19719,N_15180,N_17069);
nor U19720 (N_19720,N_16603,N_15696);
nor U19721 (N_19721,N_17327,N_16913);
and U19722 (N_19722,N_17096,N_15633);
xnor U19723 (N_19723,N_17304,N_17582);
or U19724 (N_19724,N_16893,N_15770);
nor U19725 (N_19725,N_16335,N_15049);
xor U19726 (N_19726,N_15289,N_17855);
xnor U19727 (N_19727,N_16413,N_16332);
xor U19728 (N_19728,N_15067,N_16431);
nor U19729 (N_19729,N_16993,N_15405);
or U19730 (N_19730,N_17975,N_16220);
xor U19731 (N_19731,N_17663,N_15651);
nand U19732 (N_19732,N_15634,N_16310);
and U19733 (N_19733,N_17690,N_17061);
or U19734 (N_19734,N_17898,N_15787);
nand U19735 (N_19735,N_16487,N_17698);
and U19736 (N_19736,N_16707,N_15373);
nand U19737 (N_19737,N_16433,N_16745);
nor U19738 (N_19738,N_15008,N_17657);
nand U19739 (N_19739,N_17039,N_16562);
and U19740 (N_19740,N_16427,N_15223);
xnor U19741 (N_19741,N_17347,N_16434);
nand U19742 (N_19742,N_15185,N_15403);
and U19743 (N_19743,N_17229,N_15709);
nand U19744 (N_19744,N_16385,N_17961);
xnor U19745 (N_19745,N_15721,N_15470);
nand U19746 (N_19746,N_15099,N_17232);
or U19747 (N_19747,N_16225,N_15521);
xor U19748 (N_19748,N_17792,N_15738);
xor U19749 (N_19749,N_16089,N_17062);
nor U19750 (N_19750,N_17537,N_15807);
xnor U19751 (N_19751,N_16812,N_17700);
nor U19752 (N_19752,N_15016,N_17376);
and U19753 (N_19753,N_17010,N_16769);
nand U19754 (N_19754,N_16665,N_17808);
and U19755 (N_19755,N_16524,N_16342);
nor U19756 (N_19756,N_17173,N_16886);
xnor U19757 (N_19757,N_15905,N_15907);
nor U19758 (N_19758,N_15476,N_17925);
nor U19759 (N_19759,N_15611,N_17785);
nor U19760 (N_19760,N_16964,N_15442);
nand U19761 (N_19761,N_16343,N_15323);
and U19762 (N_19762,N_17485,N_17053);
nor U19763 (N_19763,N_15527,N_17063);
nand U19764 (N_19764,N_17629,N_16644);
xnor U19765 (N_19765,N_16427,N_17124);
nor U19766 (N_19766,N_17986,N_16622);
and U19767 (N_19767,N_15392,N_15362);
nand U19768 (N_19768,N_15987,N_17965);
and U19769 (N_19769,N_17032,N_17884);
xnor U19770 (N_19770,N_17105,N_15503);
or U19771 (N_19771,N_16591,N_16083);
xor U19772 (N_19772,N_15672,N_17849);
xnor U19773 (N_19773,N_16119,N_15577);
nand U19774 (N_19774,N_17032,N_15962);
and U19775 (N_19775,N_16739,N_17381);
nand U19776 (N_19776,N_15348,N_15293);
xnor U19777 (N_19777,N_16023,N_17140);
nor U19778 (N_19778,N_17487,N_17353);
and U19779 (N_19779,N_17102,N_17392);
or U19780 (N_19780,N_17888,N_17518);
or U19781 (N_19781,N_17144,N_17137);
or U19782 (N_19782,N_15781,N_15810);
nand U19783 (N_19783,N_15174,N_15389);
or U19784 (N_19784,N_17555,N_16431);
or U19785 (N_19785,N_16462,N_16821);
and U19786 (N_19786,N_15461,N_16534);
or U19787 (N_19787,N_17768,N_17083);
xor U19788 (N_19788,N_17862,N_15538);
xnor U19789 (N_19789,N_15716,N_16488);
nor U19790 (N_19790,N_16124,N_17151);
xnor U19791 (N_19791,N_16458,N_15398);
or U19792 (N_19792,N_17510,N_17760);
and U19793 (N_19793,N_15715,N_17366);
and U19794 (N_19794,N_16591,N_15485);
nor U19795 (N_19795,N_16734,N_15237);
and U19796 (N_19796,N_17852,N_17414);
and U19797 (N_19797,N_16592,N_17211);
nor U19798 (N_19798,N_16313,N_17056);
nand U19799 (N_19799,N_17201,N_15672);
xnor U19800 (N_19800,N_16272,N_15651);
nor U19801 (N_19801,N_16333,N_15224);
xor U19802 (N_19802,N_17435,N_16267);
nor U19803 (N_19803,N_15282,N_16533);
or U19804 (N_19804,N_16945,N_15552);
and U19805 (N_19805,N_15098,N_15877);
nand U19806 (N_19806,N_17779,N_17945);
and U19807 (N_19807,N_17558,N_15843);
and U19808 (N_19808,N_16459,N_15922);
or U19809 (N_19809,N_15809,N_17879);
nor U19810 (N_19810,N_16904,N_17766);
or U19811 (N_19811,N_16803,N_17056);
xor U19812 (N_19812,N_17372,N_17669);
xor U19813 (N_19813,N_16482,N_15116);
nor U19814 (N_19814,N_15922,N_17472);
nor U19815 (N_19815,N_17875,N_16140);
xnor U19816 (N_19816,N_17167,N_15629);
xnor U19817 (N_19817,N_17853,N_16441);
or U19818 (N_19818,N_17720,N_16129);
nor U19819 (N_19819,N_16955,N_17100);
nand U19820 (N_19820,N_15726,N_15403);
nor U19821 (N_19821,N_15885,N_17845);
xor U19822 (N_19822,N_16764,N_17170);
nand U19823 (N_19823,N_17515,N_15804);
or U19824 (N_19824,N_16590,N_15801);
nor U19825 (N_19825,N_17745,N_15897);
nand U19826 (N_19826,N_15579,N_16775);
nand U19827 (N_19827,N_15342,N_17093);
nor U19828 (N_19828,N_17327,N_16167);
or U19829 (N_19829,N_16809,N_15675);
nand U19830 (N_19830,N_16373,N_17612);
nor U19831 (N_19831,N_16274,N_15318);
or U19832 (N_19832,N_15831,N_15982);
and U19833 (N_19833,N_16628,N_17768);
nand U19834 (N_19834,N_16575,N_17291);
or U19835 (N_19835,N_17235,N_16620);
and U19836 (N_19836,N_15255,N_15600);
or U19837 (N_19837,N_17601,N_15072);
nand U19838 (N_19838,N_17681,N_17028);
nor U19839 (N_19839,N_15893,N_16687);
and U19840 (N_19840,N_16637,N_15829);
and U19841 (N_19841,N_17167,N_16088);
nand U19842 (N_19842,N_16755,N_17253);
xor U19843 (N_19843,N_17280,N_15898);
nand U19844 (N_19844,N_17249,N_15751);
and U19845 (N_19845,N_15330,N_16912);
nand U19846 (N_19846,N_17943,N_16312);
or U19847 (N_19847,N_17090,N_15947);
and U19848 (N_19848,N_15758,N_15262);
and U19849 (N_19849,N_16913,N_15825);
nand U19850 (N_19850,N_16370,N_16173);
nor U19851 (N_19851,N_16427,N_16547);
nand U19852 (N_19852,N_17787,N_16818);
xnor U19853 (N_19853,N_17246,N_15446);
or U19854 (N_19854,N_15128,N_17979);
and U19855 (N_19855,N_16606,N_15348);
nand U19856 (N_19856,N_17461,N_17246);
or U19857 (N_19857,N_15451,N_16982);
nand U19858 (N_19858,N_17506,N_16966);
and U19859 (N_19859,N_17258,N_17999);
or U19860 (N_19860,N_16253,N_16405);
or U19861 (N_19861,N_17571,N_17744);
xor U19862 (N_19862,N_16543,N_15831);
or U19863 (N_19863,N_16035,N_17348);
xnor U19864 (N_19864,N_16696,N_16855);
or U19865 (N_19865,N_16766,N_17920);
nor U19866 (N_19866,N_17042,N_15562);
nand U19867 (N_19867,N_15005,N_15360);
and U19868 (N_19868,N_17243,N_17865);
or U19869 (N_19869,N_17048,N_15245);
and U19870 (N_19870,N_17463,N_16467);
xor U19871 (N_19871,N_16928,N_17033);
or U19872 (N_19872,N_15623,N_15006);
nand U19873 (N_19873,N_15193,N_16329);
or U19874 (N_19874,N_17471,N_16628);
xor U19875 (N_19875,N_17147,N_15678);
and U19876 (N_19876,N_15427,N_17676);
nor U19877 (N_19877,N_17559,N_15143);
or U19878 (N_19878,N_17501,N_16885);
nor U19879 (N_19879,N_17560,N_16861);
xnor U19880 (N_19880,N_15245,N_15473);
nand U19881 (N_19881,N_17677,N_15587);
xnor U19882 (N_19882,N_16986,N_16057);
and U19883 (N_19883,N_15940,N_17316);
nor U19884 (N_19884,N_16473,N_15589);
nand U19885 (N_19885,N_16907,N_15533);
or U19886 (N_19886,N_15455,N_15888);
xnor U19887 (N_19887,N_17509,N_17557);
xor U19888 (N_19888,N_16050,N_15776);
nor U19889 (N_19889,N_17166,N_15840);
xor U19890 (N_19890,N_17527,N_16158);
nor U19891 (N_19891,N_17900,N_17344);
xnor U19892 (N_19892,N_17970,N_17380);
nor U19893 (N_19893,N_17815,N_16107);
or U19894 (N_19894,N_15287,N_17309);
or U19895 (N_19895,N_15378,N_15497);
nand U19896 (N_19896,N_15808,N_15489);
nand U19897 (N_19897,N_15102,N_17283);
nand U19898 (N_19898,N_16584,N_17539);
and U19899 (N_19899,N_15098,N_17411);
or U19900 (N_19900,N_17415,N_17466);
xnor U19901 (N_19901,N_16089,N_17042);
and U19902 (N_19902,N_16656,N_15176);
nand U19903 (N_19903,N_16741,N_16273);
and U19904 (N_19904,N_17850,N_15854);
xor U19905 (N_19905,N_17073,N_16062);
nor U19906 (N_19906,N_15338,N_16260);
and U19907 (N_19907,N_16225,N_17498);
and U19908 (N_19908,N_15701,N_16648);
nor U19909 (N_19909,N_15090,N_16527);
or U19910 (N_19910,N_15858,N_17935);
xor U19911 (N_19911,N_16882,N_15789);
nand U19912 (N_19912,N_15612,N_15624);
nor U19913 (N_19913,N_16410,N_15946);
nand U19914 (N_19914,N_17422,N_15764);
xnor U19915 (N_19915,N_15806,N_15415);
or U19916 (N_19916,N_17529,N_17532);
and U19917 (N_19917,N_17233,N_15155);
nor U19918 (N_19918,N_16913,N_15972);
or U19919 (N_19919,N_15426,N_16495);
and U19920 (N_19920,N_17021,N_15670);
nor U19921 (N_19921,N_16378,N_16070);
and U19922 (N_19922,N_16058,N_16161);
nor U19923 (N_19923,N_15110,N_16697);
and U19924 (N_19924,N_17015,N_15811);
or U19925 (N_19925,N_17112,N_15628);
and U19926 (N_19926,N_16090,N_17160);
or U19927 (N_19927,N_17614,N_16853);
or U19928 (N_19928,N_16898,N_16710);
xnor U19929 (N_19929,N_17443,N_16109);
or U19930 (N_19930,N_17077,N_17004);
or U19931 (N_19931,N_16688,N_16821);
or U19932 (N_19932,N_17120,N_17149);
or U19933 (N_19933,N_15894,N_15341);
or U19934 (N_19934,N_17521,N_16013);
or U19935 (N_19935,N_16679,N_15381);
xnor U19936 (N_19936,N_15859,N_15679);
or U19937 (N_19937,N_17754,N_16384);
or U19938 (N_19938,N_17128,N_17714);
or U19939 (N_19939,N_17500,N_16992);
nand U19940 (N_19940,N_15005,N_16725);
nor U19941 (N_19941,N_17375,N_16771);
or U19942 (N_19942,N_15275,N_15871);
xor U19943 (N_19943,N_15027,N_17657);
and U19944 (N_19944,N_16634,N_17330);
and U19945 (N_19945,N_17511,N_16924);
nand U19946 (N_19946,N_17943,N_16103);
nand U19947 (N_19947,N_16408,N_15131);
nor U19948 (N_19948,N_17404,N_15284);
or U19949 (N_19949,N_16162,N_17700);
nor U19950 (N_19950,N_16140,N_16998);
nand U19951 (N_19951,N_17521,N_17160);
xnor U19952 (N_19952,N_15152,N_17141);
and U19953 (N_19953,N_15627,N_15787);
nor U19954 (N_19954,N_17304,N_16217);
nor U19955 (N_19955,N_15754,N_15918);
or U19956 (N_19956,N_15955,N_15032);
nand U19957 (N_19957,N_17929,N_17197);
or U19958 (N_19958,N_15383,N_15136);
xor U19959 (N_19959,N_15669,N_16324);
nor U19960 (N_19960,N_16833,N_17660);
nand U19961 (N_19961,N_17369,N_16595);
xnor U19962 (N_19962,N_15638,N_16973);
nor U19963 (N_19963,N_15404,N_15057);
nor U19964 (N_19964,N_15961,N_15156);
xor U19965 (N_19965,N_17136,N_15797);
nand U19966 (N_19966,N_16930,N_16994);
nand U19967 (N_19967,N_15833,N_17750);
nor U19968 (N_19968,N_16392,N_15032);
or U19969 (N_19969,N_15671,N_15097);
nand U19970 (N_19970,N_17219,N_16380);
or U19971 (N_19971,N_16531,N_15595);
xor U19972 (N_19972,N_17854,N_16464);
and U19973 (N_19973,N_15959,N_17913);
nor U19974 (N_19974,N_17574,N_15570);
nor U19975 (N_19975,N_17251,N_16642);
or U19976 (N_19976,N_16398,N_17065);
nand U19977 (N_19977,N_17368,N_17448);
and U19978 (N_19978,N_16106,N_16367);
xor U19979 (N_19979,N_16702,N_16422);
and U19980 (N_19980,N_15525,N_15374);
nor U19981 (N_19981,N_17160,N_16527);
nand U19982 (N_19982,N_17600,N_16351);
xor U19983 (N_19983,N_16620,N_17368);
nand U19984 (N_19984,N_16752,N_17153);
nand U19985 (N_19985,N_17866,N_15138);
nor U19986 (N_19986,N_16252,N_17468);
and U19987 (N_19987,N_16888,N_15974);
nand U19988 (N_19988,N_16036,N_16637);
nor U19989 (N_19989,N_15713,N_17760);
and U19990 (N_19990,N_15936,N_17888);
xor U19991 (N_19991,N_15244,N_17567);
xor U19992 (N_19992,N_17289,N_15563);
and U19993 (N_19993,N_16469,N_17153);
or U19994 (N_19994,N_15785,N_16290);
and U19995 (N_19995,N_16352,N_16225);
and U19996 (N_19996,N_16872,N_17553);
nor U19997 (N_19997,N_16937,N_15069);
xor U19998 (N_19998,N_15215,N_17943);
nor U19999 (N_19999,N_16576,N_15324);
nor U20000 (N_20000,N_15050,N_17086);
or U20001 (N_20001,N_16946,N_15341);
xor U20002 (N_20002,N_17969,N_17587);
nand U20003 (N_20003,N_15253,N_17585);
xnor U20004 (N_20004,N_16042,N_15667);
xor U20005 (N_20005,N_17248,N_16765);
nand U20006 (N_20006,N_15677,N_17629);
or U20007 (N_20007,N_16053,N_16067);
nor U20008 (N_20008,N_17436,N_17663);
nand U20009 (N_20009,N_15383,N_17865);
and U20010 (N_20010,N_16039,N_16048);
or U20011 (N_20011,N_16864,N_16908);
and U20012 (N_20012,N_15890,N_16162);
or U20013 (N_20013,N_15518,N_16206);
xnor U20014 (N_20014,N_17773,N_17774);
or U20015 (N_20015,N_17782,N_16631);
and U20016 (N_20016,N_17891,N_17241);
or U20017 (N_20017,N_15797,N_16890);
or U20018 (N_20018,N_15850,N_17082);
or U20019 (N_20019,N_17245,N_15770);
and U20020 (N_20020,N_17121,N_15852);
or U20021 (N_20021,N_17139,N_16890);
or U20022 (N_20022,N_17015,N_16493);
nor U20023 (N_20023,N_16944,N_17786);
or U20024 (N_20024,N_16456,N_15138);
nand U20025 (N_20025,N_17904,N_16401);
nand U20026 (N_20026,N_17763,N_17992);
and U20027 (N_20027,N_16664,N_17742);
nor U20028 (N_20028,N_16276,N_17086);
and U20029 (N_20029,N_16146,N_16269);
nand U20030 (N_20030,N_15087,N_17682);
or U20031 (N_20031,N_16863,N_15364);
or U20032 (N_20032,N_15759,N_17976);
or U20033 (N_20033,N_15328,N_15258);
or U20034 (N_20034,N_17774,N_17520);
or U20035 (N_20035,N_17750,N_17916);
nand U20036 (N_20036,N_16226,N_17781);
or U20037 (N_20037,N_15399,N_17527);
or U20038 (N_20038,N_15999,N_16363);
nand U20039 (N_20039,N_15578,N_15311);
xor U20040 (N_20040,N_15623,N_17370);
nor U20041 (N_20041,N_15321,N_15093);
nor U20042 (N_20042,N_17496,N_15951);
nand U20043 (N_20043,N_15641,N_16944);
nand U20044 (N_20044,N_16100,N_17663);
xor U20045 (N_20045,N_17935,N_16357);
nor U20046 (N_20046,N_15941,N_17735);
or U20047 (N_20047,N_15398,N_17767);
nor U20048 (N_20048,N_15637,N_16109);
xor U20049 (N_20049,N_17342,N_16108);
nand U20050 (N_20050,N_15078,N_17637);
or U20051 (N_20051,N_15091,N_17944);
nor U20052 (N_20052,N_15416,N_17974);
and U20053 (N_20053,N_15321,N_16609);
xnor U20054 (N_20054,N_17253,N_16439);
or U20055 (N_20055,N_17165,N_16406);
nor U20056 (N_20056,N_17689,N_15583);
and U20057 (N_20057,N_17831,N_17221);
and U20058 (N_20058,N_16806,N_16313);
or U20059 (N_20059,N_17929,N_16410);
nor U20060 (N_20060,N_17348,N_17226);
nand U20061 (N_20061,N_17978,N_17210);
and U20062 (N_20062,N_16003,N_16315);
nand U20063 (N_20063,N_17436,N_16355);
nand U20064 (N_20064,N_15889,N_15071);
and U20065 (N_20065,N_16967,N_17010);
and U20066 (N_20066,N_16483,N_15323);
or U20067 (N_20067,N_17074,N_15113);
or U20068 (N_20068,N_15531,N_16777);
or U20069 (N_20069,N_17147,N_15718);
nand U20070 (N_20070,N_16279,N_15589);
or U20071 (N_20071,N_15198,N_17154);
and U20072 (N_20072,N_15766,N_16934);
nor U20073 (N_20073,N_15794,N_15679);
xnor U20074 (N_20074,N_17153,N_16422);
and U20075 (N_20075,N_17609,N_17937);
nor U20076 (N_20076,N_15011,N_15437);
xor U20077 (N_20077,N_15276,N_16095);
nand U20078 (N_20078,N_16981,N_15340);
nor U20079 (N_20079,N_15618,N_16729);
or U20080 (N_20080,N_17460,N_16993);
nand U20081 (N_20081,N_17570,N_15434);
xor U20082 (N_20082,N_15984,N_17799);
xor U20083 (N_20083,N_15286,N_15566);
xnor U20084 (N_20084,N_15537,N_17853);
xor U20085 (N_20085,N_15987,N_15276);
nor U20086 (N_20086,N_15574,N_16176);
or U20087 (N_20087,N_15685,N_15217);
nand U20088 (N_20088,N_16984,N_17784);
nand U20089 (N_20089,N_17461,N_15155);
xnor U20090 (N_20090,N_17272,N_15291);
nand U20091 (N_20091,N_15728,N_16669);
and U20092 (N_20092,N_17134,N_15888);
or U20093 (N_20093,N_17898,N_15854);
and U20094 (N_20094,N_17643,N_17079);
nand U20095 (N_20095,N_15285,N_16577);
nor U20096 (N_20096,N_16068,N_17961);
nand U20097 (N_20097,N_16489,N_16495);
nand U20098 (N_20098,N_15878,N_16047);
nand U20099 (N_20099,N_15333,N_16725);
and U20100 (N_20100,N_17407,N_17042);
or U20101 (N_20101,N_17321,N_16061);
and U20102 (N_20102,N_17530,N_16477);
xnor U20103 (N_20103,N_17368,N_17728);
nand U20104 (N_20104,N_16956,N_17875);
nor U20105 (N_20105,N_16983,N_15715);
nor U20106 (N_20106,N_16800,N_15108);
nor U20107 (N_20107,N_15607,N_15610);
and U20108 (N_20108,N_16228,N_16874);
or U20109 (N_20109,N_16520,N_16438);
xnor U20110 (N_20110,N_15135,N_16508);
and U20111 (N_20111,N_17565,N_15607);
xor U20112 (N_20112,N_17129,N_15021);
or U20113 (N_20113,N_17901,N_17078);
nand U20114 (N_20114,N_16917,N_16403);
nor U20115 (N_20115,N_15840,N_15876);
or U20116 (N_20116,N_17455,N_17564);
or U20117 (N_20117,N_17388,N_16171);
xnor U20118 (N_20118,N_17316,N_17350);
or U20119 (N_20119,N_15983,N_16590);
nor U20120 (N_20120,N_15849,N_15729);
xnor U20121 (N_20121,N_17898,N_16038);
nor U20122 (N_20122,N_16102,N_17550);
xor U20123 (N_20123,N_15229,N_17262);
xor U20124 (N_20124,N_16818,N_16250);
and U20125 (N_20125,N_17007,N_15882);
and U20126 (N_20126,N_17367,N_15400);
or U20127 (N_20127,N_17586,N_16387);
or U20128 (N_20128,N_17727,N_15558);
and U20129 (N_20129,N_17375,N_16803);
nor U20130 (N_20130,N_16364,N_17409);
nand U20131 (N_20131,N_17172,N_15398);
and U20132 (N_20132,N_15102,N_16461);
nor U20133 (N_20133,N_17214,N_15822);
or U20134 (N_20134,N_16905,N_16752);
xnor U20135 (N_20135,N_15750,N_17791);
nand U20136 (N_20136,N_17600,N_17601);
xor U20137 (N_20137,N_16556,N_17400);
nand U20138 (N_20138,N_17403,N_17694);
nand U20139 (N_20139,N_16690,N_17667);
nand U20140 (N_20140,N_17932,N_16144);
nor U20141 (N_20141,N_15987,N_15057);
xor U20142 (N_20142,N_15265,N_17595);
and U20143 (N_20143,N_15923,N_15870);
nor U20144 (N_20144,N_16900,N_16718);
and U20145 (N_20145,N_17475,N_16965);
xnor U20146 (N_20146,N_16799,N_17235);
or U20147 (N_20147,N_16654,N_16912);
and U20148 (N_20148,N_16441,N_15575);
nand U20149 (N_20149,N_16029,N_15853);
nand U20150 (N_20150,N_17651,N_17731);
xnor U20151 (N_20151,N_16976,N_17439);
xnor U20152 (N_20152,N_17436,N_16378);
nor U20153 (N_20153,N_17820,N_15587);
or U20154 (N_20154,N_15972,N_16259);
or U20155 (N_20155,N_17696,N_17665);
nor U20156 (N_20156,N_16124,N_17045);
nand U20157 (N_20157,N_17570,N_16436);
nor U20158 (N_20158,N_15941,N_15470);
or U20159 (N_20159,N_16883,N_17197);
nand U20160 (N_20160,N_17349,N_16168);
or U20161 (N_20161,N_16641,N_15282);
xnor U20162 (N_20162,N_17299,N_15799);
xor U20163 (N_20163,N_15673,N_16971);
or U20164 (N_20164,N_15917,N_15440);
nand U20165 (N_20165,N_16021,N_17401);
nand U20166 (N_20166,N_15231,N_16077);
xnor U20167 (N_20167,N_16401,N_16771);
nand U20168 (N_20168,N_17825,N_16874);
nor U20169 (N_20169,N_16519,N_16046);
xor U20170 (N_20170,N_16809,N_16194);
nand U20171 (N_20171,N_16398,N_17509);
or U20172 (N_20172,N_16077,N_15593);
xnor U20173 (N_20173,N_17973,N_15108);
or U20174 (N_20174,N_16391,N_16252);
and U20175 (N_20175,N_16725,N_15286);
and U20176 (N_20176,N_17093,N_16313);
nor U20177 (N_20177,N_15414,N_15537);
and U20178 (N_20178,N_16436,N_16605);
or U20179 (N_20179,N_15767,N_16555);
nand U20180 (N_20180,N_16610,N_16162);
nor U20181 (N_20181,N_15569,N_16330);
nor U20182 (N_20182,N_16625,N_17528);
nand U20183 (N_20183,N_16435,N_16277);
or U20184 (N_20184,N_17144,N_15912);
or U20185 (N_20185,N_17508,N_16615);
xnor U20186 (N_20186,N_17110,N_16408);
and U20187 (N_20187,N_17691,N_16648);
or U20188 (N_20188,N_17050,N_16557);
nor U20189 (N_20189,N_16852,N_17502);
nor U20190 (N_20190,N_16836,N_17738);
xnor U20191 (N_20191,N_16507,N_16640);
nand U20192 (N_20192,N_15889,N_15021);
and U20193 (N_20193,N_16799,N_16740);
nand U20194 (N_20194,N_15462,N_16206);
nor U20195 (N_20195,N_17636,N_16760);
xnor U20196 (N_20196,N_16051,N_17207);
nand U20197 (N_20197,N_17757,N_16361);
nor U20198 (N_20198,N_17734,N_17599);
nand U20199 (N_20199,N_16111,N_15925);
nor U20200 (N_20200,N_17002,N_17208);
nor U20201 (N_20201,N_17001,N_15590);
and U20202 (N_20202,N_17613,N_16227);
or U20203 (N_20203,N_17168,N_17968);
nor U20204 (N_20204,N_16611,N_16761);
nor U20205 (N_20205,N_17466,N_16879);
xor U20206 (N_20206,N_15506,N_17096);
or U20207 (N_20207,N_16979,N_16981);
xor U20208 (N_20208,N_15832,N_16444);
nor U20209 (N_20209,N_15866,N_17122);
nand U20210 (N_20210,N_15946,N_16098);
nand U20211 (N_20211,N_17516,N_15790);
nand U20212 (N_20212,N_16983,N_15850);
xnor U20213 (N_20213,N_16761,N_16298);
nand U20214 (N_20214,N_15338,N_17928);
xor U20215 (N_20215,N_15802,N_16953);
nor U20216 (N_20216,N_15755,N_17589);
nor U20217 (N_20217,N_16897,N_15972);
nand U20218 (N_20218,N_17436,N_17124);
and U20219 (N_20219,N_17320,N_17681);
or U20220 (N_20220,N_15677,N_16462);
or U20221 (N_20221,N_15389,N_17246);
xnor U20222 (N_20222,N_15618,N_16224);
xor U20223 (N_20223,N_16244,N_15212);
or U20224 (N_20224,N_17321,N_15893);
nor U20225 (N_20225,N_17289,N_15408);
or U20226 (N_20226,N_16891,N_15536);
xnor U20227 (N_20227,N_15592,N_16518);
nor U20228 (N_20228,N_15711,N_17545);
and U20229 (N_20229,N_17049,N_16528);
nand U20230 (N_20230,N_15435,N_17990);
xor U20231 (N_20231,N_17065,N_16412);
or U20232 (N_20232,N_15022,N_15656);
nand U20233 (N_20233,N_17642,N_16683);
or U20234 (N_20234,N_16614,N_16952);
nor U20235 (N_20235,N_15837,N_16327);
nand U20236 (N_20236,N_17180,N_16644);
and U20237 (N_20237,N_17790,N_16110);
nor U20238 (N_20238,N_15952,N_15170);
nor U20239 (N_20239,N_17856,N_17702);
and U20240 (N_20240,N_15706,N_17274);
xor U20241 (N_20241,N_16488,N_17124);
and U20242 (N_20242,N_16399,N_15212);
xor U20243 (N_20243,N_16396,N_16471);
nor U20244 (N_20244,N_16904,N_17693);
or U20245 (N_20245,N_16198,N_17870);
xor U20246 (N_20246,N_15106,N_15874);
xor U20247 (N_20247,N_16034,N_15906);
xor U20248 (N_20248,N_15132,N_15729);
xnor U20249 (N_20249,N_16367,N_17390);
nor U20250 (N_20250,N_17264,N_15167);
nand U20251 (N_20251,N_16655,N_17414);
and U20252 (N_20252,N_15670,N_15266);
xnor U20253 (N_20253,N_16347,N_15153);
nand U20254 (N_20254,N_16998,N_17763);
nand U20255 (N_20255,N_17561,N_16870);
or U20256 (N_20256,N_15573,N_17123);
and U20257 (N_20257,N_17080,N_17078);
nor U20258 (N_20258,N_16949,N_16173);
and U20259 (N_20259,N_16412,N_17234);
nand U20260 (N_20260,N_17825,N_17537);
and U20261 (N_20261,N_16638,N_15752);
and U20262 (N_20262,N_15865,N_16450);
and U20263 (N_20263,N_16949,N_16417);
xor U20264 (N_20264,N_17377,N_16457);
xor U20265 (N_20265,N_16861,N_16384);
or U20266 (N_20266,N_17101,N_16869);
nand U20267 (N_20267,N_17127,N_16167);
and U20268 (N_20268,N_15822,N_16604);
xnor U20269 (N_20269,N_17094,N_16707);
nand U20270 (N_20270,N_16404,N_15737);
or U20271 (N_20271,N_15742,N_16294);
nor U20272 (N_20272,N_17593,N_16530);
xor U20273 (N_20273,N_16110,N_15278);
xor U20274 (N_20274,N_15592,N_17775);
and U20275 (N_20275,N_16104,N_16381);
xor U20276 (N_20276,N_17947,N_16686);
and U20277 (N_20277,N_15923,N_15289);
xnor U20278 (N_20278,N_17597,N_15543);
nand U20279 (N_20279,N_17013,N_17683);
nand U20280 (N_20280,N_16538,N_17783);
and U20281 (N_20281,N_16789,N_17377);
nor U20282 (N_20282,N_16200,N_17762);
xor U20283 (N_20283,N_17666,N_17896);
or U20284 (N_20284,N_17036,N_16409);
xnor U20285 (N_20285,N_15829,N_16011);
xnor U20286 (N_20286,N_17788,N_15301);
xor U20287 (N_20287,N_17226,N_17330);
and U20288 (N_20288,N_17239,N_17000);
and U20289 (N_20289,N_16990,N_17983);
nand U20290 (N_20290,N_17932,N_15011);
or U20291 (N_20291,N_17383,N_17678);
nor U20292 (N_20292,N_15494,N_15407);
nand U20293 (N_20293,N_16815,N_15568);
nand U20294 (N_20294,N_15590,N_15146);
and U20295 (N_20295,N_16652,N_16324);
and U20296 (N_20296,N_17482,N_17750);
and U20297 (N_20297,N_16254,N_16007);
and U20298 (N_20298,N_16455,N_16638);
nand U20299 (N_20299,N_17232,N_17057);
or U20300 (N_20300,N_15480,N_15449);
nor U20301 (N_20301,N_15366,N_16914);
nand U20302 (N_20302,N_17817,N_16718);
or U20303 (N_20303,N_17593,N_15654);
nand U20304 (N_20304,N_15058,N_15784);
or U20305 (N_20305,N_16210,N_16806);
and U20306 (N_20306,N_17776,N_16226);
xnor U20307 (N_20307,N_16400,N_16985);
nor U20308 (N_20308,N_15763,N_17197);
nor U20309 (N_20309,N_15876,N_15885);
nand U20310 (N_20310,N_15067,N_15606);
nor U20311 (N_20311,N_17637,N_16902);
nor U20312 (N_20312,N_16685,N_15080);
nor U20313 (N_20313,N_16355,N_15071);
xnor U20314 (N_20314,N_16878,N_15226);
nand U20315 (N_20315,N_16941,N_16561);
xnor U20316 (N_20316,N_16977,N_17598);
nor U20317 (N_20317,N_17295,N_15665);
or U20318 (N_20318,N_17712,N_15409);
nand U20319 (N_20319,N_17803,N_17925);
xnor U20320 (N_20320,N_16965,N_15581);
or U20321 (N_20321,N_16158,N_15752);
or U20322 (N_20322,N_16561,N_16070);
or U20323 (N_20323,N_17420,N_16405);
nand U20324 (N_20324,N_17967,N_17141);
nor U20325 (N_20325,N_15403,N_17008);
xor U20326 (N_20326,N_16051,N_17858);
and U20327 (N_20327,N_15785,N_17372);
xnor U20328 (N_20328,N_15955,N_16105);
nor U20329 (N_20329,N_17097,N_15396);
or U20330 (N_20330,N_16526,N_16662);
nand U20331 (N_20331,N_16684,N_15774);
nor U20332 (N_20332,N_16748,N_17310);
and U20333 (N_20333,N_17255,N_17854);
nand U20334 (N_20334,N_16480,N_15743);
or U20335 (N_20335,N_16049,N_16598);
nand U20336 (N_20336,N_16935,N_16506);
nor U20337 (N_20337,N_15256,N_17220);
nor U20338 (N_20338,N_15637,N_17425);
or U20339 (N_20339,N_15698,N_16442);
or U20340 (N_20340,N_17684,N_17111);
or U20341 (N_20341,N_17874,N_15002);
or U20342 (N_20342,N_17871,N_17180);
nor U20343 (N_20343,N_16479,N_15920);
nand U20344 (N_20344,N_15307,N_16173);
nor U20345 (N_20345,N_15902,N_17043);
nand U20346 (N_20346,N_16429,N_16978);
nand U20347 (N_20347,N_17870,N_17176);
and U20348 (N_20348,N_15973,N_15225);
nor U20349 (N_20349,N_17962,N_16682);
nor U20350 (N_20350,N_15879,N_17276);
or U20351 (N_20351,N_15466,N_17065);
nor U20352 (N_20352,N_16900,N_17144);
or U20353 (N_20353,N_15766,N_16384);
and U20354 (N_20354,N_15995,N_17344);
nor U20355 (N_20355,N_16058,N_15233);
xor U20356 (N_20356,N_17243,N_17929);
nor U20357 (N_20357,N_17721,N_15550);
xor U20358 (N_20358,N_17665,N_15296);
or U20359 (N_20359,N_16566,N_15564);
or U20360 (N_20360,N_16244,N_15737);
or U20361 (N_20361,N_16081,N_16751);
and U20362 (N_20362,N_15674,N_15945);
nand U20363 (N_20363,N_15439,N_15666);
or U20364 (N_20364,N_16609,N_15573);
or U20365 (N_20365,N_17519,N_17196);
nand U20366 (N_20366,N_16423,N_17065);
nor U20367 (N_20367,N_17125,N_16656);
xnor U20368 (N_20368,N_16168,N_16008);
xnor U20369 (N_20369,N_16034,N_15561);
and U20370 (N_20370,N_16186,N_15394);
nand U20371 (N_20371,N_15713,N_16276);
xor U20372 (N_20372,N_15321,N_15772);
xnor U20373 (N_20373,N_17663,N_17993);
or U20374 (N_20374,N_16585,N_16184);
and U20375 (N_20375,N_17423,N_16536);
and U20376 (N_20376,N_16621,N_15163);
nand U20377 (N_20377,N_16148,N_16781);
nand U20378 (N_20378,N_17487,N_17474);
and U20379 (N_20379,N_16055,N_16735);
xnor U20380 (N_20380,N_16116,N_15793);
and U20381 (N_20381,N_16819,N_17961);
nand U20382 (N_20382,N_15183,N_17681);
nor U20383 (N_20383,N_16876,N_16245);
and U20384 (N_20384,N_15157,N_16949);
xnor U20385 (N_20385,N_17035,N_16633);
nor U20386 (N_20386,N_16772,N_16106);
nand U20387 (N_20387,N_15517,N_17176);
nand U20388 (N_20388,N_15590,N_15857);
xor U20389 (N_20389,N_17166,N_15370);
nor U20390 (N_20390,N_17706,N_17236);
and U20391 (N_20391,N_15138,N_16933);
xor U20392 (N_20392,N_16280,N_16733);
and U20393 (N_20393,N_15895,N_17314);
or U20394 (N_20394,N_15991,N_16856);
nand U20395 (N_20395,N_15635,N_16270);
nand U20396 (N_20396,N_16542,N_17412);
xnor U20397 (N_20397,N_16777,N_16657);
nor U20398 (N_20398,N_16082,N_16133);
or U20399 (N_20399,N_16951,N_15027);
nor U20400 (N_20400,N_15560,N_15375);
nor U20401 (N_20401,N_16013,N_16566);
and U20402 (N_20402,N_17958,N_17304);
or U20403 (N_20403,N_17968,N_15288);
and U20404 (N_20404,N_16634,N_15208);
xnor U20405 (N_20405,N_15991,N_17368);
and U20406 (N_20406,N_15249,N_17655);
xor U20407 (N_20407,N_16259,N_17644);
xnor U20408 (N_20408,N_17081,N_17725);
xnor U20409 (N_20409,N_16706,N_15984);
nand U20410 (N_20410,N_15439,N_17518);
nor U20411 (N_20411,N_17435,N_15226);
nand U20412 (N_20412,N_16044,N_17953);
or U20413 (N_20413,N_16932,N_17085);
nor U20414 (N_20414,N_15933,N_17400);
or U20415 (N_20415,N_16694,N_15425);
or U20416 (N_20416,N_16463,N_15146);
and U20417 (N_20417,N_15617,N_17219);
xor U20418 (N_20418,N_16277,N_17667);
nand U20419 (N_20419,N_16901,N_17789);
xor U20420 (N_20420,N_16663,N_15461);
xor U20421 (N_20421,N_17506,N_15052);
xor U20422 (N_20422,N_15943,N_16510);
nand U20423 (N_20423,N_17340,N_15501);
xnor U20424 (N_20424,N_17258,N_16435);
xnor U20425 (N_20425,N_17661,N_16879);
or U20426 (N_20426,N_16701,N_17195);
and U20427 (N_20427,N_15426,N_16588);
xnor U20428 (N_20428,N_15940,N_17098);
nand U20429 (N_20429,N_16566,N_17721);
nand U20430 (N_20430,N_17345,N_17144);
or U20431 (N_20431,N_16909,N_15912);
nor U20432 (N_20432,N_17971,N_16770);
xor U20433 (N_20433,N_15942,N_17131);
nor U20434 (N_20434,N_17686,N_17843);
nand U20435 (N_20435,N_15597,N_15520);
nand U20436 (N_20436,N_16991,N_15210);
xnor U20437 (N_20437,N_16945,N_16234);
nor U20438 (N_20438,N_16561,N_15946);
nor U20439 (N_20439,N_17010,N_17101);
nor U20440 (N_20440,N_16771,N_16335);
or U20441 (N_20441,N_15597,N_16023);
nand U20442 (N_20442,N_16180,N_17278);
nand U20443 (N_20443,N_15773,N_17852);
and U20444 (N_20444,N_16360,N_15001);
nor U20445 (N_20445,N_17782,N_17184);
nand U20446 (N_20446,N_15537,N_17679);
nor U20447 (N_20447,N_16460,N_17790);
or U20448 (N_20448,N_17245,N_16120);
and U20449 (N_20449,N_17574,N_15247);
and U20450 (N_20450,N_17803,N_15623);
nand U20451 (N_20451,N_17784,N_17018);
xor U20452 (N_20452,N_17271,N_15762);
and U20453 (N_20453,N_15359,N_17965);
nand U20454 (N_20454,N_15162,N_17594);
or U20455 (N_20455,N_16552,N_17759);
xor U20456 (N_20456,N_17127,N_15195);
xor U20457 (N_20457,N_15016,N_16680);
xnor U20458 (N_20458,N_15569,N_17150);
nand U20459 (N_20459,N_17954,N_16820);
and U20460 (N_20460,N_15050,N_17018);
xnor U20461 (N_20461,N_17066,N_16954);
or U20462 (N_20462,N_17520,N_17591);
nor U20463 (N_20463,N_17841,N_17420);
or U20464 (N_20464,N_17676,N_17371);
and U20465 (N_20465,N_16360,N_17388);
and U20466 (N_20466,N_15472,N_16860);
nor U20467 (N_20467,N_15331,N_16509);
xor U20468 (N_20468,N_15895,N_15571);
nand U20469 (N_20469,N_16668,N_17902);
nand U20470 (N_20470,N_16942,N_16948);
or U20471 (N_20471,N_17972,N_15881);
or U20472 (N_20472,N_15125,N_16212);
nand U20473 (N_20473,N_17304,N_17707);
and U20474 (N_20474,N_16102,N_15356);
xor U20475 (N_20475,N_17200,N_15420);
or U20476 (N_20476,N_16854,N_16244);
nor U20477 (N_20477,N_16555,N_17007);
or U20478 (N_20478,N_17506,N_15154);
xor U20479 (N_20479,N_17038,N_16712);
nand U20480 (N_20480,N_15636,N_16531);
nor U20481 (N_20481,N_17343,N_15390);
or U20482 (N_20482,N_15903,N_17111);
nor U20483 (N_20483,N_17755,N_17496);
nor U20484 (N_20484,N_15568,N_16821);
and U20485 (N_20485,N_17628,N_16880);
and U20486 (N_20486,N_15728,N_16307);
xor U20487 (N_20487,N_16067,N_15548);
and U20488 (N_20488,N_17588,N_16346);
nor U20489 (N_20489,N_17422,N_17609);
and U20490 (N_20490,N_17953,N_15281);
nand U20491 (N_20491,N_17042,N_17226);
xor U20492 (N_20492,N_15897,N_16769);
or U20493 (N_20493,N_15945,N_16608);
and U20494 (N_20494,N_15267,N_15782);
and U20495 (N_20495,N_15321,N_16894);
and U20496 (N_20496,N_17959,N_16248);
or U20497 (N_20497,N_16177,N_16525);
nand U20498 (N_20498,N_17283,N_17831);
nor U20499 (N_20499,N_17567,N_17275);
and U20500 (N_20500,N_15683,N_16178);
and U20501 (N_20501,N_17453,N_15830);
nor U20502 (N_20502,N_16001,N_15482);
nand U20503 (N_20503,N_17534,N_17302);
and U20504 (N_20504,N_16317,N_15271);
nand U20505 (N_20505,N_17669,N_16252);
nand U20506 (N_20506,N_15445,N_17495);
xnor U20507 (N_20507,N_17908,N_16759);
and U20508 (N_20508,N_15046,N_15731);
xor U20509 (N_20509,N_16031,N_16059);
xor U20510 (N_20510,N_15675,N_17132);
xnor U20511 (N_20511,N_16582,N_15334);
or U20512 (N_20512,N_17891,N_17661);
nand U20513 (N_20513,N_15598,N_15138);
nand U20514 (N_20514,N_15844,N_16853);
xnor U20515 (N_20515,N_16426,N_17747);
and U20516 (N_20516,N_15962,N_15169);
and U20517 (N_20517,N_16866,N_17800);
and U20518 (N_20518,N_15172,N_17468);
xor U20519 (N_20519,N_16919,N_17321);
nor U20520 (N_20520,N_16207,N_17342);
xnor U20521 (N_20521,N_17624,N_17547);
nor U20522 (N_20522,N_15896,N_15401);
nor U20523 (N_20523,N_15591,N_15882);
nand U20524 (N_20524,N_17757,N_16763);
or U20525 (N_20525,N_17370,N_15939);
nor U20526 (N_20526,N_15438,N_16179);
and U20527 (N_20527,N_15972,N_17704);
or U20528 (N_20528,N_16474,N_15914);
xor U20529 (N_20529,N_15999,N_16500);
or U20530 (N_20530,N_17479,N_17575);
or U20531 (N_20531,N_15540,N_17330);
nand U20532 (N_20532,N_16981,N_15996);
nor U20533 (N_20533,N_17527,N_17856);
or U20534 (N_20534,N_16907,N_17299);
or U20535 (N_20535,N_15323,N_16459);
xor U20536 (N_20536,N_17946,N_16397);
or U20537 (N_20537,N_17634,N_17418);
nand U20538 (N_20538,N_17726,N_15033);
nor U20539 (N_20539,N_15589,N_16792);
nand U20540 (N_20540,N_15518,N_15285);
nand U20541 (N_20541,N_15665,N_17939);
xor U20542 (N_20542,N_16007,N_16340);
and U20543 (N_20543,N_15824,N_17643);
nand U20544 (N_20544,N_15123,N_16401);
and U20545 (N_20545,N_16050,N_16398);
nor U20546 (N_20546,N_15578,N_15188);
and U20547 (N_20547,N_16852,N_17794);
nor U20548 (N_20548,N_16310,N_17273);
nor U20549 (N_20549,N_15247,N_17049);
or U20550 (N_20550,N_17124,N_16833);
xnor U20551 (N_20551,N_16609,N_16602);
xnor U20552 (N_20552,N_16880,N_16128);
and U20553 (N_20553,N_16203,N_16917);
and U20554 (N_20554,N_17721,N_17402);
xor U20555 (N_20555,N_15403,N_15169);
nand U20556 (N_20556,N_16908,N_15541);
and U20557 (N_20557,N_15870,N_17424);
nand U20558 (N_20558,N_17494,N_16729);
or U20559 (N_20559,N_16850,N_16660);
and U20560 (N_20560,N_17966,N_17687);
nor U20561 (N_20561,N_15857,N_15826);
or U20562 (N_20562,N_16235,N_16708);
or U20563 (N_20563,N_15661,N_16841);
or U20564 (N_20564,N_15643,N_17729);
and U20565 (N_20565,N_17623,N_17778);
nor U20566 (N_20566,N_16304,N_16338);
or U20567 (N_20567,N_16377,N_17618);
xnor U20568 (N_20568,N_16979,N_15410);
nand U20569 (N_20569,N_16436,N_17133);
and U20570 (N_20570,N_17034,N_16461);
xor U20571 (N_20571,N_16239,N_17707);
nand U20572 (N_20572,N_15903,N_15923);
nand U20573 (N_20573,N_15553,N_15632);
nand U20574 (N_20574,N_17176,N_16872);
nor U20575 (N_20575,N_16228,N_17141);
xnor U20576 (N_20576,N_17385,N_17513);
nand U20577 (N_20577,N_16680,N_16892);
xnor U20578 (N_20578,N_17662,N_17307);
nor U20579 (N_20579,N_15628,N_15087);
and U20580 (N_20580,N_15877,N_15554);
nor U20581 (N_20581,N_16537,N_17651);
nor U20582 (N_20582,N_15948,N_15248);
and U20583 (N_20583,N_15847,N_15734);
nor U20584 (N_20584,N_16803,N_17068);
nor U20585 (N_20585,N_17623,N_17774);
and U20586 (N_20586,N_17268,N_17668);
and U20587 (N_20587,N_15350,N_17155);
or U20588 (N_20588,N_15105,N_15121);
or U20589 (N_20589,N_16122,N_15009);
xor U20590 (N_20590,N_16897,N_16216);
nand U20591 (N_20591,N_16916,N_15642);
or U20592 (N_20592,N_15729,N_17095);
and U20593 (N_20593,N_16800,N_17529);
nand U20594 (N_20594,N_15653,N_15949);
or U20595 (N_20595,N_16704,N_15079);
xnor U20596 (N_20596,N_17794,N_15694);
and U20597 (N_20597,N_15209,N_17221);
or U20598 (N_20598,N_17349,N_17180);
nand U20599 (N_20599,N_17958,N_17650);
nor U20600 (N_20600,N_15791,N_16939);
nand U20601 (N_20601,N_15170,N_16502);
nand U20602 (N_20602,N_16439,N_15427);
and U20603 (N_20603,N_17792,N_17357);
and U20604 (N_20604,N_15106,N_17615);
nor U20605 (N_20605,N_17452,N_17492);
and U20606 (N_20606,N_16899,N_17581);
xor U20607 (N_20607,N_15823,N_15167);
xnor U20608 (N_20608,N_17539,N_17758);
and U20609 (N_20609,N_15766,N_15174);
nor U20610 (N_20610,N_15832,N_16059);
or U20611 (N_20611,N_15625,N_16381);
nand U20612 (N_20612,N_15365,N_16972);
nor U20613 (N_20613,N_16745,N_17312);
or U20614 (N_20614,N_16776,N_15979);
xnor U20615 (N_20615,N_15124,N_15032);
nand U20616 (N_20616,N_17320,N_15169);
or U20617 (N_20617,N_16552,N_15601);
and U20618 (N_20618,N_15533,N_15126);
nor U20619 (N_20619,N_16947,N_17688);
nor U20620 (N_20620,N_17771,N_17829);
or U20621 (N_20621,N_16471,N_17499);
or U20622 (N_20622,N_15156,N_15424);
nand U20623 (N_20623,N_17889,N_16077);
xnor U20624 (N_20624,N_17274,N_16950);
nand U20625 (N_20625,N_16980,N_17410);
or U20626 (N_20626,N_16541,N_17186);
xnor U20627 (N_20627,N_17417,N_15417);
xnor U20628 (N_20628,N_16834,N_15430);
xnor U20629 (N_20629,N_17816,N_17995);
or U20630 (N_20630,N_16466,N_15865);
nand U20631 (N_20631,N_17168,N_17655);
or U20632 (N_20632,N_16104,N_15341);
nand U20633 (N_20633,N_15003,N_17216);
and U20634 (N_20634,N_16679,N_15430);
xor U20635 (N_20635,N_17056,N_16055);
nand U20636 (N_20636,N_17085,N_17022);
xor U20637 (N_20637,N_17747,N_17206);
or U20638 (N_20638,N_17280,N_17988);
or U20639 (N_20639,N_15817,N_16520);
xor U20640 (N_20640,N_16272,N_16259);
nor U20641 (N_20641,N_17959,N_15743);
or U20642 (N_20642,N_17621,N_15691);
nor U20643 (N_20643,N_17884,N_17489);
xnor U20644 (N_20644,N_17039,N_16655);
xnor U20645 (N_20645,N_16177,N_15671);
nand U20646 (N_20646,N_17742,N_17984);
nand U20647 (N_20647,N_15426,N_15944);
nor U20648 (N_20648,N_16808,N_17452);
nand U20649 (N_20649,N_16417,N_17240);
nor U20650 (N_20650,N_15400,N_15831);
xor U20651 (N_20651,N_15813,N_16644);
or U20652 (N_20652,N_16648,N_17922);
and U20653 (N_20653,N_15757,N_15447);
xor U20654 (N_20654,N_17368,N_17158);
or U20655 (N_20655,N_17247,N_16555);
and U20656 (N_20656,N_17792,N_15018);
xor U20657 (N_20657,N_17208,N_16845);
xor U20658 (N_20658,N_15403,N_16682);
and U20659 (N_20659,N_16586,N_17086);
nand U20660 (N_20660,N_15933,N_17737);
xor U20661 (N_20661,N_17929,N_15753);
nand U20662 (N_20662,N_17558,N_16289);
or U20663 (N_20663,N_17982,N_17119);
xor U20664 (N_20664,N_17065,N_17041);
nor U20665 (N_20665,N_15612,N_16233);
nor U20666 (N_20666,N_15270,N_15447);
and U20667 (N_20667,N_17307,N_16717);
and U20668 (N_20668,N_16642,N_15819);
nand U20669 (N_20669,N_17373,N_17751);
xnor U20670 (N_20670,N_17755,N_16213);
xor U20671 (N_20671,N_17837,N_15806);
nor U20672 (N_20672,N_15989,N_16506);
nor U20673 (N_20673,N_16845,N_17953);
nor U20674 (N_20674,N_16848,N_15967);
nand U20675 (N_20675,N_16658,N_15399);
and U20676 (N_20676,N_16407,N_15021);
and U20677 (N_20677,N_16330,N_16263);
xor U20678 (N_20678,N_16611,N_17363);
or U20679 (N_20679,N_16847,N_16729);
nor U20680 (N_20680,N_16528,N_15826);
nor U20681 (N_20681,N_15885,N_15171);
or U20682 (N_20682,N_16962,N_15565);
nor U20683 (N_20683,N_15865,N_17258);
nor U20684 (N_20684,N_16359,N_15463);
nor U20685 (N_20685,N_16134,N_15885);
and U20686 (N_20686,N_15201,N_17071);
or U20687 (N_20687,N_15255,N_15456);
nand U20688 (N_20688,N_17785,N_16595);
nand U20689 (N_20689,N_15600,N_15221);
nor U20690 (N_20690,N_17572,N_15473);
or U20691 (N_20691,N_15213,N_17236);
xor U20692 (N_20692,N_15021,N_16868);
xnor U20693 (N_20693,N_15262,N_15756);
nor U20694 (N_20694,N_15173,N_17642);
xor U20695 (N_20695,N_16856,N_16187);
nand U20696 (N_20696,N_17464,N_16846);
and U20697 (N_20697,N_16866,N_16128);
and U20698 (N_20698,N_15556,N_16644);
xnor U20699 (N_20699,N_17717,N_15671);
xnor U20700 (N_20700,N_17806,N_15851);
xor U20701 (N_20701,N_17422,N_17717);
or U20702 (N_20702,N_16148,N_16094);
nand U20703 (N_20703,N_16331,N_16525);
nand U20704 (N_20704,N_17109,N_15353);
nor U20705 (N_20705,N_15747,N_16530);
xnor U20706 (N_20706,N_15861,N_17260);
and U20707 (N_20707,N_15608,N_15266);
xnor U20708 (N_20708,N_17462,N_15459);
nor U20709 (N_20709,N_17884,N_16130);
nand U20710 (N_20710,N_16355,N_17701);
nor U20711 (N_20711,N_16100,N_15786);
and U20712 (N_20712,N_15154,N_16852);
and U20713 (N_20713,N_17130,N_15373);
nand U20714 (N_20714,N_17956,N_16054);
or U20715 (N_20715,N_15992,N_15045);
or U20716 (N_20716,N_17837,N_16771);
xor U20717 (N_20717,N_16799,N_16922);
xor U20718 (N_20718,N_17512,N_16746);
nand U20719 (N_20719,N_17879,N_15842);
xor U20720 (N_20720,N_16386,N_15730);
or U20721 (N_20721,N_17752,N_15492);
xnor U20722 (N_20722,N_17683,N_16269);
and U20723 (N_20723,N_17428,N_17534);
or U20724 (N_20724,N_15150,N_15908);
nor U20725 (N_20725,N_15573,N_17284);
nand U20726 (N_20726,N_17594,N_17935);
xor U20727 (N_20727,N_17424,N_16131);
nor U20728 (N_20728,N_17733,N_16890);
nor U20729 (N_20729,N_15120,N_17079);
nor U20730 (N_20730,N_16661,N_16752);
nand U20731 (N_20731,N_15084,N_17992);
and U20732 (N_20732,N_17437,N_15198);
or U20733 (N_20733,N_16854,N_17053);
and U20734 (N_20734,N_17516,N_17435);
xnor U20735 (N_20735,N_17428,N_16494);
xor U20736 (N_20736,N_16410,N_15686);
or U20737 (N_20737,N_15310,N_16633);
or U20738 (N_20738,N_15365,N_17823);
or U20739 (N_20739,N_16268,N_16451);
xnor U20740 (N_20740,N_17032,N_15049);
and U20741 (N_20741,N_16040,N_15793);
nor U20742 (N_20742,N_15763,N_16016);
nand U20743 (N_20743,N_16593,N_15063);
nor U20744 (N_20744,N_15731,N_17196);
and U20745 (N_20745,N_16837,N_16546);
and U20746 (N_20746,N_17999,N_16757);
xnor U20747 (N_20747,N_15178,N_16304);
and U20748 (N_20748,N_15513,N_17789);
xnor U20749 (N_20749,N_16169,N_17828);
xnor U20750 (N_20750,N_15311,N_16400);
nand U20751 (N_20751,N_16682,N_17297);
nand U20752 (N_20752,N_17821,N_16418);
and U20753 (N_20753,N_16402,N_17684);
nand U20754 (N_20754,N_15425,N_15468);
or U20755 (N_20755,N_16323,N_17813);
nor U20756 (N_20756,N_16797,N_15786);
xnor U20757 (N_20757,N_15680,N_17612);
nand U20758 (N_20758,N_16528,N_17667);
xor U20759 (N_20759,N_15227,N_15500);
nor U20760 (N_20760,N_16048,N_16173);
nor U20761 (N_20761,N_17422,N_17092);
nand U20762 (N_20762,N_15569,N_15897);
nor U20763 (N_20763,N_17835,N_17580);
and U20764 (N_20764,N_16283,N_17999);
and U20765 (N_20765,N_17526,N_16496);
xnor U20766 (N_20766,N_15589,N_17472);
nand U20767 (N_20767,N_17824,N_15465);
nor U20768 (N_20768,N_16913,N_16316);
and U20769 (N_20769,N_16723,N_17231);
xnor U20770 (N_20770,N_17445,N_16956);
nor U20771 (N_20771,N_16050,N_16672);
and U20772 (N_20772,N_16373,N_16756);
nor U20773 (N_20773,N_17782,N_16660);
and U20774 (N_20774,N_16786,N_17920);
nor U20775 (N_20775,N_15967,N_15143);
or U20776 (N_20776,N_15162,N_16363);
xnor U20777 (N_20777,N_16583,N_16163);
nand U20778 (N_20778,N_17267,N_15653);
xnor U20779 (N_20779,N_17546,N_15988);
nand U20780 (N_20780,N_17728,N_17082);
and U20781 (N_20781,N_15725,N_15580);
nor U20782 (N_20782,N_15096,N_15368);
and U20783 (N_20783,N_17466,N_17861);
nor U20784 (N_20784,N_16031,N_15516);
nor U20785 (N_20785,N_15995,N_15106);
nand U20786 (N_20786,N_17525,N_15609);
and U20787 (N_20787,N_15775,N_16684);
nor U20788 (N_20788,N_16123,N_17332);
and U20789 (N_20789,N_17079,N_16634);
or U20790 (N_20790,N_15320,N_15072);
and U20791 (N_20791,N_15728,N_16549);
and U20792 (N_20792,N_16144,N_17842);
nor U20793 (N_20793,N_17199,N_16332);
nand U20794 (N_20794,N_17706,N_17458);
nor U20795 (N_20795,N_17813,N_15930);
or U20796 (N_20796,N_15782,N_17285);
nand U20797 (N_20797,N_16826,N_17321);
nor U20798 (N_20798,N_15523,N_16668);
or U20799 (N_20799,N_15013,N_17992);
nand U20800 (N_20800,N_15274,N_17206);
and U20801 (N_20801,N_16474,N_15000);
nor U20802 (N_20802,N_15736,N_16951);
nand U20803 (N_20803,N_15708,N_15956);
or U20804 (N_20804,N_17460,N_16126);
or U20805 (N_20805,N_15162,N_15713);
xor U20806 (N_20806,N_16970,N_16183);
nand U20807 (N_20807,N_15812,N_16117);
and U20808 (N_20808,N_17493,N_17208);
nand U20809 (N_20809,N_15973,N_16458);
nor U20810 (N_20810,N_16624,N_16241);
nand U20811 (N_20811,N_15560,N_17134);
nand U20812 (N_20812,N_16294,N_16064);
nand U20813 (N_20813,N_15650,N_17324);
xnor U20814 (N_20814,N_16149,N_17532);
xnor U20815 (N_20815,N_15136,N_17809);
or U20816 (N_20816,N_17292,N_17112);
nand U20817 (N_20817,N_16036,N_17418);
nand U20818 (N_20818,N_16816,N_17137);
nand U20819 (N_20819,N_16894,N_16037);
xnor U20820 (N_20820,N_15912,N_17223);
or U20821 (N_20821,N_15302,N_15583);
nor U20822 (N_20822,N_16600,N_16241);
and U20823 (N_20823,N_15039,N_16479);
nand U20824 (N_20824,N_16828,N_17256);
xnor U20825 (N_20825,N_17030,N_17321);
and U20826 (N_20826,N_16314,N_17222);
nor U20827 (N_20827,N_15178,N_17113);
xnor U20828 (N_20828,N_16231,N_15031);
and U20829 (N_20829,N_15602,N_15087);
nor U20830 (N_20830,N_15620,N_15612);
or U20831 (N_20831,N_16990,N_16644);
or U20832 (N_20832,N_15136,N_17401);
nand U20833 (N_20833,N_17465,N_17369);
nor U20834 (N_20834,N_17113,N_16044);
or U20835 (N_20835,N_17141,N_16579);
xor U20836 (N_20836,N_17282,N_17363);
xnor U20837 (N_20837,N_15112,N_17417);
or U20838 (N_20838,N_17974,N_17156);
and U20839 (N_20839,N_15902,N_16547);
nor U20840 (N_20840,N_17034,N_16526);
nor U20841 (N_20841,N_16544,N_15060);
xnor U20842 (N_20842,N_15824,N_16213);
and U20843 (N_20843,N_17558,N_15039);
xnor U20844 (N_20844,N_17162,N_17878);
and U20845 (N_20845,N_16330,N_15791);
or U20846 (N_20846,N_16172,N_17961);
nor U20847 (N_20847,N_16757,N_17916);
xor U20848 (N_20848,N_15262,N_16683);
nor U20849 (N_20849,N_16078,N_16729);
xor U20850 (N_20850,N_17975,N_17285);
nand U20851 (N_20851,N_16288,N_16077);
nand U20852 (N_20852,N_15204,N_16052);
xor U20853 (N_20853,N_16041,N_16610);
nor U20854 (N_20854,N_16427,N_17462);
xor U20855 (N_20855,N_16933,N_17667);
nand U20856 (N_20856,N_16517,N_17131);
xor U20857 (N_20857,N_15748,N_15092);
nand U20858 (N_20858,N_17713,N_16361);
or U20859 (N_20859,N_16397,N_15032);
or U20860 (N_20860,N_16300,N_17779);
nor U20861 (N_20861,N_17479,N_16744);
nor U20862 (N_20862,N_15866,N_17864);
and U20863 (N_20863,N_17887,N_15827);
and U20864 (N_20864,N_17777,N_16530);
and U20865 (N_20865,N_15874,N_16012);
nand U20866 (N_20866,N_15871,N_15551);
and U20867 (N_20867,N_15010,N_17980);
nand U20868 (N_20868,N_15686,N_15492);
and U20869 (N_20869,N_15007,N_17137);
nand U20870 (N_20870,N_16740,N_16514);
nand U20871 (N_20871,N_16241,N_15140);
or U20872 (N_20872,N_15272,N_16497);
xor U20873 (N_20873,N_15977,N_15402);
nor U20874 (N_20874,N_16700,N_16009);
or U20875 (N_20875,N_16567,N_17076);
and U20876 (N_20876,N_15958,N_17250);
xor U20877 (N_20877,N_16308,N_16507);
or U20878 (N_20878,N_17350,N_16346);
nand U20879 (N_20879,N_16325,N_17858);
nand U20880 (N_20880,N_17404,N_16469);
xnor U20881 (N_20881,N_17179,N_16659);
and U20882 (N_20882,N_15314,N_15746);
nand U20883 (N_20883,N_15732,N_17955);
and U20884 (N_20884,N_17798,N_17968);
or U20885 (N_20885,N_17026,N_16714);
nand U20886 (N_20886,N_16223,N_15400);
nand U20887 (N_20887,N_15545,N_16649);
nor U20888 (N_20888,N_17356,N_17023);
nor U20889 (N_20889,N_15414,N_15686);
and U20890 (N_20890,N_16695,N_15026);
nand U20891 (N_20891,N_17921,N_15027);
or U20892 (N_20892,N_15854,N_17824);
or U20893 (N_20893,N_16475,N_16394);
and U20894 (N_20894,N_17032,N_15530);
or U20895 (N_20895,N_15818,N_15867);
nor U20896 (N_20896,N_15722,N_17953);
or U20897 (N_20897,N_17456,N_17913);
or U20898 (N_20898,N_16302,N_17904);
nand U20899 (N_20899,N_16057,N_15432);
xnor U20900 (N_20900,N_17378,N_15057);
nor U20901 (N_20901,N_17269,N_16374);
nor U20902 (N_20902,N_15172,N_15849);
and U20903 (N_20903,N_17396,N_15944);
or U20904 (N_20904,N_15489,N_17540);
nand U20905 (N_20905,N_15391,N_16993);
nor U20906 (N_20906,N_16379,N_17953);
and U20907 (N_20907,N_17351,N_15996);
nor U20908 (N_20908,N_16255,N_17070);
and U20909 (N_20909,N_17097,N_15848);
nor U20910 (N_20910,N_16384,N_15442);
nor U20911 (N_20911,N_17837,N_16379);
and U20912 (N_20912,N_15912,N_15701);
or U20913 (N_20913,N_16500,N_17709);
and U20914 (N_20914,N_16603,N_15098);
xnor U20915 (N_20915,N_17464,N_15983);
xnor U20916 (N_20916,N_17011,N_16768);
and U20917 (N_20917,N_17345,N_15995);
nand U20918 (N_20918,N_17142,N_16152);
and U20919 (N_20919,N_16007,N_16128);
nand U20920 (N_20920,N_17667,N_15368);
xor U20921 (N_20921,N_15820,N_16809);
nor U20922 (N_20922,N_16928,N_15084);
nor U20923 (N_20923,N_16258,N_16470);
xor U20924 (N_20924,N_16391,N_15205);
nand U20925 (N_20925,N_16197,N_17989);
or U20926 (N_20926,N_17767,N_15577);
or U20927 (N_20927,N_16948,N_15821);
or U20928 (N_20928,N_15787,N_16044);
nand U20929 (N_20929,N_16055,N_15746);
xor U20930 (N_20930,N_17870,N_15569);
and U20931 (N_20931,N_17501,N_17776);
and U20932 (N_20932,N_16790,N_17075);
and U20933 (N_20933,N_17058,N_16883);
nor U20934 (N_20934,N_16229,N_16300);
nand U20935 (N_20935,N_16301,N_17136);
or U20936 (N_20936,N_17343,N_15965);
and U20937 (N_20937,N_15151,N_17101);
or U20938 (N_20938,N_16854,N_16151);
nor U20939 (N_20939,N_15087,N_16127);
xor U20940 (N_20940,N_17003,N_15786);
or U20941 (N_20941,N_16584,N_17892);
or U20942 (N_20942,N_17392,N_17033);
xnor U20943 (N_20943,N_17241,N_17697);
nor U20944 (N_20944,N_15765,N_15566);
nand U20945 (N_20945,N_15252,N_16260);
xnor U20946 (N_20946,N_15137,N_17857);
xor U20947 (N_20947,N_16068,N_15790);
and U20948 (N_20948,N_16554,N_17909);
nor U20949 (N_20949,N_16224,N_16103);
and U20950 (N_20950,N_15084,N_17951);
or U20951 (N_20951,N_16225,N_15500);
nor U20952 (N_20952,N_17241,N_16830);
and U20953 (N_20953,N_15064,N_16309);
nor U20954 (N_20954,N_17831,N_15792);
and U20955 (N_20955,N_15967,N_16404);
and U20956 (N_20956,N_15676,N_16527);
and U20957 (N_20957,N_16341,N_15229);
nand U20958 (N_20958,N_15787,N_15348);
and U20959 (N_20959,N_16735,N_16106);
nand U20960 (N_20960,N_17424,N_16103);
xnor U20961 (N_20961,N_17133,N_16137);
nand U20962 (N_20962,N_16165,N_17001);
nand U20963 (N_20963,N_15418,N_17997);
and U20964 (N_20964,N_17135,N_17957);
nor U20965 (N_20965,N_17082,N_17140);
or U20966 (N_20966,N_17050,N_16026);
or U20967 (N_20967,N_15117,N_17820);
or U20968 (N_20968,N_17899,N_17278);
xnor U20969 (N_20969,N_15200,N_16166);
nand U20970 (N_20970,N_17332,N_17254);
nand U20971 (N_20971,N_15516,N_15257);
xnor U20972 (N_20972,N_17542,N_17649);
nor U20973 (N_20973,N_16419,N_17271);
and U20974 (N_20974,N_15647,N_16990);
nand U20975 (N_20975,N_15193,N_17242);
and U20976 (N_20976,N_17669,N_17381);
or U20977 (N_20977,N_17622,N_16076);
or U20978 (N_20978,N_15616,N_15194);
nand U20979 (N_20979,N_16568,N_16565);
and U20980 (N_20980,N_17958,N_17723);
or U20981 (N_20981,N_15214,N_17232);
or U20982 (N_20982,N_15882,N_15563);
or U20983 (N_20983,N_16278,N_17554);
nand U20984 (N_20984,N_16561,N_16838);
and U20985 (N_20985,N_16753,N_15769);
and U20986 (N_20986,N_16125,N_17956);
nor U20987 (N_20987,N_17000,N_16012);
xor U20988 (N_20988,N_17127,N_17172);
nand U20989 (N_20989,N_15143,N_15314);
or U20990 (N_20990,N_16098,N_16794);
xnor U20991 (N_20991,N_17112,N_17234);
nor U20992 (N_20992,N_17184,N_17680);
nand U20993 (N_20993,N_16235,N_15767);
or U20994 (N_20994,N_16062,N_15496);
nor U20995 (N_20995,N_17322,N_17173);
nand U20996 (N_20996,N_15598,N_15893);
and U20997 (N_20997,N_16552,N_15108);
xnor U20998 (N_20998,N_15808,N_17439);
xor U20999 (N_20999,N_15125,N_17608);
and U21000 (N_21000,N_18103,N_18039);
nand U21001 (N_21001,N_19190,N_19885);
xnor U21002 (N_21002,N_18737,N_19102);
nand U21003 (N_21003,N_20557,N_18053);
or U21004 (N_21004,N_18303,N_18160);
xor U21005 (N_21005,N_19693,N_18150);
or U21006 (N_21006,N_20031,N_20820);
and U21007 (N_21007,N_19501,N_18345);
or U21008 (N_21008,N_20607,N_18609);
nand U21009 (N_21009,N_19762,N_20996);
or U21010 (N_21010,N_20774,N_19840);
nor U21011 (N_21011,N_20162,N_19870);
nor U21012 (N_21012,N_19780,N_19775);
or U21013 (N_21013,N_20102,N_19084);
or U21014 (N_21014,N_19291,N_20450);
or U21015 (N_21015,N_19467,N_19619);
and U21016 (N_21016,N_19558,N_18661);
nand U21017 (N_21017,N_18066,N_18251);
nor U21018 (N_21018,N_18229,N_19822);
and U21019 (N_21019,N_20616,N_18076);
and U21020 (N_21020,N_20794,N_20378);
nand U21021 (N_21021,N_18439,N_19782);
and U21022 (N_21022,N_19734,N_20214);
and U21023 (N_21023,N_19400,N_20166);
nand U21024 (N_21024,N_18391,N_20491);
or U21025 (N_21025,N_18759,N_19014);
or U21026 (N_21026,N_20165,N_20237);
nor U21027 (N_21027,N_18557,N_18811);
xor U21028 (N_21028,N_19614,N_20457);
nor U21029 (N_21029,N_20662,N_18402);
or U21030 (N_21030,N_18506,N_20984);
nor U21031 (N_21031,N_18443,N_20257);
or U21032 (N_21032,N_20228,N_20098);
and U21033 (N_21033,N_19224,N_19328);
or U21034 (N_21034,N_19142,N_19674);
nor U21035 (N_21035,N_18314,N_20970);
and U21036 (N_21036,N_20396,N_20928);
nor U21037 (N_21037,N_20184,N_20028);
nor U21038 (N_21038,N_20536,N_18952);
nor U21039 (N_21039,N_20534,N_18726);
xor U21040 (N_21040,N_20916,N_20974);
and U21041 (N_21041,N_19903,N_20387);
nand U21042 (N_21042,N_19069,N_19237);
and U21043 (N_21043,N_18179,N_18429);
nand U21044 (N_21044,N_19352,N_19834);
and U21045 (N_21045,N_18889,N_20760);
nand U21046 (N_21046,N_19108,N_20007);
or U21047 (N_21047,N_20138,N_18919);
or U21048 (N_21048,N_18285,N_18264);
nor U21049 (N_21049,N_18817,N_20330);
nand U21050 (N_21050,N_20555,N_18754);
xor U21051 (N_21051,N_20510,N_18398);
nor U21052 (N_21052,N_19781,N_19563);
nor U21053 (N_21053,N_20342,N_19138);
xor U21054 (N_21054,N_20122,N_18981);
nor U21055 (N_21055,N_20883,N_20005);
nor U21056 (N_21056,N_19180,N_19009);
xor U21057 (N_21057,N_18549,N_20741);
or U21058 (N_21058,N_19523,N_19499);
nand U21059 (N_21059,N_20596,N_18756);
nor U21060 (N_21060,N_18108,N_18680);
or U21061 (N_21061,N_19880,N_20965);
or U21062 (N_21062,N_20952,N_20525);
xnor U21063 (N_21063,N_20429,N_19074);
or U21064 (N_21064,N_19318,N_20010);
and U21065 (N_21065,N_18449,N_20282);
nand U21066 (N_21066,N_18579,N_18789);
nand U21067 (N_21067,N_19412,N_19613);
or U21068 (N_21068,N_18724,N_18115);
or U21069 (N_21069,N_18276,N_19065);
nand U21070 (N_21070,N_19347,N_20989);
or U21071 (N_21071,N_19493,N_20489);
nand U21072 (N_21072,N_20754,N_20658);
xnor U21073 (N_21073,N_20068,N_20971);
xnor U21074 (N_21074,N_18640,N_19123);
xnor U21075 (N_21075,N_18750,N_19199);
nand U21076 (N_21076,N_18050,N_20905);
or U21077 (N_21077,N_19383,N_19579);
nor U21078 (N_21078,N_19437,N_20030);
xor U21079 (N_21079,N_19882,N_18931);
and U21080 (N_21080,N_19802,N_19760);
or U21081 (N_21081,N_20393,N_19238);
xnor U21082 (N_21082,N_18036,N_20618);
nor U21083 (N_21083,N_20594,N_18797);
nand U21084 (N_21084,N_19496,N_19322);
xor U21085 (N_21085,N_18232,N_19092);
and U21086 (N_21086,N_19675,N_18929);
nor U21087 (N_21087,N_19557,N_20020);
xnor U21088 (N_21088,N_19958,N_18978);
nand U21089 (N_21089,N_20535,N_20561);
nor U21090 (N_21090,N_18798,N_19485);
nand U21091 (N_21091,N_19051,N_20983);
nor U21092 (N_21092,N_19677,N_18683);
and U21093 (N_21093,N_18823,N_18074);
and U21094 (N_21094,N_19228,N_20035);
or U21095 (N_21095,N_20145,N_19505);
nor U21096 (N_21096,N_18942,N_19214);
xnor U21097 (N_21097,N_20714,N_18643);
and U21098 (N_21098,N_19171,N_18589);
nor U21099 (N_21099,N_19964,N_20551);
nand U21100 (N_21100,N_19516,N_18832);
xor U21101 (N_21101,N_18484,N_20625);
and U21102 (N_21102,N_19995,N_20968);
and U21103 (N_21103,N_20933,N_20624);
nand U21104 (N_21104,N_18227,N_18930);
or U21105 (N_21105,N_20384,N_18564);
nor U21106 (N_21106,N_20829,N_18289);
nor U21107 (N_21107,N_20982,N_20261);
nand U21108 (N_21108,N_18511,N_20372);
nand U21109 (N_21109,N_20630,N_19386);
nor U21110 (N_21110,N_19810,N_18901);
xnor U21111 (N_21111,N_19332,N_20918);
xor U21112 (N_21112,N_20783,N_19210);
or U21113 (N_21113,N_20921,N_18497);
nand U21114 (N_21114,N_18524,N_20678);
and U21115 (N_21115,N_18476,N_18025);
and U21116 (N_21116,N_19312,N_18385);
or U21117 (N_21117,N_19284,N_18733);
xor U21118 (N_21118,N_20546,N_19152);
or U21119 (N_21119,N_18051,N_18732);
xor U21120 (N_21120,N_18461,N_18877);
nand U21121 (N_21121,N_18742,N_20067);
nand U21122 (N_21122,N_19444,N_19851);
xor U21123 (N_21123,N_19435,N_18153);
nand U21124 (N_21124,N_19181,N_18453);
or U21125 (N_21125,N_19307,N_18745);
xnor U21126 (N_21126,N_19356,N_18651);
and U21127 (N_21127,N_18447,N_19226);
or U21128 (N_21128,N_18711,N_18793);
xnor U21129 (N_21129,N_20558,N_18974);
or U21130 (N_21130,N_18093,N_20744);
or U21131 (N_21131,N_20338,N_18863);
and U21132 (N_21132,N_18090,N_20549);
nor U21133 (N_21133,N_20751,N_20591);
nand U21134 (N_21134,N_20705,N_18342);
and U21135 (N_21135,N_19543,N_19567);
and U21136 (N_21136,N_20115,N_18715);
or U21137 (N_21137,N_20963,N_19776);
and U21138 (N_21138,N_18613,N_18082);
or U21139 (N_21139,N_18917,N_18202);
nor U21140 (N_21140,N_18329,N_19304);
and U21141 (N_21141,N_18037,N_18184);
or U21142 (N_21142,N_19736,N_19542);
nand U21143 (N_21143,N_19119,N_20936);
nand U21144 (N_21144,N_19861,N_19537);
nor U21145 (N_21145,N_20483,N_19263);
or U21146 (N_21146,N_18464,N_18213);
and U21147 (N_21147,N_18922,N_18309);
nor U21148 (N_21148,N_20879,N_20268);
nor U21149 (N_21149,N_20542,N_20692);
or U21150 (N_21150,N_20071,N_18993);
nand U21151 (N_21151,N_19478,N_20127);
and U21152 (N_21152,N_20740,N_20422);
and U21153 (N_21153,N_20597,N_20888);
or U21154 (N_21154,N_18915,N_18809);
nor U21155 (N_21155,N_19276,N_18189);
nand U21156 (N_21156,N_19544,N_18801);
or U21157 (N_21157,N_20109,N_18512);
nor U21158 (N_21158,N_20926,N_18923);
or U21159 (N_21159,N_18158,N_19118);
and U21160 (N_21160,N_19739,N_18765);
nand U21161 (N_21161,N_19256,N_20836);
or U21162 (N_21162,N_18344,N_19551);
nand U21163 (N_21163,N_19218,N_19770);
nor U21164 (N_21164,N_19335,N_18525);
and U21165 (N_21165,N_20240,N_19745);
nand U21166 (N_21166,N_18538,N_18070);
and U21167 (N_21167,N_18253,N_18011);
xnor U21168 (N_21168,N_19044,N_18612);
or U21169 (N_21169,N_19716,N_18768);
xnor U21170 (N_21170,N_18846,N_18162);
or U21171 (N_21171,N_18723,N_19337);
xnor U21172 (N_21172,N_19932,N_19911);
nand U21173 (N_21173,N_20685,N_19592);
nor U21174 (N_21174,N_18106,N_20840);
xor U21175 (N_21175,N_20497,N_19906);
or U21176 (N_21176,N_19589,N_20275);
xnor U21177 (N_21177,N_19868,N_18426);
xnor U21178 (N_21178,N_19758,N_20648);
nor U21179 (N_21179,N_19003,N_20684);
nand U21180 (N_21180,N_18654,N_20395);
nor U21181 (N_21181,N_19225,N_18495);
and U21182 (N_21182,N_19990,N_18896);
nand U21183 (N_21183,N_20319,N_20503);
nand U21184 (N_21184,N_19007,N_20643);
or U21185 (N_21185,N_19919,N_18941);
nor U21186 (N_21186,N_20262,N_19659);
and U21187 (N_21187,N_18337,N_20391);
nand U21188 (N_21188,N_18933,N_18294);
nor U21189 (N_21189,N_18097,N_19380);
or U21190 (N_21190,N_19853,N_19524);
nand U21191 (N_21191,N_18433,N_20215);
nor U21192 (N_21192,N_18114,N_18825);
and U21193 (N_21193,N_19683,N_20801);
nor U21194 (N_21194,N_20107,N_18033);
nor U21195 (N_21195,N_18280,N_19024);
xnor U21196 (N_21196,N_18713,N_18781);
xnor U21197 (N_21197,N_19050,N_19873);
and U21198 (N_21198,N_20925,N_18436);
or U21199 (N_21199,N_20029,N_19114);
and U21200 (N_21200,N_19616,N_18698);
nor U21201 (N_21201,N_20248,N_18190);
nand U21202 (N_21202,N_19654,N_18297);
or U21203 (N_21203,N_19983,N_19141);
or U21204 (N_21204,N_18568,N_18792);
and U21205 (N_21205,N_18081,N_20346);
and U21206 (N_21206,N_18007,N_18971);
xnor U21207 (N_21207,N_19136,N_18682);
nand U21208 (N_21208,N_20134,N_19531);
nand U21209 (N_21209,N_19689,N_18346);
xor U21210 (N_21210,N_18427,N_18092);
and U21211 (N_21211,N_19464,N_19976);
and U21212 (N_21212,N_18984,N_20697);
nand U21213 (N_21213,N_19872,N_18945);
xnor U21214 (N_21214,N_20825,N_20465);
nand U21215 (N_21215,N_19888,N_20039);
nand U21216 (N_21216,N_19247,N_20582);
nor U21217 (N_21217,N_18445,N_19188);
xnor U21218 (N_21218,N_20386,N_18902);
and U21219 (N_21219,N_19429,N_18003);
nand U21220 (N_21220,N_19294,N_19470);
nand U21221 (N_21221,N_20218,N_20779);
and U21222 (N_21222,N_18614,N_20514);
nor U21223 (N_21223,N_18181,N_18747);
nand U21224 (N_21224,N_18590,N_19269);
or U21225 (N_21225,N_18363,N_18250);
and U21226 (N_21226,N_19167,N_20564);
xor U21227 (N_21227,N_20075,N_19859);
nor U21228 (N_21228,N_18204,N_20588);
or U21229 (N_21229,N_19764,N_18618);
xnor U21230 (N_21230,N_18415,N_18943);
xor U21231 (N_21231,N_19841,N_19268);
and U21232 (N_21232,N_19825,N_20893);
nor U21233 (N_21233,N_20287,N_18166);
nand U21234 (N_21234,N_19771,N_20889);
nand U21235 (N_21235,N_19133,N_18205);
nand U21236 (N_21236,N_19800,N_19785);
nor U21237 (N_21237,N_18621,N_18073);
and U21238 (N_21238,N_20946,N_20575);
or U21239 (N_21239,N_18404,N_19765);
xor U21240 (N_21240,N_18606,N_18513);
or U21241 (N_21241,N_18881,N_19267);
xor U21242 (N_21242,N_19070,N_20043);
xor U21243 (N_21243,N_20259,N_20802);
and U21244 (N_21244,N_18110,N_19498);
or U21245 (N_21245,N_18061,N_20357);
xnor U21246 (N_21246,N_19178,N_18982);
nor U21247 (N_21247,N_18430,N_19809);
or U21248 (N_21248,N_19608,N_19850);
or U21249 (N_21249,N_18043,N_20998);
and U21250 (N_21250,N_19609,N_19313);
or U21251 (N_21251,N_20222,N_19362);
nor U21252 (N_21252,N_20583,N_20609);
xor U21253 (N_21253,N_19820,N_18821);
nor U21254 (N_21254,N_20307,N_18178);
xor U21255 (N_21255,N_20305,N_18975);
nand U21256 (N_21256,N_20745,N_18355);
or U21257 (N_21257,N_18968,N_19160);
nand U21258 (N_21258,N_18005,N_18559);
or U21259 (N_21259,N_18466,N_19077);
nand U21260 (N_21260,N_18826,N_20788);
xor U21261 (N_21261,N_18602,N_19292);
or U21262 (N_21262,N_20688,N_19909);
nor U21263 (N_21263,N_19460,N_18318);
nand U21264 (N_21264,N_20221,N_18326);
or U21265 (N_21265,N_19651,N_18718);
nand U21266 (N_21266,N_19988,N_19475);
or U21267 (N_21267,N_20477,N_18552);
nand U21268 (N_21268,N_20621,N_18248);
or U21269 (N_21269,N_18639,N_20593);
or U21270 (N_21270,N_19623,N_19363);
nor U21271 (N_21271,N_19961,N_20377);
nor U21272 (N_21272,N_19129,N_19144);
nor U21273 (N_21273,N_19733,N_20508);
xnor U21274 (N_21274,N_18660,N_20193);
nor U21275 (N_21275,N_19150,N_19031);
and U21276 (N_21276,N_18479,N_18959);
nand U21277 (N_21277,N_19038,N_19585);
nand U21278 (N_21278,N_18242,N_18585);
nand U21279 (N_21279,N_19692,N_19638);
nand U21280 (N_21280,N_18725,N_18164);
nand U21281 (N_21281,N_20041,N_18866);
xnor U21282 (N_21282,N_19185,N_20174);
and U21283 (N_21283,N_19408,N_18152);
xor U21284 (N_21284,N_19679,N_20047);
and U21285 (N_21285,N_18695,N_18799);
nand U21286 (N_21286,N_19720,N_19886);
and U21287 (N_21287,N_19884,N_18521);
xnor U21288 (N_21288,N_20279,N_20859);
and U21289 (N_21289,N_20762,N_18261);
or U21290 (N_21290,N_18234,N_18627);
nor U21291 (N_21291,N_19857,N_20947);
nand U21292 (N_21292,N_18482,N_18022);
nand U21293 (N_21293,N_18296,N_19486);
nand U21294 (N_21294,N_19342,N_20490);
xnor U21295 (N_21295,N_19830,N_19507);
and U21296 (N_21296,N_19447,N_19472);
nor U21297 (N_21297,N_18493,N_18702);
or U21298 (N_21298,N_20547,N_19580);
xnor U21299 (N_21299,N_18068,N_20425);
nand U21300 (N_21300,N_20877,N_20163);
and U21301 (N_21301,N_18534,N_18839);
or U21302 (N_21302,N_20834,N_20018);
xnor U21303 (N_21303,N_19135,N_19071);
nor U21304 (N_21304,N_18182,N_20169);
and U21305 (N_21305,N_19459,N_20985);
nand U21306 (N_21306,N_19948,N_20301);
xnor U21307 (N_21307,N_20224,N_18225);
nand U21308 (N_21308,N_19099,N_19871);
or U21309 (N_21309,N_18485,N_18794);
and U21310 (N_21310,N_19628,N_18616);
nand U21311 (N_21311,N_20254,N_18716);
nor U21312 (N_21312,N_20734,N_19404);
xor U21313 (N_21313,N_19900,N_20792);
and U21314 (N_21314,N_18584,N_18657);
or U21315 (N_21315,N_19049,N_19713);
nand U21316 (N_21316,N_18838,N_20781);
nand U21317 (N_21317,N_18491,N_18274);
xnor U21318 (N_21318,N_20747,N_18746);
nor U21319 (N_21319,N_20296,N_20696);
nor U21320 (N_21320,N_20175,N_18540);
and U21321 (N_21321,N_20113,N_18617);
xnor U21322 (N_21322,N_20894,N_19956);
or U21323 (N_21323,N_20638,N_18057);
and U21324 (N_21324,N_19917,N_20845);
nor U21325 (N_21325,N_18912,N_19430);
and U21326 (N_21326,N_19673,N_18649);
nand U21327 (N_21327,N_19721,N_20267);
nand U21328 (N_21328,N_18875,N_19938);
nand U21329 (N_21329,N_20430,N_19790);
xor U21330 (N_21330,N_19254,N_19803);
xor U21331 (N_21331,N_20511,N_19833);
and U21332 (N_21332,N_20008,N_20649);
and U21333 (N_21333,N_20798,N_20937);
or U21334 (N_21334,N_19371,N_18401);
nor U21335 (N_21335,N_20351,N_18079);
nor U21336 (N_21336,N_18516,N_18372);
and U21337 (N_21337,N_19743,N_19740);
xnor U21338 (N_21338,N_20938,N_18282);
nor U21339 (N_21339,N_20243,N_20456);
nand U21340 (N_21340,N_20335,N_20474);
nor U21341 (N_21341,N_19305,N_18995);
nor U21342 (N_21342,N_19055,N_18128);
and U21343 (N_21343,N_19174,N_20049);
or U21344 (N_21344,N_18174,N_18454);
or U21345 (N_21345,N_18947,N_18937);
xnor U21346 (N_21346,N_19105,N_19281);
or U21347 (N_21347,N_20683,N_20167);
and U21348 (N_21348,N_18013,N_18690);
and U21349 (N_21349,N_18562,N_20013);
nand U21350 (N_21350,N_20178,N_18463);
nor U21351 (N_21351,N_19510,N_20809);
or U21352 (N_21352,N_20331,N_19481);
and U21353 (N_21353,N_19388,N_19937);
nor U21354 (N_21354,N_20880,N_20862);
or U21355 (N_21355,N_20444,N_19583);
and U21356 (N_21356,N_18591,N_19367);
nor U21357 (N_21357,N_18381,N_18490);
and U21358 (N_21358,N_20196,N_19346);
or U21359 (N_21359,N_18900,N_18558);
xnor U21360 (N_21360,N_18842,N_19378);
xnor U21361 (N_21361,N_18503,N_19212);
xnor U21362 (N_21362,N_20874,N_20439);
and U21363 (N_21363,N_20091,N_19590);
and U21364 (N_21364,N_19904,N_20229);
or U21365 (N_21365,N_19663,N_19054);
nor U21366 (N_21366,N_20325,N_18655);
or U21367 (N_21367,N_20294,N_18547);
and U21368 (N_21368,N_19252,N_19541);
nand U21369 (N_21369,N_20464,N_19495);
xnor U21370 (N_21370,N_20955,N_20731);
xnor U21371 (N_21371,N_18743,N_18176);
and U21372 (N_21372,N_19595,N_18536);
and U21373 (N_21373,N_19093,N_19933);
or U21374 (N_21374,N_20164,N_20080);
xnor U21375 (N_21375,N_20716,N_19366);
and U21376 (N_21376,N_19710,N_19999);
or U21377 (N_21377,N_20981,N_18125);
nand U21378 (N_21378,N_20799,N_20467);
and U21379 (N_21379,N_19219,N_19097);
or U21380 (N_21380,N_18383,N_19593);
xnor U21381 (N_21381,N_20277,N_19647);
xnor U21382 (N_21382,N_18069,N_19814);
xnor U21383 (N_21383,N_20896,N_18543);
and U21384 (N_21384,N_19568,N_19082);
or U21385 (N_21385,N_19662,N_18327);
or U21386 (N_21386,N_20202,N_18456);
and U21387 (N_21387,N_20934,N_20390);
xor U21388 (N_21388,N_18641,N_19508);
or U21389 (N_21389,N_19601,N_20088);
nor U21390 (N_21390,N_18177,N_19161);
xor U21391 (N_21391,N_18884,N_19839);
and U21392 (N_21392,N_20930,N_19432);
and U21393 (N_21393,N_20757,N_19644);
xor U21394 (N_21394,N_18841,N_19407);
or U21395 (N_21395,N_19694,N_18548);
and U21396 (N_21396,N_20753,N_18451);
and U21397 (N_21397,N_18131,N_18015);
or U21398 (N_21398,N_19629,N_20204);
nor U21399 (N_21399,N_18324,N_19334);
and U21400 (N_21400,N_18173,N_18736);
or U21401 (N_21401,N_20964,N_19582);
or U21402 (N_21402,N_18494,N_18962);
xor U21403 (N_21403,N_19927,N_18669);
or U21404 (N_21404,N_18258,N_18361);
xor U21405 (N_21405,N_20646,N_18629);
or U21406 (N_21406,N_19311,N_19828);
xor U21407 (N_21407,N_18196,N_18388);
xor U21408 (N_21408,N_18950,N_18241);
nand U21409 (N_21409,N_20923,N_20598);
and U21410 (N_21410,N_19515,N_20038);
nand U21411 (N_21411,N_18500,N_19293);
and U21412 (N_21412,N_18951,N_20001);
nor U21413 (N_21413,N_19610,N_19032);
or U21414 (N_21414,N_19902,N_19977);
nor U21415 (N_21415,N_19971,N_19182);
nand U21416 (N_21416,N_20117,N_19309);
xnor U21417 (N_21417,N_20283,N_18940);
nand U21418 (N_21418,N_19239,N_19455);
nand U21419 (N_21419,N_19746,N_19474);
or U21420 (N_21420,N_19419,N_19344);
or U21421 (N_21421,N_18619,N_18008);
xor U21422 (N_21422,N_18899,N_20654);
or U21423 (N_21423,N_20852,N_18185);
xor U21424 (N_21424,N_20314,N_20176);
nor U21425 (N_21425,N_20150,N_20362);
xnor U21426 (N_21426,N_20994,N_20562);
nand U21427 (N_21427,N_20704,N_20327);
nor U21428 (N_21428,N_19148,N_18916);
or U21429 (N_21429,N_20375,N_20260);
and U21430 (N_21430,N_19805,N_18851);
xnor U21431 (N_21431,N_20940,N_18769);
nor U21432 (N_21432,N_18973,N_20942);
xnor U21433 (N_21433,N_20012,N_20345);
xor U21434 (N_21434,N_18065,N_20363);
nand U21435 (N_21435,N_19921,N_20146);
nand U21436 (N_21436,N_18257,N_18624);
nor U21437 (N_21437,N_18002,N_18366);
and U21438 (N_21438,N_18990,N_18136);
nor U21439 (N_21439,N_18628,N_19206);
nand U21440 (N_21440,N_18934,N_20710);
or U21441 (N_21441,N_18567,N_20585);
nor U21442 (N_21442,N_18928,N_19243);
and U21443 (N_21443,N_20881,N_20604);
xor U21444 (N_21444,N_19799,N_18860);
and U21445 (N_21445,N_18829,N_18281);
nor U21446 (N_21446,N_18802,N_19630);
or U21447 (N_21447,N_20181,N_18104);
nor U21448 (N_21448,N_18435,N_19887);
xnor U21449 (N_21449,N_19000,N_20110);
xnor U21450 (N_21450,N_20315,N_18313);
and U21451 (N_21451,N_18906,N_20027);
or U21452 (N_21452,N_20217,N_20058);
nor U21453 (N_21453,N_18712,N_19865);
nand U21454 (N_21454,N_20272,N_19416);
nor U21455 (N_21455,N_20786,N_19203);
xnor U21456 (N_21456,N_19034,N_20208);
and U21457 (N_21457,N_19730,N_20821);
or U21458 (N_21458,N_19146,N_19046);
nor U21459 (N_21459,N_19959,N_20920);
and U21460 (N_21460,N_20784,N_20097);
and U21461 (N_21461,N_19877,N_20695);
and U21462 (N_21462,N_19624,N_19974);
and U21463 (N_21463,N_20352,N_19376);
nand U21464 (N_21464,N_19341,N_19920);
or U21465 (N_21465,N_19687,N_19027);
nand U21466 (N_21466,N_20040,N_20816);
xor U21467 (N_21467,N_20707,N_20886);
and U21468 (N_21468,N_19845,N_18216);
or U21469 (N_21469,N_20413,N_19968);
nand U21470 (N_21470,N_19021,N_18472);
and U21471 (N_21471,N_18478,N_19333);
nor U21472 (N_21472,N_18091,N_20746);
or U21473 (N_21473,N_18165,N_20470);
or U21474 (N_21474,N_18861,N_19969);
xor U21475 (N_21475,N_19175,N_18848);
xor U21476 (N_21476,N_18060,N_19354);
nand U21477 (N_21477,N_20669,N_18704);
and U21478 (N_21478,N_19671,N_18376);
nand U21479 (N_21479,N_18186,N_18199);
nand U21480 (N_21480,N_20939,N_20950);
nor U21481 (N_21481,N_20507,N_18610);
xor U21482 (N_21482,N_18301,N_19573);
or U21483 (N_21483,N_20336,N_19187);
and U21484 (N_21484,N_20833,N_20220);
nor U21485 (N_21485,N_18156,N_20092);
xor U21486 (N_21486,N_19473,N_20297);
nand U21487 (N_21487,N_20839,N_20548);
or U21488 (N_21488,N_20924,N_20311);
xnor U21489 (N_21489,N_18673,N_19786);
xor U21490 (N_21490,N_19812,N_20251);
nand U21491 (N_21491,N_19436,N_20771);
nor U21492 (N_21492,N_20046,N_20505);
nor U21493 (N_21493,N_18710,N_20817);
nor U21494 (N_21494,N_18295,N_20280);
nor U21495 (N_21495,N_18238,N_20699);
or U21496 (N_21496,N_20539,N_19015);
nand U21497 (N_21497,N_20152,N_18813);
xor U21498 (N_21498,N_18635,N_19546);
or U21499 (N_21499,N_18667,N_20528);
nand U21500 (N_21500,N_19642,N_20796);
xor U21501 (N_21501,N_19835,N_18377);
and U21502 (N_21502,N_20861,N_19327);
and U21503 (N_21503,N_18537,N_20722);
xor U21504 (N_21504,N_18546,N_19566);
and U21505 (N_21505,N_18806,N_20735);
nor U21506 (N_21506,N_18679,N_18028);
or U21507 (N_21507,N_18010,N_19120);
or U21508 (N_21508,N_18805,N_19147);
nor U21509 (N_21509,N_19403,N_18757);
xor U21510 (N_21510,N_18523,N_18927);
or U21511 (N_21511,N_18678,N_20210);
and U21512 (N_21512,N_19536,N_19350);
nor U21513 (N_21513,N_19295,N_20855);
nor U21514 (N_21514,N_19019,N_19315);
or U21515 (N_21515,N_19625,N_20635);
and U21516 (N_21516,N_19250,N_19788);
nand U21517 (N_21517,N_18254,N_19405);
and U21518 (N_21518,N_20565,N_18960);
xnor U21519 (N_21519,N_18148,N_18486);
nand U21520 (N_21520,N_20123,N_20637);
xnor U21521 (N_21521,N_18633,N_19503);
nor U21522 (N_21522,N_19216,N_19645);
xnor U21523 (N_21523,N_20633,N_19709);
nand U21524 (N_21524,N_19894,N_18207);
nand U21525 (N_21525,N_20281,N_19379);
or U21526 (N_21526,N_20440,N_20976);
and U21527 (N_21527,N_18659,N_19860);
nor U21528 (N_21528,N_18527,N_20408);
nand U21529 (N_21529,N_19300,N_18705);
nand U21530 (N_21530,N_19134,N_18259);
and U21531 (N_21531,N_20048,N_19441);
nor U21532 (N_21532,N_19384,N_20677);
nor U21533 (N_21533,N_18795,N_20659);
or U21534 (N_21534,N_20577,N_18434);
xor U21535 (N_21535,N_18406,N_20129);
and U21536 (N_21536,N_18273,N_20841);
xnor U21537 (N_21537,N_19440,N_18531);
nand U21538 (N_21538,N_20541,N_19599);
nor U21539 (N_21539,N_18738,N_19086);
xor U21540 (N_21540,N_20693,N_18029);
nor U21541 (N_21541,N_18996,N_19963);
nand U21542 (N_21542,N_18078,N_19494);
and U21543 (N_21543,N_18032,N_18810);
or U21544 (N_21544,N_18693,N_18615);
xor U21545 (N_21545,N_18421,N_20698);
nand U21546 (N_21546,N_20235,N_20728);
or U21547 (N_21547,N_20980,N_18086);
or U21548 (N_21548,N_20225,N_19987);
or U21549 (N_21549,N_19527,N_20850);
xor U21550 (N_21550,N_20851,N_20369);
nor U21551 (N_21551,N_20922,N_18226);
and U21552 (N_21552,N_18334,N_18119);
and U21553 (N_21553,N_19230,N_19774);
nand U21554 (N_21554,N_18824,N_18987);
or U21555 (N_21555,N_18142,N_18632);
xnor U21556 (N_21556,N_19041,N_18853);
nand U21557 (N_21557,N_19368,N_20530);
or U21558 (N_21558,N_19047,N_19339);
xnor U21559 (N_21559,N_18770,N_18269);
xnor U21560 (N_21560,N_20449,N_19538);
and U21561 (N_21561,N_18828,N_18072);
and U21562 (N_21562,N_18753,N_20269);
nor U21563 (N_21563,N_18570,N_18600);
xnor U21564 (N_21564,N_19088,N_18830);
xnor U21565 (N_21565,N_19637,N_18879);
nor U21566 (N_21566,N_20371,N_19402);
or U21567 (N_21567,N_20580,N_20854);
nor U21568 (N_21568,N_19991,N_18306);
xnor U21569 (N_21569,N_20533,N_19684);
nand U21570 (N_21570,N_19955,N_18442);
nor U21571 (N_21571,N_18413,N_19253);
nor U21572 (N_21572,N_19241,N_18412);
nor U21573 (N_21573,N_19445,N_18236);
xor U21574 (N_21574,N_19488,N_19351);
or U21575 (N_21575,N_19520,N_20199);
nor U21576 (N_21576,N_20787,N_20656);
or U21577 (N_21577,N_19696,N_18014);
and U21578 (N_21578,N_18653,N_20765);
xor U21579 (N_21579,N_20755,N_19940);
nor U21580 (N_21580,N_19283,N_19661);
or U21581 (N_21581,N_20446,N_18779);
nor U21582 (N_21582,N_20100,N_18530);
nor U21583 (N_21583,N_18520,N_18139);
xor U21584 (N_21584,N_19528,N_18961);
and U21585 (N_21585,N_19666,N_19761);
nor U21586 (N_21586,N_20111,N_20830);
or U21587 (N_21587,N_20858,N_19504);
nor U21588 (N_21588,N_19410,N_18154);
and U21589 (N_21589,N_20895,N_20216);
or U21590 (N_21590,N_19936,N_19749);
nor U21591 (N_21591,N_18914,N_18766);
and U21592 (N_21592,N_20663,N_18432);
nor U21593 (N_21593,N_19973,N_20128);
or U21594 (N_21594,N_20560,N_18658);
nand U21595 (N_21595,N_20749,N_18167);
nor U21596 (N_21596,N_20022,N_18353);
xor U21597 (N_21597,N_18631,N_20323);
nor U21598 (N_21598,N_20108,N_18603);
xnor U21599 (N_21599,N_20727,N_19081);
xor U21600 (N_21600,N_19686,N_18000);
nand U21601 (N_21601,N_19298,N_19754);
xor U21602 (N_21602,N_19365,N_19875);
or U21603 (N_21603,N_20559,N_20991);
xor U21604 (N_21604,N_19668,N_20600);
nor U21605 (N_21605,N_20334,N_20074);
nor U21606 (N_21606,N_19260,N_20605);
nand U21607 (N_21607,N_18517,N_18063);
and U21608 (N_21608,N_19194,N_18501);
and U21609 (N_21609,N_20943,N_19456);
or U21610 (N_21610,N_20187,N_20399);
and U21611 (N_21611,N_18807,N_18785);
and U21612 (N_21612,N_20806,N_18672);
xnor U21613 (N_21613,N_20797,N_20179);
nor U21614 (N_21614,N_19650,N_18551);
nand U21615 (N_21615,N_20299,N_19529);
xor U21616 (N_21616,N_20831,N_19571);
xnor U21617 (N_21617,N_19897,N_19057);
and U21618 (N_21618,N_19116,N_19220);
nand U21619 (N_21619,N_19796,N_19438);
nor U21620 (N_21620,N_20537,N_18118);
nand U21621 (N_21621,N_20843,N_19349);
nor U21622 (N_21622,N_20406,N_20538);
or U21623 (N_21623,N_20480,N_18514);
nor U21624 (N_21624,N_20848,N_18529);
and U21625 (N_21625,N_18820,N_19572);
nand U21626 (N_21626,N_19856,N_20584);
and U21627 (N_21627,N_20368,N_20632);
and U21628 (N_21628,N_19807,N_19452);
nor U21629 (N_21629,N_20300,N_18509);
nand U21630 (N_21630,N_18098,N_20818);
nand U21631 (N_21631,N_19676,N_19843);
xor U21632 (N_21632,N_19215,N_20403);
xor U21633 (N_21633,N_18755,N_18626);
and U21634 (N_21634,N_19569,N_19390);
or U21635 (N_21635,N_18869,N_18601);
and U21636 (N_21636,N_18569,N_20606);
nor U21637 (N_21637,N_19895,N_18024);
nand U21638 (N_21638,N_18714,N_19153);
nor U21639 (N_21639,N_19296,N_20997);
nor U21640 (N_21640,N_20661,N_20376);
and U21641 (N_21641,N_20353,N_19600);
and U21642 (N_21642,N_20782,N_19632);
or U21643 (N_21643,N_18283,N_19617);
and U21644 (N_21644,N_18387,N_19397);
and U21645 (N_21645,N_20993,N_19741);
and U21646 (N_21646,N_18317,N_18260);
xnor U21647 (N_21647,N_19424,N_18305);
or U21648 (N_21648,N_18717,N_18206);
xor U21649 (N_21649,N_18300,N_19784);
and U21650 (N_21650,N_20521,N_19945);
or U21651 (N_21651,N_19952,N_19517);
nand U21652 (N_21652,N_18099,N_20602);
nand U21653 (N_21653,N_19649,N_18431);
nand U21654 (N_21654,N_20995,N_18112);
xor U21655 (N_21655,N_20824,N_19944);
xnor U21656 (N_21656,N_18847,N_19080);
nor U21657 (N_21657,N_20545,N_18338);
and U21658 (N_21658,N_18582,N_18328);
nor U21659 (N_21659,N_19079,N_18992);
or U21660 (N_21660,N_18030,N_20509);
and U21661 (N_21661,N_20293,N_20927);
nor U21662 (N_21662,N_20434,N_19324);
or U21663 (N_21663,N_19942,N_20628);
and U21664 (N_21664,N_19646,N_18597);
xnor U21665 (N_21665,N_19972,N_18840);
or U21666 (N_21666,N_20003,N_18071);
and U21667 (N_21667,N_18358,N_18773);
nand U21668 (N_21668,N_18201,N_20773);
or U21669 (N_21669,N_19876,N_18044);
or U21670 (N_21670,N_19245,N_18854);
nand U21671 (N_21671,N_20623,N_18457);
nor U21672 (N_21672,N_20468,N_20389);
xnor U21673 (N_21673,N_19061,N_19559);
xnor U21674 (N_21674,N_19477,N_18685);
or U21675 (N_21675,N_19338,N_18587);
nand U21676 (N_21676,N_18371,N_20647);
and U21677 (N_21677,N_19483,N_19089);
or U21678 (N_21678,N_20409,N_20160);
xor U21679 (N_21679,N_19454,N_20004);
or U21680 (N_21680,N_19899,N_19753);
nand U21681 (N_21681,N_19040,N_18703);
xor U21682 (N_21682,N_18563,N_18911);
and U21683 (N_21683,N_20308,N_20844);
nor U21684 (N_21684,N_18428,N_18997);
xnor U21685 (N_21685,N_20042,N_18145);
nand U21686 (N_21686,N_19149,N_18532);
nor U21687 (N_21687,N_18581,N_20493);
and U21688 (N_21688,N_19928,N_19914);
nor U21689 (N_21689,N_19489,N_19045);
nand U21690 (N_21690,N_19425,N_20703);
nor U21691 (N_21691,N_18132,N_19013);
or U21692 (N_21692,N_20484,N_20112);
nand U21693 (N_21693,N_20155,N_18336);
and U21694 (N_21694,N_18576,N_20929);
nand U21695 (N_21695,N_19117,N_18193);
xnor U21696 (N_21696,N_18677,N_20298);
and U21697 (N_21697,N_20532,N_20884);
or U21698 (N_21698,N_20316,N_18604);
and U21699 (N_21699,N_18316,N_20158);
nand U21700 (N_21700,N_19222,N_18465);
and U21701 (N_21701,N_19635,N_19130);
or U21702 (N_21702,N_19540,N_18630);
or U21703 (N_21703,N_19555,N_18397);
nand U21704 (N_21704,N_19479,N_18335);
nor U21705 (N_21705,N_20192,N_20328);
and U21706 (N_21706,N_20239,N_20232);
nor U21707 (N_21707,N_19288,N_20832);
and U21708 (N_21708,N_18645,N_19469);
and U21709 (N_21709,N_20553,N_19862);
or U21710 (N_21710,N_18038,N_20476);
and U21711 (N_21711,N_20887,N_19487);
or U21712 (N_21712,N_18835,N_18572);
xor U21713 (N_21713,N_18708,N_20898);
or U21714 (N_21714,N_20592,N_20247);
or U21715 (N_21715,N_18855,N_20304);
nor U21716 (N_21716,N_18647,N_19036);
or U21717 (N_21717,N_20761,N_20278);
xor U21718 (N_21718,N_18217,N_19562);
and U21719 (N_21719,N_19157,N_18230);
nor U21720 (N_21720,N_20121,N_20571);
or U21721 (N_21721,N_18907,N_18488);
nor U21722 (N_21722,N_18489,N_20766);
xnor U21723 (N_21723,N_18262,N_19204);
nand U21724 (N_21724,N_20454,N_18734);
and U21725 (N_21725,N_18140,N_19023);
nor U21726 (N_21726,N_20813,N_20417);
or U21727 (N_21727,N_19223,N_20791);
xor U21728 (N_21728,N_19420,N_19231);
xor U21729 (N_21729,N_18903,N_19035);
nor U21730 (N_21730,N_19511,N_20990);
nand U21731 (N_21731,N_19392,N_18340);
and U21732 (N_21732,N_20709,N_19062);
nor U21733 (N_21733,N_18390,N_18394);
and U21734 (N_21734,N_20072,N_19221);
xnor U21735 (N_21735,N_18083,N_20867);
and U21736 (N_21736,N_18310,N_18198);
or U21737 (N_21737,N_19043,N_18067);
and U21738 (N_21738,N_19691,N_20083);
xnor U21739 (N_21739,N_19449,N_20554);
and U21740 (N_21740,N_18539,N_19139);
or U21741 (N_21741,N_20045,N_20385);
xnor U21742 (N_21742,N_18384,N_20733);
or U21743 (N_21743,N_19509,N_20322);
nand U21744 (N_21744,N_19979,N_19090);
nand U21745 (N_21745,N_19735,N_18134);
and U21746 (N_21746,N_19457,N_20212);
or U21747 (N_21747,N_20089,N_19303);
nand U21748 (N_21748,N_20726,N_18784);
or U21749 (N_21749,N_20015,N_20724);
nand U21750 (N_21750,N_19026,N_18749);
xor U21751 (N_21751,N_18575,N_18913);
or U21752 (N_21752,N_20428,N_18116);
nor U21753 (N_21753,N_20133,N_18348);
nand U21754 (N_21754,N_18596,N_18814);
nand U21755 (N_21755,N_20114,N_20689);
or U21756 (N_21756,N_19577,N_18408);
nor U21757 (N_21757,N_19905,N_18403);
and U21758 (N_21758,N_19848,N_19205);
nand U21759 (N_21759,N_18849,N_19173);
or U21760 (N_21760,N_19244,N_20932);
nor U21761 (N_21761,N_20795,N_20827);
or U21762 (N_21762,N_19866,N_19002);
xnor U21763 (N_21763,N_18341,N_18237);
and U21764 (N_21764,N_20679,N_18740);
nor U21765 (N_21765,N_19700,N_19297);
nand U21766 (N_21766,N_18623,N_18599);
xor U21767 (N_21767,N_18857,N_18735);
xor U21768 (N_21768,N_19306,N_20171);
nand U21769 (N_21769,N_19570,N_18721);
nand U21770 (N_21770,N_19576,N_19672);
and U21771 (N_21771,N_18121,N_20711);
nor U21772 (N_21772,N_20137,N_20329);
nand U21773 (N_21773,N_19950,N_20140);
xor U21774 (N_21774,N_20636,N_19030);
nor U21775 (N_21775,N_18634,N_18055);
nor U21776 (N_21776,N_19598,N_20383);
xnor U21777 (N_21777,N_18731,N_20131);
nor U21778 (N_21778,N_18856,N_18141);
nand U21779 (N_21779,N_20462,N_18646);
or U21780 (N_21780,N_20601,N_20337);
nor U21781 (N_21781,N_19832,N_18009);
nor U21782 (N_21782,N_18367,N_20566);
or U21783 (N_21783,N_18192,N_19277);
xnor U21784 (N_21784,N_20156,N_19794);
xor U21785 (N_21785,N_20266,N_18268);
nand U21786 (N_21786,N_19719,N_19058);
and U21787 (N_21787,N_19198,N_20653);
xor U21788 (N_21788,N_18058,N_19626);
nor U21789 (N_21789,N_20461,N_18507);
and U21790 (N_21790,N_19165,N_20073);
or U21791 (N_21791,N_19837,N_19262);
and U21792 (N_21792,N_19763,N_20139);
xor U21793 (N_21793,N_18373,N_19881);
and U21794 (N_21794,N_20017,N_20835);
nand U21795 (N_21795,N_20289,N_19110);
xor U21796 (N_21796,N_18417,N_18468);
or U21797 (N_21797,N_19907,N_19179);
and U21798 (N_21798,N_18016,N_18778);
nand U21799 (N_21799,N_18775,N_20614);
nand U21800 (N_21800,N_19847,N_19087);
and U21801 (N_21801,N_18304,N_18045);
nand U21802 (N_21802,N_20526,N_19759);
nand U21803 (N_21803,N_20873,N_19553);
nand U21804 (N_21804,N_20999,N_20657);
xnor U21805 (N_21805,N_18422,N_19521);
or U21806 (N_21806,N_19838,N_18012);
nor U21807 (N_21807,N_20977,N_18263);
or U21808 (N_21808,N_20617,N_18791);
xor U21809 (N_21809,N_19106,N_19707);
nand U21810 (N_21810,N_20572,N_20901);
and U21811 (N_21811,N_20397,N_20651);
nor U21812 (N_21812,N_20016,N_19712);
nand U21813 (N_21813,N_20055,N_18414);
xor U21814 (N_21814,N_18298,N_20421);
or U21815 (N_21815,N_20563,N_19931);
xor U21816 (N_21816,N_18777,N_18967);
and U21817 (N_21817,N_20737,N_20767);
and U21818 (N_21818,N_19792,N_18374);
xnor U21819 (N_21819,N_19387,N_19986);
xnor U21820 (N_21820,N_19411,N_20721);
xnor U21821 (N_21821,N_20142,N_20789);
and U21822 (N_21822,N_18686,N_20104);
and U21823 (N_21823,N_20119,N_19453);
or U21824 (N_21824,N_18885,N_20324);
nor U21825 (N_21825,N_19426,N_18194);
or U21826 (N_21826,N_19323,N_19289);
nor U21827 (N_21827,N_20076,N_20608);
nor U21828 (N_21828,N_19715,N_18034);
nand U21829 (N_21829,N_19813,N_19399);
nor U21830 (N_21830,N_18218,N_18979);
and U21831 (N_21831,N_20373,N_20495);
nand U21832 (N_21832,N_18102,N_18410);
xor U21833 (N_21833,N_19382,N_20077);
xnor U21834 (N_21834,N_18593,N_18553);
and U21835 (N_21835,N_18986,N_20034);
or U21836 (N_21836,N_20949,N_18963);
and U21837 (N_21837,N_18035,N_20668);
or U21838 (N_21838,N_19319,N_20063);
nand U21839 (N_21839,N_20944,N_20025);
nand U21840 (N_21840,N_20910,N_19326);
xnor U21841 (N_21841,N_18780,N_20332);
xor U21842 (N_21842,N_20200,N_19418);
xor U21843 (N_21843,N_19201,N_20717);
and U21844 (N_21844,N_19393,N_20790);
nand U21845 (N_21845,N_20078,N_20725);
and U21846 (N_21846,N_18460,N_18772);
or U21847 (N_21847,N_18827,N_19336);
nor U21848 (N_21848,N_20988,N_19073);
xnor U21849 (N_21849,N_18858,N_19278);
or U21850 (N_21850,N_20234,N_19795);
nor U21851 (N_21851,N_18541,N_19197);
and U21852 (N_21852,N_18450,N_20438);
nor U21853 (N_21853,N_18441,N_20700);
and U21854 (N_21854,N_19434,N_18411);
and U21855 (N_21855,N_19960,N_18275);
xor U21856 (N_21856,N_19998,N_18954);
xnor U21857 (N_21857,N_18474,N_18137);
xor U21858 (N_21858,N_20130,N_20793);
and U21859 (N_21859,N_18396,N_19688);
xor U21860 (N_21860,N_19727,N_20019);
and U21861 (N_21861,N_18966,N_19824);
or U21862 (N_21862,N_18423,N_18159);
nand U21863 (N_21863,N_18290,N_18697);
or U21864 (N_21864,N_20036,N_18595);
nor U21865 (N_21865,N_19122,N_19717);
nor U21866 (N_21866,N_19697,N_18578);
or U21867 (N_21867,N_20069,N_18921);
and U21868 (N_21868,N_18240,N_20350);
or U21869 (N_21869,N_19502,N_20909);
xnor U21870 (N_21870,N_20370,N_20227);
or U21871 (N_21871,N_20953,N_18510);
nand U21872 (N_21872,N_18146,N_19725);
and U21873 (N_21873,N_20183,N_18064);
nand U21874 (N_21874,N_20024,N_18343);
and U21875 (N_21875,N_19767,N_19417);
xnor U21876 (N_21876,N_18220,N_19091);
and U21877 (N_21877,N_19655,N_19874);
and U21878 (N_21878,N_19039,N_20958);
or U21879 (N_21879,N_20540,N_20904);
or U21880 (N_21880,N_18637,N_19996);
nor U21881 (N_21881,N_18701,N_18638);
and U21882 (N_21882,N_20492,N_20527);
nand U21883 (N_21883,N_18499,N_19029);
xnor U21884 (N_21884,N_20452,N_18356);
and U21885 (N_21885,N_19534,N_18675);
or U21886 (N_21886,N_20611,N_18935);
or U21887 (N_21887,N_19535,N_18210);
and U21888 (N_21888,N_18386,N_19127);
and U21889 (N_21889,N_20366,N_18932);
xor U21890 (N_21890,N_19615,N_20258);
and U21891 (N_21891,N_18739,N_20569);
and U21892 (N_21892,N_18994,N_20106);
nor U21893 (N_21893,N_20455,N_19648);
nand U21894 (N_21894,N_19353,N_19519);
and U21895 (N_21895,N_20407,N_18533);
nand U21896 (N_21896,N_19490,N_20579);
and U21897 (N_21897,N_18077,N_20021);
xnor U21898 (N_21898,N_18496,N_18347);
or U21899 (N_21899,N_20054,N_18666);
nand U21900 (N_21900,N_20341,N_19729);
xnor U21901 (N_21901,N_20568,N_19068);
and U21902 (N_21902,N_20520,N_19431);
nor U21903 (N_21903,N_18352,N_20211);
nand U21904 (N_21904,N_19302,N_18687);
nor U21905 (N_21905,N_20374,N_19748);
and U21906 (N_21906,N_20917,N_18052);
xor U21907 (N_21907,N_20116,N_19893);
nand U21908 (N_21908,N_19605,N_20349);
or U21909 (N_21909,N_19450,N_20382);
nand U21910 (N_21910,N_20360,N_18818);
nand U21911 (N_21911,N_20674,N_18498);
or U21912 (N_21912,N_18223,N_20567);
and U21913 (N_21913,N_20223,N_20050);
or U21914 (N_21914,N_18399,N_19232);
and U21915 (N_21915,N_18308,N_19056);
and U21916 (N_21916,N_19929,N_18650);
or U21917 (N_21917,N_19016,N_18244);
nor U21918 (N_21918,N_19169,N_20154);
xnor U21919 (N_21919,N_19274,N_20241);
nor U21920 (N_21920,N_18611,N_19299);
nand U21921 (N_21921,N_19975,N_18127);
xnor U21922 (N_21922,N_19806,N_19458);
and U21923 (N_21923,N_18893,N_18694);
nand U21924 (N_21924,N_20715,N_20878);
or U21925 (N_21925,N_18109,N_18819);
or U21926 (N_21926,N_20079,N_20141);
or U21927 (N_21927,N_19532,N_20915);
xor U21928 (N_21928,N_20686,N_18880);
nor U21929 (N_21929,N_20513,N_19193);
and U21930 (N_21930,N_20284,N_18054);
xnor U21931 (N_21931,N_20172,N_19836);
xor U21932 (N_21932,N_18320,N_20868);
nand U21933 (N_21933,N_19726,N_19176);
or U21934 (N_21934,N_20650,N_20552);
or U21935 (N_21935,N_20051,N_20009);
and U21936 (N_21936,N_19657,N_20743);
or U21937 (N_21937,N_18988,N_18999);
and U21938 (N_21938,N_18560,N_19316);
xnor U21939 (N_21939,N_18243,N_20361);
or U21940 (N_21940,N_18583,N_19308);
nand U21941 (N_21941,N_19168,N_18379);
or U21942 (N_21942,N_19131,N_20785);
nand U21943 (N_21943,N_20448,N_20729);
nor U21944 (N_21944,N_20244,N_19744);
and U21945 (N_21945,N_20180,N_18652);
nand U21946 (N_21946,N_20629,N_20132);
or U21947 (N_21947,N_20890,N_19779);
or U21948 (N_21948,N_19783,N_20478);
or U21949 (N_21949,N_19575,N_20411);
nand U21950 (N_21950,N_20972,N_20603);
nor U21951 (N_21951,N_20501,N_19934);
xnor U21952 (N_21952,N_19922,N_19702);
and U21953 (N_21953,N_19918,N_19255);
xor U21954 (N_21954,N_19398,N_18094);
nand U21955 (N_21955,N_20381,N_18416);
or U21956 (N_21956,N_18867,N_20423);
and U21957 (N_21957,N_19083,N_18252);
nand U21958 (N_21958,N_20826,N_18741);
xor U21959 (N_21959,N_18870,N_20188);
or U21960 (N_21960,N_18001,N_19653);
or U21961 (N_21961,N_18644,N_19618);
or U21962 (N_21962,N_19797,N_19183);
nand U21963 (N_21963,N_18788,N_18286);
or U21964 (N_21964,N_18891,N_19361);
nor U21965 (N_21965,N_18844,N_18625);
xnor U21966 (N_21966,N_18271,N_19389);
nand U21967 (N_21967,N_20475,N_18209);
nor U21968 (N_21968,N_18293,N_18359);
nor U21969 (N_21969,N_18664,N_20911);
or U21970 (N_21970,N_19257,N_19989);
nor U21971 (N_21971,N_19821,N_19414);
or U21972 (N_21972,N_19705,N_19556);
nand U21973 (N_21973,N_20246,N_19433);
nor U21974 (N_21974,N_20673,N_18122);
nor U21975 (N_21975,N_18437,N_20485);
or U21976 (N_21976,N_19620,N_18219);
nand U21977 (N_21977,N_18895,N_19172);
xnor U21978 (N_21978,N_20780,N_19270);
nor U21979 (N_21979,N_18728,N_20574);
or U21980 (N_21980,N_19163,N_19910);
or U21981 (N_21981,N_19500,N_19724);
nor U21982 (N_21982,N_19993,N_20667);
and U21983 (N_21983,N_18147,N_19639);
nor U21984 (N_21984,N_19060,N_19234);
xor U21985 (N_21985,N_19098,N_20230);
nand U21986 (N_21986,N_19242,N_20772);
or U21987 (N_21987,N_20061,N_19162);
and U21988 (N_21988,N_20405,N_20189);
nor U21989 (N_21989,N_18222,N_20672);
xnor U21990 (N_21990,N_19798,N_19603);
nand U21991 (N_21991,N_18852,N_18089);
or U21992 (N_21992,N_20032,N_19854);
nand U21993 (N_21993,N_19804,N_20687);
and U21994 (N_21994,N_19196,N_19578);
nor U21995 (N_21995,N_20044,N_19891);
xor U21996 (N_21996,N_19863,N_18574);
and U21997 (N_21997,N_19370,N_20857);
nor U21998 (N_21998,N_18822,N_19997);
xor U21999 (N_21999,N_20919,N_18200);
nor U22000 (N_22000,N_20931,N_20494);
and U22001 (N_22001,N_19492,N_20086);
nand U22002 (N_22002,N_19104,N_19842);
or U22003 (N_22003,N_19272,N_20276);
nand U22004 (N_22004,N_18418,N_20333);
nor U22005 (N_22005,N_18477,N_19067);
nor U22006 (N_22006,N_18168,N_19755);
nor U22007 (N_22007,N_18459,N_19913);
nor U22008 (N_22008,N_18325,N_20136);
nor U22009 (N_22009,N_20263,N_18133);
nand U22010 (N_22010,N_20908,N_18444);
xor U22011 (N_22011,N_20451,N_19670);
or U22012 (N_22012,N_18684,N_19166);
nor U22013 (N_22013,N_19451,N_20084);
or U22014 (N_22014,N_20194,N_18696);
nand U22015 (N_22015,N_20978,N_18803);
and U22016 (N_22016,N_18228,N_18448);
and U22017 (N_22017,N_19006,N_18908);
xnor U22018 (N_22018,N_20436,N_20471);
nor U22019 (N_22019,N_19935,N_20613);
nand U22020 (N_22020,N_18850,N_19612);
xor U22021 (N_22021,N_20719,N_20238);
xnor U22022 (N_22022,N_19463,N_18424);
xor U22023 (N_22023,N_20093,N_20645);
nor U22024 (N_22024,N_18886,N_19924);
or U22025 (N_22025,N_19789,N_20531);
and U22026 (N_22026,N_18031,N_19053);
xnor U22027 (N_22027,N_19391,N_19443);
nor U22028 (N_22028,N_18566,N_20713);
nor U22029 (N_22029,N_18405,N_19701);
xnor U22030 (N_22030,N_19325,N_20472);
xnor U22031 (N_22031,N_18085,N_18171);
nor U22032 (N_22032,N_18111,N_19591);
or U22033 (N_22033,N_20432,N_18047);
and U22034 (N_22034,N_20736,N_20498);
nand U22035 (N_22035,N_18017,N_20401);
or U22036 (N_22036,N_19915,N_19664);
nor U22037 (N_22037,N_19819,N_18256);
or U22038 (N_22038,N_19728,N_20147);
nand U22039 (N_22039,N_18837,N_19422);
xnor U22040 (N_22040,N_19355,N_18758);
or U22041 (N_22041,N_18620,N_19195);
and U22042 (N_22042,N_20578,N_20060);
nand U22043 (N_22043,N_20105,N_20903);
nand U22044 (N_22044,N_20011,N_19340);
or U22045 (N_22045,N_18124,N_20967);
nand U22046 (N_22046,N_20655,N_20622);
and U22047 (N_22047,N_19518,N_20945);
xor U22048 (N_22048,N_18970,N_18267);
nor U22049 (N_22049,N_19317,N_20339);
nor U22050 (N_22050,N_19703,N_18526);
nor U22051 (N_22051,N_19844,N_19137);
nor U22052 (N_22052,N_20412,N_20524);
xnor U22053 (N_22053,N_18926,N_18965);
nand U22054 (N_22054,N_18722,N_20691);
and U22055 (N_22055,N_18113,N_20037);
or U22056 (N_22056,N_18169,N_18420);
nand U22057 (N_22057,N_20312,N_19965);
and U22058 (N_22058,N_20410,N_19385);
or U22059 (N_22059,N_18330,N_19143);
or U22060 (N_22060,N_19343,N_19982);
nor U22061 (N_22061,N_18483,N_18580);
and U22062 (N_22062,N_20052,N_20466);
xnor U22063 (N_22063,N_18946,N_18438);
nor U22064 (N_22064,N_18812,N_19064);
or U22065 (N_22065,N_20550,N_18760);
nand U22066 (N_22066,N_18834,N_19471);
and U22067 (N_22067,N_18351,N_18143);
nor U22068 (N_22068,N_20094,N_18729);
and U22069 (N_22069,N_18607,N_20866);
nand U22070 (N_22070,N_19264,N_18873);
nand U22071 (N_22071,N_19533,N_19584);
or U22072 (N_22072,N_20153,N_18957);
or U22073 (N_22073,N_20522,N_20665);
nand U22074 (N_22074,N_20245,N_20706);
or U22075 (N_22075,N_19497,N_19680);
or U22076 (N_22076,N_18255,N_18360);
nor U22077 (N_22077,N_20644,N_18100);
or U22078 (N_22078,N_20576,N_18622);
xor U22079 (N_22079,N_19811,N_18452);
xor U22080 (N_22080,N_19095,N_19949);
nand U22081 (N_22081,N_20286,N_19249);
and U22082 (N_22082,N_20897,N_20441);
nor U22083 (N_22083,N_20487,N_19012);
nand U22084 (N_22084,N_19192,N_18123);
or U22085 (N_22085,N_20641,N_19132);
xor U22086 (N_22086,N_18888,N_20253);
nor U22087 (N_22087,N_19096,N_19564);
nand U22088 (N_22088,N_20948,N_18767);
nand U22089 (N_22089,N_20064,N_20846);
and U22090 (N_22090,N_20512,N_20000);
nor U22091 (N_22091,N_19552,N_20213);
nand U22092 (N_22092,N_19667,N_19817);
or U22093 (N_22093,N_19994,N_19827);
nand U22094 (N_22094,N_19829,N_19953);
and U22095 (N_22095,N_18752,N_20053);
nand U22096 (N_22096,N_20173,N_18550);
nand U22097 (N_22097,N_18467,N_19737);
and U22098 (N_22098,N_19265,N_20203);
nor U22099 (N_22099,N_18969,N_18149);
nand U22100 (N_22100,N_20863,N_19375);
nand U22101 (N_22101,N_18544,N_20882);
nand U22102 (N_22102,N_18964,N_19476);
or U22103 (N_22103,N_20118,N_18473);
xor U22104 (N_22104,N_19113,N_19548);
nand U22105 (N_22105,N_19259,N_19076);
nor U22106 (N_22106,N_20815,N_19320);
or U22107 (N_22107,N_18985,N_20087);
xor U22108 (N_22108,N_20912,N_18350);
nor U22109 (N_22109,N_18956,N_19011);
nor U22110 (N_22110,N_18369,N_20900);
or U22111 (N_22111,N_20620,N_20198);
or U22112 (N_22112,N_19778,N_19100);
nand U22113 (N_22113,N_20957,N_19992);
nor U22114 (N_22114,N_19465,N_20343);
nor U22115 (N_22115,N_20680,N_18120);
nand U22116 (N_22116,N_18535,N_18469);
nor U22117 (N_22117,N_18287,N_19506);
nor U22118 (N_22118,N_18096,N_19128);
nand U22119 (N_22119,N_20712,N_19658);
or U22120 (N_22120,N_18892,N_19699);
xor U22121 (N_22121,N_20803,N_19985);
or U22122 (N_22122,N_19751,N_20348);
and U22123 (N_22123,N_20775,N_20236);
and U22124 (N_22124,N_20899,N_18135);
nand U22125 (N_22125,N_20979,N_20309);
nor U22126 (N_22126,N_19271,N_19345);
nand U22127 (N_22127,N_20504,N_19602);
xor U22128 (N_22128,N_19448,N_20619);
xor U22129 (N_22129,N_20159,N_19151);
and U22130 (N_22130,N_19656,N_18365);
nand U22131 (N_22131,N_20907,N_19233);
nor U22132 (N_22132,N_20402,N_19275);
or U22133 (N_22133,N_18084,N_18938);
or U22134 (N_22134,N_19112,N_19200);
xnor U22135 (N_22135,N_19554,N_20306);
nand U22136 (N_22136,N_19923,N_18586);
nor U22137 (N_22137,N_19606,N_20556);
xor U22138 (N_22138,N_19413,N_19660);
nor U22139 (N_22139,N_20219,N_20481);
nor U22140 (N_22140,N_19018,N_18505);
nand U22141 (N_22141,N_19984,N_19823);
or U22142 (N_22142,N_18555,N_20065);
nor U22143 (N_22143,N_18845,N_19164);
or U22144 (N_22144,N_19109,N_19251);
and U22145 (N_22145,N_18409,N_18668);
xor U22146 (N_22146,N_18080,N_18019);
or U22147 (N_22147,N_19757,N_19022);
and U22148 (N_22148,N_20313,N_20805);
xnor U22149 (N_22149,N_19059,N_20838);
or U22150 (N_22150,N_18331,N_20249);
xnor U22151 (N_22151,N_19512,N_18871);
or U22152 (N_22152,N_20732,N_19258);
nor U22153 (N_22153,N_18144,N_18920);
and U22154 (N_22154,N_19640,N_19285);
nor U22155 (N_22155,N_18291,N_20914);
nand U22156 (N_22156,N_20759,N_18936);
xnor U22157 (N_22157,N_19867,N_18197);
xor U22158 (N_22158,N_20082,N_20869);
xnor U22159 (N_22159,N_18519,N_20205);
and U22160 (N_22160,N_20975,N_18333);
and U22161 (N_22161,N_18270,N_19816);
nor U22162 (N_22162,N_20804,N_20151);
nand U22163 (N_22163,N_20865,N_19550);
xnor U22164 (N_22164,N_19962,N_18446);
nor U22165 (N_22165,N_18730,N_19750);
nor U22166 (N_22166,N_20812,N_20469);
or U22167 (N_22167,N_20070,N_19357);
or U22168 (N_22168,N_18021,N_19678);
xor U22169 (N_22169,N_20913,N_18939);
or U22170 (N_22170,N_19622,N_19282);
nand U22171 (N_22171,N_20367,N_19772);
or U22172 (N_22172,N_19287,N_20326);
nor U22173 (N_22173,N_19189,N_19442);
and U22174 (N_22174,N_19681,N_19480);
nand U22175 (N_22175,N_18545,N_19547);
or U22176 (N_22176,N_18023,N_20473);
or U22177 (N_22177,N_19125,N_20447);
or U22178 (N_22178,N_18042,N_19428);
nor U22179 (N_22179,N_19396,N_18790);
nand U22180 (N_22180,N_18998,N_20807);
nor U22181 (N_22181,N_19731,N_20191);
and U22182 (N_22182,N_20144,N_18815);
nand U22183 (N_22183,N_20096,N_19177);
nor U22184 (N_22184,N_19240,N_20388);
nor U22185 (N_22185,N_19669,N_19939);
xnor U22186 (N_22186,N_18126,N_19581);
nand U22187 (N_22187,N_20718,N_20090);
nand U22188 (N_22188,N_18006,N_20708);
or U22189 (N_22189,N_18573,N_20103);
xnor U22190 (N_22190,N_19273,N_18887);
nand U22191 (N_22191,N_18321,N_20320);
and U22192 (N_22192,N_18909,N_18764);
nand U22193 (N_22193,N_18958,N_18265);
and U22194 (N_22194,N_20479,N_20570);
nor U22195 (N_22195,N_20864,N_18375);
nor U22196 (N_22196,N_18663,N_19423);
nand U22197 (N_22197,N_18674,N_19078);
or U22198 (N_22198,N_20099,N_18831);
xnor U22199 (N_22199,N_19207,N_19966);
nor U22200 (N_22200,N_19394,N_18380);
or U22201 (N_22201,N_19372,N_19227);
nor U22202 (N_22202,N_20274,N_18681);
xor U22203 (N_22203,N_20303,N_18247);
nand U22204 (N_22204,N_18796,N_19395);
and U22205 (N_22205,N_20810,N_18195);
xnor U22206 (N_22206,N_20627,N_18026);
or U22207 (N_22207,N_18662,N_20941);
nor U22208 (N_22208,N_20956,N_20420);
and U22209 (N_22209,N_19513,N_20394);
and U22210 (N_22210,N_18101,N_20660);
xnor U22211 (N_22211,N_18594,N_18130);
or U22212 (N_22212,N_18368,N_20292);
nand U22213 (N_22213,N_20543,N_20458);
xor U22214 (N_22214,N_19111,N_20587);
nor U22215 (N_22215,N_20207,N_20270);
and U22216 (N_22216,N_18235,N_18004);
nor U22217 (N_22217,N_19981,N_19482);
or U22218 (N_22218,N_20002,N_18706);
or U22219 (N_22219,N_18470,N_18191);
or U22220 (N_22220,N_18323,N_20355);
nor U22221 (N_22221,N_20023,N_18808);
or U22222 (N_22222,N_20101,N_18041);
or U22223 (N_22223,N_18763,N_18284);
nor U22224 (N_22224,N_18211,N_19858);
nand U22225 (N_22225,N_20681,N_18393);
xnor U22226 (N_22226,N_18105,N_19145);
or U22227 (N_22227,N_18214,N_20095);
xnor U22228 (N_22228,N_18874,N_19052);
nand U22229 (N_22229,N_19970,N_20872);
xor U22230 (N_22230,N_18049,N_18872);
or U22231 (N_22231,N_20443,N_18231);
and U22232 (N_22232,N_18203,N_18157);
xor U22233 (N_22233,N_20414,N_18059);
and U22234 (N_22234,N_20177,N_20344);
xor U22235 (N_22235,N_18382,N_18605);
nor U22236 (N_22236,N_18315,N_20364);
and U22237 (N_22237,N_20502,N_18095);
or U22238 (N_22238,N_20347,N_20986);
and U22239 (N_22239,N_20317,N_19831);
or U22240 (N_22240,N_20482,N_19738);
nand U22241 (N_22241,N_19747,N_19594);
xor U22242 (N_22242,N_20206,N_19266);
or U22243 (N_22243,N_18056,N_20756);
or U22244 (N_22244,N_18949,N_19846);
or U22245 (N_22245,N_19978,N_18188);
or U22246 (N_22246,N_19665,N_20768);
nor U22247 (N_22247,N_19348,N_19607);
nand U22248 (N_22248,N_20496,N_20285);
nor U22249 (N_22249,N_18786,N_19170);
nand U22250 (N_22250,N_18862,N_18400);
nor U22251 (N_22251,N_19063,N_19752);
or U22252 (N_22252,N_18608,N_20026);
nor U22253 (N_22253,N_20664,N_20415);
and U22254 (N_22254,N_20057,N_18299);
nand U22255 (N_22255,N_20066,N_18868);
and U22256 (N_22256,N_20723,N_19010);
nand U22257 (N_22257,N_18087,N_19290);
nand U22258 (N_22258,N_20959,N_19826);
xor U22259 (N_22259,N_18278,N_19186);
nor U22260 (N_22260,N_19560,N_20427);
nand U22261 (N_22261,N_20233,N_18357);
or U22262 (N_22262,N_19633,N_18339);
or U22263 (N_22263,N_18804,N_20271);
and U22264 (N_22264,N_20748,N_19901);
xnor U22265 (N_22265,N_19967,N_18288);
or U22266 (N_22266,N_19439,N_20885);
nor U22267 (N_22267,N_19072,N_19191);
and U22268 (N_22268,N_20033,N_20488);
nor U22269 (N_22269,N_18481,N_18370);
xnor U22270 (N_22270,N_19954,N_20252);
nand U22271 (N_22271,N_20250,N_20358);
nor U22272 (N_22272,N_19462,N_18161);
and U22273 (N_22273,N_20742,N_18138);
or U22274 (N_22274,N_20463,N_20288);
nor U22275 (N_22275,N_18040,N_20256);
xor U22276 (N_22276,N_19756,N_20380);
xor U22277 (N_22277,N_19154,N_20290);
or U22278 (N_22278,N_19466,N_19037);
or U22279 (N_22279,N_19156,N_18864);
nor U22280 (N_22280,N_20318,N_20702);
or U22281 (N_22281,N_20777,N_19732);
nor U22282 (N_22282,N_19849,N_18692);
and U22283 (N_22283,N_20544,N_20190);
xnor U22284 (N_22284,N_20517,N_20365);
nor U22285 (N_22285,N_20871,N_20310);
nand U22286 (N_22286,N_19075,N_19314);
or U22287 (N_22287,N_18163,N_19714);
xor U22288 (N_22288,N_20860,N_20392);
or U22289 (N_22289,N_18492,N_19421);
nor U22290 (N_22290,N_20738,N_18208);
xnor U22291 (N_22291,N_20870,N_18224);
nor U22292 (N_22292,N_20499,N_19925);
nor U22293 (N_22293,N_18719,N_20902);
xnor U22294 (N_22294,N_19048,N_18075);
xnor U22295 (N_22295,N_20157,N_19852);
and U22296 (N_22296,N_18894,N_18487);
and U22297 (N_22297,N_18129,N_19229);
and U22298 (N_22298,N_19001,N_20125);
xor U22299 (N_22299,N_19261,N_18508);
nand U22300 (N_22300,N_18897,N_18665);
nand U22301 (N_22301,N_20515,N_18953);
nand U22302 (N_22302,N_19468,N_20962);
or U22303 (N_22303,N_19530,N_18392);
nor U22304 (N_22304,N_19358,N_19373);
xor U22305 (N_22305,N_19706,N_20642);
nand U22306 (N_22306,N_18948,N_20853);
xor U22307 (N_22307,N_18239,N_18898);
or U22308 (N_22308,N_20437,N_18859);
nor U22309 (N_22309,N_20671,N_20404);
xnor U22310 (N_22310,N_19246,N_18748);
xnor U22311 (N_22311,N_19020,N_18419);
nor U22312 (N_22312,N_19484,N_19279);
nand U22313 (N_22313,N_19539,N_18172);
nand U22314 (N_22314,N_18925,N_19545);
or U22315 (N_22315,N_19773,N_20185);
nor U22316 (N_22316,N_19898,N_18676);
or U22317 (N_22317,N_19124,N_20892);
nor U22318 (N_22318,N_19912,N_18910);
or U22319 (N_22319,N_19008,N_19208);
nand U22320 (N_22320,N_19695,N_19791);
nand U22321 (N_22321,N_20168,N_18455);
nand U22322 (N_22322,N_19321,N_19793);
nand U22323 (N_22323,N_18175,N_19107);
nand U22324 (N_22324,N_19374,N_18107);
nand U22325 (N_22325,N_19415,N_19946);
xor U22326 (N_22326,N_18364,N_18245);
nand U22327 (N_22327,N_20453,N_18989);
and U22328 (N_22328,N_18155,N_18462);
nor U22329 (N_22329,N_19236,N_20445);
xnor U22330 (N_22330,N_18395,N_18699);
nand U22331 (N_22331,N_18918,N_20500);
and U22332 (N_22332,N_19631,N_19310);
nor U22333 (N_22333,N_20639,N_19235);
and U22334 (N_22334,N_19409,N_19301);
xnor U22335 (N_22335,N_20954,N_18117);
nand U22336 (N_22336,N_20764,N_20701);
xor U22337 (N_22337,N_20599,N_18233);
nor U22338 (N_22338,N_18955,N_19980);
or U22339 (N_22339,N_20442,N_18833);
xor U22340 (N_22340,N_20085,N_19115);
nand U22341 (N_22341,N_19280,N_19514);
xor U22342 (N_22342,N_20586,N_19930);
nand U22343 (N_22343,N_18561,N_18279);
or U22344 (N_22344,N_18636,N_19211);
and U22345 (N_22345,N_20730,N_19028);
xor U22346 (N_22346,N_19121,N_19908);
and U22347 (N_22347,N_19682,N_20182);
nor U22348 (N_22348,N_19066,N_20581);
nand U22349 (N_22349,N_18709,N_18319);
nor U22350 (N_22350,N_20966,N_19209);
xnor U22351 (N_22351,N_19377,N_19604);
xnor U22352 (N_22352,N_19406,N_19777);
and U22353 (N_22353,N_20056,N_18571);
nor U22354 (N_22354,N_19202,N_20987);
or U22355 (N_22355,N_20973,N_18565);
and U22356 (N_22356,N_20951,N_18689);
and U22357 (N_22357,N_20808,N_18843);
nand U22358 (N_22358,N_18046,N_18151);
nand U22359 (N_22359,N_20615,N_18592);
nand U22360 (N_22360,N_20842,N_19085);
xnor U22361 (N_22361,N_19916,N_18062);
or U22362 (N_22362,N_20906,N_18588);
or U22363 (N_22363,N_18322,N_19217);
or U22364 (N_22364,N_19364,N_18700);
and U22365 (N_22365,N_20778,N_18980);
nor U22366 (N_22366,N_19766,N_18471);
and U22367 (N_22367,N_20226,N_20143);
and U22368 (N_22368,N_20295,N_19634);
nand U22369 (N_22369,N_19926,N_19033);
nand U22370 (N_22370,N_20426,N_20856);
xnor U22371 (N_22371,N_18292,N_20961);
nand U22372 (N_22372,N_19330,N_18475);
nor U22373 (N_22373,N_18458,N_19004);
nand U22374 (N_22374,N_18688,N_20519);
nor U22375 (N_22375,N_18720,N_20135);
xor U22376 (N_22376,N_18215,N_18904);
or U22377 (N_22377,N_20291,N_20837);
nand U22378 (N_22378,N_19140,N_18522);
xor U22379 (N_22379,N_20769,N_19025);
nor U22380 (N_22380,N_20770,N_20875);
xor U22381 (N_22381,N_18311,N_20523);
nand U22382 (N_22382,N_20460,N_20209);
or U22383 (N_22383,N_18944,N_18656);
or U22384 (N_22384,N_18554,N_20197);
nor U22385 (N_22385,N_19526,N_19711);
and U22386 (N_22386,N_18187,N_20170);
and U22387 (N_22387,N_20321,N_20935);
and U22388 (N_22388,N_20416,N_20819);
xor U22389 (N_22389,N_18670,N_18876);
or U22390 (N_22390,N_18836,N_18407);
and U22391 (N_22391,N_18502,N_18883);
and U22392 (N_22392,N_19641,N_18480);
nand U22393 (N_22393,N_20969,N_19587);
xnor U22394 (N_22394,N_20242,N_18972);
or U22395 (N_22395,N_20148,N_19815);
and U22396 (N_22396,N_20631,N_20354);
nor U22397 (N_22397,N_20758,N_19286);
xor U22398 (N_22398,N_19864,N_20595);
nand U22399 (N_22399,N_19101,N_20800);
and U22400 (N_22400,N_18800,N_19329);
and U22401 (N_22401,N_18272,N_19597);
nor U22402 (N_22402,N_18924,N_18312);
nand U22403 (N_22403,N_18354,N_18362);
or U22404 (N_22404,N_19574,N_19401);
nor U22405 (N_22405,N_20516,N_18865);
nand U22406 (N_22406,N_20652,N_19596);
xnor U22407 (N_22407,N_19690,N_18221);
nor U22408 (N_22408,N_19718,N_20814);
and U22409 (N_22409,N_18878,N_19941);
nand U22410 (N_22410,N_18389,N_19017);
nor U22411 (N_22411,N_19042,N_18425);
nor U22412 (N_22412,N_18991,N_18577);
xnor U22413 (N_22413,N_18349,N_19787);
or U22414 (N_22414,N_19957,N_20823);
nand U22415 (N_22415,N_20694,N_19769);
xor U22416 (N_22416,N_18018,N_19005);
xnor U22417 (N_22417,N_18518,N_20626);
xor U22418 (N_22418,N_18691,N_19627);
xnor U22419 (N_22419,N_18816,N_20419);
or U22420 (N_22420,N_19094,N_20690);
nand U22421 (N_22421,N_20161,N_20059);
xor U22422 (N_22422,N_20529,N_20822);
nor U22423 (N_22423,N_20124,N_20518);
nor U22424 (N_22424,N_19768,N_18170);
nor U22425 (N_22425,N_18783,N_18504);
nor U22426 (N_22426,N_19427,N_18642);
xnor U22427 (N_22427,N_18302,N_18976);
nor U22428 (N_22428,N_19878,N_20891);
and U22429 (N_22429,N_19943,N_18212);
nand U22430 (N_22430,N_19588,N_19565);
nand U22431 (N_22431,N_18183,N_20265);
xnor U22432 (N_22432,N_19491,N_20640);
nor U22433 (N_22433,N_19446,N_18440);
and U22434 (N_22434,N_19892,N_19126);
xnor U22435 (N_22435,N_20418,N_19213);
xnor U22436 (N_22436,N_20424,N_18751);
xnor U22437 (N_22437,N_18782,N_18515);
xnor U22438 (N_22438,N_20302,N_18266);
nor U22439 (N_22439,N_18977,N_18020);
xor U22440 (N_22440,N_19621,N_18727);
and U22441 (N_22441,N_20231,N_19643);
xor U22442 (N_22442,N_19889,N_20876);
and U22443 (N_22443,N_20682,N_20610);
nor U22444 (N_22444,N_18598,N_20126);
xnor U22445 (N_22445,N_18246,N_20273);
or U22446 (N_22446,N_20255,N_19742);
and U22447 (N_22447,N_19722,N_19951);
nand U22448 (N_22448,N_18671,N_19155);
nor U22449 (N_22449,N_20081,N_19158);
nand U22450 (N_22450,N_20763,N_20398);
xor U22451 (N_22451,N_19611,N_20359);
xor U22452 (N_22452,N_20400,N_20847);
xor U22453 (N_22453,N_20589,N_20828);
xor U22454 (N_22454,N_19549,N_20435);
or U22455 (N_22455,N_20676,N_19947);
xnor U22456 (N_22456,N_19184,N_18761);
or U22457 (N_22457,N_20006,N_19896);
nor U22458 (N_22458,N_20720,N_20195);
xnor U22459 (N_22459,N_18771,N_19704);
xor U22460 (N_22460,N_20960,N_19561);
nand U22461 (N_22461,N_18542,N_20750);
and U22462 (N_22462,N_18027,N_19855);
nor U22463 (N_22463,N_19103,N_18528);
nand U22464 (N_22464,N_20776,N_19652);
nor U22465 (N_22465,N_19869,N_19369);
and U22466 (N_22466,N_18556,N_19522);
and U22467 (N_22467,N_20634,N_20811);
xor U22468 (N_22468,N_20506,N_19698);
or U22469 (N_22469,N_18088,N_20264);
xnor U22470 (N_22470,N_20739,N_18707);
nand U22471 (N_22471,N_18905,N_18249);
xnor U22472 (N_22472,N_20666,N_19801);
or U22473 (N_22473,N_18776,N_18762);
nand U22474 (N_22474,N_18307,N_20590);
or U22475 (N_22475,N_20670,N_19723);
nor U22476 (N_22476,N_19461,N_19636);
xnor U22477 (N_22477,N_20431,N_20149);
nand U22478 (N_22478,N_18744,N_19685);
and U22479 (N_22479,N_19708,N_18048);
xnor U22480 (N_22480,N_18648,N_20752);
nor U22481 (N_22481,N_19879,N_18983);
nand U22482 (N_22482,N_18277,N_18882);
nand U22483 (N_22483,N_20356,N_20186);
or U22484 (N_22484,N_20612,N_19381);
and U22485 (N_22485,N_18787,N_19331);
and U22486 (N_22486,N_20062,N_19525);
and U22487 (N_22487,N_19818,N_20379);
and U22488 (N_22488,N_18180,N_19808);
nor U22489 (N_22489,N_20573,N_19360);
xor U22490 (N_22490,N_20849,N_19359);
xnor U22491 (N_22491,N_19883,N_20459);
nand U22492 (N_22492,N_20120,N_20675);
nand U22493 (N_22493,N_19586,N_19248);
nand U22494 (N_22494,N_18378,N_20201);
or U22495 (N_22495,N_18774,N_19890);
and U22496 (N_22496,N_18890,N_20992);
nand U22497 (N_22497,N_19159,N_20433);
and U22498 (N_22498,N_20486,N_20340);
nor U22499 (N_22499,N_18332,N_20014);
and U22500 (N_22500,N_20992,N_18857);
xnor U22501 (N_22501,N_18034,N_18480);
xor U22502 (N_22502,N_19590,N_20892);
and U22503 (N_22503,N_19585,N_19767);
nand U22504 (N_22504,N_18822,N_19449);
and U22505 (N_22505,N_19644,N_20326);
nand U22506 (N_22506,N_19942,N_19624);
nor U22507 (N_22507,N_18287,N_18305);
nand U22508 (N_22508,N_18232,N_19829);
xor U22509 (N_22509,N_18782,N_18099);
xor U22510 (N_22510,N_18361,N_20920);
xor U22511 (N_22511,N_20666,N_20980);
nor U22512 (N_22512,N_19845,N_20738);
nand U22513 (N_22513,N_18581,N_18056);
and U22514 (N_22514,N_18375,N_19131);
nand U22515 (N_22515,N_19283,N_20400);
nor U22516 (N_22516,N_18187,N_20743);
nand U22517 (N_22517,N_19573,N_19755);
nand U22518 (N_22518,N_18250,N_19667);
nor U22519 (N_22519,N_18333,N_20562);
xnor U22520 (N_22520,N_18903,N_19478);
or U22521 (N_22521,N_19258,N_20676);
or U22522 (N_22522,N_18537,N_18329);
xor U22523 (N_22523,N_20860,N_18754);
nor U22524 (N_22524,N_18326,N_19606);
and U22525 (N_22525,N_18868,N_20302);
nand U22526 (N_22526,N_19364,N_19480);
and U22527 (N_22527,N_18501,N_20322);
and U22528 (N_22528,N_18005,N_20345);
and U22529 (N_22529,N_18971,N_18218);
and U22530 (N_22530,N_19468,N_20073);
and U22531 (N_22531,N_20919,N_19370);
or U22532 (N_22532,N_18304,N_18337);
or U22533 (N_22533,N_19128,N_18899);
nand U22534 (N_22534,N_20068,N_18515);
xnor U22535 (N_22535,N_20036,N_20700);
nor U22536 (N_22536,N_19216,N_20703);
nand U22537 (N_22537,N_20565,N_20230);
or U22538 (N_22538,N_20984,N_20047);
xnor U22539 (N_22539,N_20998,N_20516);
nand U22540 (N_22540,N_19569,N_20453);
nand U22541 (N_22541,N_19720,N_18454);
nor U22542 (N_22542,N_19620,N_18548);
and U22543 (N_22543,N_20658,N_18068);
nor U22544 (N_22544,N_18258,N_18279);
or U22545 (N_22545,N_18088,N_19374);
or U22546 (N_22546,N_18918,N_20101);
nand U22547 (N_22547,N_20896,N_18517);
nand U22548 (N_22548,N_18669,N_20230);
or U22549 (N_22549,N_19795,N_20468);
or U22550 (N_22550,N_19123,N_20386);
xor U22551 (N_22551,N_19011,N_18675);
nand U22552 (N_22552,N_18522,N_18731);
nand U22553 (N_22553,N_20989,N_19640);
xor U22554 (N_22554,N_20067,N_20127);
or U22555 (N_22555,N_18708,N_19433);
nor U22556 (N_22556,N_18275,N_19855);
xnor U22557 (N_22557,N_20701,N_19164);
nor U22558 (N_22558,N_18761,N_19560);
or U22559 (N_22559,N_20301,N_19204);
xnor U22560 (N_22560,N_19308,N_19169);
or U22561 (N_22561,N_19585,N_20096);
nand U22562 (N_22562,N_18916,N_20606);
xnor U22563 (N_22563,N_20080,N_20417);
nand U22564 (N_22564,N_18786,N_20782);
or U22565 (N_22565,N_20289,N_18108);
nand U22566 (N_22566,N_20135,N_18451);
or U22567 (N_22567,N_19979,N_18437);
nand U22568 (N_22568,N_19286,N_20932);
nor U22569 (N_22569,N_20131,N_18729);
nand U22570 (N_22570,N_18238,N_19152);
nor U22571 (N_22571,N_18079,N_20002);
and U22572 (N_22572,N_20143,N_18025);
xor U22573 (N_22573,N_18522,N_20090);
or U22574 (N_22574,N_19237,N_19493);
and U22575 (N_22575,N_18759,N_20501);
xor U22576 (N_22576,N_20139,N_18733);
or U22577 (N_22577,N_19752,N_19780);
nand U22578 (N_22578,N_20182,N_18337);
and U22579 (N_22579,N_20430,N_20116);
and U22580 (N_22580,N_20038,N_20695);
xnor U22581 (N_22581,N_18887,N_20041);
and U22582 (N_22582,N_19563,N_18792);
and U22583 (N_22583,N_20688,N_19853);
nand U22584 (N_22584,N_19519,N_20499);
nand U22585 (N_22585,N_18390,N_19863);
xnor U22586 (N_22586,N_20181,N_20855);
xnor U22587 (N_22587,N_20814,N_19741);
nor U22588 (N_22588,N_19749,N_20435);
and U22589 (N_22589,N_20961,N_20212);
xnor U22590 (N_22590,N_18842,N_20175);
nand U22591 (N_22591,N_20069,N_18122);
nor U22592 (N_22592,N_20639,N_18074);
and U22593 (N_22593,N_19589,N_19112);
nand U22594 (N_22594,N_19318,N_19569);
xor U22595 (N_22595,N_18317,N_20756);
or U22596 (N_22596,N_19726,N_19212);
and U22597 (N_22597,N_20246,N_20200);
nor U22598 (N_22598,N_20893,N_18087);
xor U22599 (N_22599,N_18269,N_18143);
xnor U22600 (N_22600,N_20458,N_18622);
and U22601 (N_22601,N_19686,N_19847);
xnor U22602 (N_22602,N_20064,N_19626);
nand U22603 (N_22603,N_19584,N_18776);
nand U22604 (N_22604,N_18640,N_20057);
nor U22605 (N_22605,N_19267,N_19862);
or U22606 (N_22606,N_20201,N_19073);
and U22607 (N_22607,N_18969,N_18562);
nor U22608 (N_22608,N_19697,N_18270);
xor U22609 (N_22609,N_18697,N_19144);
nor U22610 (N_22610,N_20938,N_20875);
nor U22611 (N_22611,N_20587,N_19456);
nor U22612 (N_22612,N_18177,N_18712);
or U22613 (N_22613,N_18807,N_18630);
xor U22614 (N_22614,N_20843,N_20459);
nand U22615 (N_22615,N_18203,N_19421);
or U22616 (N_22616,N_20593,N_18682);
or U22617 (N_22617,N_20853,N_19634);
nand U22618 (N_22618,N_20705,N_19520);
or U22619 (N_22619,N_19461,N_18892);
xnor U22620 (N_22620,N_19228,N_19694);
xnor U22621 (N_22621,N_18308,N_20437);
and U22622 (N_22622,N_19965,N_20030);
and U22623 (N_22623,N_20860,N_20493);
or U22624 (N_22624,N_19518,N_18122);
or U22625 (N_22625,N_19497,N_18058);
or U22626 (N_22626,N_18376,N_20648);
xnor U22627 (N_22627,N_19795,N_20905);
or U22628 (N_22628,N_18546,N_20187);
nand U22629 (N_22629,N_19929,N_18785);
xnor U22630 (N_22630,N_18068,N_20835);
or U22631 (N_22631,N_20909,N_18184);
or U22632 (N_22632,N_20842,N_20910);
nand U22633 (N_22633,N_18677,N_20208);
nor U22634 (N_22634,N_19864,N_20382);
and U22635 (N_22635,N_19065,N_18451);
xor U22636 (N_22636,N_19285,N_20805);
nand U22637 (N_22637,N_19214,N_20393);
nand U22638 (N_22638,N_20124,N_19864);
nor U22639 (N_22639,N_18391,N_20292);
and U22640 (N_22640,N_18305,N_19333);
nor U22641 (N_22641,N_20975,N_19149);
nand U22642 (N_22642,N_20984,N_18559);
and U22643 (N_22643,N_20185,N_18360);
and U22644 (N_22644,N_19662,N_18404);
xnor U22645 (N_22645,N_18953,N_18617);
xnor U22646 (N_22646,N_18635,N_19300);
nor U22647 (N_22647,N_20334,N_20285);
and U22648 (N_22648,N_19305,N_18379);
nor U22649 (N_22649,N_19695,N_19303);
nand U22650 (N_22650,N_20913,N_20511);
nand U22651 (N_22651,N_19248,N_20757);
nor U22652 (N_22652,N_18727,N_19789);
nor U22653 (N_22653,N_18658,N_20038);
xor U22654 (N_22654,N_19905,N_20504);
nor U22655 (N_22655,N_20753,N_19286);
nor U22656 (N_22656,N_18401,N_20482);
and U22657 (N_22657,N_20472,N_18513);
nand U22658 (N_22658,N_18344,N_19217);
xnor U22659 (N_22659,N_18977,N_19644);
nand U22660 (N_22660,N_20747,N_20617);
nor U22661 (N_22661,N_20386,N_18044);
nor U22662 (N_22662,N_18747,N_18855);
nor U22663 (N_22663,N_20169,N_18137);
and U22664 (N_22664,N_18987,N_18739);
and U22665 (N_22665,N_19090,N_18440);
xnor U22666 (N_22666,N_20439,N_20281);
nor U22667 (N_22667,N_19820,N_19837);
and U22668 (N_22668,N_19497,N_19099);
or U22669 (N_22669,N_18498,N_19669);
and U22670 (N_22670,N_19728,N_20808);
and U22671 (N_22671,N_20462,N_19919);
or U22672 (N_22672,N_19327,N_20879);
nand U22673 (N_22673,N_20202,N_18019);
xnor U22674 (N_22674,N_19041,N_18300);
nor U22675 (N_22675,N_19137,N_19592);
xor U22676 (N_22676,N_18853,N_18631);
xnor U22677 (N_22677,N_19077,N_20150);
and U22678 (N_22678,N_18294,N_19729);
xor U22679 (N_22679,N_20238,N_19827);
nor U22680 (N_22680,N_19508,N_18450);
xor U22681 (N_22681,N_19133,N_18428);
and U22682 (N_22682,N_18874,N_18000);
nor U22683 (N_22683,N_18121,N_19066);
nand U22684 (N_22684,N_19198,N_18035);
and U22685 (N_22685,N_19604,N_19508);
xnor U22686 (N_22686,N_18397,N_18335);
or U22687 (N_22687,N_19278,N_20351);
xnor U22688 (N_22688,N_18825,N_18860);
and U22689 (N_22689,N_19483,N_18302);
and U22690 (N_22690,N_20712,N_18065);
nor U22691 (N_22691,N_20126,N_20662);
nor U22692 (N_22692,N_19335,N_20823);
nand U22693 (N_22693,N_20209,N_20385);
and U22694 (N_22694,N_20086,N_18983);
or U22695 (N_22695,N_18986,N_20676);
nand U22696 (N_22696,N_19742,N_18746);
nor U22697 (N_22697,N_18471,N_20271);
or U22698 (N_22698,N_18963,N_19229);
xnor U22699 (N_22699,N_19244,N_19002);
and U22700 (N_22700,N_19823,N_19103);
and U22701 (N_22701,N_20277,N_20214);
or U22702 (N_22702,N_18166,N_20198);
or U22703 (N_22703,N_19126,N_19719);
and U22704 (N_22704,N_20389,N_20320);
and U22705 (N_22705,N_19061,N_20047);
and U22706 (N_22706,N_19014,N_18985);
and U22707 (N_22707,N_20011,N_20729);
xor U22708 (N_22708,N_18080,N_18885);
nor U22709 (N_22709,N_19610,N_18025);
nand U22710 (N_22710,N_19343,N_18429);
nand U22711 (N_22711,N_19228,N_18003);
nand U22712 (N_22712,N_19211,N_19303);
and U22713 (N_22713,N_18505,N_19984);
nand U22714 (N_22714,N_18935,N_18552);
nand U22715 (N_22715,N_19645,N_20601);
xor U22716 (N_22716,N_18317,N_18588);
nand U22717 (N_22717,N_18345,N_18380);
nand U22718 (N_22718,N_20663,N_20110);
nor U22719 (N_22719,N_18374,N_18318);
xnor U22720 (N_22720,N_20149,N_18552);
nand U22721 (N_22721,N_19110,N_20532);
xor U22722 (N_22722,N_19968,N_20602);
or U22723 (N_22723,N_19152,N_20998);
and U22724 (N_22724,N_20067,N_19252);
or U22725 (N_22725,N_18935,N_19858);
xor U22726 (N_22726,N_20756,N_18478);
nand U22727 (N_22727,N_20465,N_20020);
xor U22728 (N_22728,N_19885,N_19284);
or U22729 (N_22729,N_18966,N_20846);
and U22730 (N_22730,N_19534,N_20584);
or U22731 (N_22731,N_18233,N_20508);
xor U22732 (N_22732,N_19784,N_19483);
nor U22733 (N_22733,N_19243,N_18366);
and U22734 (N_22734,N_20769,N_19951);
or U22735 (N_22735,N_18944,N_20550);
and U22736 (N_22736,N_19373,N_19450);
nand U22737 (N_22737,N_19735,N_20520);
nand U22738 (N_22738,N_19255,N_18628);
or U22739 (N_22739,N_18457,N_20965);
xor U22740 (N_22740,N_20275,N_19585);
or U22741 (N_22741,N_20375,N_19835);
and U22742 (N_22742,N_20176,N_18345);
nor U22743 (N_22743,N_18591,N_18193);
and U22744 (N_22744,N_19875,N_18212);
nor U22745 (N_22745,N_18641,N_19237);
xnor U22746 (N_22746,N_20110,N_20104);
nor U22747 (N_22747,N_19666,N_19735);
or U22748 (N_22748,N_19159,N_19443);
nor U22749 (N_22749,N_20835,N_18914);
nand U22750 (N_22750,N_20610,N_20305);
or U22751 (N_22751,N_18160,N_20113);
and U22752 (N_22752,N_19590,N_18918);
and U22753 (N_22753,N_19014,N_18168);
or U22754 (N_22754,N_19297,N_19954);
nor U22755 (N_22755,N_20183,N_20871);
and U22756 (N_22756,N_19845,N_18143);
xor U22757 (N_22757,N_19569,N_18877);
and U22758 (N_22758,N_20199,N_18941);
and U22759 (N_22759,N_20626,N_18861);
nor U22760 (N_22760,N_20905,N_20545);
or U22761 (N_22761,N_20419,N_18880);
xor U22762 (N_22762,N_20337,N_19394);
xnor U22763 (N_22763,N_19712,N_20633);
nand U22764 (N_22764,N_19977,N_19734);
and U22765 (N_22765,N_20603,N_18641);
and U22766 (N_22766,N_20424,N_18916);
or U22767 (N_22767,N_19240,N_18106);
and U22768 (N_22768,N_20685,N_18783);
nor U22769 (N_22769,N_18969,N_19668);
xnor U22770 (N_22770,N_19035,N_18068);
xnor U22771 (N_22771,N_18265,N_19622);
or U22772 (N_22772,N_19753,N_18570);
or U22773 (N_22773,N_19408,N_18983);
nand U22774 (N_22774,N_20879,N_18032);
xor U22775 (N_22775,N_18623,N_18966);
nor U22776 (N_22776,N_18753,N_20273);
nor U22777 (N_22777,N_19733,N_18659);
nor U22778 (N_22778,N_19427,N_19525);
and U22779 (N_22779,N_20363,N_19245);
or U22780 (N_22780,N_18796,N_20848);
nand U22781 (N_22781,N_18888,N_20292);
nand U22782 (N_22782,N_20149,N_18328);
and U22783 (N_22783,N_18051,N_19868);
or U22784 (N_22784,N_18935,N_18272);
nand U22785 (N_22785,N_19917,N_20315);
xnor U22786 (N_22786,N_19781,N_20565);
xor U22787 (N_22787,N_18969,N_19223);
or U22788 (N_22788,N_19273,N_19392);
and U22789 (N_22789,N_19159,N_19901);
nand U22790 (N_22790,N_19339,N_19892);
nor U22791 (N_22791,N_18652,N_20300);
and U22792 (N_22792,N_20234,N_18098);
or U22793 (N_22793,N_18345,N_20946);
nor U22794 (N_22794,N_19462,N_19878);
nand U22795 (N_22795,N_20218,N_18275);
and U22796 (N_22796,N_19369,N_19502);
nor U22797 (N_22797,N_18824,N_19265);
nor U22798 (N_22798,N_20127,N_20933);
xor U22799 (N_22799,N_19568,N_20837);
or U22800 (N_22800,N_20880,N_20501);
nand U22801 (N_22801,N_20786,N_20193);
xnor U22802 (N_22802,N_20709,N_20229);
nor U22803 (N_22803,N_19955,N_20780);
xnor U22804 (N_22804,N_19273,N_19420);
xor U22805 (N_22805,N_18318,N_20894);
nor U22806 (N_22806,N_20313,N_18392);
or U22807 (N_22807,N_19290,N_20643);
and U22808 (N_22808,N_19681,N_19589);
xnor U22809 (N_22809,N_19348,N_20162);
and U22810 (N_22810,N_18042,N_18018);
or U22811 (N_22811,N_19267,N_18810);
xor U22812 (N_22812,N_20903,N_20301);
nor U22813 (N_22813,N_19123,N_19672);
or U22814 (N_22814,N_19129,N_18293);
or U22815 (N_22815,N_19459,N_19953);
and U22816 (N_22816,N_18807,N_18166);
nand U22817 (N_22817,N_20667,N_19073);
xor U22818 (N_22818,N_18633,N_19631);
or U22819 (N_22819,N_20026,N_20206);
nor U22820 (N_22820,N_18226,N_20193);
xor U22821 (N_22821,N_19534,N_19617);
xor U22822 (N_22822,N_20078,N_18862);
nor U22823 (N_22823,N_19948,N_19777);
nor U22824 (N_22824,N_19918,N_18847);
nor U22825 (N_22825,N_18913,N_20916);
or U22826 (N_22826,N_19940,N_20675);
or U22827 (N_22827,N_20834,N_18506);
or U22828 (N_22828,N_20453,N_18455);
nand U22829 (N_22829,N_20054,N_19665);
xor U22830 (N_22830,N_19827,N_18295);
nand U22831 (N_22831,N_18707,N_18022);
and U22832 (N_22832,N_19431,N_19384);
nand U22833 (N_22833,N_19675,N_18275);
nand U22834 (N_22834,N_19510,N_18163);
nand U22835 (N_22835,N_20315,N_18175);
nor U22836 (N_22836,N_19114,N_20039);
and U22837 (N_22837,N_18950,N_18954);
nor U22838 (N_22838,N_20906,N_18696);
xnor U22839 (N_22839,N_19341,N_19996);
xor U22840 (N_22840,N_18205,N_19976);
nor U22841 (N_22841,N_18134,N_19840);
nor U22842 (N_22842,N_20164,N_18113);
nand U22843 (N_22843,N_19319,N_20032);
and U22844 (N_22844,N_20692,N_20787);
nor U22845 (N_22845,N_20294,N_20478);
nand U22846 (N_22846,N_18566,N_19584);
xor U22847 (N_22847,N_18524,N_18919);
and U22848 (N_22848,N_18766,N_18961);
and U22849 (N_22849,N_20446,N_20331);
xor U22850 (N_22850,N_18162,N_20177);
and U22851 (N_22851,N_18325,N_18896);
or U22852 (N_22852,N_19596,N_19232);
or U22853 (N_22853,N_19536,N_18630);
and U22854 (N_22854,N_20210,N_19460);
nor U22855 (N_22855,N_18588,N_18902);
nor U22856 (N_22856,N_18710,N_20187);
nor U22857 (N_22857,N_19169,N_20237);
xor U22858 (N_22858,N_18920,N_19919);
nand U22859 (N_22859,N_18302,N_18416);
xnor U22860 (N_22860,N_20731,N_19350);
or U22861 (N_22861,N_19978,N_19882);
nand U22862 (N_22862,N_20866,N_20347);
or U22863 (N_22863,N_20349,N_20660);
nand U22864 (N_22864,N_18962,N_19882);
xnor U22865 (N_22865,N_18982,N_18050);
nand U22866 (N_22866,N_18112,N_20910);
nand U22867 (N_22867,N_20619,N_19294);
xnor U22868 (N_22868,N_18884,N_19540);
nand U22869 (N_22869,N_20708,N_20152);
or U22870 (N_22870,N_19563,N_18406);
and U22871 (N_22871,N_18372,N_19910);
nand U22872 (N_22872,N_18386,N_19061);
or U22873 (N_22873,N_20048,N_19821);
nand U22874 (N_22874,N_19226,N_19523);
xor U22875 (N_22875,N_20379,N_20629);
nor U22876 (N_22876,N_18681,N_20075);
xnor U22877 (N_22877,N_19725,N_18114);
xor U22878 (N_22878,N_18781,N_19380);
nand U22879 (N_22879,N_20696,N_20721);
and U22880 (N_22880,N_20646,N_18445);
or U22881 (N_22881,N_20266,N_19954);
or U22882 (N_22882,N_20448,N_20885);
nor U22883 (N_22883,N_18477,N_19249);
nand U22884 (N_22884,N_18091,N_18331);
and U22885 (N_22885,N_18114,N_20201);
nand U22886 (N_22886,N_20540,N_18998);
or U22887 (N_22887,N_18233,N_19074);
xnor U22888 (N_22888,N_19481,N_20838);
nor U22889 (N_22889,N_19768,N_19851);
and U22890 (N_22890,N_18613,N_18558);
or U22891 (N_22891,N_18325,N_18681);
nand U22892 (N_22892,N_18390,N_20234);
or U22893 (N_22893,N_19131,N_20529);
nor U22894 (N_22894,N_18951,N_19480);
xnor U22895 (N_22895,N_18153,N_20163);
or U22896 (N_22896,N_20202,N_20661);
nand U22897 (N_22897,N_19874,N_18828);
xor U22898 (N_22898,N_19010,N_18194);
nor U22899 (N_22899,N_18777,N_19677);
nor U22900 (N_22900,N_19223,N_19676);
or U22901 (N_22901,N_19782,N_20275);
or U22902 (N_22902,N_18608,N_20903);
and U22903 (N_22903,N_18062,N_20373);
nor U22904 (N_22904,N_18563,N_19639);
nand U22905 (N_22905,N_19069,N_19955);
nor U22906 (N_22906,N_19745,N_19961);
nand U22907 (N_22907,N_19667,N_19446);
nand U22908 (N_22908,N_18758,N_20722);
nand U22909 (N_22909,N_18917,N_20885);
nand U22910 (N_22910,N_20345,N_20095);
and U22911 (N_22911,N_18589,N_20970);
xor U22912 (N_22912,N_19688,N_19059);
and U22913 (N_22913,N_18747,N_19783);
or U22914 (N_22914,N_18731,N_20391);
xnor U22915 (N_22915,N_20198,N_18986);
or U22916 (N_22916,N_19388,N_19655);
nor U22917 (N_22917,N_20060,N_19515);
nor U22918 (N_22918,N_20390,N_18245);
nor U22919 (N_22919,N_19753,N_18109);
xor U22920 (N_22920,N_18133,N_20111);
or U22921 (N_22921,N_20044,N_18113);
nor U22922 (N_22922,N_20639,N_19470);
or U22923 (N_22923,N_19418,N_20812);
xor U22924 (N_22924,N_19094,N_18879);
nand U22925 (N_22925,N_18437,N_18345);
or U22926 (N_22926,N_18008,N_19121);
xnor U22927 (N_22927,N_20703,N_20484);
xor U22928 (N_22928,N_19284,N_19012);
xnor U22929 (N_22929,N_19285,N_19621);
or U22930 (N_22930,N_20339,N_18552);
nand U22931 (N_22931,N_18645,N_20907);
nand U22932 (N_22932,N_18136,N_18818);
xor U22933 (N_22933,N_18321,N_20354);
nand U22934 (N_22934,N_18703,N_20813);
nor U22935 (N_22935,N_19838,N_18400);
and U22936 (N_22936,N_19923,N_18143);
xor U22937 (N_22937,N_20528,N_20300);
nor U22938 (N_22938,N_20991,N_19436);
and U22939 (N_22939,N_19560,N_19399);
or U22940 (N_22940,N_18060,N_18869);
and U22941 (N_22941,N_18137,N_18321);
nor U22942 (N_22942,N_20131,N_19660);
xnor U22943 (N_22943,N_19545,N_19769);
nor U22944 (N_22944,N_20447,N_18657);
xor U22945 (N_22945,N_20716,N_18113);
xnor U22946 (N_22946,N_20401,N_20545);
nand U22947 (N_22947,N_20935,N_19939);
or U22948 (N_22948,N_19086,N_18485);
xor U22949 (N_22949,N_19043,N_20528);
nand U22950 (N_22950,N_19915,N_19294);
nor U22951 (N_22951,N_18202,N_19831);
and U22952 (N_22952,N_20710,N_20149);
xnor U22953 (N_22953,N_19428,N_18586);
and U22954 (N_22954,N_18191,N_18325);
nor U22955 (N_22955,N_19737,N_19394);
xor U22956 (N_22956,N_20670,N_18508);
xor U22957 (N_22957,N_19019,N_19646);
nand U22958 (N_22958,N_20742,N_19718);
xor U22959 (N_22959,N_19516,N_19905);
nand U22960 (N_22960,N_19687,N_19084);
xnor U22961 (N_22961,N_18892,N_19735);
nor U22962 (N_22962,N_19065,N_20636);
xor U22963 (N_22963,N_18068,N_18343);
nand U22964 (N_22964,N_19535,N_19987);
or U22965 (N_22965,N_18899,N_19415);
xnor U22966 (N_22966,N_18787,N_19978);
xor U22967 (N_22967,N_18126,N_19929);
xnor U22968 (N_22968,N_18907,N_20670);
and U22969 (N_22969,N_19647,N_19604);
and U22970 (N_22970,N_18637,N_19250);
and U22971 (N_22971,N_20800,N_19888);
xor U22972 (N_22972,N_19079,N_18388);
nand U22973 (N_22973,N_18645,N_18878);
or U22974 (N_22974,N_20453,N_19261);
and U22975 (N_22975,N_19626,N_18430);
nor U22976 (N_22976,N_20801,N_18258);
nor U22977 (N_22977,N_18569,N_19843);
xnor U22978 (N_22978,N_18569,N_18191);
nand U22979 (N_22979,N_18567,N_19399);
xor U22980 (N_22980,N_18273,N_20798);
xnor U22981 (N_22981,N_18425,N_19272);
nor U22982 (N_22982,N_18067,N_18602);
and U22983 (N_22983,N_19271,N_20894);
or U22984 (N_22984,N_20851,N_19794);
or U22985 (N_22985,N_20711,N_18182);
and U22986 (N_22986,N_20657,N_20696);
or U22987 (N_22987,N_20093,N_20802);
nand U22988 (N_22988,N_18788,N_19860);
xnor U22989 (N_22989,N_18042,N_19537);
and U22990 (N_22990,N_19043,N_18903);
nand U22991 (N_22991,N_19639,N_18842);
nand U22992 (N_22992,N_20174,N_19703);
nand U22993 (N_22993,N_18417,N_18066);
xor U22994 (N_22994,N_18266,N_18377);
nand U22995 (N_22995,N_18214,N_20908);
and U22996 (N_22996,N_20546,N_19967);
and U22997 (N_22997,N_18560,N_20527);
nand U22998 (N_22998,N_20052,N_19294);
xor U22999 (N_22999,N_18972,N_18684);
and U23000 (N_23000,N_19189,N_20988);
xor U23001 (N_23001,N_20170,N_19355);
nand U23002 (N_23002,N_19041,N_20857);
and U23003 (N_23003,N_20019,N_18986);
or U23004 (N_23004,N_19177,N_19687);
and U23005 (N_23005,N_18771,N_19061);
nand U23006 (N_23006,N_19333,N_18438);
xnor U23007 (N_23007,N_19164,N_20898);
nor U23008 (N_23008,N_19287,N_20968);
or U23009 (N_23009,N_19950,N_18108);
or U23010 (N_23010,N_20563,N_20801);
and U23011 (N_23011,N_20082,N_20516);
nor U23012 (N_23012,N_18112,N_20669);
nor U23013 (N_23013,N_19914,N_18721);
and U23014 (N_23014,N_20315,N_18186);
and U23015 (N_23015,N_19164,N_19619);
and U23016 (N_23016,N_19862,N_20630);
nand U23017 (N_23017,N_18211,N_19948);
xnor U23018 (N_23018,N_19401,N_18070);
and U23019 (N_23019,N_19720,N_18465);
nor U23020 (N_23020,N_20377,N_18161);
or U23021 (N_23021,N_19212,N_18450);
nand U23022 (N_23022,N_18628,N_18671);
nor U23023 (N_23023,N_19259,N_20260);
nand U23024 (N_23024,N_20074,N_19614);
xor U23025 (N_23025,N_19590,N_20219);
xor U23026 (N_23026,N_20712,N_19004);
xnor U23027 (N_23027,N_19469,N_18923);
and U23028 (N_23028,N_18939,N_19031);
nor U23029 (N_23029,N_20994,N_20381);
and U23030 (N_23030,N_18388,N_19208);
and U23031 (N_23031,N_19027,N_18639);
nor U23032 (N_23032,N_19359,N_20564);
nand U23033 (N_23033,N_19567,N_18782);
nor U23034 (N_23034,N_18271,N_20172);
xor U23035 (N_23035,N_19932,N_19259);
or U23036 (N_23036,N_19137,N_20928);
xnor U23037 (N_23037,N_20487,N_20546);
and U23038 (N_23038,N_20914,N_19752);
nor U23039 (N_23039,N_20477,N_19508);
nand U23040 (N_23040,N_19797,N_20917);
nand U23041 (N_23041,N_20280,N_19349);
xor U23042 (N_23042,N_18320,N_20109);
and U23043 (N_23043,N_19551,N_18076);
nand U23044 (N_23044,N_18380,N_18978);
and U23045 (N_23045,N_19508,N_18653);
nand U23046 (N_23046,N_19058,N_20414);
nand U23047 (N_23047,N_18908,N_20251);
xor U23048 (N_23048,N_18569,N_19926);
and U23049 (N_23049,N_18375,N_20901);
nand U23050 (N_23050,N_20210,N_19075);
and U23051 (N_23051,N_18771,N_18705);
xnor U23052 (N_23052,N_20066,N_20630);
nand U23053 (N_23053,N_20085,N_20262);
and U23054 (N_23054,N_20892,N_20634);
or U23055 (N_23055,N_18092,N_20548);
or U23056 (N_23056,N_18405,N_20012);
and U23057 (N_23057,N_20845,N_20172);
nor U23058 (N_23058,N_19745,N_19277);
and U23059 (N_23059,N_19818,N_18612);
nand U23060 (N_23060,N_19257,N_20574);
and U23061 (N_23061,N_18544,N_18794);
xor U23062 (N_23062,N_18592,N_18511);
nand U23063 (N_23063,N_18983,N_20002);
or U23064 (N_23064,N_20541,N_18628);
xor U23065 (N_23065,N_18406,N_19385);
xor U23066 (N_23066,N_18969,N_18117);
nor U23067 (N_23067,N_18798,N_20476);
nand U23068 (N_23068,N_18184,N_19925);
or U23069 (N_23069,N_18888,N_18645);
xnor U23070 (N_23070,N_18700,N_19851);
or U23071 (N_23071,N_18361,N_20903);
or U23072 (N_23072,N_20649,N_18746);
or U23073 (N_23073,N_19394,N_18403);
nor U23074 (N_23074,N_20532,N_18187);
or U23075 (N_23075,N_19530,N_19678);
nor U23076 (N_23076,N_18863,N_19954);
nand U23077 (N_23077,N_20075,N_18829);
xor U23078 (N_23078,N_18479,N_20909);
xnor U23079 (N_23079,N_20456,N_18744);
nand U23080 (N_23080,N_20033,N_19906);
nor U23081 (N_23081,N_20461,N_19456);
xor U23082 (N_23082,N_18931,N_18076);
and U23083 (N_23083,N_18740,N_18948);
or U23084 (N_23084,N_20231,N_19347);
and U23085 (N_23085,N_18883,N_19781);
xnor U23086 (N_23086,N_18513,N_18461);
nand U23087 (N_23087,N_19990,N_18210);
and U23088 (N_23088,N_18326,N_18321);
xnor U23089 (N_23089,N_20983,N_20894);
or U23090 (N_23090,N_20025,N_20832);
xor U23091 (N_23091,N_18220,N_18615);
and U23092 (N_23092,N_18587,N_20346);
and U23093 (N_23093,N_20092,N_19462);
nor U23094 (N_23094,N_18371,N_18231);
nand U23095 (N_23095,N_18611,N_18685);
nand U23096 (N_23096,N_18120,N_18996);
xnor U23097 (N_23097,N_20232,N_19286);
xor U23098 (N_23098,N_19119,N_19567);
or U23099 (N_23099,N_18227,N_19063);
nor U23100 (N_23100,N_18358,N_19377);
nor U23101 (N_23101,N_20977,N_18384);
and U23102 (N_23102,N_18666,N_19093);
nor U23103 (N_23103,N_19822,N_20329);
nor U23104 (N_23104,N_18106,N_18160);
or U23105 (N_23105,N_20927,N_19371);
or U23106 (N_23106,N_20267,N_19737);
xnor U23107 (N_23107,N_20604,N_19632);
or U23108 (N_23108,N_20034,N_20628);
xnor U23109 (N_23109,N_19324,N_20799);
and U23110 (N_23110,N_18019,N_18786);
and U23111 (N_23111,N_18523,N_18283);
nor U23112 (N_23112,N_19304,N_19229);
xnor U23113 (N_23113,N_18017,N_18069);
nand U23114 (N_23114,N_20880,N_19816);
or U23115 (N_23115,N_19214,N_19563);
nand U23116 (N_23116,N_20554,N_19517);
nor U23117 (N_23117,N_20807,N_18817);
nand U23118 (N_23118,N_19726,N_20862);
xnor U23119 (N_23119,N_19946,N_20258);
nor U23120 (N_23120,N_18958,N_18229);
xnor U23121 (N_23121,N_19445,N_18712);
and U23122 (N_23122,N_18677,N_18016);
and U23123 (N_23123,N_18449,N_19684);
nor U23124 (N_23124,N_18963,N_20154);
nand U23125 (N_23125,N_19292,N_19673);
nand U23126 (N_23126,N_18588,N_19182);
nand U23127 (N_23127,N_19682,N_19914);
xor U23128 (N_23128,N_20585,N_19667);
and U23129 (N_23129,N_18817,N_18995);
and U23130 (N_23130,N_18133,N_20153);
and U23131 (N_23131,N_20098,N_19129);
nand U23132 (N_23132,N_18002,N_18956);
and U23133 (N_23133,N_18690,N_20732);
or U23134 (N_23134,N_20837,N_20098);
and U23135 (N_23135,N_18415,N_20166);
nand U23136 (N_23136,N_20061,N_19201);
and U23137 (N_23137,N_18933,N_19299);
and U23138 (N_23138,N_19187,N_19246);
and U23139 (N_23139,N_20695,N_20743);
xor U23140 (N_23140,N_18040,N_18664);
and U23141 (N_23141,N_18541,N_19579);
xnor U23142 (N_23142,N_19095,N_20534);
and U23143 (N_23143,N_20544,N_18719);
or U23144 (N_23144,N_19237,N_18774);
and U23145 (N_23145,N_20470,N_18821);
nor U23146 (N_23146,N_19134,N_18813);
xor U23147 (N_23147,N_18647,N_20133);
nand U23148 (N_23148,N_18005,N_19633);
nand U23149 (N_23149,N_18724,N_19663);
xnor U23150 (N_23150,N_20861,N_19889);
and U23151 (N_23151,N_19803,N_20693);
nand U23152 (N_23152,N_19965,N_18986);
nand U23153 (N_23153,N_19719,N_20244);
and U23154 (N_23154,N_18454,N_20037);
xor U23155 (N_23155,N_19134,N_20214);
xnor U23156 (N_23156,N_19860,N_19863);
nand U23157 (N_23157,N_20648,N_20611);
xnor U23158 (N_23158,N_19069,N_19372);
nand U23159 (N_23159,N_19714,N_20856);
or U23160 (N_23160,N_19303,N_18557);
or U23161 (N_23161,N_18908,N_18243);
nor U23162 (N_23162,N_20642,N_19798);
xor U23163 (N_23163,N_19594,N_19216);
or U23164 (N_23164,N_19373,N_19323);
nand U23165 (N_23165,N_19519,N_20772);
xnor U23166 (N_23166,N_19105,N_19569);
or U23167 (N_23167,N_18436,N_18085);
xor U23168 (N_23168,N_20656,N_20523);
nand U23169 (N_23169,N_20432,N_19068);
xnor U23170 (N_23170,N_18931,N_19948);
or U23171 (N_23171,N_20494,N_18188);
nor U23172 (N_23172,N_19935,N_19108);
and U23173 (N_23173,N_19617,N_19976);
nand U23174 (N_23174,N_18319,N_19585);
or U23175 (N_23175,N_18275,N_19804);
nand U23176 (N_23176,N_20226,N_20505);
nor U23177 (N_23177,N_18656,N_19629);
nor U23178 (N_23178,N_18721,N_19741);
xor U23179 (N_23179,N_19859,N_20649);
xor U23180 (N_23180,N_19961,N_20729);
or U23181 (N_23181,N_20846,N_19247);
nor U23182 (N_23182,N_18309,N_18539);
nand U23183 (N_23183,N_20198,N_20536);
nor U23184 (N_23184,N_19831,N_18189);
or U23185 (N_23185,N_20717,N_20831);
xnor U23186 (N_23186,N_20033,N_19798);
xnor U23187 (N_23187,N_19065,N_18548);
or U23188 (N_23188,N_18956,N_18162);
xnor U23189 (N_23189,N_19293,N_19796);
xor U23190 (N_23190,N_18014,N_18898);
or U23191 (N_23191,N_20060,N_20985);
and U23192 (N_23192,N_18695,N_18430);
or U23193 (N_23193,N_20626,N_19736);
xor U23194 (N_23194,N_20329,N_20984);
or U23195 (N_23195,N_20449,N_18037);
nor U23196 (N_23196,N_18368,N_18587);
nor U23197 (N_23197,N_20283,N_18243);
xnor U23198 (N_23198,N_19047,N_19204);
or U23199 (N_23199,N_19592,N_19480);
nand U23200 (N_23200,N_20121,N_19777);
nor U23201 (N_23201,N_19795,N_20509);
nor U23202 (N_23202,N_20068,N_20490);
or U23203 (N_23203,N_18594,N_19216);
or U23204 (N_23204,N_20964,N_20937);
and U23205 (N_23205,N_19179,N_19266);
and U23206 (N_23206,N_20488,N_20114);
or U23207 (N_23207,N_18819,N_18052);
or U23208 (N_23208,N_20607,N_18410);
xor U23209 (N_23209,N_18901,N_19273);
or U23210 (N_23210,N_19796,N_19103);
nor U23211 (N_23211,N_20070,N_18113);
nor U23212 (N_23212,N_18423,N_19180);
xnor U23213 (N_23213,N_18625,N_20349);
and U23214 (N_23214,N_18080,N_18560);
nor U23215 (N_23215,N_19274,N_20342);
and U23216 (N_23216,N_19041,N_20998);
nand U23217 (N_23217,N_20619,N_20275);
nor U23218 (N_23218,N_19709,N_19863);
or U23219 (N_23219,N_20370,N_18907);
nor U23220 (N_23220,N_18341,N_18711);
and U23221 (N_23221,N_20266,N_18300);
nand U23222 (N_23222,N_19715,N_19437);
and U23223 (N_23223,N_18450,N_20377);
xor U23224 (N_23224,N_20467,N_18426);
and U23225 (N_23225,N_19377,N_18025);
or U23226 (N_23226,N_18869,N_19963);
xor U23227 (N_23227,N_20206,N_20680);
nor U23228 (N_23228,N_20097,N_20958);
nor U23229 (N_23229,N_18778,N_19271);
and U23230 (N_23230,N_18115,N_18876);
nand U23231 (N_23231,N_18799,N_20799);
or U23232 (N_23232,N_18002,N_20851);
nand U23233 (N_23233,N_20839,N_19963);
nor U23234 (N_23234,N_20652,N_18024);
nand U23235 (N_23235,N_19349,N_20780);
nand U23236 (N_23236,N_18049,N_19418);
or U23237 (N_23237,N_18046,N_18232);
nand U23238 (N_23238,N_20514,N_18525);
xor U23239 (N_23239,N_19408,N_20942);
xnor U23240 (N_23240,N_19521,N_19130);
xor U23241 (N_23241,N_19155,N_20151);
and U23242 (N_23242,N_18828,N_18032);
xor U23243 (N_23243,N_18590,N_20965);
nand U23244 (N_23244,N_20607,N_18608);
nand U23245 (N_23245,N_19410,N_20750);
nor U23246 (N_23246,N_18001,N_20460);
and U23247 (N_23247,N_19670,N_20104);
nand U23248 (N_23248,N_19911,N_18731);
nor U23249 (N_23249,N_18895,N_18147);
nor U23250 (N_23250,N_20219,N_20882);
nor U23251 (N_23251,N_19033,N_20553);
nand U23252 (N_23252,N_20692,N_19785);
nor U23253 (N_23253,N_20743,N_18374);
nand U23254 (N_23254,N_19902,N_19726);
nor U23255 (N_23255,N_18115,N_20318);
nor U23256 (N_23256,N_20469,N_18512);
and U23257 (N_23257,N_18883,N_20677);
nor U23258 (N_23258,N_20763,N_18140);
or U23259 (N_23259,N_19251,N_19768);
and U23260 (N_23260,N_19316,N_20131);
nor U23261 (N_23261,N_20046,N_20861);
xor U23262 (N_23262,N_18374,N_18522);
xnor U23263 (N_23263,N_18428,N_18972);
nand U23264 (N_23264,N_20232,N_20936);
and U23265 (N_23265,N_19797,N_18630);
nor U23266 (N_23266,N_20219,N_20855);
nand U23267 (N_23267,N_20726,N_20028);
nand U23268 (N_23268,N_19204,N_20658);
nor U23269 (N_23269,N_18883,N_18060);
nand U23270 (N_23270,N_19861,N_19716);
nor U23271 (N_23271,N_20569,N_19392);
xnor U23272 (N_23272,N_18456,N_19075);
xnor U23273 (N_23273,N_19514,N_18232);
and U23274 (N_23274,N_19430,N_19969);
xor U23275 (N_23275,N_20829,N_19690);
xnor U23276 (N_23276,N_18778,N_20921);
or U23277 (N_23277,N_18456,N_18232);
nand U23278 (N_23278,N_20045,N_20026);
nor U23279 (N_23279,N_20283,N_19741);
nor U23280 (N_23280,N_20706,N_20651);
xor U23281 (N_23281,N_19178,N_18768);
and U23282 (N_23282,N_19948,N_18297);
and U23283 (N_23283,N_20811,N_18590);
and U23284 (N_23284,N_18347,N_18657);
nand U23285 (N_23285,N_19080,N_20798);
nor U23286 (N_23286,N_20753,N_20636);
xnor U23287 (N_23287,N_20032,N_20614);
xor U23288 (N_23288,N_20041,N_19078);
and U23289 (N_23289,N_20810,N_20739);
and U23290 (N_23290,N_18436,N_20233);
xnor U23291 (N_23291,N_18979,N_18845);
or U23292 (N_23292,N_19802,N_19933);
nor U23293 (N_23293,N_19886,N_19153);
xnor U23294 (N_23294,N_18624,N_19709);
nand U23295 (N_23295,N_20691,N_19617);
nor U23296 (N_23296,N_20275,N_18761);
or U23297 (N_23297,N_18464,N_19002);
or U23298 (N_23298,N_20088,N_20206);
nand U23299 (N_23299,N_20376,N_20542);
or U23300 (N_23300,N_18295,N_18695);
nor U23301 (N_23301,N_18415,N_20045);
and U23302 (N_23302,N_18772,N_20884);
nor U23303 (N_23303,N_19284,N_19673);
or U23304 (N_23304,N_18164,N_20831);
xor U23305 (N_23305,N_18256,N_20944);
or U23306 (N_23306,N_19855,N_19807);
xnor U23307 (N_23307,N_20502,N_18308);
nor U23308 (N_23308,N_18501,N_19905);
xnor U23309 (N_23309,N_19980,N_19222);
xor U23310 (N_23310,N_19783,N_19718);
and U23311 (N_23311,N_19887,N_18314);
or U23312 (N_23312,N_19976,N_20105);
nand U23313 (N_23313,N_19309,N_19022);
and U23314 (N_23314,N_18213,N_18667);
nor U23315 (N_23315,N_20888,N_18806);
or U23316 (N_23316,N_18832,N_18242);
xor U23317 (N_23317,N_18466,N_18670);
and U23318 (N_23318,N_18279,N_19001);
nand U23319 (N_23319,N_20504,N_19156);
nor U23320 (N_23320,N_20293,N_20727);
nand U23321 (N_23321,N_20224,N_18024);
nand U23322 (N_23322,N_19617,N_19584);
or U23323 (N_23323,N_19698,N_20583);
nor U23324 (N_23324,N_18865,N_18429);
xnor U23325 (N_23325,N_20092,N_18297);
xnor U23326 (N_23326,N_20009,N_20522);
nand U23327 (N_23327,N_20968,N_19220);
xor U23328 (N_23328,N_19035,N_18801);
nor U23329 (N_23329,N_18666,N_18858);
or U23330 (N_23330,N_19050,N_20578);
and U23331 (N_23331,N_20471,N_20734);
nand U23332 (N_23332,N_20703,N_18067);
and U23333 (N_23333,N_20848,N_18766);
nor U23334 (N_23334,N_18102,N_20502);
nor U23335 (N_23335,N_19547,N_19505);
nand U23336 (N_23336,N_19069,N_19016);
and U23337 (N_23337,N_20983,N_19082);
or U23338 (N_23338,N_18423,N_19856);
nand U23339 (N_23339,N_20038,N_18815);
and U23340 (N_23340,N_19719,N_20482);
nand U23341 (N_23341,N_19162,N_18276);
and U23342 (N_23342,N_19769,N_18282);
nor U23343 (N_23343,N_18384,N_18913);
nand U23344 (N_23344,N_18455,N_19266);
nor U23345 (N_23345,N_20459,N_20671);
nand U23346 (N_23346,N_20232,N_20275);
and U23347 (N_23347,N_18890,N_19430);
or U23348 (N_23348,N_20948,N_20213);
and U23349 (N_23349,N_19081,N_19189);
xor U23350 (N_23350,N_20699,N_18821);
xor U23351 (N_23351,N_18275,N_19861);
nor U23352 (N_23352,N_18177,N_20947);
or U23353 (N_23353,N_18935,N_18017);
and U23354 (N_23354,N_20391,N_18696);
nand U23355 (N_23355,N_19668,N_19758);
xnor U23356 (N_23356,N_20414,N_18814);
and U23357 (N_23357,N_20240,N_19432);
nand U23358 (N_23358,N_19776,N_20383);
or U23359 (N_23359,N_18404,N_20477);
nand U23360 (N_23360,N_18388,N_19660);
xor U23361 (N_23361,N_19437,N_20364);
or U23362 (N_23362,N_20083,N_19363);
and U23363 (N_23363,N_20430,N_19544);
or U23364 (N_23364,N_18643,N_19055);
xnor U23365 (N_23365,N_18908,N_18857);
nor U23366 (N_23366,N_19558,N_20984);
nand U23367 (N_23367,N_18111,N_18145);
nor U23368 (N_23368,N_18022,N_20524);
and U23369 (N_23369,N_20505,N_19212);
and U23370 (N_23370,N_18071,N_20501);
xor U23371 (N_23371,N_18117,N_20186);
or U23372 (N_23372,N_18042,N_19945);
nor U23373 (N_23373,N_20283,N_19592);
xnor U23374 (N_23374,N_19425,N_20111);
nor U23375 (N_23375,N_18560,N_19482);
and U23376 (N_23376,N_19780,N_19485);
and U23377 (N_23377,N_19603,N_18529);
or U23378 (N_23378,N_20963,N_19797);
and U23379 (N_23379,N_19835,N_20293);
and U23380 (N_23380,N_19022,N_19479);
nand U23381 (N_23381,N_20110,N_20582);
nor U23382 (N_23382,N_18662,N_19888);
xor U23383 (N_23383,N_18785,N_19059);
nor U23384 (N_23384,N_19822,N_19190);
xnor U23385 (N_23385,N_19965,N_18446);
nand U23386 (N_23386,N_18430,N_20018);
nor U23387 (N_23387,N_19508,N_20806);
xnor U23388 (N_23388,N_18076,N_18406);
xnor U23389 (N_23389,N_20679,N_20114);
xnor U23390 (N_23390,N_18250,N_20876);
and U23391 (N_23391,N_19593,N_19620);
and U23392 (N_23392,N_18640,N_18962);
or U23393 (N_23393,N_20171,N_20617);
nand U23394 (N_23394,N_18476,N_19079);
nor U23395 (N_23395,N_19531,N_18976);
or U23396 (N_23396,N_18032,N_20297);
or U23397 (N_23397,N_20963,N_18288);
and U23398 (N_23398,N_20829,N_20746);
and U23399 (N_23399,N_18387,N_20664);
or U23400 (N_23400,N_19934,N_18438);
nand U23401 (N_23401,N_18392,N_19698);
and U23402 (N_23402,N_19997,N_18535);
or U23403 (N_23403,N_18381,N_20370);
nor U23404 (N_23404,N_18673,N_19926);
nand U23405 (N_23405,N_18047,N_20257);
nand U23406 (N_23406,N_20650,N_20992);
or U23407 (N_23407,N_19750,N_18481);
and U23408 (N_23408,N_18798,N_19352);
and U23409 (N_23409,N_19891,N_20973);
and U23410 (N_23410,N_20553,N_18849);
and U23411 (N_23411,N_20657,N_19796);
nand U23412 (N_23412,N_20800,N_19791);
nand U23413 (N_23413,N_18468,N_18353);
and U23414 (N_23414,N_19379,N_19303);
and U23415 (N_23415,N_18258,N_18045);
or U23416 (N_23416,N_18952,N_19519);
xor U23417 (N_23417,N_20663,N_20561);
nor U23418 (N_23418,N_20105,N_18210);
or U23419 (N_23419,N_20618,N_18957);
and U23420 (N_23420,N_18802,N_20371);
nor U23421 (N_23421,N_20526,N_19801);
nand U23422 (N_23422,N_20790,N_19796);
or U23423 (N_23423,N_18233,N_20721);
nand U23424 (N_23424,N_18640,N_20359);
nor U23425 (N_23425,N_19537,N_20787);
xnor U23426 (N_23426,N_20741,N_19640);
nor U23427 (N_23427,N_19843,N_18119);
and U23428 (N_23428,N_20745,N_20568);
or U23429 (N_23429,N_19465,N_20499);
or U23430 (N_23430,N_19095,N_20101);
or U23431 (N_23431,N_20771,N_19638);
nor U23432 (N_23432,N_19723,N_20381);
nor U23433 (N_23433,N_18635,N_19315);
nand U23434 (N_23434,N_20269,N_20402);
or U23435 (N_23435,N_20413,N_20860);
and U23436 (N_23436,N_18166,N_18130);
or U23437 (N_23437,N_20410,N_20956);
xor U23438 (N_23438,N_18369,N_20495);
and U23439 (N_23439,N_18542,N_18425);
or U23440 (N_23440,N_19642,N_18384);
or U23441 (N_23441,N_18599,N_19543);
nor U23442 (N_23442,N_19870,N_19102);
or U23443 (N_23443,N_19983,N_19427);
or U23444 (N_23444,N_18648,N_20629);
nor U23445 (N_23445,N_18945,N_18159);
and U23446 (N_23446,N_18584,N_20546);
nor U23447 (N_23447,N_19953,N_20465);
or U23448 (N_23448,N_18042,N_19824);
nor U23449 (N_23449,N_19835,N_20106);
and U23450 (N_23450,N_19978,N_20354);
nor U23451 (N_23451,N_18534,N_18490);
nand U23452 (N_23452,N_20384,N_18109);
or U23453 (N_23453,N_19858,N_19383);
nor U23454 (N_23454,N_20399,N_20001);
nor U23455 (N_23455,N_18696,N_20313);
nand U23456 (N_23456,N_19141,N_19061);
nand U23457 (N_23457,N_20846,N_18874);
or U23458 (N_23458,N_20106,N_19986);
nor U23459 (N_23459,N_19986,N_18137);
nor U23460 (N_23460,N_18029,N_18357);
and U23461 (N_23461,N_20022,N_20293);
nand U23462 (N_23462,N_19694,N_19430);
and U23463 (N_23463,N_19652,N_19786);
nand U23464 (N_23464,N_20438,N_20425);
or U23465 (N_23465,N_20734,N_20170);
nand U23466 (N_23466,N_18858,N_19553);
nand U23467 (N_23467,N_19576,N_18975);
nand U23468 (N_23468,N_20337,N_19127);
nor U23469 (N_23469,N_18991,N_19038);
xnor U23470 (N_23470,N_18446,N_20674);
nand U23471 (N_23471,N_19809,N_20910);
and U23472 (N_23472,N_20621,N_19375);
xnor U23473 (N_23473,N_18052,N_20873);
xor U23474 (N_23474,N_20439,N_19153);
nor U23475 (N_23475,N_20980,N_20540);
xor U23476 (N_23476,N_20926,N_20867);
and U23477 (N_23477,N_18229,N_18840);
nor U23478 (N_23478,N_19023,N_20638);
xnor U23479 (N_23479,N_18308,N_18649);
nand U23480 (N_23480,N_20497,N_20420);
xnor U23481 (N_23481,N_19975,N_20899);
nor U23482 (N_23482,N_20013,N_19073);
xnor U23483 (N_23483,N_20971,N_20947);
xnor U23484 (N_23484,N_19906,N_19216);
nand U23485 (N_23485,N_19290,N_19493);
and U23486 (N_23486,N_20034,N_18090);
xor U23487 (N_23487,N_19557,N_18413);
nand U23488 (N_23488,N_20071,N_18617);
and U23489 (N_23489,N_20931,N_18072);
or U23490 (N_23490,N_20884,N_20028);
or U23491 (N_23491,N_19705,N_18136);
nand U23492 (N_23492,N_20221,N_18412);
or U23493 (N_23493,N_20620,N_18000);
xor U23494 (N_23494,N_18279,N_20046);
nand U23495 (N_23495,N_20412,N_20184);
nand U23496 (N_23496,N_18557,N_20548);
xnor U23497 (N_23497,N_20043,N_20505);
nor U23498 (N_23498,N_20434,N_19755);
or U23499 (N_23499,N_19931,N_19534);
nand U23500 (N_23500,N_19162,N_18031);
xnor U23501 (N_23501,N_18594,N_20512);
nand U23502 (N_23502,N_18574,N_20174);
and U23503 (N_23503,N_20757,N_20417);
nor U23504 (N_23504,N_18196,N_19621);
xor U23505 (N_23505,N_19791,N_19356);
xnor U23506 (N_23506,N_18798,N_18891);
xor U23507 (N_23507,N_20447,N_19443);
and U23508 (N_23508,N_19115,N_20018);
or U23509 (N_23509,N_18126,N_19803);
xnor U23510 (N_23510,N_20584,N_19935);
or U23511 (N_23511,N_20722,N_19957);
or U23512 (N_23512,N_20339,N_20574);
nor U23513 (N_23513,N_19937,N_20985);
nor U23514 (N_23514,N_19576,N_18996);
nand U23515 (N_23515,N_19717,N_19214);
and U23516 (N_23516,N_18696,N_20277);
nand U23517 (N_23517,N_18022,N_20189);
nand U23518 (N_23518,N_19459,N_19079);
nand U23519 (N_23519,N_20346,N_19800);
nor U23520 (N_23520,N_19462,N_19505);
or U23521 (N_23521,N_20370,N_20103);
nand U23522 (N_23522,N_20560,N_18459);
and U23523 (N_23523,N_20573,N_19544);
and U23524 (N_23524,N_18880,N_19187);
xnor U23525 (N_23525,N_18313,N_19538);
and U23526 (N_23526,N_19142,N_18337);
nand U23527 (N_23527,N_20135,N_20346);
xnor U23528 (N_23528,N_18554,N_20357);
nand U23529 (N_23529,N_18127,N_20116);
nor U23530 (N_23530,N_18603,N_19726);
xnor U23531 (N_23531,N_19390,N_19753);
nor U23532 (N_23532,N_19242,N_19349);
or U23533 (N_23533,N_18143,N_18770);
xnor U23534 (N_23534,N_19762,N_20228);
xor U23535 (N_23535,N_18032,N_18312);
nor U23536 (N_23536,N_19754,N_19622);
xor U23537 (N_23537,N_19512,N_20059);
and U23538 (N_23538,N_18972,N_19992);
nand U23539 (N_23539,N_19103,N_20572);
xnor U23540 (N_23540,N_19328,N_18974);
and U23541 (N_23541,N_20936,N_20558);
nand U23542 (N_23542,N_20701,N_18619);
xnor U23543 (N_23543,N_20798,N_19460);
nor U23544 (N_23544,N_20853,N_20318);
nand U23545 (N_23545,N_19275,N_20896);
or U23546 (N_23546,N_20771,N_18001);
nor U23547 (N_23547,N_18697,N_18120);
or U23548 (N_23548,N_20785,N_20612);
and U23549 (N_23549,N_20662,N_19336);
nor U23550 (N_23550,N_19471,N_18632);
nand U23551 (N_23551,N_18217,N_19476);
or U23552 (N_23552,N_19487,N_18481);
or U23553 (N_23553,N_20086,N_20272);
and U23554 (N_23554,N_18072,N_18037);
xor U23555 (N_23555,N_19802,N_18593);
nor U23556 (N_23556,N_18784,N_20790);
xnor U23557 (N_23557,N_19564,N_19176);
and U23558 (N_23558,N_18376,N_18686);
and U23559 (N_23559,N_20918,N_19585);
and U23560 (N_23560,N_19732,N_20925);
xnor U23561 (N_23561,N_18123,N_20272);
or U23562 (N_23562,N_18703,N_19683);
nand U23563 (N_23563,N_18591,N_20711);
or U23564 (N_23564,N_18693,N_18356);
nand U23565 (N_23565,N_20538,N_18248);
nand U23566 (N_23566,N_20930,N_20319);
nand U23567 (N_23567,N_20659,N_19855);
nand U23568 (N_23568,N_19049,N_18889);
nand U23569 (N_23569,N_20860,N_19864);
nand U23570 (N_23570,N_19177,N_19596);
nor U23571 (N_23571,N_19085,N_20542);
xnor U23572 (N_23572,N_20534,N_18805);
nor U23573 (N_23573,N_19036,N_18127);
or U23574 (N_23574,N_19537,N_19673);
nor U23575 (N_23575,N_19121,N_18552);
nor U23576 (N_23576,N_18984,N_20828);
xor U23577 (N_23577,N_20228,N_20237);
xnor U23578 (N_23578,N_18710,N_18811);
xor U23579 (N_23579,N_18683,N_18203);
nand U23580 (N_23580,N_18377,N_19954);
nand U23581 (N_23581,N_20983,N_18635);
nand U23582 (N_23582,N_20972,N_19325);
nand U23583 (N_23583,N_19346,N_20911);
and U23584 (N_23584,N_18862,N_19224);
xnor U23585 (N_23585,N_18692,N_18720);
xnor U23586 (N_23586,N_18147,N_19715);
and U23587 (N_23587,N_20017,N_20758);
and U23588 (N_23588,N_18907,N_20997);
or U23589 (N_23589,N_18678,N_18008);
and U23590 (N_23590,N_20560,N_19338);
nand U23591 (N_23591,N_20098,N_19549);
and U23592 (N_23592,N_20321,N_20624);
xnor U23593 (N_23593,N_20275,N_19471);
nor U23594 (N_23594,N_18106,N_20167);
nand U23595 (N_23595,N_18571,N_19445);
and U23596 (N_23596,N_18641,N_20347);
xnor U23597 (N_23597,N_20079,N_19615);
nor U23598 (N_23598,N_20355,N_18283);
or U23599 (N_23599,N_18192,N_20993);
and U23600 (N_23600,N_18746,N_18511);
or U23601 (N_23601,N_20622,N_18904);
xor U23602 (N_23602,N_19397,N_20595);
xor U23603 (N_23603,N_18411,N_20779);
nor U23604 (N_23604,N_19077,N_19981);
or U23605 (N_23605,N_18648,N_20885);
nand U23606 (N_23606,N_19840,N_19469);
nor U23607 (N_23607,N_18571,N_20834);
and U23608 (N_23608,N_20228,N_19862);
or U23609 (N_23609,N_19072,N_19643);
nor U23610 (N_23610,N_19345,N_19262);
and U23611 (N_23611,N_18303,N_19504);
or U23612 (N_23612,N_20708,N_18821);
and U23613 (N_23613,N_20798,N_20786);
and U23614 (N_23614,N_18242,N_20551);
or U23615 (N_23615,N_20958,N_19316);
xor U23616 (N_23616,N_19115,N_19406);
and U23617 (N_23617,N_20152,N_20933);
or U23618 (N_23618,N_20121,N_19528);
and U23619 (N_23619,N_19096,N_20715);
xnor U23620 (N_23620,N_18429,N_20503);
and U23621 (N_23621,N_19771,N_18081);
and U23622 (N_23622,N_20461,N_18655);
nor U23623 (N_23623,N_19387,N_20160);
and U23624 (N_23624,N_19633,N_20723);
nand U23625 (N_23625,N_20663,N_18713);
nand U23626 (N_23626,N_20607,N_18070);
nor U23627 (N_23627,N_20297,N_18586);
nand U23628 (N_23628,N_19783,N_20807);
and U23629 (N_23629,N_18221,N_20067);
nor U23630 (N_23630,N_18523,N_20422);
and U23631 (N_23631,N_18159,N_18683);
or U23632 (N_23632,N_20830,N_20912);
xor U23633 (N_23633,N_20692,N_18603);
and U23634 (N_23634,N_19900,N_19561);
nand U23635 (N_23635,N_18052,N_18858);
nor U23636 (N_23636,N_19869,N_19534);
and U23637 (N_23637,N_18211,N_20462);
and U23638 (N_23638,N_20470,N_19230);
or U23639 (N_23639,N_19847,N_19947);
and U23640 (N_23640,N_20960,N_19275);
nand U23641 (N_23641,N_20959,N_20306);
nand U23642 (N_23642,N_18260,N_20643);
or U23643 (N_23643,N_18217,N_19869);
nand U23644 (N_23644,N_18907,N_18574);
xnor U23645 (N_23645,N_18750,N_19636);
or U23646 (N_23646,N_20804,N_18449);
nand U23647 (N_23647,N_20959,N_18164);
or U23648 (N_23648,N_19903,N_18306);
and U23649 (N_23649,N_19361,N_20301);
nand U23650 (N_23650,N_19971,N_18669);
and U23651 (N_23651,N_19296,N_18056);
xor U23652 (N_23652,N_19146,N_18593);
and U23653 (N_23653,N_20422,N_19332);
and U23654 (N_23654,N_20817,N_18871);
nand U23655 (N_23655,N_20390,N_18391);
and U23656 (N_23656,N_19232,N_20572);
or U23657 (N_23657,N_18576,N_20371);
nand U23658 (N_23658,N_19460,N_20729);
or U23659 (N_23659,N_20686,N_20627);
nand U23660 (N_23660,N_19770,N_19118);
or U23661 (N_23661,N_18482,N_18918);
and U23662 (N_23662,N_18385,N_20136);
nand U23663 (N_23663,N_20951,N_19101);
or U23664 (N_23664,N_20925,N_20028);
nor U23665 (N_23665,N_20697,N_20193);
and U23666 (N_23666,N_19696,N_18661);
nor U23667 (N_23667,N_18800,N_20005);
nor U23668 (N_23668,N_19645,N_18960);
nor U23669 (N_23669,N_18785,N_20317);
and U23670 (N_23670,N_20360,N_19708);
and U23671 (N_23671,N_19838,N_18572);
and U23672 (N_23672,N_20741,N_19938);
or U23673 (N_23673,N_19307,N_19844);
xor U23674 (N_23674,N_18964,N_18448);
nand U23675 (N_23675,N_20425,N_20057);
nor U23676 (N_23676,N_20459,N_20360);
nor U23677 (N_23677,N_19977,N_19724);
or U23678 (N_23678,N_20068,N_19381);
or U23679 (N_23679,N_19292,N_20022);
and U23680 (N_23680,N_18299,N_19120);
or U23681 (N_23681,N_20734,N_19381);
and U23682 (N_23682,N_19321,N_20784);
nor U23683 (N_23683,N_18429,N_19687);
and U23684 (N_23684,N_19846,N_18208);
nand U23685 (N_23685,N_19115,N_20945);
or U23686 (N_23686,N_20069,N_18238);
nand U23687 (N_23687,N_18399,N_18181);
nand U23688 (N_23688,N_18815,N_18995);
nand U23689 (N_23689,N_20855,N_19171);
xor U23690 (N_23690,N_20428,N_18753);
or U23691 (N_23691,N_19894,N_19288);
and U23692 (N_23692,N_20902,N_19183);
and U23693 (N_23693,N_20007,N_18031);
nor U23694 (N_23694,N_19990,N_19283);
or U23695 (N_23695,N_19897,N_20117);
xor U23696 (N_23696,N_19922,N_19917);
nand U23697 (N_23697,N_18674,N_20146);
xnor U23698 (N_23698,N_20212,N_19977);
nor U23699 (N_23699,N_20845,N_19444);
xnor U23700 (N_23700,N_20840,N_19728);
and U23701 (N_23701,N_20436,N_19545);
and U23702 (N_23702,N_19457,N_19309);
nand U23703 (N_23703,N_20530,N_18395);
xnor U23704 (N_23704,N_20700,N_18536);
or U23705 (N_23705,N_19808,N_18406);
or U23706 (N_23706,N_18698,N_20155);
nor U23707 (N_23707,N_18071,N_18835);
xor U23708 (N_23708,N_19404,N_18559);
or U23709 (N_23709,N_18301,N_20387);
or U23710 (N_23710,N_20340,N_18229);
or U23711 (N_23711,N_19013,N_19308);
xnor U23712 (N_23712,N_19240,N_19355);
nand U23713 (N_23713,N_20092,N_20926);
or U23714 (N_23714,N_20053,N_20878);
xor U23715 (N_23715,N_20907,N_18788);
and U23716 (N_23716,N_20885,N_19179);
xor U23717 (N_23717,N_20131,N_19989);
nor U23718 (N_23718,N_18128,N_20534);
and U23719 (N_23719,N_19304,N_19746);
nor U23720 (N_23720,N_19337,N_19303);
nand U23721 (N_23721,N_20239,N_18084);
or U23722 (N_23722,N_20323,N_19110);
nand U23723 (N_23723,N_18502,N_19864);
nand U23724 (N_23724,N_19599,N_18750);
xor U23725 (N_23725,N_18551,N_20934);
xor U23726 (N_23726,N_20031,N_18219);
and U23727 (N_23727,N_18282,N_18626);
and U23728 (N_23728,N_20729,N_20936);
nand U23729 (N_23729,N_20226,N_19151);
and U23730 (N_23730,N_18523,N_20377);
and U23731 (N_23731,N_18518,N_20397);
nand U23732 (N_23732,N_19723,N_19236);
or U23733 (N_23733,N_20899,N_20375);
nor U23734 (N_23734,N_18408,N_20037);
xor U23735 (N_23735,N_20735,N_18100);
or U23736 (N_23736,N_20705,N_18595);
and U23737 (N_23737,N_20392,N_19033);
or U23738 (N_23738,N_19799,N_18300);
and U23739 (N_23739,N_19506,N_20625);
xnor U23740 (N_23740,N_18526,N_18170);
and U23741 (N_23741,N_20044,N_20629);
xnor U23742 (N_23742,N_19689,N_18487);
nor U23743 (N_23743,N_19172,N_18437);
and U23744 (N_23744,N_18441,N_20348);
or U23745 (N_23745,N_20430,N_20208);
and U23746 (N_23746,N_19490,N_18814);
xor U23747 (N_23747,N_20609,N_20866);
and U23748 (N_23748,N_18692,N_20690);
and U23749 (N_23749,N_20055,N_18060);
nand U23750 (N_23750,N_20649,N_19306);
and U23751 (N_23751,N_18300,N_20602);
nand U23752 (N_23752,N_20018,N_20996);
nand U23753 (N_23753,N_18009,N_19994);
nor U23754 (N_23754,N_20067,N_18442);
or U23755 (N_23755,N_18778,N_19045);
nor U23756 (N_23756,N_19334,N_20417);
or U23757 (N_23757,N_18150,N_20759);
nand U23758 (N_23758,N_20460,N_20657);
and U23759 (N_23759,N_18081,N_20073);
or U23760 (N_23760,N_20223,N_18189);
xnor U23761 (N_23761,N_20923,N_18447);
nand U23762 (N_23762,N_20331,N_20301);
nand U23763 (N_23763,N_20065,N_18934);
and U23764 (N_23764,N_20139,N_19992);
nor U23765 (N_23765,N_18514,N_18598);
xnor U23766 (N_23766,N_19685,N_19290);
and U23767 (N_23767,N_18021,N_18471);
and U23768 (N_23768,N_19214,N_19855);
and U23769 (N_23769,N_18768,N_19238);
nor U23770 (N_23770,N_18531,N_18163);
xnor U23771 (N_23771,N_20290,N_18804);
xor U23772 (N_23772,N_20177,N_19396);
xnor U23773 (N_23773,N_18893,N_18601);
or U23774 (N_23774,N_19038,N_18920);
nand U23775 (N_23775,N_18627,N_18358);
nor U23776 (N_23776,N_19867,N_18550);
or U23777 (N_23777,N_20577,N_18815);
nand U23778 (N_23778,N_18812,N_19548);
and U23779 (N_23779,N_20076,N_18977);
nor U23780 (N_23780,N_19444,N_20491);
nor U23781 (N_23781,N_20114,N_19407);
nor U23782 (N_23782,N_18540,N_18059);
and U23783 (N_23783,N_18966,N_18429);
or U23784 (N_23784,N_18233,N_19463);
nor U23785 (N_23785,N_20965,N_20821);
or U23786 (N_23786,N_18521,N_18316);
and U23787 (N_23787,N_18517,N_19980);
xnor U23788 (N_23788,N_18495,N_20900);
xnor U23789 (N_23789,N_18727,N_18788);
xor U23790 (N_23790,N_20380,N_20215);
nand U23791 (N_23791,N_20533,N_20683);
and U23792 (N_23792,N_20057,N_18337);
or U23793 (N_23793,N_20985,N_18534);
and U23794 (N_23794,N_18383,N_20166);
or U23795 (N_23795,N_20704,N_18221);
or U23796 (N_23796,N_18240,N_18620);
nand U23797 (N_23797,N_19059,N_19524);
or U23798 (N_23798,N_19783,N_18923);
nand U23799 (N_23799,N_19185,N_19419);
nor U23800 (N_23800,N_20512,N_20016);
nand U23801 (N_23801,N_18967,N_18857);
or U23802 (N_23802,N_18017,N_18740);
nand U23803 (N_23803,N_20276,N_20087);
nand U23804 (N_23804,N_19405,N_18814);
xor U23805 (N_23805,N_20221,N_19287);
xor U23806 (N_23806,N_19434,N_18855);
nand U23807 (N_23807,N_20191,N_20845);
or U23808 (N_23808,N_18629,N_19941);
nand U23809 (N_23809,N_19766,N_18388);
nand U23810 (N_23810,N_19512,N_19704);
or U23811 (N_23811,N_19780,N_19326);
xor U23812 (N_23812,N_18803,N_18868);
xnor U23813 (N_23813,N_20457,N_18521);
and U23814 (N_23814,N_19030,N_18886);
xnor U23815 (N_23815,N_18048,N_20377);
nand U23816 (N_23816,N_20765,N_20620);
nand U23817 (N_23817,N_18461,N_18787);
nand U23818 (N_23818,N_19489,N_19705);
and U23819 (N_23819,N_19704,N_20498);
nor U23820 (N_23820,N_18594,N_19413);
and U23821 (N_23821,N_20619,N_18440);
xnor U23822 (N_23822,N_20584,N_19131);
and U23823 (N_23823,N_19081,N_20684);
and U23824 (N_23824,N_18216,N_20501);
nor U23825 (N_23825,N_20778,N_20692);
nand U23826 (N_23826,N_18091,N_19289);
nor U23827 (N_23827,N_20810,N_18283);
or U23828 (N_23828,N_20557,N_20601);
and U23829 (N_23829,N_18307,N_20295);
and U23830 (N_23830,N_18940,N_18664);
nand U23831 (N_23831,N_20692,N_19300);
and U23832 (N_23832,N_19420,N_20760);
and U23833 (N_23833,N_19789,N_19524);
nor U23834 (N_23834,N_20096,N_18555);
nor U23835 (N_23835,N_19671,N_18643);
or U23836 (N_23836,N_20767,N_18992);
nor U23837 (N_23837,N_19431,N_18675);
nor U23838 (N_23838,N_20687,N_20510);
nor U23839 (N_23839,N_20666,N_20540);
xor U23840 (N_23840,N_20829,N_20838);
and U23841 (N_23841,N_19810,N_20576);
nand U23842 (N_23842,N_18547,N_20854);
nor U23843 (N_23843,N_19151,N_19949);
xnor U23844 (N_23844,N_18990,N_18963);
and U23845 (N_23845,N_19943,N_18038);
nor U23846 (N_23846,N_18516,N_18711);
nor U23847 (N_23847,N_20221,N_19990);
xnor U23848 (N_23848,N_19598,N_19229);
nand U23849 (N_23849,N_19984,N_18862);
xnor U23850 (N_23850,N_19804,N_19627);
xnor U23851 (N_23851,N_18403,N_20660);
or U23852 (N_23852,N_18030,N_20685);
xor U23853 (N_23853,N_20709,N_20235);
nor U23854 (N_23854,N_18098,N_18668);
and U23855 (N_23855,N_20388,N_19347);
nor U23856 (N_23856,N_19871,N_19912);
nand U23857 (N_23857,N_20949,N_19410);
nor U23858 (N_23858,N_18761,N_18292);
nor U23859 (N_23859,N_19758,N_19136);
and U23860 (N_23860,N_20005,N_19147);
xor U23861 (N_23861,N_19798,N_19321);
nand U23862 (N_23862,N_18044,N_18910);
or U23863 (N_23863,N_20732,N_19183);
and U23864 (N_23864,N_19043,N_19633);
nor U23865 (N_23865,N_20976,N_19997);
nor U23866 (N_23866,N_19194,N_18770);
nand U23867 (N_23867,N_20637,N_18809);
or U23868 (N_23868,N_20808,N_19095);
xnor U23869 (N_23869,N_19391,N_18520);
xnor U23870 (N_23870,N_20372,N_19954);
nand U23871 (N_23871,N_19541,N_18736);
nand U23872 (N_23872,N_18214,N_19480);
nor U23873 (N_23873,N_20860,N_20625);
nand U23874 (N_23874,N_20223,N_20493);
or U23875 (N_23875,N_20875,N_18411);
or U23876 (N_23876,N_19573,N_19241);
and U23877 (N_23877,N_18334,N_18172);
nor U23878 (N_23878,N_19299,N_20719);
nor U23879 (N_23879,N_18887,N_19823);
nand U23880 (N_23880,N_19161,N_18282);
nand U23881 (N_23881,N_19969,N_20403);
or U23882 (N_23882,N_20214,N_20895);
nor U23883 (N_23883,N_19145,N_19299);
and U23884 (N_23884,N_18099,N_19273);
and U23885 (N_23885,N_19726,N_18283);
and U23886 (N_23886,N_20122,N_18495);
nor U23887 (N_23887,N_19247,N_19972);
xnor U23888 (N_23888,N_20915,N_19202);
nand U23889 (N_23889,N_18320,N_20491);
nor U23890 (N_23890,N_20893,N_20708);
or U23891 (N_23891,N_19003,N_18074);
nor U23892 (N_23892,N_18408,N_18035);
nand U23893 (N_23893,N_18487,N_18010);
and U23894 (N_23894,N_20200,N_19302);
xnor U23895 (N_23895,N_20471,N_20253);
or U23896 (N_23896,N_19419,N_19913);
nand U23897 (N_23897,N_18634,N_19346);
or U23898 (N_23898,N_20474,N_19385);
or U23899 (N_23899,N_18425,N_19811);
xor U23900 (N_23900,N_20193,N_20923);
and U23901 (N_23901,N_19642,N_19557);
xnor U23902 (N_23902,N_20010,N_20837);
xnor U23903 (N_23903,N_19803,N_20060);
nand U23904 (N_23904,N_19999,N_18992);
nor U23905 (N_23905,N_18584,N_19576);
xnor U23906 (N_23906,N_20421,N_18888);
or U23907 (N_23907,N_18199,N_20377);
or U23908 (N_23908,N_20535,N_19606);
nor U23909 (N_23909,N_20641,N_18059);
or U23910 (N_23910,N_18923,N_19530);
or U23911 (N_23911,N_19933,N_19659);
nor U23912 (N_23912,N_19450,N_18132);
nand U23913 (N_23913,N_19512,N_18140);
nand U23914 (N_23914,N_19797,N_18971);
xor U23915 (N_23915,N_19519,N_19186);
xnor U23916 (N_23916,N_19569,N_18777);
and U23917 (N_23917,N_18603,N_18060);
nand U23918 (N_23918,N_20761,N_18920);
nand U23919 (N_23919,N_19519,N_18533);
and U23920 (N_23920,N_18136,N_20967);
nand U23921 (N_23921,N_20822,N_20226);
and U23922 (N_23922,N_18983,N_19042);
or U23923 (N_23923,N_18242,N_20236);
and U23924 (N_23924,N_18599,N_19053);
or U23925 (N_23925,N_18648,N_18045);
nand U23926 (N_23926,N_20282,N_19562);
nor U23927 (N_23927,N_19171,N_19656);
and U23928 (N_23928,N_20027,N_18103);
nand U23929 (N_23929,N_20829,N_18672);
nor U23930 (N_23930,N_19932,N_19873);
nand U23931 (N_23931,N_20140,N_19261);
and U23932 (N_23932,N_20071,N_19670);
nand U23933 (N_23933,N_20289,N_19645);
and U23934 (N_23934,N_18500,N_18199);
and U23935 (N_23935,N_18045,N_18319);
and U23936 (N_23936,N_19922,N_19308);
or U23937 (N_23937,N_19217,N_20742);
nand U23938 (N_23938,N_18120,N_19121);
and U23939 (N_23939,N_20641,N_19367);
nor U23940 (N_23940,N_20075,N_18937);
nand U23941 (N_23941,N_19229,N_19485);
or U23942 (N_23942,N_18133,N_18917);
nor U23943 (N_23943,N_18677,N_19799);
nor U23944 (N_23944,N_19268,N_18137);
nand U23945 (N_23945,N_19223,N_18909);
nor U23946 (N_23946,N_19922,N_18866);
or U23947 (N_23947,N_19997,N_19322);
xnor U23948 (N_23948,N_19234,N_20209);
or U23949 (N_23949,N_19583,N_18984);
nor U23950 (N_23950,N_20303,N_18729);
nor U23951 (N_23951,N_19502,N_18327);
and U23952 (N_23952,N_20261,N_20880);
nand U23953 (N_23953,N_19604,N_18699);
or U23954 (N_23954,N_19764,N_18184);
xor U23955 (N_23955,N_18803,N_19324);
nor U23956 (N_23956,N_20863,N_20915);
xnor U23957 (N_23957,N_18399,N_19921);
xor U23958 (N_23958,N_19143,N_19409);
nand U23959 (N_23959,N_19631,N_18572);
or U23960 (N_23960,N_20626,N_19659);
nand U23961 (N_23961,N_18914,N_19278);
or U23962 (N_23962,N_19988,N_20482);
or U23963 (N_23963,N_19466,N_20615);
and U23964 (N_23964,N_20180,N_19722);
xnor U23965 (N_23965,N_19825,N_18788);
or U23966 (N_23966,N_19297,N_19920);
xor U23967 (N_23967,N_18732,N_20551);
or U23968 (N_23968,N_20591,N_19334);
nor U23969 (N_23969,N_18336,N_18043);
or U23970 (N_23970,N_19548,N_19435);
nor U23971 (N_23971,N_19911,N_18015);
or U23972 (N_23972,N_18308,N_20323);
and U23973 (N_23973,N_18068,N_20076);
nor U23974 (N_23974,N_20035,N_20688);
or U23975 (N_23975,N_20532,N_19306);
nand U23976 (N_23976,N_18439,N_18713);
or U23977 (N_23977,N_20761,N_19799);
xor U23978 (N_23978,N_20898,N_19860);
nand U23979 (N_23979,N_19523,N_19639);
or U23980 (N_23980,N_20730,N_18117);
nand U23981 (N_23981,N_19084,N_18701);
nor U23982 (N_23982,N_18336,N_19499);
and U23983 (N_23983,N_20970,N_19549);
nand U23984 (N_23984,N_18381,N_20217);
xor U23985 (N_23985,N_18140,N_19433);
or U23986 (N_23986,N_18827,N_18493);
xor U23987 (N_23987,N_19677,N_18040);
xor U23988 (N_23988,N_18411,N_20611);
or U23989 (N_23989,N_20265,N_19332);
nor U23990 (N_23990,N_18516,N_19767);
nor U23991 (N_23991,N_19586,N_18986);
nand U23992 (N_23992,N_20330,N_18939);
nor U23993 (N_23993,N_18758,N_19109);
xnor U23994 (N_23994,N_20208,N_18121);
or U23995 (N_23995,N_18029,N_20316);
nand U23996 (N_23996,N_20420,N_19424);
nand U23997 (N_23997,N_18314,N_20453);
or U23998 (N_23998,N_19899,N_19602);
and U23999 (N_23999,N_19437,N_19808);
xnor U24000 (N_24000,N_23621,N_21984);
nor U24001 (N_24001,N_22763,N_23952);
xor U24002 (N_24002,N_23410,N_23988);
xor U24003 (N_24003,N_21365,N_23237);
and U24004 (N_24004,N_23830,N_22084);
nor U24005 (N_24005,N_21171,N_21946);
or U24006 (N_24006,N_22679,N_23177);
xnor U24007 (N_24007,N_22955,N_21545);
or U24008 (N_24008,N_23438,N_22009);
and U24009 (N_24009,N_22116,N_23972);
and U24010 (N_24010,N_22282,N_21113);
nand U24011 (N_24011,N_22767,N_23366);
or U24012 (N_24012,N_22622,N_21093);
or U24013 (N_24013,N_21190,N_22978);
xnor U24014 (N_24014,N_23453,N_22214);
nor U24015 (N_24015,N_22958,N_22405);
nor U24016 (N_24016,N_23036,N_21947);
or U24017 (N_24017,N_23164,N_23877);
and U24018 (N_24018,N_21852,N_23535);
nand U24019 (N_24019,N_23662,N_22764);
nand U24020 (N_24020,N_23484,N_22965);
nand U24021 (N_24021,N_23132,N_22065);
xnor U24022 (N_24022,N_23476,N_21998);
nand U24023 (N_24023,N_22204,N_21121);
nand U24024 (N_24024,N_21359,N_21868);
and U24025 (N_24025,N_23914,N_23992);
nand U24026 (N_24026,N_22423,N_21301);
nor U24027 (N_24027,N_21576,N_22926);
and U24028 (N_24028,N_21245,N_22010);
nand U24029 (N_24029,N_21367,N_23383);
and U24030 (N_24030,N_22143,N_21199);
xnor U24031 (N_24031,N_23031,N_22513);
nand U24032 (N_24032,N_22520,N_21765);
xor U24033 (N_24033,N_22480,N_22422);
nor U24034 (N_24034,N_22177,N_22355);
nand U24035 (N_24035,N_21914,N_21202);
nor U24036 (N_24036,N_22671,N_21858);
xor U24037 (N_24037,N_22791,N_23214);
nand U24038 (N_24038,N_22979,N_21971);
xnor U24039 (N_24039,N_21102,N_21944);
nand U24040 (N_24040,N_22882,N_21471);
nor U24041 (N_24041,N_22085,N_21683);
nand U24042 (N_24042,N_23599,N_23794);
nor U24043 (N_24043,N_21494,N_23879);
or U24044 (N_24044,N_21784,N_21414);
and U24045 (N_24045,N_22318,N_21303);
and U24046 (N_24046,N_21571,N_23720);
or U24047 (N_24047,N_21737,N_22505);
nor U24048 (N_24048,N_22275,N_21641);
nor U24049 (N_24049,N_21867,N_21838);
nand U24050 (N_24050,N_21486,N_22596);
nor U24051 (N_24051,N_22139,N_22709);
and U24052 (N_24052,N_22160,N_23334);
or U24053 (N_24053,N_21442,N_21011);
and U24054 (N_24054,N_23417,N_23895);
and U24055 (N_24055,N_21636,N_23746);
nand U24056 (N_24056,N_22225,N_23270);
nand U24057 (N_24057,N_22776,N_21297);
or U24058 (N_24058,N_21279,N_23550);
nor U24059 (N_24059,N_22155,N_21770);
or U24060 (N_24060,N_21813,N_21862);
xor U24061 (N_24061,N_23886,N_23773);
xnor U24062 (N_24062,N_22723,N_21308);
nor U24063 (N_24063,N_23816,N_21273);
xnor U24064 (N_24064,N_23595,N_21752);
xor U24065 (N_24065,N_21083,N_22019);
and U24066 (N_24066,N_21272,N_23456);
nor U24067 (N_24067,N_22445,N_22238);
and U24068 (N_24068,N_23306,N_21440);
and U24069 (N_24069,N_22687,N_22025);
or U24070 (N_24070,N_22855,N_22852);
nor U24071 (N_24071,N_22298,N_21022);
or U24072 (N_24072,N_22525,N_21699);
nand U24073 (N_24073,N_23011,N_23931);
xnor U24074 (N_24074,N_23087,N_23471);
or U24075 (N_24075,N_22583,N_21812);
nand U24076 (N_24076,N_22031,N_23154);
and U24077 (N_24077,N_23806,N_22786);
or U24078 (N_24078,N_23543,N_23465);
xor U24079 (N_24079,N_22384,N_21969);
xor U24080 (N_24080,N_21695,N_22839);
and U24081 (N_24081,N_22293,N_21747);
xor U24082 (N_24082,N_23677,N_23867);
nand U24083 (N_24083,N_22798,N_22544);
and U24084 (N_24084,N_21891,N_22416);
xor U24085 (N_24085,N_21778,N_21403);
nand U24086 (N_24086,N_23586,N_22655);
nand U24087 (N_24087,N_22317,N_22372);
nor U24088 (N_24088,N_22195,N_21415);
nor U24089 (N_24089,N_23745,N_23754);
and U24090 (N_24090,N_23212,N_23182);
xor U24091 (N_24091,N_23887,N_23752);
nand U24092 (N_24092,N_23812,N_21251);
xnor U24093 (N_24093,N_23184,N_23292);
or U24094 (N_24094,N_21192,N_21108);
nor U24095 (N_24095,N_23810,N_23198);
and U24096 (N_24096,N_23430,N_23679);
and U24097 (N_24097,N_23285,N_23555);
or U24098 (N_24098,N_21532,N_22280);
xor U24099 (N_24099,N_22847,N_23847);
or U24100 (N_24100,N_22610,N_21421);
nand U24101 (N_24101,N_23315,N_23638);
and U24102 (N_24102,N_23670,N_23842);
or U24103 (N_24103,N_23829,N_23160);
or U24104 (N_24104,N_21012,N_22913);
nor U24105 (N_24105,N_22130,N_23464);
nand U24106 (N_24106,N_23788,N_21363);
nor U24107 (N_24107,N_21933,N_23710);
and U24108 (N_24108,N_23560,N_23910);
or U24109 (N_24109,N_23678,N_21227);
xnor U24110 (N_24110,N_23071,N_23823);
nor U24111 (N_24111,N_23900,N_22600);
xor U24112 (N_24112,N_22069,N_23561);
xnor U24113 (N_24113,N_21476,N_23461);
nor U24114 (N_24114,N_22050,N_22620);
or U24115 (N_24115,N_22093,N_23520);
or U24116 (N_24116,N_23050,N_21943);
or U24117 (N_24117,N_21579,N_21934);
nor U24118 (N_24118,N_23103,N_23717);
nand U24119 (N_24119,N_21529,N_22587);
nor U24120 (N_24120,N_21470,N_23431);
nand U24121 (N_24121,N_21617,N_23674);
nand U24122 (N_24122,N_22234,N_21066);
and U24123 (N_24123,N_21963,N_22412);
nor U24124 (N_24124,N_21788,N_22098);
or U24125 (N_24125,N_23331,N_22346);
nand U24126 (N_24126,N_21473,N_23147);
nand U24127 (N_24127,N_21268,N_21509);
or U24128 (N_24128,N_22117,N_21091);
nand U24129 (N_24129,N_23015,N_23848);
or U24130 (N_24130,N_23739,N_23922);
nand U24131 (N_24131,N_21352,N_22656);
xor U24132 (N_24132,N_21131,N_22083);
xor U24133 (N_24133,N_23094,N_23001);
and U24134 (N_24134,N_22780,N_23907);
and U24135 (N_24135,N_23322,N_23409);
or U24136 (N_24136,N_21158,N_23042);
or U24137 (N_24137,N_23023,N_22636);
xor U24138 (N_24138,N_23018,N_23704);
xnor U24139 (N_24139,N_23281,N_22023);
or U24140 (N_24140,N_23296,N_23457);
nor U24141 (N_24141,N_22758,N_22621);
xor U24142 (N_24142,N_22945,N_22518);
and U24143 (N_24143,N_23188,N_22822);
and U24144 (N_24144,N_22411,N_23753);
xor U24145 (N_24145,N_22503,N_22916);
and U24146 (N_24146,N_23303,N_21446);
xnor U24147 (N_24147,N_21300,N_22331);
nor U24148 (N_24148,N_21334,N_22987);
or U24149 (N_24149,N_21890,N_23379);
and U24150 (N_24150,N_21089,N_21926);
or U24151 (N_24151,N_23722,N_22438);
xnor U24152 (N_24152,N_21003,N_22894);
nand U24153 (N_24153,N_23013,N_22850);
and U24154 (N_24154,N_22860,N_22435);
nand U24155 (N_24155,N_21389,N_23458);
xor U24156 (N_24156,N_22296,N_23712);
and U24157 (N_24157,N_22733,N_23882);
xor U24158 (N_24158,N_23008,N_23658);
and U24159 (N_24159,N_21733,N_23771);
nand U24160 (N_24160,N_22256,N_23192);
and U24161 (N_24161,N_23064,N_21793);
xor U24162 (N_24162,N_22768,N_23928);
xnor U24163 (N_24163,N_23267,N_21729);
xor U24164 (N_24164,N_22419,N_21225);
nand U24165 (N_24165,N_21647,N_21217);
or U24166 (N_24166,N_23191,N_23761);
nand U24167 (N_24167,N_23868,N_23028);
nand U24168 (N_24168,N_21327,N_22012);
nand U24169 (N_24169,N_21013,N_23547);
or U24170 (N_24170,N_23994,N_21981);
nand U24171 (N_24171,N_23261,N_23903);
and U24172 (N_24172,N_23479,N_21357);
xnor U24173 (N_24173,N_22273,N_21704);
nor U24174 (N_24174,N_23120,N_23143);
or U24175 (N_24175,N_22429,N_21856);
or U24176 (N_24176,N_21652,N_21205);
nor U24177 (N_24177,N_23259,N_21060);
nor U24178 (N_24178,N_23901,N_22404);
xor U24179 (N_24179,N_21761,N_21086);
or U24180 (N_24180,N_22255,N_21696);
nand U24181 (N_24181,N_22936,N_22581);
nor U24182 (N_24182,N_22672,N_23571);
xnor U24183 (N_24183,N_21691,N_23386);
nor U24184 (N_24184,N_23568,N_23302);
and U24185 (N_24185,N_21407,N_21062);
nor U24186 (N_24186,N_21372,N_21749);
nor U24187 (N_24187,N_21449,N_23148);
nor U24188 (N_24188,N_23528,N_21458);
nand U24189 (N_24189,N_21193,N_23820);
nand U24190 (N_24190,N_22848,N_23396);
and U24191 (N_24191,N_21700,N_22729);
nand U24192 (N_24192,N_23022,N_22568);
or U24193 (N_24193,N_22585,N_23956);
or U24194 (N_24194,N_22618,N_22719);
nor U24195 (N_24195,N_21275,N_22030);
nor U24196 (N_24196,N_21779,N_23858);
xor U24197 (N_24197,N_23387,N_23144);
xnor U24198 (N_24198,N_21750,N_22515);
xnor U24199 (N_24199,N_22543,N_23522);
xor U24200 (N_24200,N_21094,N_22647);
and U24201 (N_24201,N_21680,N_23740);
nor U24202 (N_24202,N_21951,N_21924);
or U24203 (N_24203,N_22036,N_23973);
or U24204 (N_24204,N_22260,N_23989);
and U24205 (N_24205,N_21855,N_21870);
nor U24206 (N_24206,N_22232,N_22113);
nor U24207 (N_24207,N_23365,N_22292);
or U24208 (N_24208,N_23680,N_22247);
and U24209 (N_24209,N_21212,N_22872);
and U24210 (N_24210,N_22315,N_22111);
and U24211 (N_24211,N_22027,N_21075);
nand U24212 (N_24212,N_22675,N_22920);
or U24213 (N_24213,N_21754,N_22481);
and U24214 (N_24214,N_21850,N_22948);
nand U24215 (N_24215,N_22836,N_22013);
or U24216 (N_24216,N_23216,N_22588);
xnor U24217 (N_24217,N_21625,N_23054);
and U24218 (N_24218,N_23240,N_22076);
nor U24219 (N_24219,N_22316,N_22952);
xor U24220 (N_24220,N_21716,N_23169);
nor U24221 (N_24221,N_22365,N_22577);
and U24222 (N_24222,N_23519,N_22519);
nor U24223 (N_24223,N_21533,N_22179);
or U24224 (N_24224,N_23570,N_23004);
nand U24225 (N_24225,N_22566,N_23363);
and U24226 (N_24226,N_22330,N_23529);
nor U24227 (N_24227,N_23787,N_23616);
nand U24228 (N_24228,N_21026,N_23539);
nand U24229 (N_24229,N_21954,N_23057);
and U24230 (N_24230,N_21336,N_21377);
xnor U24231 (N_24231,N_21459,N_22099);
xnor U24232 (N_24232,N_23220,N_21031);
or U24233 (N_24233,N_21499,N_22248);
xnor U24234 (N_24234,N_23055,N_22349);
nor U24235 (N_24235,N_22388,N_23052);
and U24236 (N_24236,N_21172,N_22614);
and U24237 (N_24237,N_22212,N_21772);
and U24238 (N_24238,N_23935,N_22998);
xor U24239 (N_24239,N_22601,N_23357);
nor U24240 (N_24240,N_21077,N_21601);
nor U24241 (N_24241,N_23927,N_21953);
nor U24242 (N_24242,N_21775,N_23501);
nand U24243 (N_24243,N_22259,N_23633);
and U24244 (N_24244,N_23862,N_21823);
nor U24245 (N_24245,N_22989,N_22868);
and U24246 (N_24246,N_23659,N_22569);
and U24247 (N_24247,N_22068,N_23970);
nor U24248 (N_24248,N_21834,N_22639);
xnor U24249 (N_24249,N_21719,N_21874);
nand U24250 (N_24250,N_23853,N_23174);
or U24251 (N_24251,N_22340,N_21540);
or U24252 (N_24252,N_22761,N_23872);
xor U24253 (N_24253,N_23737,N_21903);
nor U24254 (N_24254,N_21628,N_22714);
or U24255 (N_24255,N_21827,N_22870);
nand U24256 (N_24256,N_22443,N_23514);
nor U24257 (N_24257,N_22550,N_22322);
and U24258 (N_24258,N_23137,N_21718);
or U24259 (N_24259,N_23354,N_21991);
nand U24260 (N_24260,N_21067,N_21826);
and U24261 (N_24261,N_22348,N_21059);
or U24262 (N_24262,N_21349,N_22706);
and U24263 (N_24263,N_21546,N_21049);
or U24264 (N_24264,N_22746,N_23647);
or U24265 (N_24265,N_22563,N_21288);
nand U24266 (N_24266,N_22556,N_22135);
or U24267 (N_24267,N_21338,N_21588);
or U24268 (N_24268,N_21201,N_23286);
xor U24269 (N_24269,N_22575,N_23653);
nand U24270 (N_24270,N_22022,N_23832);
or U24271 (N_24271,N_23950,N_23074);
or U24272 (N_24272,N_21203,N_23005);
xor U24273 (N_24273,N_23797,N_21892);
xnor U24274 (N_24274,N_23609,N_21679);
nor U24275 (N_24275,N_23178,N_23038);
and U24276 (N_24276,N_22903,N_23685);
or U24277 (N_24277,N_23891,N_22444);
xor U24278 (N_24278,N_21702,N_22721);
nor U24279 (N_24279,N_23238,N_22873);
xnor U24280 (N_24280,N_21516,N_22686);
and U24281 (N_24281,N_23089,N_21005);
xnor U24282 (N_24282,N_23949,N_23146);
nor U24283 (N_24283,N_21046,N_23345);
or U24284 (N_24284,N_22536,N_21405);
or U24285 (N_24285,N_21237,N_22364);
nand U24286 (N_24286,N_21585,N_22947);
nor U24287 (N_24287,N_21606,N_23530);
nor U24288 (N_24288,N_21803,N_23093);
xnor U24289 (N_24289,N_21575,N_22222);
nor U24290 (N_24290,N_21910,N_23881);
xor U24291 (N_24291,N_22096,N_23524);
nand U24292 (N_24292,N_22199,N_22421);
or U24293 (N_24293,N_22912,N_23266);
and U24294 (N_24294,N_23051,N_21469);
nand U24295 (N_24295,N_22814,N_21942);
nor U24296 (N_24296,N_22984,N_21339);
nor U24297 (N_24297,N_23835,N_22000);
and U24298 (N_24298,N_23268,N_21810);
nand U24299 (N_24299,N_22172,N_23667);
nand U24300 (N_24300,N_21580,N_21880);
or U24301 (N_24301,N_22261,N_22194);
and U24302 (N_24302,N_22838,N_22286);
xnor U24303 (N_24303,N_21615,N_23111);
or U24304 (N_24304,N_23825,N_21952);
and U24305 (N_24305,N_22593,N_23860);
nor U24306 (N_24306,N_23559,N_21650);
or U24307 (N_24307,N_23580,N_23855);
xnor U24308 (N_24308,N_23598,N_22991);
or U24309 (N_24309,N_21124,N_21298);
nand U24310 (N_24310,N_23567,N_22127);
nor U24311 (N_24311,N_23367,N_21391);
and U24312 (N_24312,N_21731,N_22402);
nor U24313 (N_24313,N_21116,N_21343);
nand U24314 (N_24314,N_22613,N_22967);
nand U24315 (N_24315,N_21786,N_23518);
and U24316 (N_24316,N_23579,N_22149);
or U24317 (N_24317,N_22227,N_23690);
and U24318 (N_24318,N_23236,N_22919);
xor U24319 (N_24319,N_23856,N_22245);
nand U24320 (N_24320,N_22157,N_23772);
and U24321 (N_24321,N_23557,N_21655);
nand U24322 (N_24322,N_22762,N_21692);
nor U24323 (N_24323,N_21309,N_23516);
nor U24324 (N_24324,N_21590,N_21767);
xnor U24325 (N_24325,N_22694,N_23702);
or U24326 (N_24326,N_22980,N_21435);
xnor U24327 (N_24327,N_21474,N_22026);
xnor U24328 (N_24328,N_23705,N_21422);
nand U24329 (N_24329,N_22506,N_21787);
or U24330 (N_24330,N_22399,N_23817);
and U24331 (N_24331,N_23070,N_23328);
and U24332 (N_24332,N_22934,N_22333);
or U24333 (N_24333,N_23030,N_21229);
and U24334 (N_24334,N_21222,N_22005);
nand U24335 (N_24335,N_22815,N_22643);
nand U24336 (N_24336,N_23415,N_23210);
and U24337 (N_24337,N_21063,N_21829);
or U24338 (N_24338,N_22409,N_23003);
nand U24339 (N_24339,N_21353,N_22570);
xor U24340 (N_24340,N_23946,N_23061);
and U24341 (N_24341,N_22307,N_22832);
and U24342 (N_24342,N_22862,N_21137);
or U24343 (N_24343,N_22203,N_22477);
xor U24344 (N_24344,N_22864,N_22827);
and U24345 (N_24345,N_23181,N_22207);
and U24346 (N_24346,N_21697,N_22299);
or U24347 (N_24347,N_22757,N_21189);
and U24348 (N_24348,N_23116,N_23246);
or U24349 (N_24349,N_23814,N_22810);
or U24350 (N_24350,N_21672,N_21748);
nor U24351 (N_24351,N_23955,N_23156);
or U24352 (N_24352,N_21634,N_22304);
and U24353 (N_24353,N_21538,N_23346);
nor U24354 (N_24354,N_23958,N_23122);
or U24355 (N_24355,N_23002,N_23876);
xnor U24356 (N_24356,N_21651,N_22526);
nor U24357 (N_24357,N_23280,N_23849);
nand U24358 (N_24358,N_23977,N_22779);
or U24359 (N_24359,N_21935,N_23779);
xor U24360 (N_24360,N_23091,N_23092);
nor U24361 (N_24361,N_22849,N_22262);
nand U24362 (N_24362,N_22028,N_23587);
and U24363 (N_24363,N_21569,N_21746);
nor U24364 (N_24364,N_22996,N_21751);
nor U24365 (N_24365,N_23827,N_22825);
nand U24366 (N_24366,N_23399,N_21381);
nand U24367 (N_24367,N_23698,N_22181);
or U24368 (N_24368,N_21004,N_21883);
nand U24369 (N_24369,N_23209,N_21147);
nand U24370 (N_24370,N_23460,N_23324);
xnor U24371 (N_24371,N_22042,N_21138);
nand U24372 (N_24372,N_23067,N_22734);
and U24373 (N_24373,N_21281,N_22020);
nand U24374 (N_24374,N_21399,N_22890);
nand U24375 (N_24375,N_23026,N_21962);
or U24376 (N_24376,N_21082,N_22125);
and U24377 (N_24377,N_21148,N_21564);
or U24378 (N_24378,N_21648,N_21658);
xor U24379 (N_24379,N_22001,N_21785);
and U24380 (N_24380,N_21987,N_23128);
or U24381 (N_24381,N_21909,N_22521);
xor U24382 (N_24382,N_22535,N_22724);
and U24383 (N_24383,N_21286,N_22871);
xor U24384 (N_24384,N_23252,N_22564);
nand U24385 (N_24385,N_21065,N_23890);
or U24386 (N_24386,N_21197,N_21837);
xor U24387 (N_24387,N_21736,N_22403);
nor U24388 (N_24388,N_23839,N_22891);
xor U24389 (N_24389,N_21875,N_23158);
nand U24390 (N_24390,N_22442,N_23938);
nor U24391 (N_24391,N_21491,N_23371);
or U24392 (N_24392,N_22052,N_21493);
nor U24393 (N_24393,N_22830,N_23919);
or U24394 (N_24394,N_22252,N_23079);
xnor U24395 (N_24395,N_22151,N_22276);
nand U24396 (N_24396,N_22866,N_21815);
nor U24397 (N_24397,N_21774,N_22743);
or U24398 (N_24398,N_22347,N_23358);
nor U24399 (N_24399,N_21295,N_22059);
and U24400 (N_24400,N_21723,N_21234);
xor U24401 (N_24401,N_22705,N_22358);
nand U24402 (N_24402,N_22826,N_21743);
and U24403 (N_24403,N_21503,N_21966);
or U24404 (N_24404,N_21605,N_22617);
xnor U24405 (N_24405,N_23414,N_23153);
or U24406 (N_24406,N_23791,N_21356);
nor U24407 (N_24407,N_22278,N_22962);
xnor U24408 (N_24408,N_23392,N_22385);
nand U24409 (N_24409,N_22792,N_22156);
nor U24410 (N_24410,N_21355,N_21574);
or U24411 (N_24411,N_22797,N_21110);
or U24412 (N_24412,N_22677,N_22327);
and U24413 (N_24413,N_23707,N_21956);
or U24414 (N_24414,N_23000,N_23024);
nand U24415 (N_24415,N_23470,N_21671);
and U24416 (N_24416,N_22021,N_23915);
or U24417 (N_24417,N_22611,N_23715);
nand U24418 (N_24418,N_23778,N_22586);
xor U24419 (N_24419,N_23614,N_23059);
nor U24420 (N_24420,N_23044,N_22073);
nand U24421 (N_24421,N_21000,N_22641);
xor U24422 (N_24422,N_23603,N_21805);
nand U24423 (N_24423,N_23673,N_22562);
nor U24424 (N_24424,N_21687,N_21006);
nor U24425 (N_24425,N_23504,N_22484);
xnor U24426 (N_24426,N_23100,N_21475);
nor U24427 (N_24427,N_22904,N_23606);
or U24428 (N_24428,N_22942,N_21587);
xor U24429 (N_24429,N_23506,N_23749);
nand U24430 (N_24430,N_23736,N_21163);
nor U24431 (N_24431,N_21889,N_23083);
nand U24432 (N_24432,N_21453,N_23796);
nand U24433 (N_24433,N_22367,N_23462);
and U24434 (N_24434,N_23581,N_21487);
nand U24435 (N_24435,N_21975,N_23766);
or U24436 (N_24436,N_22909,N_21835);
and U24437 (N_24437,N_22753,N_21328);
and U24438 (N_24438,N_21708,N_22279);
and U24439 (N_24439,N_22966,N_22198);
and U24440 (N_24440,N_22615,N_23645);
or U24441 (N_24441,N_22314,N_23343);
nor U24442 (N_24442,N_21174,N_23339);
or U24443 (N_24443,N_22141,N_23811);
nor U24444 (N_24444,N_21782,N_23951);
nand U24445 (N_24445,N_22329,N_21264);
nand U24446 (N_24446,N_21964,N_22071);
nor U24447 (N_24447,N_23552,N_22213);
or U24448 (N_24448,N_21017,N_21550);
or U24449 (N_24449,N_22311,N_23250);
nand U24450 (N_24450,N_23841,N_22016);
nand U24451 (N_24451,N_22136,N_21807);
nand U24452 (N_24452,N_23403,N_21167);
nand U24453 (N_24453,N_22108,N_22253);
xnor U24454 (N_24454,N_21982,N_22538);
nand U24455 (N_24455,N_22750,N_23434);
or U24456 (N_24456,N_22537,N_21893);
and U24457 (N_24457,N_22788,N_23774);
or U24458 (N_24458,N_23219,N_23613);
xnor U24459 (N_24459,N_22977,N_21836);
nor U24460 (N_24460,N_23545,N_21477);
and U24461 (N_24461,N_22877,N_21076);
and U24462 (N_24462,N_21958,N_21123);
and U24463 (N_24463,N_23300,N_22995);
nand U24464 (N_24464,N_22271,N_21613);
and U24465 (N_24465,N_22993,N_22634);
nand U24466 (N_24466,N_21898,N_21512);
nand U24467 (N_24467,N_23313,N_21895);
xor U24468 (N_24468,N_23892,N_22932);
xnor U24469 (N_24469,N_23009,N_21930);
and U24470 (N_24470,N_21115,N_22407);
nand U24471 (N_24471,N_23831,N_22501);
nand U24472 (N_24472,N_21348,N_22772);
xnor U24473 (N_24473,N_22003,N_21183);
nor U24474 (N_24474,N_22024,N_21596);
nor U24475 (N_24475,N_21515,N_22922);
xor U24476 (N_24476,N_23819,N_22376);
nand U24477 (N_24477,N_23447,N_21467);
nor U24478 (N_24478,N_22353,N_22215);
or U24479 (N_24479,N_21420,N_22997);
or U24480 (N_24480,N_21443,N_23728);
nand U24481 (N_24481,N_23969,N_23025);
xor U24482 (N_24482,N_21358,N_23218);
xnor U24483 (N_24483,N_23290,N_22661);
nor U24484 (N_24484,N_22992,N_22488);
and U24485 (N_24485,N_23764,N_23062);
nor U24486 (N_24486,N_21244,N_21848);
nand U24487 (N_24487,N_22453,N_23641);
nand U24488 (N_24488,N_21151,N_23512);
nand U24489 (N_24489,N_21559,N_23960);
nor U24490 (N_24490,N_22369,N_22976);
or U24491 (N_24491,N_21781,N_23584);
xor U24492 (N_24492,N_22756,N_23997);
nor U24493 (N_24493,N_22863,N_23205);
or U24494 (N_24494,N_22469,N_23375);
nor U24495 (N_24495,N_23523,N_21081);
or U24496 (N_24496,N_22164,N_21098);
or U24497 (N_24497,N_23897,N_23807);
nand U24498 (N_24498,N_22487,N_22133);
nor U24499 (N_24499,N_23691,N_22693);
or U24500 (N_24500,N_23724,N_21830);
and U24501 (N_24501,N_22389,N_21794);
or U24502 (N_24502,N_22580,N_22554);
or U24503 (N_24503,N_23077,N_22209);
nand U24504 (N_24504,N_21941,N_21053);
or U24505 (N_24505,N_23789,N_23213);
nor U24506 (N_24506,N_21937,N_21092);
nor U24507 (N_24507,N_21665,N_22146);
or U24508 (N_24508,N_22107,N_22841);
xnor U24509 (N_24509,N_23199,N_23696);
nand U24510 (N_24510,N_22165,N_21607);
or U24511 (N_24511,N_23006,N_21329);
and U24512 (N_24512,N_22783,N_23427);
xnor U24513 (N_24513,N_23834,N_21085);
or U24514 (N_24514,N_23634,N_21888);
nor U24515 (N_24515,N_22582,N_23335);
or U24516 (N_24516,N_23118,N_23232);
nor U24517 (N_24517,N_22040,N_23047);
xor U24518 (N_24518,N_22387,N_22637);
nor U24519 (N_24519,N_22599,N_22778);
and U24520 (N_24520,N_21287,N_21999);
or U24521 (N_24521,N_23262,N_22785);
nor U24522 (N_24522,N_21169,N_22594);
nor U24523 (N_24523,N_23196,N_22152);
xnor U24524 (N_24524,N_22303,N_22801);
nand U24525 (N_24525,N_23119,N_21361);
nor U24526 (N_24526,N_21997,N_21056);
or U24527 (N_24527,N_23944,N_23107);
xor U24528 (N_24528,N_21530,N_21196);
or U24529 (N_24529,N_22674,N_21931);
nand U24530 (N_24530,N_21404,N_21134);
or U24531 (N_24531,N_22789,N_22450);
and U24532 (N_24532,N_21425,N_23364);
or U24533 (N_24533,N_22735,N_21160);
nand U24534 (N_24534,N_21236,N_21445);
xnor U24535 (N_24535,N_22845,N_23656);
or U24536 (N_24536,N_21316,N_23287);
nand U24537 (N_24537,N_23368,N_22478);
xor U24538 (N_24538,N_21143,N_23362);
or U24539 (N_24539,N_22631,N_22459);
or U24540 (N_24540,N_22185,N_22337);
and U24541 (N_24541,N_21438,N_23253);
nor U24542 (N_24542,N_22342,N_21468);
nor U24543 (N_24543,N_22288,N_21911);
nor U24544 (N_24544,N_23920,N_23846);
nor U24545 (N_24545,N_23359,N_23991);
or U24546 (N_24546,N_23433,N_22999);
or U24547 (N_24547,N_22041,N_21542);
or U24548 (N_24548,N_23808,N_21945);
nor U24549 (N_24549,N_21289,N_22471);
and U24550 (N_24550,N_21500,N_22887);
and U24551 (N_24551,N_22448,N_23592);
nand U24552 (N_24552,N_22857,N_21757);
nor U24553 (N_24553,N_21375,N_21632);
xor U24554 (N_24554,N_21908,N_23755);
nor U24555 (N_24555,N_22070,N_23953);
nand U24556 (N_24556,N_22014,N_22603);
or U24557 (N_24557,N_21208,N_21317);
xor U24558 (N_24558,N_21025,N_21675);
nand U24559 (N_24559,N_22885,N_22092);
or U24560 (N_24560,N_22738,N_21084);
or U24561 (N_24561,N_23845,N_21379);
or U24562 (N_24562,N_21497,N_22170);
and U24563 (N_24563,N_22032,N_22306);
and U24564 (N_24564,N_23747,N_22229);
or U24565 (N_24565,N_21221,N_21258);
or U24566 (N_24566,N_21795,N_22716);
or U24567 (N_24567,N_22906,N_21551);
nor U24568 (N_24568,N_23481,N_21558);
or U24569 (N_24569,N_22162,N_21248);
or U24570 (N_24570,N_22168,N_21010);
xnor U24571 (N_24571,N_21881,N_21955);
or U24572 (N_24572,N_22095,N_21256);
nor U24573 (N_24573,N_23485,N_22530);
and U24574 (N_24574,N_23500,N_23859);
or U24575 (N_24575,N_23454,N_21432);
nand U24576 (N_24576,N_22228,N_23027);
nand U24577 (N_24577,N_23301,N_23619);
xor U24578 (N_24578,N_22274,N_23016);
and U24579 (N_24579,N_22378,N_23637);
or U24580 (N_24580,N_21247,N_22954);
nand U24581 (N_24581,N_23642,N_21218);
nor U24582 (N_24582,N_21127,N_22775);
nor U24583 (N_24583,N_23600,N_22382);
or U24584 (N_24584,N_21598,N_23542);
and U24585 (N_24585,N_23532,N_23675);
nor U24586 (N_24586,N_23693,N_22119);
and U24587 (N_24587,N_21142,N_22251);
or U24588 (N_24588,N_21001,N_22426);
or U24589 (N_24589,N_23097,N_21078);
nand U24590 (N_24590,N_21114,N_22673);
or U24591 (N_24591,N_21396,N_23578);
xor U24592 (N_24592,N_22874,N_21326);
nand U24593 (N_24593,N_21041,N_21904);
nor U24594 (N_24594,N_21433,N_23923);
xnor U24595 (N_24595,N_21260,N_22496);
nor U24596 (N_24596,N_23437,N_23502);
or U24597 (N_24597,N_22676,N_23271);
and U24598 (N_24598,N_23323,N_21412);
nor U24599 (N_24599,N_21577,N_21548);
and U24600 (N_24600,N_22428,N_22557);
xnor U24601 (N_24601,N_21364,N_23703);
xor U24602 (N_24602,N_21369,N_21839);
and U24603 (N_24603,N_23496,N_21649);
and U24604 (N_24604,N_22844,N_22802);
and U24605 (N_24605,N_22663,N_23668);
nand U24606 (N_24606,N_22499,N_23215);
nor U24607 (N_24607,N_22502,N_21684);
nor U24608 (N_24608,N_21024,N_22334);
nand U24609 (N_24609,N_22191,N_22974);
nor U24610 (N_24610,N_21293,N_22698);
xor U24611 (N_24611,N_21175,N_21922);
nand U24612 (N_24612,N_21463,N_23727);
nor U24613 (N_24613,N_21411,N_22846);
or U24614 (N_24614,N_22142,N_21517);
xnor U24615 (N_24615,N_23446,N_21866);
nor U24616 (N_24616,N_22865,N_23330);
nor U24617 (N_24617,N_22559,N_21821);
nor U24618 (N_24618,N_21586,N_22470);
or U24619 (N_24619,N_23185,N_21156);
or U24620 (N_24620,N_22701,N_21007);
nor U24621 (N_24621,N_21016,N_22745);
nand U24622 (N_24622,N_22140,N_21630);
and U24623 (N_24623,N_23961,N_23971);
nand U24624 (N_24624,N_21825,N_23305);
nand U24625 (N_24625,N_23426,N_23167);
nand U24626 (N_24626,N_22938,N_23491);
nand U24627 (N_24627,N_23684,N_22138);
xnor U24628 (N_24628,N_22605,N_21032);
nand U24629 (N_24629,N_21583,N_21662);
or U24630 (N_24630,N_21323,N_23078);
and U24631 (N_24631,N_23152,N_22988);
or U24632 (N_24632,N_23439,N_23594);
xnor U24633 (N_24633,N_21796,N_21802);
and U24634 (N_24634,N_21990,N_21811);
and U24635 (N_24635,N_22268,N_23204);
nand U24636 (N_24636,N_21178,N_22077);
and U24637 (N_24637,N_22858,N_21734);
nand U24638 (N_24638,N_21029,N_22546);
nor U24639 (N_24639,N_23913,N_21070);
or U24640 (N_24640,N_21290,N_23505);
xor U24641 (N_24641,N_22751,N_23499);
nor U24642 (N_24642,N_22283,N_23942);
nand U24643 (N_24643,N_21527,N_22472);
xnor U24644 (N_24644,N_23828,N_22876);
nand U24645 (N_24645,N_21100,N_21074);
nand U24646 (N_24646,N_23309,N_23983);
nor U24647 (N_24647,N_23173,N_21153);
xnor U24648 (N_24648,N_21557,N_21136);
xor U24649 (N_24649,N_22956,N_23593);
and U24650 (N_24650,N_23799,N_21507);
xnor U24651 (N_24651,N_22047,N_21616);
nor U24652 (N_24652,N_21831,N_23615);
or U24653 (N_24653,N_21745,N_22824);
and U24654 (N_24654,N_22508,N_23957);
or U24655 (N_24655,N_21028,N_23477);
nor U24656 (N_24656,N_23276,N_21840);
xnor U24657 (N_24657,N_23565,N_21872);
and U24658 (N_24658,N_23577,N_22455);
and U24659 (N_24659,N_22354,N_23655);
xnor U24660 (N_24660,N_21664,N_22662);
and U24661 (N_24661,N_21900,N_21413);
xor U24662 (N_24662,N_21553,N_21383);
nand U24663 (N_24663,N_22178,N_22175);
nor U24664 (N_24664,N_21194,N_22061);
xor U24665 (N_24665,N_21635,N_23947);
xor U24666 (N_24666,N_23360,N_21573);
or U24667 (N_24667,N_21537,N_21619);
or U24668 (N_24668,N_22608,N_23106);
or U24669 (N_24669,N_22795,N_23189);
and U24670 (N_24670,N_23084,N_21970);
xor U24671 (N_24671,N_21242,N_21885);
and U24672 (N_24672,N_23272,N_22081);
and U24673 (N_24673,N_22773,N_22737);
nor U24674 (N_24674,N_23423,N_21656);
xor U24675 (N_24675,N_23202,N_22592);
and U24676 (N_24676,N_23194,N_21139);
nand U24677 (N_24677,N_23894,N_21832);
or U24678 (N_24678,N_23474,N_23917);
nand U24679 (N_24679,N_22118,N_22063);
xnor U24680 (N_24680,N_23497,N_22366);
nand U24681 (N_24681,N_23381,N_23332);
nand U24682 (N_24682,N_21209,N_22267);
xnor U24683 (N_24683,N_23697,N_23629);
or U24684 (N_24684,N_21071,N_23975);
and U24685 (N_24685,N_23984,N_21820);
nor U24686 (N_24686,N_23758,N_21531);
and U24687 (N_24687,N_23792,N_22653);
nor U24688 (N_24688,N_21478,N_22907);
or U24689 (N_24689,N_21995,N_21430);
and U24690 (N_24690,N_22831,N_21986);
or U24691 (N_24691,N_23932,N_23982);
or U24692 (N_24692,N_22297,N_23622);
nor U24693 (N_24693,N_23709,N_22835);
nor U24694 (N_24694,N_23384,N_23793);
xnor U24695 (N_24695,N_21129,N_21018);
xnor U24696 (N_24696,N_21155,N_21916);
or U24697 (N_24697,N_23436,N_21567);
xnor U24698 (N_24698,N_23802,N_23076);
xnor U24699 (N_24699,N_23289,N_21246);
xnor U24700 (N_24700,N_22668,N_23790);
xnor U24701 (N_24701,N_21498,N_22390);
nor U24702 (N_24702,N_21373,N_22100);
nor U24703 (N_24703,N_21220,N_23569);
nor U24704 (N_24704,N_23010,N_21602);
or U24705 (N_24705,N_22635,N_23782);
and U24706 (N_24706,N_23007,N_22739);
nand U24707 (N_24707,N_23780,N_21170);
or U24708 (N_24708,N_22823,N_22878);
or U24709 (N_24709,N_22398,N_22043);
nor U24710 (N_24710,N_21618,N_23875);
xnor U24711 (N_24711,N_21912,N_23843);
nor U24712 (N_24712,N_22167,N_22057);
nor U24713 (N_24713,N_21777,N_21261);
or U24714 (N_24714,N_23034,N_22491);
xnor U24715 (N_24715,N_22144,N_21693);
or U24716 (N_24716,N_23311,N_21873);
and U24717 (N_24717,N_23818,N_22432);
xor U24718 (N_24718,N_21690,N_21660);
nor U24719 (N_24719,N_23170,N_22363);
and U24720 (N_24720,N_22727,N_22468);
nor U24721 (N_24721,N_23597,N_22102);
xnor U24722 (N_24722,N_23822,N_22744);
and U24723 (N_24723,N_23291,N_22717);
or U24724 (N_24724,N_22964,N_21185);
and U24725 (N_24725,N_22211,N_22834);
nand U24726 (N_24726,N_22627,N_22290);
and U24727 (N_24727,N_22796,N_22931);
nor U24728 (N_24728,N_22441,N_22715);
xnor U24729 (N_24729,N_23589,N_21818);
nand U24730 (N_24730,N_22218,N_21448);
nand U24731 (N_24731,N_23596,N_21132);
nor U24732 (N_24732,N_21378,N_23750);
and U24733 (N_24733,N_21382,N_21927);
and U24734 (N_24734,N_23411,N_23566);
and U24735 (N_24735,N_22893,N_22134);
xnor U24736 (N_24736,N_21401,N_21522);
or U24737 (N_24737,N_21960,N_22731);
nand U24738 (N_24738,N_23726,N_23244);
nor U24739 (N_24739,N_21713,N_23911);
or U24740 (N_24740,N_23155,N_22532);
or U24741 (N_24741,N_21508,N_22633);
nand U24742 (N_24742,N_23242,N_21393);
nand U24743 (N_24743,N_21644,N_23711);
nand U24744 (N_24744,N_21058,N_23651);
nor U24745 (N_24745,N_22579,N_23068);
nand U24746 (N_24746,N_22046,N_22196);
or U24747 (N_24747,N_22029,N_22254);
xor U24748 (N_24748,N_23043,N_22373);
or U24749 (N_24749,N_22192,N_22345);
nand U24750 (N_24750,N_21681,N_23352);
xnor U24751 (N_24751,N_23388,N_21073);
nand U24752 (N_24752,N_21627,N_22033);
nand U24753 (N_24753,N_23563,N_23896);
xor U24754 (N_24754,N_23288,N_22558);
and U24755 (N_24755,N_23671,N_22049);
and U24756 (N_24756,N_22434,N_23325);
nand U24757 (N_24757,N_21019,N_23161);
and U24758 (N_24758,N_22524,N_23646);
nand U24759 (N_24759,N_22174,N_22258);
nor U24760 (N_24760,N_23265,N_22094);
nor U24761 (N_24761,N_21489,N_22759);
nand U24762 (N_24762,N_22129,N_22681);
nor U24763 (N_24763,N_23733,N_22380);
and U24764 (N_24764,N_21582,N_21790);
nor U24765 (N_24765,N_22090,N_22700);
nor U24766 (N_24766,N_23666,N_22567);
and U24767 (N_24767,N_21461,N_21721);
and U24768 (N_24768,N_21140,N_22702);
nor U24769 (N_24769,N_21667,N_21801);
nor U24770 (N_24770,N_22418,N_23398);
nand U24771 (N_24771,N_21107,N_23800);
nor U24772 (N_24772,N_22408,N_22208);
nor U24773 (N_24773,N_21936,N_21054);
nand U24774 (N_24774,N_23039,N_21313);
and U24775 (N_24775,N_21861,N_23195);
nor U24776 (N_24776,N_21565,N_21384);
or U24777 (N_24777,N_23233,N_23838);
nor U24778 (N_24778,N_21847,N_22576);
nor U24779 (N_24779,N_23730,N_21099);
nand U24780 (N_24780,N_21720,N_21233);
xnor U24781 (N_24781,N_21306,N_22697);
nor U24782 (N_24782,N_21330,N_21452);
nand U24783 (N_24783,N_21186,N_23451);
xor U24784 (N_24784,N_21715,N_23234);
and U24785 (N_24785,N_21145,N_22305);
nor U24786 (N_24786,N_23304,N_21701);
nor U24787 (N_24787,N_22774,N_22350);
xor U24788 (N_24788,N_22666,N_22625);
and U24789 (N_24789,N_23448,N_22859);
and U24790 (N_24790,N_22393,N_21481);
nand U24791 (N_24791,N_21210,N_22180);
and U24792 (N_24792,N_23889,N_22946);
or U24793 (N_24793,N_22748,N_21033);
nand U24794 (N_24794,N_21431,N_21195);
xnor U24795 (N_24795,N_22154,N_21771);
and U24796 (N_24796,N_22079,N_23225);
nor U24797 (N_24797,N_21591,N_22578);
nand U24798 (N_24798,N_22205,N_22713);
nor U24799 (N_24799,N_22902,N_21485);
and U24800 (N_24800,N_22612,N_23759);
and U24801 (N_24801,N_22335,N_23489);
nand U24802 (N_24802,N_22264,N_22362);
and U24803 (N_24803,N_23625,N_21228);
nor U24804 (N_24804,N_21224,N_21968);
nor U24805 (N_24805,N_23190,N_23959);
xor U24806 (N_24806,N_22089,N_21161);
xnor U24807 (N_24807,N_22602,N_23527);
and U24808 (N_24808,N_21180,N_21057);
and U24809 (N_24809,N_21637,N_23418);
or U24810 (N_24810,N_22794,N_21524);
nor U24811 (N_24811,N_22854,N_22510);
xor U24812 (N_24812,N_21090,N_21623);
nand U24813 (N_24813,N_23264,N_21521);
nand U24814 (N_24814,N_22121,N_21739);
xor U24815 (N_24815,N_22414,N_22534);
nand U24816 (N_24816,N_22494,N_23980);
or U24817 (N_24817,N_23372,N_21096);
and U24818 (N_24818,N_21111,N_23714);
xnor U24819 (N_24819,N_22541,N_22285);
or U24820 (N_24820,N_22861,N_21614);
and U24821 (N_24821,N_23987,N_23916);
nor U24822 (N_24822,N_22332,N_23507);
xnor U24823 (N_24823,N_22137,N_23588);
nand U24824 (N_24824,N_22875,N_23777);
xor U24825 (N_24825,N_22632,N_22514);
nor U24826 (N_24826,N_22482,N_21816);
or U24827 (N_24827,N_22106,N_23206);
xor U24828 (N_24828,N_22324,N_22840);
or U24829 (N_24829,N_21302,N_23072);
or U24830 (N_24830,N_23075,N_23544);
and U24831 (N_24831,N_21689,N_21216);
nor U24832 (N_24832,N_22752,N_21572);
xnor U24833 (N_24833,N_23429,N_22806);
xor U24834 (N_24834,N_21899,N_23729);
and U24835 (N_24835,N_22629,N_22712);
or U24836 (N_24836,N_22120,N_23385);
or U24837 (N_24837,N_23105,N_23377);
nor U24838 (N_24838,N_22295,N_23966);
and U24839 (N_24839,N_22527,N_22037);
and U24840 (N_24840,N_21267,N_22928);
xnor U24841 (N_24841,N_21204,N_22216);
and U24842 (N_24842,N_21488,N_23549);
nor U24843 (N_24843,N_23525,N_22960);
nor U24844 (N_24844,N_23933,N_23435);
or U24845 (N_24845,N_21918,N_22466);
or U24846 (N_24846,N_22901,N_22383);
nor U24847 (N_24847,N_21726,N_22386);
nand U24848 (N_24848,N_23664,N_22131);
xnor U24849 (N_24849,N_22781,N_21913);
or U24850 (N_24850,N_21525,N_23117);
and U24851 (N_24851,N_22821,N_23548);
xnor U24852 (N_24852,N_21162,N_21368);
or U24853 (N_24853,N_22201,N_23934);
nor U24854 (N_24854,N_22457,N_21423);
and U24855 (N_24855,N_22711,N_21257);
or U24856 (N_24856,N_23086,N_23734);
and U24857 (N_24857,N_23467,N_21597);
xor U24858 (N_24858,N_21639,N_21514);
nor U24859 (N_24859,N_22011,N_23487);
nor U24860 (N_24860,N_21502,N_22742);
and U24861 (N_24861,N_22226,N_21337);
or U24862 (N_24862,N_21159,N_22547);
nand U24863 (N_24863,N_22911,N_22881);
nor U24864 (N_24864,N_23443,N_22054);
nor U24865 (N_24865,N_21959,N_22344);
nor U24866 (N_24866,N_21240,N_23344);
xnor U24867 (N_24867,N_22939,N_22684);
or U24868 (N_24868,N_21042,N_23798);
xnor U24869 (N_24869,N_21249,N_21051);
and U24870 (N_24870,N_22820,N_21322);
nand U24871 (N_24871,N_21050,N_22193);
xor U24872 (N_24872,N_22374,N_23676);
or U24873 (N_24873,N_21472,N_23297);
or U24874 (N_24874,N_22272,N_21080);
nor U24875 (N_24875,N_23201,N_22007);
or U24876 (N_24876,N_22004,N_21387);
nor U24877 (N_24877,N_21611,N_21274);
xor U24878 (N_24878,N_23230,N_21284);
nand U24879 (N_24879,N_22495,N_21119);
nor U24880 (N_24880,N_23307,N_23186);
nand U24881 (N_24881,N_23999,N_21484);
nand U24882 (N_24882,N_23141,N_21462);
or U24883 (N_24883,N_21950,N_21118);
nand U24884 (N_24884,N_23748,N_22308);
xnor U24885 (N_24885,N_22640,N_21230);
xor U24886 (N_24886,N_21009,N_23687);
nand U24887 (N_24887,N_23945,N_22359);
and U24888 (N_24888,N_23058,N_22128);
nor U24889 (N_24889,N_22078,N_21657);
xor U24890 (N_24890,N_21865,N_23475);
nand U24891 (N_24891,N_21495,N_22424);
and U24892 (N_24892,N_22720,N_23870);
or U24893 (N_24893,N_22963,N_23056);
nand U24894 (N_24894,N_22941,N_21263);
nand U24895 (N_24895,N_21674,N_23706);
or U24896 (N_24896,N_22689,N_22182);
nor U24897 (N_24897,N_23163,N_21902);
xor U24898 (N_24898,N_23391,N_22927);
or U24899 (N_24899,N_23590,N_21666);
nand U24900 (N_24900,N_23906,N_21321);
nor U24901 (N_24901,N_23166,N_21417);
xor U24902 (N_24902,N_21511,N_21504);
or U24903 (N_24903,N_21465,N_23045);
nor U24904 (N_24904,N_23929,N_22528);
xnor U24905 (N_24905,N_21780,N_23871);
xor U24906 (N_24906,N_22161,N_23531);
xnor U24907 (N_24907,N_23993,N_21318);
xnor U24908 (N_24908,N_22328,N_23627);
nand U24909 (N_24909,N_22699,N_21426);
xnor U24910 (N_24910,N_21633,N_23492);
nand U24911 (N_24911,N_21030,N_22055);
xor U24912 (N_24912,N_22458,N_23221);
nand U24913 (N_24913,N_21101,N_23382);
and U24914 (N_24914,N_22242,N_21709);
and U24915 (N_24915,N_23786,N_23912);
nor U24916 (N_24916,N_21120,N_21126);
and U24917 (N_24917,N_22500,N_22985);
and U24918 (N_24918,N_22417,N_22233);
or U24919 (N_24919,N_22277,N_22726);
xnor U24920 (N_24920,N_21397,N_21520);
xor U24921 (N_24921,N_23483,N_22289);
nor U24922 (N_24922,N_23632,N_21506);
nor U24923 (N_24923,N_23974,N_23245);
nand U24924 (N_24924,N_23510,N_22765);
nand U24925 (N_24925,N_21897,N_22235);
xnor U24926 (N_24926,N_23361,N_22760);
or U24927 (N_24927,N_23327,N_22053);
or U24928 (N_24928,N_21350,N_21859);
and U24929 (N_24929,N_23540,N_22951);
xor U24930 (N_24930,N_21677,N_23440);
nor U24931 (N_24931,N_22708,N_21534);
or U24932 (N_24932,N_22669,N_23142);
or U24933 (N_24933,N_23251,N_22571);
xor U24934 (N_24934,N_21766,N_21768);
xnor U24935 (N_24935,N_21406,N_21157);
nor U24936 (N_24936,N_22665,N_23405);
xor U24937 (N_24937,N_22219,N_21165);
and U24938 (N_24938,N_22790,N_23157);
nand U24939 (N_24939,N_21603,N_22449);
xor U24940 (N_24940,N_22153,N_21996);
nand U24941 (N_24941,N_21663,N_21460);
and U24942 (N_24942,N_21271,N_22646);
xnor U24943 (N_24943,N_21622,N_21394);
and U24944 (N_24944,N_23864,N_23425);
and U24945 (N_24945,N_21940,N_23355);
or U24946 (N_24946,N_22843,N_22813);
or U24947 (N_24947,N_22310,N_23905);
and U24948 (N_24948,N_23321,N_21266);
xnor U24949 (N_24949,N_21371,N_22595);
nand U24950 (N_24950,N_23582,N_22112);
nand U24951 (N_24951,N_21211,N_23573);
nor U24952 (N_24952,N_21447,N_21360);
nand U24953 (N_24953,N_23450,N_22410);
nor U24954 (N_24954,N_21769,N_22413);
nor U24955 (N_24955,N_21668,N_23217);
xor U24956 (N_24956,N_21544,N_23976);
or U24957 (N_24957,N_22725,N_21842);
nand U24958 (N_24958,N_22045,N_23962);
or U24959 (N_24959,N_23115,N_22659);
xnor U24960 (N_24960,N_23121,N_22949);
nor U24961 (N_24961,N_22497,N_23630);
nor U24962 (N_24962,N_22935,N_23863);
xnor U24963 (N_24963,N_23416,N_23318);
nor U24964 (N_24964,N_23021,N_21418);
xor U24965 (N_24965,N_22375,N_23854);
and U24966 (N_24966,N_23762,N_21021);
nand U24967 (N_24967,N_22452,N_21038);
and U24968 (N_24968,N_21252,N_22427);
nand U24969 (N_24969,N_22109,N_23908);
and U24970 (N_24970,N_22644,N_21505);
xor U24971 (N_24971,N_22787,N_23338);
nand U24972 (N_24972,N_23247,N_22607);
xor U24973 (N_24973,N_21390,N_22490);
or U24974 (N_24974,N_21688,N_23610);
and U24975 (N_24975,N_23114,N_21044);
or U24976 (N_24976,N_22169,N_22048);
or U24977 (N_24977,N_21416,N_23449);
xnor U24978 (N_24978,N_23861,N_23104);
nand U24979 (N_24979,N_21896,N_21173);
nor U24980 (N_24980,N_21055,N_21061);
nand U24981 (N_24981,N_23493,N_22718);
and U24982 (N_24982,N_22101,N_23053);
nand U24983 (N_24983,N_21039,N_23256);
xnor U24984 (N_24984,N_21654,N_22420);
or U24985 (N_24985,N_23784,N_22326);
and U24986 (N_24986,N_21455,N_23986);
or U24987 (N_24987,N_22058,N_21844);
and U24988 (N_24988,N_21798,N_23769);
and U24989 (N_24989,N_22391,N_21562);
nor U24990 (N_24990,N_22250,N_22246);
or U24991 (N_24991,N_22339,N_23102);
nand U24992 (N_24992,N_22628,N_22529);
xnor U24993 (N_24993,N_21262,N_22467);
nor U24994 (N_24994,N_22728,N_23612);
and U24995 (N_24995,N_23572,N_22937);
nor U24996 (N_24996,N_21604,N_23326);
or U24997 (N_24997,N_22809,N_22561);
or U24998 (N_24998,N_22200,N_21168);
and U24999 (N_24999,N_22454,N_23918);
nand U25000 (N_25000,N_21424,N_22892);
nand U25001 (N_25001,N_23090,N_23312);
or U25002 (N_25002,N_21882,N_23511);
xnor U25003 (N_25003,N_21640,N_21753);
xnor U25004 (N_25004,N_21014,N_23775);
and U25005 (N_25005,N_21276,N_23241);
nor U25006 (N_25006,N_23413,N_23401);
and U25007 (N_25007,N_22392,N_22923);
or U25008 (N_25008,N_22189,N_23995);
and U25009 (N_25009,N_23888,N_23657);
nor U25010 (N_25010,N_21223,N_22741);
nand U25011 (N_25011,N_21929,N_23224);
xnor U25012 (N_25012,N_21549,N_23080);
or U25013 (N_25013,N_21919,N_22231);
and U25014 (N_25014,N_21386,N_22190);
and U25015 (N_25015,N_21589,N_23165);
and U25016 (N_25016,N_23258,N_23130);
and U25017 (N_25017,N_23490,N_21402);
or U25018 (N_25018,N_21109,N_22747);
nor U25019 (N_25019,N_22159,N_21841);
nand U25020 (N_25020,N_21905,N_23473);
and U25021 (N_25021,N_23099,N_22243);
or U25022 (N_25022,N_22929,N_22301);
nor U25023 (N_25023,N_23725,N_23228);
or U25024 (N_25024,N_21543,N_22670);
nor U25025 (N_25025,N_23785,N_23428);
or U25026 (N_25026,N_22682,N_21706);
and U25027 (N_25027,N_22291,N_23636);
nor U25028 (N_25028,N_21993,N_21294);
xor U25029 (N_25029,N_23562,N_22982);
nor U25030 (N_25030,N_22722,N_23336);
nor U25031 (N_25031,N_22898,N_23954);
or U25032 (N_25032,N_22512,N_22066);
or U25033 (N_25033,N_21762,N_22451);
nor U25034 (N_25034,N_21133,N_23294);
xnor U25035 (N_25035,N_22188,N_23649);
nand U25036 (N_25036,N_21806,N_23274);
nor U25037 (N_25037,N_23412,N_22645);
xnor U25038 (N_25038,N_21626,N_21048);
and U25039 (N_25039,N_23127,N_23468);
and U25040 (N_25040,N_21226,N_23941);
nand U25041 (N_25041,N_23498,N_22703);
and U25042 (N_25042,N_22396,N_23112);
or U25043 (N_25043,N_23110,N_22397);
nor U25044 (N_25044,N_22370,N_22433);
or U25045 (N_25045,N_22184,N_23688);
xor U25046 (N_25046,N_21351,N_22691);
xor U25047 (N_25047,N_23873,N_21215);
xnor U25048 (N_25048,N_22660,N_21670);
nand U25049 (N_25049,N_21988,N_21849);
nor U25050 (N_25050,N_23626,N_21291);
nor U25051 (N_25051,N_22736,N_21965);
xnor U25052 (N_25052,N_21187,N_21207);
nor U25053 (N_25053,N_22509,N_22953);
xor U25054 (N_25054,N_21219,N_21198);
nand U25055 (N_25055,N_22202,N_21980);
xnor U25056 (N_25056,N_21106,N_22969);
nor U25057 (N_25057,N_22884,N_21181);
and U25058 (N_25058,N_21104,N_23669);
or U25059 (N_25059,N_23591,N_23803);
nand U25060 (N_25060,N_23295,N_23731);
nor U25061 (N_25061,N_21141,N_23538);
and U25062 (N_25062,N_22173,N_21255);
nor U25063 (N_25063,N_23098,N_23073);
nor U25064 (N_25064,N_22828,N_22943);
nand U25065 (N_25065,N_21112,N_21730);
or U25066 (N_25066,N_22236,N_23179);
nor U25067 (N_25067,N_23254,N_22623);
or U25068 (N_25068,N_21869,N_21035);
and U25069 (N_25069,N_22807,N_22220);
nand U25070 (N_25070,N_21740,N_21985);
or U25071 (N_25071,N_22800,N_22244);
and U25072 (N_25072,N_22975,N_22560);
and U25073 (N_25073,N_22899,N_21776);
nor U25074 (N_25074,N_23376,N_21243);
nor U25075 (N_25075,N_21860,N_21184);
and U25076 (N_25076,N_22343,N_22777);
xor U25077 (N_25077,N_23175,N_22654);
or U25078 (N_25078,N_21682,N_23378);
nand U25079 (N_25079,N_22973,N_22097);
nor U25080 (N_25080,N_23686,N_22680);
and U25081 (N_25081,N_23223,N_22269);
or U25082 (N_25082,N_22522,N_22517);
nor U25083 (N_25083,N_22223,N_21324);
or U25084 (N_25084,N_23644,N_22658);
and U25085 (N_25085,N_21333,N_23159);
xor U25086 (N_25086,N_23937,N_22908);
or U25087 (N_25087,N_23035,N_23940);
nand U25088 (N_25088,N_22320,N_21282);
xnor U25089 (N_25089,N_22379,N_22368);
and U25090 (N_25090,N_22690,N_22970);
or U25091 (N_25091,N_23723,N_23756);
xnor U25092 (N_25092,N_23314,N_23964);
nor U25093 (N_25093,N_23537,N_23692);
nand U25094 (N_25094,N_22122,N_22539);
or U25095 (N_25095,N_23836,N_23904);
xor U25096 (N_25096,N_23689,N_21434);
nand U25097 (N_25097,N_21354,N_23229);
or U25098 (N_25098,N_21698,N_22018);
or U25099 (N_25099,N_23020,N_23207);
or U25100 (N_25100,N_22394,N_21722);
or U25101 (N_25101,N_23340,N_21312);
nor U25102 (N_25102,N_21015,N_21814);
and U25103 (N_25103,N_22657,N_21064);
and U25104 (N_25104,N_23795,N_21122);
xor U25105 (N_25105,N_22166,N_22381);
nor U25106 (N_25106,N_23948,N_23640);
nor U25107 (N_25107,N_22148,N_22425);
or U25108 (N_25108,N_21214,N_23546);
and U25109 (N_25109,N_23380,N_22067);
nand U25110 (N_25110,N_23063,N_21510);
and U25111 (N_25111,N_22035,N_22545);
xnor U25112 (N_25112,N_23996,N_21270);
nor U25113 (N_25113,N_22377,N_21593);
xnor U25114 (N_25114,N_23012,N_22755);
xnor U25115 (N_25115,N_22704,N_22082);
xor U25116 (N_25116,N_23395,N_23033);
and U25117 (N_25117,N_21932,N_23402);
xor U25118 (N_25118,N_21901,N_22707);
or U25119 (N_25119,N_23564,N_21166);
or U25120 (N_25120,N_21072,N_21182);
nand U25121 (N_25121,N_23299,N_23554);
xor U25122 (N_25122,N_21428,N_21555);
nand U25123 (N_25123,N_22456,N_23936);
xnor U25124 (N_25124,N_21388,N_22087);
nor U25125 (N_25125,N_23235,N_23065);
nand U25126 (N_25126,N_21864,N_21915);
and U25127 (N_25127,N_22474,N_23652);
xnor U25128 (N_25128,N_21717,N_21200);
nor U25129 (N_25129,N_22784,N_22695);
nor U25130 (N_25130,N_22511,N_23310);
and U25131 (N_25131,N_23445,N_21961);
or U25132 (N_25132,N_21146,N_22944);
and U25133 (N_25133,N_22240,N_23095);
xnor U25134 (N_25134,N_21427,N_23695);
xor U25135 (N_25135,N_23124,N_21232);
and U25136 (N_25136,N_22950,N_21299);
nor U25137 (N_25137,N_21105,N_22360);
or U25138 (N_25138,N_23208,N_23422);
and U25139 (N_25139,N_23041,N_21342);
xnor U25140 (N_25140,N_22361,N_22483);
nand U25141 (N_25141,N_22217,N_21763);
or U25142 (N_25142,N_22325,N_23732);
or U25143 (N_25143,N_22312,N_23665);
nand U25144 (N_25144,N_22678,N_22921);
nor U25145 (N_25145,N_23869,N_23719);
or U25146 (N_25146,N_21370,N_22114);
nor U25147 (N_25147,N_22309,N_22688);
nor U25148 (N_25148,N_23017,N_22088);
nand U25149 (N_25149,N_23123,N_21917);
xor U25150 (N_25150,N_23273,N_21341);
nand U25151 (N_25151,N_23601,N_21304);
xor U25152 (N_25152,N_22479,N_23060);
or U25153 (N_25153,N_21385,N_21760);
nor U25154 (N_25154,N_21037,N_21600);
nand U25155 (N_25155,N_22300,N_23660);
nor U25156 (N_25156,N_23136,N_22124);
nand U25157 (N_25157,N_23113,N_21566);
or U25158 (N_25158,N_21707,N_21560);
or U25159 (N_25159,N_22239,N_23459);
nor U25160 (N_25160,N_22008,N_21989);
or U25161 (N_25161,N_21191,N_21346);
nand U25162 (N_25162,N_23926,N_21408);
or U25163 (N_25163,N_21335,N_23751);
nand U25164 (N_25164,N_22817,N_23874);
and U25165 (N_25165,N_23503,N_21034);
xor U25166 (N_25166,N_21278,N_23048);
and U25167 (N_25167,N_21973,N_23985);
nor U25168 (N_25168,N_23407,N_22983);
nand U25169 (N_25169,N_23700,N_23200);
or U25170 (N_25170,N_21150,N_23187);
xnor U25171 (N_25171,N_22492,N_23408);
xnor U25172 (N_25172,N_22981,N_23283);
or U25173 (N_25173,N_21259,N_21479);
nand U25174 (N_25174,N_21887,N_23432);
nand U25175 (N_25175,N_21097,N_22933);
nor U25176 (N_25176,N_21612,N_23998);
xnor U25177 (N_25177,N_22889,N_21797);
nor U25178 (N_25178,N_23770,N_21992);
nor U25179 (N_25179,N_22968,N_22437);
and U25180 (N_25180,N_22461,N_22572);
nor U25181 (N_25181,N_22842,N_22171);
nor U25182 (N_25182,N_23419,N_21967);
or U25183 (N_25183,N_23902,N_21002);
and U25184 (N_25184,N_21645,N_23611);
nand U25185 (N_25185,N_23488,N_22516);
nor U25186 (N_25186,N_22918,N_22504);
nor U25187 (N_25187,N_22574,N_22851);
and U25188 (N_25188,N_23337,N_21599);
xnor U25189 (N_25189,N_22091,N_23708);
or U25190 (N_25190,N_23203,N_22287);
nor U25191 (N_25191,N_23421,N_21496);
nand U25192 (N_25192,N_21957,N_23193);
or U25193 (N_25193,N_21315,N_23574);
xnor U25194 (N_25194,N_23319,N_22683);
and U25195 (N_25195,N_23515,N_21876);
nand U25196 (N_25196,N_23096,N_22266);
xnor U25197 (N_25197,N_22351,N_22044);
or U25198 (N_25198,N_21974,N_21456);
nor U25199 (N_25199,N_23833,N_23968);
and U25200 (N_25200,N_23138,N_21631);
or U25201 (N_25201,N_21325,N_21079);
nor U25202 (N_25202,N_23032,N_22498);
and U25203 (N_25203,N_23049,N_23369);
nand U25204 (N_25204,N_23909,N_22017);
or U25205 (N_25205,N_23231,N_23180);
nand U25206 (N_25206,N_22914,N_23374);
nand U25207 (N_25207,N_22888,N_21925);
nand U25208 (N_25208,N_21344,N_22589);
nand U25209 (N_25209,N_21676,N_22060);
nand U25210 (N_25210,N_22804,N_23885);
and U25211 (N_25211,N_22692,N_22132);
and U25212 (N_25212,N_23298,N_21238);
nor U25213 (N_25213,N_23081,N_23508);
and U25214 (N_25214,N_23617,N_21164);
and U25215 (N_25215,N_23509,N_22880);
and U25216 (N_25216,N_22619,N_23151);
nand U25217 (N_25217,N_21920,N_21808);
xnor U25218 (N_25218,N_21239,N_23618);
nand U25219 (N_25219,N_23140,N_23257);
or U25220 (N_25220,N_23046,N_21653);
nor U25221 (N_25221,N_22533,N_21659);
nand U25222 (N_25222,N_21135,N_23226);
or U25223 (N_25223,N_23131,N_23767);
nor U25224 (N_25224,N_23347,N_23424);
xnor U25225 (N_25225,N_23480,N_22206);
and U25226 (N_25226,N_23541,N_22710);
nor U25227 (N_25227,N_22990,N_23040);
or U25228 (N_25228,N_21800,N_21994);
or U25229 (N_25229,N_21792,N_21027);
nand U25230 (N_25230,N_21592,N_23878);
xor U25231 (N_25231,N_23851,N_22476);
and U25232 (N_25232,N_21020,N_23893);
nand U25233 (N_25233,N_22341,N_21450);
xnor U25234 (N_25234,N_21419,N_23624);
xor U25235 (N_25235,N_22961,N_21755);
or U25236 (N_25236,N_23883,N_22696);
nand U25237 (N_25237,N_22905,N_21728);
nor U25238 (N_25238,N_21492,N_21789);
or U25239 (N_25239,N_23558,N_22856);
and U25240 (N_25240,N_21556,N_23126);
or U25241 (N_25241,N_23444,N_22464);
xor U25242 (N_25242,N_23222,N_22187);
and U25243 (N_25243,N_23350,N_22565);
and U25244 (N_25244,N_21878,N_22648);
and U25245 (N_25245,N_21087,N_21409);
nor U25246 (N_25246,N_21149,N_23320);
xnor U25247 (N_25247,N_23275,N_23899);
and U25248 (N_25248,N_22064,N_22323);
and U25249 (N_25249,N_21128,N_22606);
or U25250 (N_25250,N_23880,N_23672);
nand U25251 (N_25251,N_22263,N_23526);
or U25252 (N_25252,N_22357,N_22624);
xnor U25253 (N_25253,N_22638,N_21853);
nand U25254 (N_25254,N_22431,N_21519);
or U25255 (N_25255,N_23783,N_23585);
nand U25256 (N_25256,N_21457,N_21877);
xnor U25257 (N_25257,N_21362,N_22158);
and U25258 (N_25258,N_23643,N_22769);
nor U25259 (N_25259,N_23694,N_21144);
nor U25260 (N_25260,N_23329,N_22869);
nor U25261 (N_25261,N_21526,N_23308);
xnor U25262 (N_25262,N_21578,N_21117);
xnor U25263 (N_25263,N_21480,N_21285);
and U25264 (N_25264,N_23735,N_22086);
and U25265 (N_25265,N_22924,N_21483);
xnor U25266 (N_25266,N_21732,N_23837);
nor U25267 (N_25267,N_22626,N_21621);
nand U25268 (N_25268,N_21906,N_22110);
nor U25269 (N_25269,N_21735,N_22667);
xnor U25270 (N_25270,N_21296,N_23939);
and U25271 (N_25271,N_22080,N_22313);
or U25272 (N_25272,N_21206,N_21976);
xnor U25273 (N_25273,N_22805,N_21742);
nor U25274 (N_25274,N_22371,N_21314);
and U25275 (N_25275,N_21250,N_22270);
and U25276 (N_25276,N_23243,N_22910);
nor U25277 (N_25277,N_21436,N_22833);
nand U25278 (N_25278,N_23930,N_22163);
xor U25279 (N_25279,N_23466,N_23716);
nor U25280 (N_25280,N_23620,N_21871);
and U25281 (N_25281,N_23149,N_23813);
or U25282 (N_25282,N_23682,N_21879);
nor U25283 (N_25283,N_22548,N_21518);
nand U25284 (N_25284,N_22002,N_22754);
or U25285 (N_25285,N_23168,N_22473);
and U25286 (N_25286,N_22651,N_22284);
and U25287 (N_25287,N_22038,N_22819);
or U25288 (N_25288,N_23551,N_23763);
or U25289 (N_25289,N_21023,N_23400);
xnor U25290 (N_25290,N_23353,N_22732);
and U25291 (N_25291,N_21177,N_21398);
xnor U25292 (N_25292,N_23840,N_22531);
nand U25293 (N_25293,N_21241,N_21340);
xor U25294 (N_25294,N_22338,N_21712);
or U25295 (N_25295,N_21305,N_22356);
or U25296 (N_25296,N_21819,N_22486);
or U25297 (N_25297,N_23101,N_21646);
xor U25298 (N_25298,N_21380,N_21783);
nand U25299 (N_25299,N_23990,N_22740);
and U25300 (N_25300,N_21444,N_23279);
nor U25301 (N_25301,N_21972,N_23742);
nor U25302 (N_25302,N_23943,N_21629);
nand U25303 (N_25303,N_21724,N_21277);
or U25304 (N_25304,N_21886,N_23455);
nand U25305 (N_25305,N_22237,N_23082);
and U25306 (N_25306,N_23513,N_23277);
nor U25307 (N_25307,N_21764,N_21678);
and U25308 (N_25308,N_23260,N_21711);
and U25309 (N_25309,N_22446,N_21638);
and U25310 (N_25310,N_21983,N_23316);
nand U25311 (N_25311,N_21410,N_21609);
nand U25312 (N_25312,N_22650,N_23134);
nor U25313 (N_25313,N_22957,N_22039);
nand U25314 (N_25314,N_23495,N_21741);
or U25315 (N_25315,N_22523,N_22994);
and U25316 (N_25316,N_21833,N_22115);
or U25317 (N_25317,N_22616,N_21554);
or U25318 (N_25318,N_21978,N_22766);
nor U25319 (N_25319,N_23014,N_21437);
xor U25320 (N_25320,N_21799,N_22104);
or U25321 (N_25321,N_23227,N_23269);
and U25322 (N_25322,N_21938,N_22879);
or U25323 (N_25323,N_22493,N_22818);
xnor U25324 (N_25324,N_22186,N_23865);
or U25325 (N_25325,N_22590,N_21152);
nand U25326 (N_25326,N_23139,N_22883);
nor U25327 (N_25327,N_22224,N_23171);
nand U25328 (N_25328,N_22799,N_21523);
nor U25329 (N_25329,N_21366,N_22210);
or U25330 (N_25330,N_22915,N_23069);
or U25331 (N_25331,N_23393,N_22183);
or U25332 (N_25332,N_23172,N_21125);
nor U25333 (N_25333,N_21176,N_23921);
nor U25334 (N_25334,N_23967,N_22925);
nand U25335 (N_25335,N_23133,N_22971);
nand U25336 (N_25336,N_22542,N_21643);
xnor U25337 (N_25337,N_23575,N_23317);
and U25338 (N_25338,N_23469,N_22415);
nor U25339 (N_25339,N_21095,N_23824);
nor U25340 (N_25340,N_21454,N_21863);
or U25341 (N_25341,N_22230,N_23741);
nor U25342 (N_25342,N_23129,N_23608);
xor U25343 (N_25343,N_22460,N_22265);
xnor U25344 (N_25344,N_23701,N_22986);
xnor U25345 (N_25345,N_23866,N_22406);
nor U25346 (N_25346,N_23721,N_22221);
xor U25347 (N_25347,N_23341,N_21694);
nand U25348 (N_25348,N_22642,N_21594);
xor U25349 (N_25349,N_23650,N_22816);
or U25350 (N_25350,N_21846,N_21703);
nor U25351 (N_25351,N_23135,N_21547);
nor U25352 (N_25352,N_22436,N_21539);
xnor U25353 (N_25353,N_21466,N_21705);
nand U25354 (N_25354,N_23394,N_23125);
and U25355 (N_25355,N_21727,N_21332);
and U25356 (N_25356,N_21213,N_21809);
nor U25357 (N_25357,N_23348,N_22917);
nand U25358 (N_25358,N_21642,N_21843);
nor U25359 (N_25359,N_23804,N_23333);
and U25360 (N_25360,N_21154,N_21036);
nand U25361 (N_25361,N_21307,N_23801);
or U25362 (N_25362,N_22051,N_21103);
and U25363 (N_25363,N_22319,N_23183);
xor U25364 (N_25364,N_23963,N_22463);
nand U25365 (N_25365,N_23482,N_21347);
xnor U25366 (N_25366,N_21395,N_23420);
xnor U25367 (N_25367,N_22930,N_23370);
xnor U25368 (N_25368,N_21828,N_23494);
nand U25369 (N_25369,N_21857,N_22015);
xnor U25370 (N_25370,N_21490,N_21269);
or U25371 (N_25371,N_21374,N_22811);
nand U25372 (N_25372,N_23282,N_23898);
xor U25373 (N_25373,N_21939,N_22540);
nor U25374 (N_25374,N_23463,N_22895);
nand U25375 (N_25375,N_21008,N_23852);
and U25376 (N_25376,N_22896,N_23534);
and U25377 (N_25377,N_21845,N_23351);
and U25378 (N_25378,N_23263,N_22401);
nand U25379 (N_25379,N_22147,N_23850);
or U25380 (N_25380,N_22609,N_21824);
or U25381 (N_25381,N_23713,N_21235);
nor U25382 (N_25382,N_22972,N_23397);
nand U25383 (N_25383,N_23844,N_21725);
or U25384 (N_25384,N_22150,N_23576);
or U25385 (N_25385,N_23604,N_22395);
or U25386 (N_25386,N_21948,N_23925);
and U25387 (N_25387,N_23635,N_22465);
xnor U25388 (N_25388,N_21541,N_21710);
nor U25389 (N_25389,N_21441,N_23699);
nor U25390 (N_25390,N_21513,N_22145);
xnor U25391 (N_25391,N_23718,N_22430);
nand U25392 (N_25392,N_23607,N_23145);
and U25393 (N_25393,N_22056,N_23356);
xor U25394 (N_25394,N_22072,N_23805);
and U25395 (N_25395,N_23472,N_21283);
and U25396 (N_25396,N_22549,N_22439);
or U25397 (N_25397,N_21804,N_21254);
or U25398 (N_25398,N_23857,N_21043);
nand U25399 (N_25399,N_23605,N_22837);
nor U25400 (N_25400,N_22886,N_21907);
or U25401 (N_25401,N_23821,N_23776);
or U25402 (N_25402,N_21265,N_21758);
nor U25403 (N_25403,N_23517,N_21624);
nand U25404 (N_25404,N_21535,N_22034);
xnor U25405 (N_25405,N_21570,N_22940);
nor U25406 (N_25406,N_21528,N_23683);
and U25407 (N_25407,N_21331,N_21320);
xor U25408 (N_25408,N_21977,N_21620);
nand U25409 (N_25409,N_23744,N_22123);
nor U25410 (N_25410,N_21744,N_21451);
and U25411 (N_25411,N_23743,N_23278);
xnor U25412 (N_25412,N_23757,N_22793);
or U25413 (N_25413,N_23631,N_23654);
xnor U25414 (N_25414,N_22630,N_23809);
xnor U25415 (N_25415,N_22352,N_21536);
nand U25416 (N_25416,N_21345,N_22249);
nand U25417 (N_25417,N_23924,N_23373);
nand U25418 (N_25418,N_22552,N_23533);
xor U25419 (N_25419,N_23197,N_21311);
nand U25420 (N_25420,N_23760,N_21179);
or U25421 (N_25421,N_22475,N_21759);
nand U25422 (N_25422,N_22074,N_23981);
nand U25423 (N_25423,N_21894,N_23255);
and U25424 (N_25424,N_21052,N_22321);
or U25425 (N_25425,N_22598,N_23583);
nand U25426 (N_25426,N_21392,N_23681);
nor U25427 (N_25427,N_22400,N_21756);
nor U25428 (N_25428,N_22105,N_21822);
or U25429 (N_25429,N_22808,N_23826);
nand U25430 (N_25430,N_21568,N_23478);
xnor U25431 (N_25431,N_23781,N_21501);
nor U25432 (N_25432,N_23108,N_23248);
xnor U25433 (N_25433,N_23239,N_23556);
and U25434 (N_25434,N_21979,N_23815);
or U25435 (N_25435,N_21584,N_22803);
or U25436 (N_25436,N_22664,N_23404);
and U25437 (N_25437,N_22555,N_21045);
or U25438 (N_25438,N_23965,N_21231);
and U25439 (N_25439,N_23088,N_21552);
and U25440 (N_25440,N_21319,N_23109);
nor U25441 (N_25441,N_21923,N_23249);
nor U25442 (N_25442,N_22197,N_21464);
nand U25443 (N_25443,N_21088,N_22281);
nor U25444 (N_25444,N_21130,N_21400);
and U25445 (N_25445,N_23037,N_23628);
or U25446 (N_25446,N_21280,N_23019);
xor U25447 (N_25447,N_23342,N_22241);
or U25448 (N_25448,N_21673,N_23066);
nand U25449 (N_25449,N_21429,N_21817);
or U25450 (N_25450,N_22829,N_23452);
or U25451 (N_25451,N_21253,N_23623);
or U25452 (N_25452,N_21188,N_23284);
nand U25453 (N_25453,N_22584,N_23648);
or U25454 (N_25454,N_23765,N_23536);
and U25455 (N_25455,N_22853,N_22649);
nand U25456 (N_25456,N_23162,N_22447);
xor U25457 (N_25457,N_23293,N_22489);
or U25458 (N_25458,N_21563,N_22006);
and U25459 (N_25459,N_23390,N_21292);
or U25460 (N_25460,N_23389,N_23406);
xnor U25461 (N_25461,N_21773,N_22302);
and U25462 (N_25462,N_21561,N_21669);
nor U25463 (N_25463,N_21921,N_22812);
and U25464 (N_25464,N_22900,N_22294);
nor U25465 (N_25465,N_23176,N_21047);
or U25466 (N_25466,N_22604,N_21482);
or U25467 (N_25467,N_23639,N_21851);
and U25468 (N_25468,N_21595,N_23486);
xnor U25469 (N_25469,N_23661,N_22553);
nor U25470 (N_25470,N_23979,N_22103);
nand U25471 (N_25471,N_22440,N_23768);
and U25472 (N_25472,N_21714,N_21884);
or U25473 (N_25473,N_22551,N_22770);
xnor U25474 (N_25474,N_22485,N_21686);
nand U25475 (N_25475,N_22652,N_23602);
xor U25476 (N_25476,N_21854,N_21661);
and U25477 (N_25477,N_22126,N_21439);
and U25478 (N_25478,N_21738,N_22336);
xnor U25479 (N_25479,N_23738,N_22867);
and U25480 (N_25480,N_23150,N_22176);
nand U25481 (N_25481,N_22897,N_21040);
or U25482 (N_25482,N_21791,N_22782);
or U25483 (N_25483,N_23553,N_22507);
and U25484 (N_25484,N_23521,N_21610);
and U25485 (N_25485,N_22075,N_23029);
and U25486 (N_25486,N_22771,N_21068);
xnor U25487 (N_25487,N_21608,N_23884);
and U25488 (N_25488,N_23349,N_21069);
xnor U25489 (N_25489,N_21581,N_23442);
and U25490 (N_25490,N_22685,N_21685);
or U25491 (N_25491,N_21949,N_23085);
nand U25492 (N_25492,N_22257,N_21310);
nand U25493 (N_25493,N_21376,N_22462);
or U25494 (N_25494,N_22591,N_21928);
and U25495 (N_25495,N_23441,N_22597);
or U25496 (N_25496,N_22062,N_22573);
and U25497 (N_25497,N_22730,N_23211);
xnor U25498 (N_25498,N_22959,N_22749);
or U25499 (N_25499,N_23978,N_23663);
nor U25500 (N_25500,N_22795,N_22177);
nand U25501 (N_25501,N_23912,N_23254);
nand U25502 (N_25502,N_23585,N_23838);
or U25503 (N_25503,N_21173,N_22927);
and U25504 (N_25504,N_21339,N_22382);
nand U25505 (N_25505,N_22131,N_23001);
or U25506 (N_25506,N_23607,N_21878);
nand U25507 (N_25507,N_22631,N_21080);
xor U25508 (N_25508,N_21230,N_23491);
and U25509 (N_25509,N_21918,N_23761);
nand U25510 (N_25510,N_22182,N_22040);
nand U25511 (N_25511,N_23930,N_23349);
xor U25512 (N_25512,N_22266,N_21710);
nand U25513 (N_25513,N_23541,N_22474);
nor U25514 (N_25514,N_23389,N_21782);
xor U25515 (N_25515,N_22480,N_23712);
xnor U25516 (N_25516,N_22130,N_23587);
and U25517 (N_25517,N_23773,N_22174);
xor U25518 (N_25518,N_22652,N_21258);
and U25519 (N_25519,N_22957,N_21167);
nand U25520 (N_25520,N_21242,N_22010);
and U25521 (N_25521,N_22573,N_22773);
and U25522 (N_25522,N_23762,N_23302);
xor U25523 (N_25523,N_21584,N_22044);
or U25524 (N_25524,N_22062,N_22996);
nand U25525 (N_25525,N_22702,N_23749);
or U25526 (N_25526,N_21348,N_22042);
xor U25527 (N_25527,N_22421,N_21136);
nand U25528 (N_25528,N_23723,N_23488);
and U25529 (N_25529,N_23363,N_21399);
nor U25530 (N_25530,N_21488,N_23934);
nor U25531 (N_25531,N_23432,N_23334);
and U25532 (N_25532,N_21682,N_21606);
and U25533 (N_25533,N_21616,N_21135);
nor U25534 (N_25534,N_21786,N_21221);
or U25535 (N_25535,N_22264,N_22236);
xnor U25536 (N_25536,N_21859,N_22971);
nand U25537 (N_25537,N_22800,N_22729);
or U25538 (N_25538,N_23903,N_22540);
nand U25539 (N_25539,N_22413,N_23929);
and U25540 (N_25540,N_23979,N_22287);
or U25541 (N_25541,N_23409,N_22153);
xor U25542 (N_25542,N_21482,N_23551);
xor U25543 (N_25543,N_22380,N_23661);
nand U25544 (N_25544,N_23549,N_22878);
xnor U25545 (N_25545,N_21023,N_22464);
and U25546 (N_25546,N_23543,N_21779);
nor U25547 (N_25547,N_23351,N_22089);
nor U25548 (N_25548,N_21309,N_23756);
nand U25549 (N_25549,N_22879,N_21902);
and U25550 (N_25550,N_22428,N_22549);
nor U25551 (N_25551,N_22476,N_23537);
and U25552 (N_25552,N_22554,N_22005);
nor U25553 (N_25553,N_21096,N_21916);
nand U25554 (N_25554,N_21896,N_22392);
or U25555 (N_25555,N_23048,N_22095);
xnor U25556 (N_25556,N_21310,N_22895);
nor U25557 (N_25557,N_21835,N_23128);
nor U25558 (N_25558,N_22782,N_23912);
xor U25559 (N_25559,N_22015,N_22882);
xor U25560 (N_25560,N_21895,N_21653);
or U25561 (N_25561,N_22332,N_23783);
nand U25562 (N_25562,N_21551,N_22705);
or U25563 (N_25563,N_22516,N_22446);
and U25564 (N_25564,N_22578,N_21934);
nor U25565 (N_25565,N_21439,N_23641);
or U25566 (N_25566,N_23174,N_22513);
nand U25567 (N_25567,N_21561,N_22588);
nor U25568 (N_25568,N_23905,N_22184);
nor U25569 (N_25569,N_22861,N_21718);
xnor U25570 (N_25570,N_23211,N_21666);
and U25571 (N_25571,N_22453,N_23136);
nand U25572 (N_25572,N_23284,N_21565);
or U25573 (N_25573,N_23613,N_23527);
nand U25574 (N_25574,N_23396,N_23725);
nor U25575 (N_25575,N_22244,N_23191);
xnor U25576 (N_25576,N_23660,N_23567);
nor U25577 (N_25577,N_23150,N_23314);
nand U25578 (N_25578,N_21093,N_22944);
and U25579 (N_25579,N_22956,N_23854);
or U25580 (N_25580,N_23814,N_21215);
nor U25581 (N_25581,N_23750,N_22488);
and U25582 (N_25582,N_23244,N_21260);
nor U25583 (N_25583,N_23831,N_23923);
nor U25584 (N_25584,N_22678,N_23859);
or U25585 (N_25585,N_22602,N_23982);
nor U25586 (N_25586,N_21312,N_21169);
nor U25587 (N_25587,N_21301,N_21077);
xnor U25588 (N_25588,N_23770,N_22567);
nand U25589 (N_25589,N_23948,N_23592);
nand U25590 (N_25590,N_22210,N_23922);
and U25591 (N_25591,N_22214,N_22962);
or U25592 (N_25592,N_22365,N_21789);
nor U25593 (N_25593,N_21871,N_22168);
and U25594 (N_25594,N_21626,N_23318);
nand U25595 (N_25595,N_23414,N_21865);
nor U25596 (N_25596,N_21905,N_22723);
nor U25597 (N_25597,N_21086,N_23528);
or U25598 (N_25598,N_21054,N_21868);
and U25599 (N_25599,N_23090,N_22122);
nand U25600 (N_25600,N_22339,N_22594);
and U25601 (N_25601,N_22992,N_21502);
nor U25602 (N_25602,N_21978,N_21280);
nand U25603 (N_25603,N_23273,N_22172);
and U25604 (N_25604,N_22608,N_21841);
and U25605 (N_25605,N_22167,N_21616);
nand U25606 (N_25606,N_22802,N_21095);
xor U25607 (N_25607,N_22219,N_23065);
nand U25608 (N_25608,N_21153,N_21369);
and U25609 (N_25609,N_21828,N_22395);
xor U25610 (N_25610,N_23600,N_23014);
and U25611 (N_25611,N_21204,N_22573);
xnor U25612 (N_25612,N_21752,N_22305);
nand U25613 (N_25613,N_21819,N_21942);
xnor U25614 (N_25614,N_23431,N_22897);
and U25615 (N_25615,N_22901,N_21838);
nor U25616 (N_25616,N_23773,N_21334);
or U25617 (N_25617,N_23438,N_23328);
nor U25618 (N_25618,N_21268,N_22346);
and U25619 (N_25619,N_23569,N_22578);
nor U25620 (N_25620,N_23167,N_21694);
or U25621 (N_25621,N_22776,N_21745);
nor U25622 (N_25622,N_22934,N_22546);
or U25623 (N_25623,N_22727,N_21030);
and U25624 (N_25624,N_21313,N_22697);
and U25625 (N_25625,N_21580,N_22208);
nand U25626 (N_25626,N_23810,N_23586);
and U25627 (N_25627,N_22683,N_23325);
nand U25628 (N_25628,N_21866,N_23700);
xor U25629 (N_25629,N_23609,N_21465);
nor U25630 (N_25630,N_21942,N_23409);
nor U25631 (N_25631,N_23507,N_23479);
and U25632 (N_25632,N_21544,N_22593);
nor U25633 (N_25633,N_23505,N_23619);
nand U25634 (N_25634,N_21535,N_21143);
nand U25635 (N_25635,N_22324,N_21479);
nor U25636 (N_25636,N_23420,N_21676);
nand U25637 (N_25637,N_23115,N_22957);
xor U25638 (N_25638,N_21784,N_22698);
xor U25639 (N_25639,N_21867,N_21272);
and U25640 (N_25640,N_23578,N_23321);
xor U25641 (N_25641,N_23021,N_23409);
xnor U25642 (N_25642,N_23393,N_23413);
and U25643 (N_25643,N_21077,N_23597);
nor U25644 (N_25644,N_22652,N_22830);
xor U25645 (N_25645,N_23271,N_21609);
nand U25646 (N_25646,N_21288,N_21118);
nand U25647 (N_25647,N_22278,N_22759);
nor U25648 (N_25648,N_22246,N_21843);
xor U25649 (N_25649,N_21815,N_21902);
xor U25650 (N_25650,N_23285,N_21279);
nor U25651 (N_25651,N_22212,N_21348);
and U25652 (N_25652,N_22442,N_21623);
nor U25653 (N_25653,N_21166,N_21836);
or U25654 (N_25654,N_22728,N_23380);
nand U25655 (N_25655,N_22871,N_21869);
nor U25656 (N_25656,N_22494,N_22069);
nand U25657 (N_25657,N_21065,N_22835);
and U25658 (N_25658,N_21167,N_23088);
nor U25659 (N_25659,N_22194,N_22404);
xor U25660 (N_25660,N_21417,N_22548);
nor U25661 (N_25661,N_22939,N_22252);
or U25662 (N_25662,N_21919,N_23649);
nand U25663 (N_25663,N_21324,N_23475);
and U25664 (N_25664,N_21800,N_22394);
nor U25665 (N_25665,N_22909,N_21730);
nor U25666 (N_25666,N_22484,N_21395);
xnor U25667 (N_25667,N_23024,N_22665);
xnor U25668 (N_25668,N_21283,N_21531);
and U25669 (N_25669,N_22849,N_23398);
nor U25670 (N_25670,N_22177,N_22160);
xor U25671 (N_25671,N_21528,N_22987);
or U25672 (N_25672,N_23659,N_21486);
nor U25673 (N_25673,N_21867,N_21384);
nand U25674 (N_25674,N_21542,N_21732);
nand U25675 (N_25675,N_23240,N_21667);
and U25676 (N_25676,N_21221,N_22847);
or U25677 (N_25677,N_23600,N_23502);
xor U25678 (N_25678,N_22490,N_23478);
nor U25679 (N_25679,N_21832,N_23077);
xnor U25680 (N_25680,N_22001,N_23198);
or U25681 (N_25681,N_23614,N_22137);
or U25682 (N_25682,N_22722,N_21835);
xnor U25683 (N_25683,N_22367,N_21707);
nor U25684 (N_25684,N_21037,N_22976);
nand U25685 (N_25685,N_22316,N_21520);
nand U25686 (N_25686,N_22488,N_21298);
or U25687 (N_25687,N_23104,N_21305);
and U25688 (N_25688,N_21257,N_22311);
nor U25689 (N_25689,N_21995,N_22253);
and U25690 (N_25690,N_23517,N_21318);
or U25691 (N_25691,N_23535,N_21008);
nand U25692 (N_25692,N_22536,N_21373);
or U25693 (N_25693,N_21163,N_22312);
nand U25694 (N_25694,N_22013,N_21688);
nand U25695 (N_25695,N_22866,N_21695);
or U25696 (N_25696,N_23544,N_22367);
and U25697 (N_25697,N_23245,N_22225);
nand U25698 (N_25698,N_22503,N_22265);
and U25699 (N_25699,N_23225,N_21804);
nor U25700 (N_25700,N_23458,N_22592);
xnor U25701 (N_25701,N_22279,N_21366);
nor U25702 (N_25702,N_23427,N_22455);
xnor U25703 (N_25703,N_21511,N_22397);
xnor U25704 (N_25704,N_21559,N_23550);
and U25705 (N_25705,N_21174,N_23985);
nor U25706 (N_25706,N_21208,N_22495);
nand U25707 (N_25707,N_23323,N_21943);
and U25708 (N_25708,N_22077,N_23156);
nor U25709 (N_25709,N_21471,N_22673);
nor U25710 (N_25710,N_23262,N_21055);
or U25711 (N_25711,N_21261,N_22114);
nor U25712 (N_25712,N_21742,N_21855);
or U25713 (N_25713,N_23170,N_23760);
nor U25714 (N_25714,N_22608,N_23894);
xnor U25715 (N_25715,N_22216,N_22601);
or U25716 (N_25716,N_23207,N_23091);
nor U25717 (N_25717,N_23646,N_21590);
nand U25718 (N_25718,N_22690,N_21204);
or U25719 (N_25719,N_23224,N_21665);
or U25720 (N_25720,N_21608,N_22744);
and U25721 (N_25721,N_22747,N_23979);
or U25722 (N_25722,N_22390,N_21423);
and U25723 (N_25723,N_22006,N_21154);
and U25724 (N_25724,N_22009,N_21891);
nand U25725 (N_25725,N_22347,N_23300);
xnor U25726 (N_25726,N_21433,N_22107);
nand U25727 (N_25727,N_23326,N_21322);
or U25728 (N_25728,N_22150,N_21052);
xnor U25729 (N_25729,N_21276,N_21305);
nor U25730 (N_25730,N_23908,N_23387);
and U25731 (N_25731,N_22740,N_22993);
xor U25732 (N_25732,N_22695,N_21021);
and U25733 (N_25733,N_21514,N_21712);
xnor U25734 (N_25734,N_23813,N_21132);
nor U25735 (N_25735,N_21603,N_23320);
nand U25736 (N_25736,N_21285,N_23279);
xnor U25737 (N_25737,N_22301,N_23408);
nor U25738 (N_25738,N_22344,N_21520);
or U25739 (N_25739,N_21315,N_21427);
and U25740 (N_25740,N_23693,N_23530);
nand U25741 (N_25741,N_21956,N_21988);
xnor U25742 (N_25742,N_22215,N_21314);
and U25743 (N_25743,N_23576,N_23654);
xnor U25744 (N_25744,N_22554,N_21574);
nand U25745 (N_25745,N_23892,N_23206);
nand U25746 (N_25746,N_23144,N_23204);
or U25747 (N_25747,N_22873,N_22721);
or U25748 (N_25748,N_23133,N_21509);
nand U25749 (N_25749,N_22662,N_21360);
nor U25750 (N_25750,N_22293,N_21139);
or U25751 (N_25751,N_23426,N_23352);
or U25752 (N_25752,N_23590,N_23970);
nand U25753 (N_25753,N_22084,N_22287);
nor U25754 (N_25754,N_21060,N_23737);
and U25755 (N_25755,N_23290,N_23238);
xor U25756 (N_25756,N_21649,N_21700);
and U25757 (N_25757,N_21161,N_21780);
nor U25758 (N_25758,N_23602,N_23971);
nand U25759 (N_25759,N_22993,N_21988);
or U25760 (N_25760,N_21681,N_21800);
and U25761 (N_25761,N_23760,N_21770);
xnor U25762 (N_25762,N_21004,N_23455);
xnor U25763 (N_25763,N_23498,N_22698);
and U25764 (N_25764,N_23586,N_22724);
nand U25765 (N_25765,N_21268,N_22076);
or U25766 (N_25766,N_21131,N_21285);
and U25767 (N_25767,N_23230,N_23844);
nand U25768 (N_25768,N_22977,N_22316);
xnor U25769 (N_25769,N_22616,N_21444);
and U25770 (N_25770,N_22429,N_22562);
nand U25771 (N_25771,N_23024,N_22279);
nand U25772 (N_25772,N_22365,N_22741);
nor U25773 (N_25773,N_22343,N_22228);
and U25774 (N_25774,N_21575,N_22184);
and U25775 (N_25775,N_22944,N_21276);
xnor U25776 (N_25776,N_21834,N_23165);
or U25777 (N_25777,N_22517,N_23277);
and U25778 (N_25778,N_22383,N_22013);
nor U25779 (N_25779,N_22605,N_23811);
xnor U25780 (N_25780,N_22669,N_22993);
nand U25781 (N_25781,N_22508,N_22343);
nor U25782 (N_25782,N_23512,N_21630);
nor U25783 (N_25783,N_23811,N_23137);
nand U25784 (N_25784,N_23064,N_23051);
nor U25785 (N_25785,N_21799,N_21424);
xnor U25786 (N_25786,N_23076,N_22191);
xnor U25787 (N_25787,N_22798,N_23221);
nor U25788 (N_25788,N_21950,N_23870);
nand U25789 (N_25789,N_23203,N_22532);
nor U25790 (N_25790,N_21127,N_23264);
xor U25791 (N_25791,N_21193,N_22228);
nor U25792 (N_25792,N_23962,N_21151);
or U25793 (N_25793,N_21501,N_22504);
and U25794 (N_25794,N_23138,N_23080);
nand U25795 (N_25795,N_23167,N_21370);
nor U25796 (N_25796,N_22029,N_21926);
xor U25797 (N_25797,N_23241,N_23826);
nor U25798 (N_25798,N_21545,N_21055);
or U25799 (N_25799,N_22675,N_21615);
and U25800 (N_25800,N_23919,N_22409);
or U25801 (N_25801,N_23705,N_22423);
or U25802 (N_25802,N_21443,N_22048);
nor U25803 (N_25803,N_22331,N_22818);
or U25804 (N_25804,N_21975,N_23572);
nand U25805 (N_25805,N_23820,N_21935);
xor U25806 (N_25806,N_22398,N_23336);
and U25807 (N_25807,N_21585,N_22884);
or U25808 (N_25808,N_22314,N_22598);
or U25809 (N_25809,N_21308,N_21214);
nor U25810 (N_25810,N_22382,N_22918);
xor U25811 (N_25811,N_22161,N_21763);
nor U25812 (N_25812,N_23939,N_21294);
or U25813 (N_25813,N_22422,N_22539);
nor U25814 (N_25814,N_22244,N_21740);
nand U25815 (N_25815,N_23563,N_23782);
xor U25816 (N_25816,N_23481,N_23316);
xnor U25817 (N_25817,N_22268,N_22265);
and U25818 (N_25818,N_23114,N_22642);
nor U25819 (N_25819,N_23865,N_23635);
nand U25820 (N_25820,N_22438,N_21046);
or U25821 (N_25821,N_23791,N_22804);
xor U25822 (N_25822,N_21917,N_21765);
nor U25823 (N_25823,N_21945,N_21244);
and U25824 (N_25824,N_23850,N_23459);
and U25825 (N_25825,N_23272,N_22024);
and U25826 (N_25826,N_21560,N_21185);
or U25827 (N_25827,N_21162,N_21715);
nand U25828 (N_25828,N_22438,N_23980);
nor U25829 (N_25829,N_23505,N_22997);
and U25830 (N_25830,N_22858,N_21527);
xnor U25831 (N_25831,N_21286,N_22423);
and U25832 (N_25832,N_22090,N_21549);
xor U25833 (N_25833,N_23715,N_21179);
nand U25834 (N_25834,N_23278,N_22705);
nor U25835 (N_25835,N_23633,N_23177);
nand U25836 (N_25836,N_23251,N_22067);
or U25837 (N_25837,N_23545,N_23730);
nand U25838 (N_25838,N_23691,N_21647);
nand U25839 (N_25839,N_22798,N_23031);
nor U25840 (N_25840,N_23651,N_21409);
nor U25841 (N_25841,N_23961,N_23995);
nand U25842 (N_25842,N_23702,N_23306);
or U25843 (N_25843,N_21250,N_23049);
or U25844 (N_25844,N_23798,N_21273);
or U25845 (N_25845,N_23122,N_21731);
and U25846 (N_25846,N_22084,N_22281);
and U25847 (N_25847,N_22651,N_22177);
nand U25848 (N_25848,N_22021,N_21238);
and U25849 (N_25849,N_23166,N_22873);
nand U25850 (N_25850,N_22987,N_23816);
and U25851 (N_25851,N_22969,N_21201);
nor U25852 (N_25852,N_23016,N_23123);
xor U25853 (N_25853,N_23570,N_22305);
nor U25854 (N_25854,N_23315,N_23779);
or U25855 (N_25855,N_22574,N_21495);
and U25856 (N_25856,N_23510,N_23239);
and U25857 (N_25857,N_22221,N_21664);
nand U25858 (N_25858,N_22862,N_22104);
and U25859 (N_25859,N_23444,N_23794);
and U25860 (N_25860,N_23822,N_21867);
xnor U25861 (N_25861,N_21511,N_23651);
and U25862 (N_25862,N_22729,N_22440);
and U25863 (N_25863,N_21896,N_21042);
xnor U25864 (N_25864,N_23024,N_23683);
xor U25865 (N_25865,N_23157,N_23748);
and U25866 (N_25866,N_22762,N_21768);
or U25867 (N_25867,N_22217,N_21836);
or U25868 (N_25868,N_22206,N_22184);
and U25869 (N_25869,N_22451,N_21832);
or U25870 (N_25870,N_22367,N_23736);
nand U25871 (N_25871,N_23295,N_21743);
and U25872 (N_25872,N_21788,N_22771);
or U25873 (N_25873,N_23754,N_22508);
and U25874 (N_25874,N_21108,N_23457);
xor U25875 (N_25875,N_23301,N_23902);
nor U25876 (N_25876,N_22712,N_22804);
and U25877 (N_25877,N_21324,N_22047);
or U25878 (N_25878,N_21799,N_22267);
xnor U25879 (N_25879,N_23612,N_22695);
or U25880 (N_25880,N_22987,N_21857);
xnor U25881 (N_25881,N_21388,N_21222);
xor U25882 (N_25882,N_21970,N_23473);
xor U25883 (N_25883,N_23955,N_21289);
and U25884 (N_25884,N_23766,N_22947);
or U25885 (N_25885,N_23012,N_21827);
nand U25886 (N_25886,N_21250,N_22897);
nor U25887 (N_25887,N_23173,N_21484);
nor U25888 (N_25888,N_23024,N_21601);
nand U25889 (N_25889,N_22509,N_23299);
and U25890 (N_25890,N_23486,N_22965);
or U25891 (N_25891,N_21928,N_23200);
nand U25892 (N_25892,N_21793,N_22249);
or U25893 (N_25893,N_21078,N_23686);
xnor U25894 (N_25894,N_21267,N_22526);
nor U25895 (N_25895,N_22417,N_21557);
xor U25896 (N_25896,N_23938,N_22700);
nor U25897 (N_25897,N_23740,N_22064);
and U25898 (N_25898,N_21713,N_21469);
nor U25899 (N_25899,N_23587,N_23911);
and U25900 (N_25900,N_23543,N_23884);
xnor U25901 (N_25901,N_22418,N_22641);
xnor U25902 (N_25902,N_21292,N_21046);
and U25903 (N_25903,N_21440,N_21228);
or U25904 (N_25904,N_23850,N_22897);
xor U25905 (N_25905,N_23374,N_23643);
and U25906 (N_25906,N_22233,N_21254);
nand U25907 (N_25907,N_21618,N_23641);
xor U25908 (N_25908,N_23527,N_21832);
and U25909 (N_25909,N_21820,N_22116);
nand U25910 (N_25910,N_23682,N_22502);
and U25911 (N_25911,N_23707,N_21656);
nand U25912 (N_25912,N_23806,N_23804);
nand U25913 (N_25913,N_22111,N_21831);
nand U25914 (N_25914,N_22754,N_23224);
nand U25915 (N_25915,N_21426,N_23187);
or U25916 (N_25916,N_23035,N_22304);
nand U25917 (N_25917,N_23039,N_23816);
nand U25918 (N_25918,N_23860,N_23039);
xnor U25919 (N_25919,N_22955,N_22518);
nor U25920 (N_25920,N_21741,N_23185);
nand U25921 (N_25921,N_22340,N_21123);
nor U25922 (N_25922,N_21637,N_22098);
xor U25923 (N_25923,N_22906,N_22348);
or U25924 (N_25924,N_22621,N_22311);
nand U25925 (N_25925,N_21750,N_23013);
or U25926 (N_25926,N_21315,N_23825);
xnor U25927 (N_25927,N_21867,N_23000);
xnor U25928 (N_25928,N_21283,N_21364);
and U25929 (N_25929,N_22525,N_22770);
or U25930 (N_25930,N_21644,N_22190);
nor U25931 (N_25931,N_23685,N_22746);
and U25932 (N_25932,N_22481,N_22347);
nand U25933 (N_25933,N_21984,N_22841);
nand U25934 (N_25934,N_21499,N_23746);
xnor U25935 (N_25935,N_22796,N_22656);
and U25936 (N_25936,N_22450,N_23437);
xnor U25937 (N_25937,N_22498,N_21669);
or U25938 (N_25938,N_21106,N_22016);
or U25939 (N_25939,N_23360,N_22647);
and U25940 (N_25940,N_21101,N_23271);
or U25941 (N_25941,N_23052,N_21893);
or U25942 (N_25942,N_22508,N_22588);
nor U25943 (N_25943,N_22745,N_21611);
nand U25944 (N_25944,N_23310,N_21916);
or U25945 (N_25945,N_22200,N_22201);
or U25946 (N_25946,N_21318,N_22439);
and U25947 (N_25947,N_22235,N_21912);
nand U25948 (N_25948,N_23860,N_21075);
and U25949 (N_25949,N_21807,N_21805);
nand U25950 (N_25950,N_21343,N_21709);
nand U25951 (N_25951,N_21984,N_23088);
xnor U25952 (N_25952,N_22139,N_21071);
nor U25953 (N_25953,N_21988,N_21996);
nor U25954 (N_25954,N_23656,N_23379);
xnor U25955 (N_25955,N_23745,N_23516);
and U25956 (N_25956,N_23331,N_21386);
or U25957 (N_25957,N_23640,N_22979);
nand U25958 (N_25958,N_22634,N_23502);
and U25959 (N_25959,N_22940,N_22560);
nand U25960 (N_25960,N_21851,N_22177);
or U25961 (N_25961,N_22995,N_23805);
and U25962 (N_25962,N_22888,N_23011);
nand U25963 (N_25963,N_21997,N_23465);
or U25964 (N_25964,N_21810,N_22226);
nor U25965 (N_25965,N_21350,N_21748);
xnor U25966 (N_25966,N_21177,N_22091);
xor U25967 (N_25967,N_22052,N_23581);
nor U25968 (N_25968,N_21253,N_21283);
and U25969 (N_25969,N_22504,N_23383);
xnor U25970 (N_25970,N_22400,N_21558);
xor U25971 (N_25971,N_21519,N_21042);
or U25972 (N_25972,N_22219,N_22856);
or U25973 (N_25973,N_22443,N_21868);
nor U25974 (N_25974,N_22672,N_23296);
nand U25975 (N_25975,N_21226,N_22602);
or U25976 (N_25976,N_22373,N_21234);
or U25977 (N_25977,N_21971,N_21518);
or U25978 (N_25978,N_23451,N_22727);
nand U25979 (N_25979,N_21458,N_22444);
or U25980 (N_25980,N_23745,N_22401);
or U25981 (N_25981,N_21782,N_22272);
or U25982 (N_25982,N_23943,N_22055);
or U25983 (N_25983,N_23165,N_21014);
and U25984 (N_25984,N_22624,N_23429);
nand U25985 (N_25985,N_22207,N_21081);
or U25986 (N_25986,N_22832,N_23931);
or U25987 (N_25987,N_22093,N_21338);
nand U25988 (N_25988,N_23543,N_22597);
and U25989 (N_25989,N_23065,N_22983);
xor U25990 (N_25990,N_21278,N_21011);
nand U25991 (N_25991,N_23977,N_23991);
nand U25992 (N_25992,N_23508,N_21925);
nand U25993 (N_25993,N_21554,N_23055);
nor U25994 (N_25994,N_21530,N_21140);
xnor U25995 (N_25995,N_22924,N_21056);
xor U25996 (N_25996,N_21582,N_22534);
nor U25997 (N_25997,N_21034,N_23166);
nand U25998 (N_25998,N_23655,N_21527);
or U25999 (N_25999,N_21309,N_22986);
xor U26000 (N_26000,N_23655,N_23660);
or U26001 (N_26001,N_21560,N_21966);
nor U26002 (N_26002,N_21545,N_21482);
and U26003 (N_26003,N_23064,N_23025);
nand U26004 (N_26004,N_22727,N_23555);
nand U26005 (N_26005,N_23551,N_21361);
nand U26006 (N_26006,N_21386,N_22797);
or U26007 (N_26007,N_21126,N_21218);
nand U26008 (N_26008,N_22472,N_23426);
xnor U26009 (N_26009,N_22977,N_22877);
or U26010 (N_26010,N_23536,N_23666);
and U26011 (N_26011,N_21242,N_23075);
nor U26012 (N_26012,N_22476,N_21030);
nand U26013 (N_26013,N_21765,N_21351);
or U26014 (N_26014,N_22818,N_22905);
nor U26015 (N_26015,N_22462,N_23793);
nand U26016 (N_26016,N_21467,N_21061);
and U26017 (N_26017,N_21158,N_21034);
and U26018 (N_26018,N_22261,N_21337);
and U26019 (N_26019,N_23394,N_21834);
nor U26020 (N_26020,N_22984,N_22864);
nand U26021 (N_26021,N_21845,N_21105);
nor U26022 (N_26022,N_21360,N_23783);
nor U26023 (N_26023,N_21024,N_23125);
and U26024 (N_26024,N_21321,N_23467);
or U26025 (N_26025,N_23337,N_23126);
nand U26026 (N_26026,N_22997,N_22053);
and U26027 (N_26027,N_23718,N_21312);
or U26028 (N_26028,N_23434,N_23016);
or U26029 (N_26029,N_23521,N_23977);
and U26030 (N_26030,N_23735,N_22665);
xor U26031 (N_26031,N_22502,N_23924);
and U26032 (N_26032,N_21617,N_22827);
and U26033 (N_26033,N_23053,N_21910);
or U26034 (N_26034,N_21457,N_23484);
nor U26035 (N_26035,N_23186,N_21368);
nor U26036 (N_26036,N_23118,N_21551);
xnor U26037 (N_26037,N_22473,N_22803);
xor U26038 (N_26038,N_22143,N_23512);
or U26039 (N_26039,N_21159,N_23471);
or U26040 (N_26040,N_21725,N_23432);
nand U26041 (N_26041,N_22052,N_23443);
nor U26042 (N_26042,N_22024,N_21131);
nor U26043 (N_26043,N_21234,N_22319);
xnor U26044 (N_26044,N_22443,N_23278);
xor U26045 (N_26045,N_22276,N_23582);
and U26046 (N_26046,N_23106,N_23060);
nand U26047 (N_26047,N_22880,N_23301);
xor U26048 (N_26048,N_23323,N_23666);
and U26049 (N_26049,N_23790,N_21550);
xor U26050 (N_26050,N_21600,N_23083);
or U26051 (N_26051,N_22136,N_22005);
xnor U26052 (N_26052,N_21567,N_22976);
nand U26053 (N_26053,N_22989,N_22349);
nand U26054 (N_26054,N_22359,N_21156);
xnor U26055 (N_26055,N_22948,N_22716);
and U26056 (N_26056,N_23075,N_22345);
xnor U26057 (N_26057,N_23945,N_22669);
xnor U26058 (N_26058,N_23324,N_21565);
or U26059 (N_26059,N_21798,N_21135);
and U26060 (N_26060,N_23956,N_22470);
xor U26061 (N_26061,N_21693,N_23539);
and U26062 (N_26062,N_21334,N_21766);
nor U26063 (N_26063,N_22996,N_21288);
nand U26064 (N_26064,N_21358,N_21679);
or U26065 (N_26065,N_23312,N_22814);
nor U26066 (N_26066,N_21460,N_23672);
xnor U26067 (N_26067,N_21914,N_21205);
nand U26068 (N_26068,N_22493,N_21477);
nor U26069 (N_26069,N_21035,N_21922);
xor U26070 (N_26070,N_23059,N_23615);
nor U26071 (N_26071,N_21304,N_21228);
nor U26072 (N_26072,N_23159,N_23484);
or U26073 (N_26073,N_23246,N_22530);
nor U26074 (N_26074,N_23440,N_22453);
and U26075 (N_26075,N_21143,N_21654);
and U26076 (N_26076,N_22233,N_21456);
xnor U26077 (N_26077,N_23612,N_22724);
nor U26078 (N_26078,N_23452,N_21479);
or U26079 (N_26079,N_21539,N_23148);
nand U26080 (N_26080,N_22699,N_22467);
or U26081 (N_26081,N_21531,N_23297);
nor U26082 (N_26082,N_21910,N_22727);
and U26083 (N_26083,N_23737,N_21481);
nand U26084 (N_26084,N_23260,N_21876);
and U26085 (N_26085,N_23191,N_22988);
nor U26086 (N_26086,N_22209,N_22114);
nor U26087 (N_26087,N_21307,N_21193);
or U26088 (N_26088,N_21817,N_23575);
or U26089 (N_26089,N_23868,N_22052);
nor U26090 (N_26090,N_22978,N_21720);
nor U26091 (N_26091,N_23731,N_22648);
or U26092 (N_26092,N_22906,N_21687);
nand U26093 (N_26093,N_21542,N_22891);
or U26094 (N_26094,N_22334,N_23308);
xor U26095 (N_26095,N_22097,N_22958);
nand U26096 (N_26096,N_22635,N_23933);
and U26097 (N_26097,N_22108,N_22087);
or U26098 (N_26098,N_23065,N_23575);
nand U26099 (N_26099,N_23140,N_21778);
xor U26100 (N_26100,N_21824,N_21940);
nand U26101 (N_26101,N_22505,N_22213);
or U26102 (N_26102,N_22024,N_21261);
nand U26103 (N_26103,N_22383,N_22158);
or U26104 (N_26104,N_22733,N_21845);
or U26105 (N_26105,N_23998,N_23953);
xnor U26106 (N_26106,N_21781,N_21282);
or U26107 (N_26107,N_21687,N_23957);
xnor U26108 (N_26108,N_23202,N_23782);
and U26109 (N_26109,N_22305,N_23041);
nor U26110 (N_26110,N_21233,N_23546);
nor U26111 (N_26111,N_21664,N_21385);
or U26112 (N_26112,N_23187,N_21277);
or U26113 (N_26113,N_21895,N_23101);
xor U26114 (N_26114,N_21519,N_22658);
xnor U26115 (N_26115,N_22133,N_21688);
nor U26116 (N_26116,N_23043,N_23189);
nand U26117 (N_26117,N_22593,N_23913);
and U26118 (N_26118,N_23746,N_21892);
xnor U26119 (N_26119,N_21687,N_23515);
or U26120 (N_26120,N_22353,N_22802);
nor U26121 (N_26121,N_22276,N_23431);
nand U26122 (N_26122,N_23117,N_22381);
and U26123 (N_26123,N_22965,N_22962);
or U26124 (N_26124,N_22957,N_21407);
or U26125 (N_26125,N_22715,N_22967);
xnor U26126 (N_26126,N_23735,N_23554);
and U26127 (N_26127,N_22497,N_21362);
or U26128 (N_26128,N_21108,N_23598);
nand U26129 (N_26129,N_21734,N_22756);
and U26130 (N_26130,N_21027,N_23279);
nand U26131 (N_26131,N_21302,N_22522);
or U26132 (N_26132,N_21611,N_21050);
or U26133 (N_26133,N_22855,N_21050);
and U26134 (N_26134,N_22724,N_21457);
and U26135 (N_26135,N_21811,N_21614);
nand U26136 (N_26136,N_22528,N_21061);
xnor U26137 (N_26137,N_21357,N_23438);
or U26138 (N_26138,N_22174,N_23967);
nand U26139 (N_26139,N_21987,N_21264);
nand U26140 (N_26140,N_21474,N_23937);
or U26141 (N_26141,N_23414,N_22683);
nand U26142 (N_26142,N_21346,N_23833);
nand U26143 (N_26143,N_22809,N_22611);
nand U26144 (N_26144,N_21079,N_21630);
or U26145 (N_26145,N_22579,N_21727);
and U26146 (N_26146,N_22043,N_21383);
nor U26147 (N_26147,N_21452,N_22628);
nand U26148 (N_26148,N_22624,N_21609);
nand U26149 (N_26149,N_23911,N_23009);
xnor U26150 (N_26150,N_21017,N_23487);
or U26151 (N_26151,N_21897,N_22457);
nand U26152 (N_26152,N_22738,N_21184);
or U26153 (N_26153,N_21093,N_23633);
nand U26154 (N_26154,N_23045,N_23030);
or U26155 (N_26155,N_21959,N_22955);
and U26156 (N_26156,N_22870,N_21389);
nand U26157 (N_26157,N_23371,N_23375);
or U26158 (N_26158,N_23149,N_21011);
nor U26159 (N_26159,N_21673,N_23768);
nor U26160 (N_26160,N_21580,N_23733);
and U26161 (N_26161,N_23340,N_22919);
and U26162 (N_26162,N_22174,N_23206);
and U26163 (N_26163,N_22916,N_22734);
nand U26164 (N_26164,N_23569,N_23711);
xor U26165 (N_26165,N_23195,N_23717);
or U26166 (N_26166,N_23915,N_23226);
nor U26167 (N_26167,N_22529,N_21657);
or U26168 (N_26168,N_21171,N_22945);
or U26169 (N_26169,N_21831,N_21940);
and U26170 (N_26170,N_21850,N_21378);
xnor U26171 (N_26171,N_23473,N_22688);
nand U26172 (N_26172,N_21641,N_23091);
xnor U26173 (N_26173,N_22494,N_23602);
nor U26174 (N_26174,N_23034,N_23317);
nor U26175 (N_26175,N_23907,N_21406);
nor U26176 (N_26176,N_23404,N_22493);
nor U26177 (N_26177,N_22873,N_23314);
nand U26178 (N_26178,N_21863,N_23218);
and U26179 (N_26179,N_23110,N_23753);
nand U26180 (N_26180,N_21061,N_22871);
xor U26181 (N_26181,N_21950,N_22102);
nor U26182 (N_26182,N_21358,N_22312);
nor U26183 (N_26183,N_21307,N_22551);
xor U26184 (N_26184,N_21900,N_23019);
or U26185 (N_26185,N_23759,N_21717);
and U26186 (N_26186,N_21421,N_23967);
nand U26187 (N_26187,N_22730,N_21489);
nor U26188 (N_26188,N_21588,N_22107);
xnor U26189 (N_26189,N_22028,N_22246);
xnor U26190 (N_26190,N_21044,N_22017);
or U26191 (N_26191,N_23034,N_23841);
or U26192 (N_26192,N_23093,N_21881);
or U26193 (N_26193,N_21499,N_23723);
and U26194 (N_26194,N_22630,N_23234);
or U26195 (N_26195,N_23342,N_22767);
or U26196 (N_26196,N_23152,N_22886);
nand U26197 (N_26197,N_23903,N_21199);
and U26198 (N_26198,N_23729,N_21069);
nand U26199 (N_26199,N_23728,N_23833);
xnor U26200 (N_26200,N_23237,N_21315);
and U26201 (N_26201,N_23060,N_23546);
and U26202 (N_26202,N_23343,N_21384);
nor U26203 (N_26203,N_22678,N_22417);
or U26204 (N_26204,N_22765,N_21761);
nand U26205 (N_26205,N_21969,N_22032);
xor U26206 (N_26206,N_21041,N_21247);
nand U26207 (N_26207,N_21676,N_22012);
nor U26208 (N_26208,N_23556,N_21121);
nor U26209 (N_26209,N_23413,N_21928);
and U26210 (N_26210,N_23258,N_21640);
nor U26211 (N_26211,N_23784,N_21613);
or U26212 (N_26212,N_22612,N_22255);
xor U26213 (N_26213,N_23268,N_21842);
and U26214 (N_26214,N_23602,N_22234);
nor U26215 (N_26215,N_23730,N_21310);
or U26216 (N_26216,N_22498,N_21650);
xor U26217 (N_26217,N_22376,N_21412);
or U26218 (N_26218,N_23941,N_23743);
nand U26219 (N_26219,N_23057,N_23456);
or U26220 (N_26220,N_23492,N_22435);
nor U26221 (N_26221,N_23755,N_21379);
nor U26222 (N_26222,N_21346,N_21485);
nand U26223 (N_26223,N_22013,N_23025);
xor U26224 (N_26224,N_23757,N_22371);
nor U26225 (N_26225,N_23387,N_22871);
nand U26226 (N_26226,N_21447,N_23612);
nor U26227 (N_26227,N_21635,N_21665);
nor U26228 (N_26228,N_22206,N_22661);
and U26229 (N_26229,N_21800,N_22573);
xor U26230 (N_26230,N_21276,N_21684);
and U26231 (N_26231,N_21999,N_23388);
nand U26232 (N_26232,N_23491,N_22229);
xnor U26233 (N_26233,N_22833,N_23893);
or U26234 (N_26234,N_21661,N_22050);
nand U26235 (N_26235,N_23313,N_21748);
or U26236 (N_26236,N_23410,N_21709);
xnor U26237 (N_26237,N_21605,N_22299);
nor U26238 (N_26238,N_21389,N_23728);
and U26239 (N_26239,N_21805,N_22368);
xor U26240 (N_26240,N_22573,N_21697);
nor U26241 (N_26241,N_21226,N_21380);
nand U26242 (N_26242,N_22216,N_23941);
xnor U26243 (N_26243,N_22384,N_21587);
xnor U26244 (N_26244,N_21242,N_21746);
xnor U26245 (N_26245,N_22025,N_21609);
nand U26246 (N_26246,N_22048,N_22915);
xor U26247 (N_26247,N_21707,N_21921);
nand U26248 (N_26248,N_22209,N_21863);
xor U26249 (N_26249,N_21645,N_21768);
and U26250 (N_26250,N_22643,N_22985);
or U26251 (N_26251,N_22301,N_23597);
or U26252 (N_26252,N_23251,N_23424);
xor U26253 (N_26253,N_21927,N_23286);
or U26254 (N_26254,N_22433,N_23684);
nand U26255 (N_26255,N_23017,N_21614);
xnor U26256 (N_26256,N_21577,N_23539);
nor U26257 (N_26257,N_22080,N_22879);
or U26258 (N_26258,N_21644,N_23318);
and U26259 (N_26259,N_23069,N_21765);
and U26260 (N_26260,N_23678,N_22156);
or U26261 (N_26261,N_23424,N_22471);
or U26262 (N_26262,N_22788,N_21542);
nor U26263 (N_26263,N_22226,N_21209);
xor U26264 (N_26264,N_23947,N_22518);
nand U26265 (N_26265,N_21753,N_23793);
and U26266 (N_26266,N_22676,N_23954);
nor U26267 (N_26267,N_21851,N_22841);
or U26268 (N_26268,N_23848,N_22493);
and U26269 (N_26269,N_22615,N_21965);
nand U26270 (N_26270,N_22536,N_21218);
xnor U26271 (N_26271,N_21423,N_23390);
and U26272 (N_26272,N_23454,N_21399);
and U26273 (N_26273,N_22805,N_22465);
or U26274 (N_26274,N_22470,N_22001);
xor U26275 (N_26275,N_22939,N_21122);
or U26276 (N_26276,N_23857,N_23386);
xor U26277 (N_26277,N_22245,N_21993);
or U26278 (N_26278,N_21133,N_21617);
nand U26279 (N_26279,N_22217,N_21923);
nand U26280 (N_26280,N_21743,N_22194);
or U26281 (N_26281,N_22084,N_22080);
or U26282 (N_26282,N_21744,N_23447);
nand U26283 (N_26283,N_21632,N_21299);
nor U26284 (N_26284,N_21534,N_22170);
xor U26285 (N_26285,N_21767,N_21074);
nor U26286 (N_26286,N_21452,N_21823);
xnor U26287 (N_26287,N_21005,N_22496);
xor U26288 (N_26288,N_23232,N_21863);
or U26289 (N_26289,N_22491,N_22802);
and U26290 (N_26290,N_23035,N_23315);
nand U26291 (N_26291,N_23173,N_22986);
nand U26292 (N_26292,N_22928,N_23749);
nand U26293 (N_26293,N_21340,N_22453);
nand U26294 (N_26294,N_22667,N_21383);
nand U26295 (N_26295,N_21931,N_23498);
xnor U26296 (N_26296,N_21862,N_23916);
xor U26297 (N_26297,N_21168,N_23152);
xnor U26298 (N_26298,N_21248,N_22186);
xnor U26299 (N_26299,N_22321,N_23217);
and U26300 (N_26300,N_23830,N_22703);
nand U26301 (N_26301,N_22102,N_22611);
or U26302 (N_26302,N_22781,N_23283);
xor U26303 (N_26303,N_23838,N_21111);
nor U26304 (N_26304,N_23289,N_22008);
nor U26305 (N_26305,N_22186,N_21472);
nand U26306 (N_26306,N_21296,N_23690);
xor U26307 (N_26307,N_23822,N_22428);
or U26308 (N_26308,N_22932,N_21001);
and U26309 (N_26309,N_21253,N_21379);
and U26310 (N_26310,N_22136,N_22222);
and U26311 (N_26311,N_21402,N_21287);
xor U26312 (N_26312,N_21916,N_23398);
nand U26313 (N_26313,N_22538,N_22371);
xor U26314 (N_26314,N_23102,N_22130);
or U26315 (N_26315,N_21708,N_22076);
or U26316 (N_26316,N_22127,N_22402);
and U26317 (N_26317,N_22489,N_22588);
and U26318 (N_26318,N_21236,N_22553);
or U26319 (N_26319,N_21762,N_22998);
and U26320 (N_26320,N_23745,N_23873);
nor U26321 (N_26321,N_22790,N_23187);
nor U26322 (N_26322,N_21562,N_23335);
and U26323 (N_26323,N_23494,N_23388);
xor U26324 (N_26324,N_21855,N_22418);
nor U26325 (N_26325,N_21393,N_23987);
or U26326 (N_26326,N_21577,N_21220);
nand U26327 (N_26327,N_23469,N_22143);
and U26328 (N_26328,N_21401,N_21425);
nand U26329 (N_26329,N_21664,N_22671);
nor U26330 (N_26330,N_23417,N_22447);
or U26331 (N_26331,N_21516,N_21614);
nand U26332 (N_26332,N_22351,N_22419);
xnor U26333 (N_26333,N_23513,N_21254);
and U26334 (N_26334,N_21802,N_23328);
xnor U26335 (N_26335,N_21703,N_23557);
xnor U26336 (N_26336,N_22098,N_23895);
nand U26337 (N_26337,N_23591,N_22367);
and U26338 (N_26338,N_23633,N_22454);
xor U26339 (N_26339,N_22695,N_23473);
nor U26340 (N_26340,N_21445,N_23702);
or U26341 (N_26341,N_21563,N_21224);
nor U26342 (N_26342,N_22458,N_23947);
and U26343 (N_26343,N_21876,N_23806);
nor U26344 (N_26344,N_23867,N_22635);
nand U26345 (N_26345,N_21118,N_22534);
nor U26346 (N_26346,N_22117,N_22823);
nand U26347 (N_26347,N_21635,N_21821);
and U26348 (N_26348,N_22825,N_22360);
and U26349 (N_26349,N_23510,N_23262);
nand U26350 (N_26350,N_21124,N_22053);
xor U26351 (N_26351,N_23347,N_21602);
or U26352 (N_26352,N_22298,N_23072);
nor U26353 (N_26353,N_21659,N_22959);
xnor U26354 (N_26354,N_23723,N_23503);
or U26355 (N_26355,N_21505,N_22318);
or U26356 (N_26356,N_23839,N_22137);
nor U26357 (N_26357,N_21228,N_21839);
xnor U26358 (N_26358,N_22733,N_22082);
nor U26359 (N_26359,N_23800,N_22341);
or U26360 (N_26360,N_23013,N_23129);
nor U26361 (N_26361,N_23685,N_23935);
nor U26362 (N_26362,N_21912,N_23913);
nand U26363 (N_26363,N_23284,N_23099);
nor U26364 (N_26364,N_22684,N_22803);
and U26365 (N_26365,N_21994,N_23923);
nand U26366 (N_26366,N_21314,N_21849);
or U26367 (N_26367,N_21920,N_23348);
nor U26368 (N_26368,N_23532,N_23625);
and U26369 (N_26369,N_21769,N_23858);
or U26370 (N_26370,N_22638,N_23064);
xnor U26371 (N_26371,N_23730,N_22341);
and U26372 (N_26372,N_23165,N_23410);
nor U26373 (N_26373,N_21354,N_22081);
nand U26374 (N_26374,N_23463,N_22668);
xnor U26375 (N_26375,N_23479,N_21495);
nor U26376 (N_26376,N_23972,N_21060);
or U26377 (N_26377,N_22363,N_22935);
xnor U26378 (N_26378,N_21778,N_21072);
xnor U26379 (N_26379,N_22363,N_23926);
and U26380 (N_26380,N_23173,N_21609);
nand U26381 (N_26381,N_22635,N_22170);
and U26382 (N_26382,N_22582,N_21753);
nand U26383 (N_26383,N_22603,N_21452);
and U26384 (N_26384,N_23835,N_21392);
or U26385 (N_26385,N_23115,N_21633);
nand U26386 (N_26386,N_23843,N_21977);
or U26387 (N_26387,N_21512,N_22216);
or U26388 (N_26388,N_21602,N_21184);
or U26389 (N_26389,N_23637,N_21732);
xor U26390 (N_26390,N_22067,N_22778);
nor U26391 (N_26391,N_22351,N_21557);
nand U26392 (N_26392,N_21095,N_22795);
nand U26393 (N_26393,N_21527,N_23668);
and U26394 (N_26394,N_22587,N_21148);
and U26395 (N_26395,N_23528,N_22518);
xnor U26396 (N_26396,N_21834,N_23492);
nand U26397 (N_26397,N_21967,N_23253);
and U26398 (N_26398,N_21849,N_23649);
nor U26399 (N_26399,N_23740,N_23607);
or U26400 (N_26400,N_23828,N_22244);
nor U26401 (N_26401,N_23441,N_22133);
and U26402 (N_26402,N_21799,N_23098);
or U26403 (N_26403,N_23812,N_21427);
xor U26404 (N_26404,N_22104,N_22450);
nand U26405 (N_26405,N_22720,N_22055);
and U26406 (N_26406,N_22909,N_22326);
nand U26407 (N_26407,N_22601,N_21468);
or U26408 (N_26408,N_23340,N_22020);
nand U26409 (N_26409,N_22254,N_22131);
or U26410 (N_26410,N_22375,N_22163);
or U26411 (N_26411,N_23043,N_22974);
or U26412 (N_26412,N_23683,N_23764);
xor U26413 (N_26413,N_22750,N_23060);
or U26414 (N_26414,N_22071,N_22829);
and U26415 (N_26415,N_22766,N_22367);
nand U26416 (N_26416,N_21656,N_22789);
nand U26417 (N_26417,N_23070,N_21354);
nor U26418 (N_26418,N_23008,N_21199);
nor U26419 (N_26419,N_22307,N_22925);
or U26420 (N_26420,N_21027,N_23354);
nor U26421 (N_26421,N_23158,N_22295);
or U26422 (N_26422,N_22030,N_23417);
or U26423 (N_26423,N_23544,N_23119);
and U26424 (N_26424,N_21473,N_23104);
xnor U26425 (N_26425,N_22876,N_21278);
nand U26426 (N_26426,N_23716,N_21031);
xnor U26427 (N_26427,N_21637,N_21036);
xor U26428 (N_26428,N_21403,N_23141);
or U26429 (N_26429,N_23313,N_22609);
or U26430 (N_26430,N_23442,N_22509);
xor U26431 (N_26431,N_21410,N_23726);
or U26432 (N_26432,N_23774,N_22383);
nor U26433 (N_26433,N_23429,N_23444);
nand U26434 (N_26434,N_21958,N_23755);
nand U26435 (N_26435,N_21685,N_22574);
xor U26436 (N_26436,N_21729,N_23024);
and U26437 (N_26437,N_21335,N_23014);
xnor U26438 (N_26438,N_21031,N_22076);
nand U26439 (N_26439,N_21985,N_21755);
nand U26440 (N_26440,N_22654,N_21813);
and U26441 (N_26441,N_22302,N_21776);
or U26442 (N_26442,N_22464,N_23521);
nor U26443 (N_26443,N_23230,N_21889);
nor U26444 (N_26444,N_21802,N_23389);
xor U26445 (N_26445,N_23391,N_23745);
or U26446 (N_26446,N_23242,N_22246);
xor U26447 (N_26447,N_21889,N_23929);
nor U26448 (N_26448,N_23076,N_23992);
nor U26449 (N_26449,N_22274,N_21918);
nand U26450 (N_26450,N_23228,N_22165);
nand U26451 (N_26451,N_22504,N_22520);
or U26452 (N_26452,N_23907,N_22342);
or U26453 (N_26453,N_22254,N_21878);
nor U26454 (N_26454,N_22676,N_21933);
xnor U26455 (N_26455,N_23681,N_23682);
nand U26456 (N_26456,N_22874,N_22656);
xnor U26457 (N_26457,N_21822,N_23420);
xor U26458 (N_26458,N_23101,N_22935);
nor U26459 (N_26459,N_22585,N_23500);
nor U26460 (N_26460,N_23711,N_22901);
or U26461 (N_26461,N_23224,N_22765);
nand U26462 (N_26462,N_21135,N_22537);
nor U26463 (N_26463,N_21842,N_23703);
or U26464 (N_26464,N_21957,N_22654);
nor U26465 (N_26465,N_22599,N_22544);
xnor U26466 (N_26466,N_23233,N_23620);
xnor U26467 (N_26467,N_22178,N_23537);
nand U26468 (N_26468,N_21055,N_23063);
nor U26469 (N_26469,N_22356,N_21278);
nand U26470 (N_26470,N_23593,N_22416);
and U26471 (N_26471,N_23018,N_21660);
and U26472 (N_26472,N_22290,N_21728);
nand U26473 (N_26473,N_21006,N_21501);
nand U26474 (N_26474,N_23729,N_23494);
nand U26475 (N_26475,N_22450,N_23378);
nor U26476 (N_26476,N_23690,N_22613);
or U26477 (N_26477,N_23615,N_23790);
or U26478 (N_26478,N_21815,N_22769);
nand U26479 (N_26479,N_21221,N_23251);
nand U26480 (N_26480,N_23551,N_23123);
xnor U26481 (N_26481,N_23393,N_21059);
nor U26482 (N_26482,N_23139,N_23710);
or U26483 (N_26483,N_23293,N_22883);
nor U26484 (N_26484,N_21102,N_23177);
nand U26485 (N_26485,N_21538,N_22352);
nand U26486 (N_26486,N_23625,N_21055);
and U26487 (N_26487,N_22665,N_21671);
nor U26488 (N_26488,N_22692,N_21487);
nor U26489 (N_26489,N_21352,N_23028);
and U26490 (N_26490,N_22055,N_21097);
and U26491 (N_26491,N_23801,N_21265);
or U26492 (N_26492,N_22549,N_21291);
nor U26493 (N_26493,N_22717,N_21155);
or U26494 (N_26494,N_22240,N_21357);
and U26495 (N_26495,N_22755,N_21601);
nand U26496 (N_26496,N_22886,N_23465);
nand U26497 (N_26497,N_22116,N_22710);
and U26498 (N_26498,N_23158,N_23462);
nand U26499 (N_26499,N_23850,N_21387);
nor U26500 (N_26500,N_21718,N_21563);
xor U26501 (N_26501,N_22656,N_23065);
and U26502 (N_26502,N_23505,N_22935);
nand U26503 (N_26503,N_23355,N_22497);
nor U26504 (N_26504,N_23010,N_21939);
or U26505 (N_26505,N_22743,N_21946);
and U26506 (N_26506,N_23209,N_21868);
xnor U26507 (N_26507,N_21363,N_23776);
or U26508 (N_26508,N_21777,N_21118);
xnor U26509 (N_26509,N_22136,N_23770);
or U26510 (N_26510,N_23073,N_22826);
nand U26511 (N_26511,N_23546,N_22828);
nand U26512 (N_26512,N_23461,N_22112);
and U26513 (N_26513,N_23587,N_22046);
nor U26514 (N_26514,N_23522,N_22783);
and U26515 (N_26515,N_23165,N_22175);
nand U26516 (N_26516,N_23071,N_22613);
or U26517 (N_26517,N_21836,N_23984);
nor U26518 (N_26518,N_21238,N_22996);
nor U26519 (N_26519,N_23926,N_21574);
and U26520 (N_26520,N_21689,N_23711);
and U26521 (N_26521,N_22403,N_21284);
or U26522 (N_26522,N_21484,N_21810);
or U26523 (N_26523,N_22571,N_22114);
xor U26524 (N_26524,N_21175,N_22693);
or U26525 (N_26525,N_23804,N_21367);
nand U26526 (N_26526,N_23276,N_23377);
and U26527 (N_26527,N_22563,N_21084);
and U26528 (N_26528,N_22698,N_21689);
nand U26529 (N_26529,N_22851,N_22269);
xnor U26530 (N_26530,N_21516,N_23758);
or U26531 (N_26531,N_21289,N_22527);
or U26532 (N_26532,N_22149,N_23734);
xor U26533 (N_26533,N_21897,N_22816);
nor U26534 (N_26534,N_21890,N_21929);
nand U26535 (N_26535,N_22653,N_21829);
xnor U26536 (N_26536,N_22153,N_23862);
and U26537 (N_26537,N_22154,N_23659);
xor U26538 (N_26538,N_23662,N_21941);
and U26539 (N_26539,N_21040,N_22747);
nand U26540 (N_26540,N_22826,N_22078);
and U26541 (N_26541,N_21101,N_22280);
xor U26542 (N_26542,N_23665,N_23815);
and U26543 (N_26543,N_21111,N_21553);
or U26544 (N_26544,N_23541,N_21535);
xor U26545 (N_26545,N_22566,N_23423);
or U26546 (N_26546,N_21728,N_21443);
nor U26547 (N_26547,N_23873,N_22202);
or U26548 (N_26548,N_22228,N_21293);
and U26549 (N_26549,N_22738,N_23821);
xor U26550 (N_26550,N_23622,N_22446);
nor U26551 (N_26551,N_23858,N_21964);
nand U26552 (N_26552,N_21030,N_21068);
or U26553 (N_26553,N_23249,N_22416);
xnor U26554 (N_26554,N_22783,N_21572);
xor U26555 (N_26555,N_23508,N_21092);
nand U26556 (N_26556,N_23079,N_21555);
or U26557 (N_26557,N_22504,N_21368);
xor U26558 (N_26558,N_21625,N_23817);
xor U26559 (N_26559,N_21332,N_22626);
or U26560 (N_26560,N_21120,N_23056);
xnor U26561 (N_26561,N_22573,N_22257);
nor U26562 (N_26562,N_22475,N_21233);
nor U26563 (N_26563,N_23176,N_22787);
or U26564 (N_26564,N_21564,N_21409);
and U26565 (N_26565,N_21751,N_21264);
or U26566 (N_26566,N_23999,N_21379);
or U26567 (N_26567,N_22512,N_23618);
and U26568 (N_26568,N_21951,N_21562);
xnor U26569 (N_26569,N_21865,N_21247);
nor U26570 (N_26570,N_23649,N_22392);
nor U26571 (N_26571,N_21597,N_21695);
xor U26572 (N_26572,N_23454,N_21027);
or U26573 (N_26573,N_23381,N_23640);
nand U26574 (N_26574,N_22241,N_21830);
xnor U26575 (N_26575,N_22185,N_21106);
and U26576 (N_26576,N_21884,N_22953);
and U26577 (N_26577,N_21287,N_23246);
or U26578 (N_26578,N_21113,N_22552);
nand U26579 (N_26579,N_22465,N_21118);
xor U26580 (N_26580,N_22011,N_22304);
nor U26581 (N_26581,N_23635,N_23368);
nor U26582 (N_26582,N_22172,N_22544);
and U26583 (N_26583,N_23095,N_21120);
or U26584 (N_26584,N_23012,N_23970);
xor U26585 (N_26585,N_23048,N_23648);
xor U26586 (N_26586,N_23633,N_23001);
xnor U26587 (N_26587,N_23537,N_23390);
nand U26588 (N_26588,N_22577,N_22298);
and U26589 (N_26589,N_21031,N_23127);
or U26590 (N_26590,N_21701,N_22434);
nand U26591 (N_26591,N_21556,N_21150);
xnor U26592 (N_26592,N_23248,N_22386);
nor U26593 (N_26593,N_21947,N_23951);
xnor U26594 (N_26594,N_23832,N_22000);
nor U26595 (N_26595,N_21959,N_21322);
or U26596 (N_26596,N_22344,N_23662);
or U26597 (N_26597,N_21812,N_21159);
xor U26598 (N_26598,N_21048,N_22748);
and U26599 (N_26599,N_23222,N_23937);
and U26600 (N_26600,N_21105,N_21165);
xor U26601 (N_26601,N_22460,N_23058);
nand U26602 (N_26602,N_23906,N_22138);
and U26603 (N_26603,N_23035,N_21721);
or U26604 (N_26604,N_21894,N_21589);
nand U26605 (N_26605,N_23919,N_23897);
nand U26606 (N_26606,N_21513,N_23304);
or U26607 (N_26607,N_21569,N_21806);
or U26608 (N_26608,N_22179,N_22905);
xnor U26609 (N_26609,N_22498,N_22528);
or U26610 (N_26610,N_22054,N_22963);
xor U26611 (N_26611,N_23586,N_22729);
nand U26612 (N_26612,N_22346,N_22986);
nand U26613 (N_26613,N_21203,N_22310);
nor U26614 (N_26614,N_22458,N_21589);
or U26615 (N_26615,N_23615,N_22351);
nor U26616 (N_26616,N_22135,N_23585);
nand U26617 (N_26617,N_22088,N_23356);
or U26618 (N_26618,N_22377,N_21257);
and U26619 (N_26619,N_21351,N_21912);
xor U26620 (N_26620,N_23493,N_23036);
and U26621 (N_26621,N_21807,N_21997);
nor U26622 (N_26622,N_22850,N_21577);
and U26623 (N_26623,N_22617,N_21331);
and U26624 (N_26624,N_21198,N_23041);
or U26625 (N_26625,N_21534,N_21314);
nor U26626 (N_26626,N_23237,N_22997);
nor U26627 (N_26627,N_23043,N_23180);
nand U26628 (N_26628,N_22887,N_22508);
xor U26629 (N_26629,N_23885,N_22383);
nand U26630 (N_26630,N_22937,N_23461);
and U26631 (N_26631,N_21645,N_22876);
nor U26632 (N_26632,N_22442,N_23651);
nand U26633 (N_26633,N_21775,N_22209);
nor U26634 (N_26634,N_23910,N_23258);
nand U26635 (N_26635,N_22328,N_23474);
and U26636 (N_26636,N_22890,N_22640);
nor U26637 (N_26637,N_21530,N_22752);
xor U26638 (N_26638,N_22867,N_23601);
nand U26639 (N_26639,N_23261,N_21014);
and U26640 (N_26640,N_22747,N_22637);
or U26641 (N_26641,N_21131,N_22558);
xnor U26642 (N_26642,N_22087,N_23136);
and U26643 (N_26643,N_23936,N_21014);
and U26644 (N_26644,N_22217,N_21862);
or U26645 (N_26645,N_23065,N_23898);
nand U26646 (N_26646,N_23684,N_21619);
and U26647 (N_26647,N_22954,N_22654);
or U26648 (N_26648,N_23152,N_22364);
nand U26649 (N_26649,N_21586,N_23505);
xnor U26650 (N_26650,N_23435,N_23483);
nor U26651 (N_26651,N_21011,N_21950);
nor U26652 (N_26652,N_22121,N_21359);
or U26653 (N_26653,N_23692,N_22457);
xor U26654 (N_26654,N_22523,N_21773);
nand U26655 (N_26655,N_23058,N_21287);
xor U26656 (N_26656,N_22793,N_22264);
or U26657 (N_26657,N_22401,N_22718);
xor U26658 (N_26658,N_23913,N_22652);
xor U26659 (N_26659,N_23062,N_21263);
nand U26660 (N_26660,N_22399,N_22332);
nor U26661 (N_26661,N_22268,N_23561);
or U26662 (N_26662,N_21559,N_21262);
or U26663 (N_26663,N_22712,N_21292);
and U26664 (N_26664,N_23478,N_23160);
and U26665 (N_26665,N_23775,N_22753);
and U26666 (N_26666,N_22674,N_21581);
nor U26667 (N_26667,N_23709,N_22014);
or U26668 (N_26668,N_21548,N_22022);
and U26669 (N_26669,N_21376,N_22424);
nand U26670 (N_26670,N_23789,N_23670);
xor U26671 (N_26671,N_23008,N_23235);
and U26672 (N_26672,N_21798,N_21822);
and U26673 (N_26673,N_23189,N_21583);
nand U26674 (N_26674,N_21675,N_21537);
nor U26675 (N_26675,N_23523,N_22688);
nor U26676 (N_26676,N_22284,N_23011);
and U26677 (N_26677,N_23220,N_21225);
and U26678 (N_26678,N_23901,N_22294);
nand U26679 (N_26679,N_23245,N_23278);
nor U26680 (N_26680,N_23162,N_21056);
xnor U26681 (N_26681,N_22872,N_21770);
and U26682 (N_26682,N_21304,N_22496);
and U26683 (N_26683,N_22374,N_22986);
nor U26684 (N_26684,N_21367,N_21062);
nor U26685 (N_26685,N_21297,N_21843);
or U26686 (N_26686,N_21100,N_22568);
and U26687 (N_26687,N_21482,N_22091);
and U26688 (N_26688,N_21626,N_23319);
and U26689 (N_26689,N_23244,N_22212);
xnor U26690 (N_26690,N_23145,N_23650);
and U26691 (N_26691,N_21729,N_23345);
and U26692 (N_26692,N_23344,N_23374);
xor U26693 (N_26693,N_22726,N_21325);
or U26694 (N_26694,N_21327,N_21221);
nand U26695 (N_26695,N_23585,N_21908);
xor U26696 (N_26696,N_22795,N_23509);
or U26697 (N_26697,N_21181,N_23769);
and U26698 (N_26698,N_21841,N_21171);
nor U26699 (N_26699,N_22358,N_22747);
or U26700 (N_26700,N_21706,N_23717);
xnor U26701 (N_26701,N_22717,N_21716);
nand U26702 (N_26702,N_21920,N_23743);
nand U26703 (N_26703,N_22773,N_21633);
xnor U26704 (N_26704,N_21652,N_21546);
nor U26705 (N_26705,N_21550,N_23067);
and U26706 (N_26706,N_23380,N_23518);
or U26707 (N_26707,N_23266,N_22047);
nor U26708 (N_26708,N_23502,N_23233);
xnor U26709 (N_26709,N_22339,N_22262);
and U26710 (N_26710,N_23214,N_23518);
nor U26711 (N_26711,N_22828,N_21269);
nor U26712 (N_26712,N_22380,N_22464);
nand U26713 (N_26713,N_21328,N_21657);
or U26714 (N_26714,N_22183,N_21217);
nand U26715 (N_26715,N_23065,N_22447);
xnor U26716 (N_26716,N_21390,N_21583);
or U26717 (N_26717,N_23771,N_21060);
or U26718 (N_26718,N_22136,N_22870);
and U26719 (N_26719,N_21238,N_23299);
nor U26720 (N_26720,N_23291,N_21748);
nor U26721 (N_26721,N_21289,N_23450);
or U26722 (N_26722,N_21877,N_21183);
or U26723 (N_26723,N_21191,N_22669);
nand U26724 (N_26724,N_22516,N_21817);
nor U26725 (N_26725,N_23800,N_22401);
nor U26726 (N_26726,N_23902,N_23352);
or U26727 (N_26727,N_21942,N_23473);
xnor U26728 (N_26728,N_23214,N_21943);
nor U26729 (N_26729,N_23380,N_23927);
nand U26730 (N_26730,N_21066,N_22966);
xnor U26731 (N_26731,N_23051,N_22786);
and U26732 (N_26732,N_23522,N_22081);
nand U26733 (N_26733,N_22771,N_23670);
nand U26734 (N_26734,N_21204,N_21802);
xor U26735 (N_26735,N_23873,N_22675);
xor U26736 (N_26736,N_21441,N_21378);
and U26737 (N_26737,N_22810,N_23574);
nand U26738 (N_26738,N_21838,N_23151);
nor U26739 (N_26739,N_22786,N_21018);
nor U26740 (N_26740,N_22595,N_23504);
or U26741 (N_26741,N_22330,N_21283);
and U26742 (N_26742,N_21990,N_21191);
and U26743 (N_26743,N_21984,N_21308);
or U26744 (N_26744,N_23596,N_22147);
nand U26745 (N_26745,N_22735,N_23208);
and U26746 (N_26746,N_22612,N_23617);
xnor U26747 (N_26747,N_23472,N_21774);
nand U26748 (N_26748,N_22322,N_23857);
nor U26749 (N_26749,N_23426,N_23172);
and U26750 (N_26750,N_21946,N_23744);
or U26751 (N_26751,N_23004,N_23957);
nand U26752 (N_26752,N_22108,N_22846);
xnor U26753 (N_26753,N_22992,N_22690);
xnor U26754 (N_26754,N_22683,N_21170);
and U26755 (N_26755,N_23195,N_22976);
or U26756 (N_26756,N_23210,N_21391);
nand U26757 (N_26757,N_21847,N_22232);
and U26758 (N_26758,N_21344,N_22897);
nor U26759 (N_26759,N_22765,N_23185);
nor U26760 (N_26760,N_21921,N_22097);
or U26761 (N_26761,N_22541,N_23501);
or U26762 (N_26762,N_22579,N_23314);
nor U26763 (N_26763,N_21882,N_22740);
and U26764 (N_26764,N_23336,N_22434);
or U26765 (N_26765,N_23335,N_23840);
xnor U26766 (N_26766,N_23161,N_21277);
xnor U26767 (N_26767,N_22115,N_22420);
nor U26768 (N_26768,N_22441,N_21532);
nor U26769 (N_26769,N_23355,N_23695);
or U26770 (N_26770,N_21519,N_23691);
xnor U26771 (N_26771,N_21757,N_21536);
or U26772 (N_26772,N_21190,N_23868);
or U26773 (N_26773,N_22336,N_21727);
nor U26774 (N_26774,N_23705,N_22634);
nand U26775 (N_26775,N_21446,N_22457);
nor U26776 (N_26776,N_21912,N_21964);
xnor U26777 (N_26777,N_23795,N_21497);
nor U26778 (N_26778,N_21378,N_22842);
xnor U26779 (N_26779,N_22073,N_22335);
nor U26780 (N_26780,N_21397,N_23473);
or U26781 (N_26781,N_21979,N_21226);
and U26782 (N_26782,N_21804,N_22789);
nand U26783 (N_26783,N_21057,N_21051);
nor U26784 (N_26784,N_21594,N_22818);
and U26785 (N_26785,N_23320,N_22704);
xor U26786 (N_26786,N_23334,N_22700);
nand U26787 (N_26787,N_21220,N_22990);
nand U26788 (N_26788,N_22553,N_21180);
nand U26789 (N_26789,N_22067,N_23250);
and U26790 (N_26790,N_21083,N_21861);
xnor U26791 (N_26791,N_22627,N_23921);
or U26792 (N_26792,N_22152,N_23902);
or U26793 (N_26793,N_23006,N_21920);
nand U26794 (N_26794,N_23657,N_22752);
xnor U26795 (N_26795,N_22552,N_23684);
or U26796 (N_26796,N_22390,N_21924);
xnor U26797 (N_26797,N_21790,N_23958);
nand U26798 (N_26798,N_23661,N_22011);
xor U26799 (N_26799,N_21860,N_23557);
nor U26800 (N_26800,N_23199,N_22150);
and U26801 (N_26801,N_23082,N_23332);
and U26802 (N_26802,N_21642,N_23384);
or U26803 (N_26803,N_23020,N_22088);
nand U26804 (N_26804,N_22586,N_21379);
nor U26805 (N_26805,N_22038,N_21360);
xor U26806 (N_26806,N_21970,N_21075);
nor U26807 (N_26807,N_21685,N_21729);
xnor U26808 (N_26808,N_21977,N_22892);
nand U26809 (N_26809,N_21291,N_21968);
or U26810 (N_26810,N_22201,N_22652);
nor U26811 (N_26811,N_22613,N_21753);
or U26812 (N_26812,N_22972,N_22456);
xor U26813 (N_26813,N_21799,N_23193);
nand U26814 (N_26814,N_23318,N_21204);
nor U26815 (N_26815,N_23199,N_21003);
nand U26816 (N_26816,N_22248,N_21712);
and U26817 (N_26817,N_21522,N_21165);
nor U26818 (N_26818,N_22713,N_21549);
or U26819 (N_26819,N_23606,N_21502);
nor U26820 (N_26820,N_22097,N_22936);
nand U26821 (N_26821,N_23862,N_21871);
xnor U26822 (N_26822,N_23120,N_21408);
nand U26823 (N_26823,N_22348,N_21227);
or U26824 (N_26824,N_23690,N_21134);
and U26825 (N_26825,N_23532,N_21113);
xor U26826 (N_26826,N_22828,N_22187);
xor U26827 (N_26827,N_23456,N_22263);
nand U26828 (N_26828,N_21924,N_22025);
nand U26829 (N_26829,N_21256,N_21063);
nand U26830 (N_26830,N_22258,N_23786);
and U26831 (N_26831,N_23028,N_23922);
xor U26832 (N_26832,N_22425,N_22661);
nand U26833 (N_26833,N_21359,N_22160);
or U26834 (N_26834,N_23268,N_22099);
xor U26835 (N_26835,N_21956,N_21799);
and U26836 (N_26836,N_23401,N_21444);
nor U26837 (N_26837,N_21853,N_22198);
and U26838 (N_26838,N_22379,N_21432);
nor U26839 (N_26839,N_21764,N_23654);
and U26840 (N_26840,N_23400,N_21971);
nand U26841 (N_26841,N_21496,N_22165);
xnor U26842 (N_26842,N_22903,N_23627);
xnor U26843 (N_26843,N_21982,N_23434);
nor U26844 (N_26844,N_21806,N_23321);
nand U26845 (N_26845,N_23529,N_23936);
or U26846 (N_26846,N_21622,N_23320);
or U26847 (N_26847,N_23117,N_21488);
nand U26848 (N_26848,N_22358,N_21496);
or U26849 (N_26849,N_23221,N_21287);
and U26850 (N_26850,N_22603,N_22110);
xnor U26851 (N_26851,N_21812,N_21444);
or U26852 (N_26852,N_23525,N_23335);
xnor U26853 (N_26853,N_23146,N_21585);
nor U26854 (N_26854,N_23943,N_21726);
nor U26855 (N_26855,N_22670,N_23888);
nand U26856 (N_26856,N_23811,N_21969);
or U26857 (N_26857,N_21630,N_21716);
and U26858 (N_26858,N_23861,N_23909);
nand U26859 (N_26859,N_21969,N_22904);
and U26860 (N_26860,N_21541,N_21322);
xor U26861 (N_26861,N_21312,N_21694);
or U26862 (N_26862,N_21637,N_23384);
nand U26863 (N_26863,N_22676,N_23378);
nand U26864 (N_26864,N_22347,N_21820);
nor U26865 (N_26865,N_22946,N_22371);
nor U26866 (N_26866,N_21546,N_21734);
nor U26867 (N_26867,N_23075,N_22158);
and U26868 (N_26868,N_21880,N_21504);
and U26869 (N_26869,N_22492,N_21170);
and U26870 (N_26870,N_22212,N_22168);
or U26871 (N_26871,N_23169,N_22797);
or U26872 (N_26872,N_23854,N_22071);
and U26873 (N_26873,N_23660,N_21182);
and U26874 (N_26874,N_23358,N_23497);
nand U26875 (N_26875,N_23110,N_23549);
and U26876 (N_26876,N_23466,N_21898);
nand U26877 (N_26877,N_21347,N_22004);
or U26878 (N_26878,N_22364,N_21159);
or U26879 (N_26879,N_22852,N_21341);
xnor U26880 (N_26880,N_21159,N_21977);
nand U26881 (N_26881,N_23877,N_22187);
or U26882 (N_26882,N_23706,N_22630);
and U26883 (N_26883,N_23892,N_21885);
xnor U26884 (N_26884,N_23167,N_23241);
xnor U26885 (N_26885,N_22023,N_23667);
nand U26886 (N_26886,N_21176,N_22073);
or U26887 (N_26887,N_21664,N_21235);
and U26888 (N_26888,N_23746,N_23401);
or U26889 (N_26889,N_21974,N_22820);
or U26890 (N_26890,N_23966,N_21912);
nand U26891 (N_26891,N_23607,N_22690);
xnor U26892 (N_26892,N_22268,N_21258);
nor U26893 (N_26893,N_21920,N_21151);
or U26894 (N_26894,N_23849,N_22978);
nand U26895 (N_26895,N_21898,N_21553);
nor U26896 (N_26896,N_22824,N_22296);
and U26897 (N_26897,N_21975,N_23742);
nor U26898 (N_26898,N_23589,N_21855);
nand U26899 (N_26899,N_23154,N_21241);
or U26900 (N_26900,N_22942,N_22323);
or U26901 (N_26901,N_22869,N_23745);
xor U26902 (N_26902,N_22512,N_23415);
and U26903 (N_26903,N_22685,N_22917);
nor U26904 (N_26904,N_22331,N_21144);
nor U26905 (N_26905,N_21457,N_23676);
nor U26906 (N_26906,N_21182,N_23940);
xnor U26907 (N_26907,N_22444,N_23393);
nand U26908 (N_26908,N_22205,N_21872);
nand U26909 (N_26909,N_23128,N_23895);
and U26910 (N_26910,N_23673,N_23694);
or U26911 (N_26911,N_23720,N_22749);
and U26912 (N_26912,N_21807,N_22208);
nand U26913 (N_26913,N_21947,N_23654);
or U26914 (N_26914,N_23709,N_23755);
nor U26915 (N_26915,N_22808,N_21847);
or U26916 (N_26916,N_23950,N_22130);
nand U26917 (N_26917,N_23118,N_23322);
and U26918 (N_26918,N_21059,N_21837);
and U26919 (N_26919,N_22186,N_23502);
nand U26920 (N_26920,N_21391,N_22082);
and U26921 (N_26921,N_22468,N_22093);
nand U26922 (N_26922,N_23103,N_21801);
nand U26923 (N_26923,N_23530,N_21603);
xor U26924 (N_26924,N_23240,N_23343);
nand U26925 (N_26925,N_21618,N_21863);
xor U26926 (N_26926,N_23208,N_23383);
and U26927 (N_26927,N_23812,N_22551);
nand U26928 (N_26928,N_21062,N_23315);
or U26929 (N_26929,N_21404,N_21238);
nor U26930 (N_26930,N_21590,N_23003);
xor U26931 (N_26931,N_22267,N_21322);
nor U26932 (N_26932,N_21166,N_23883);
xnor U26933 (N_26933,N_21066,N_21402);
nand U26934 (N_26934,N_22737,N_22830);
nand U26935 (N_26935,N_21324,N_21282);
nand U26936 (N_26936,N_22861,N_21004);
nor U26937 (N_26937,N_22080,N_23206);
nand U26938 (N_26938,N_21694,N_23761);
and U26939 (N_26939,N_23022,N_23262);
or U26940 (N_26940,N_22707,N_23516);
xnor U26941 (N_26941,N_21317,N_21544);
nand U26942 (N_26942,N_22241,N_21806);
and U26943 (N_26943,N_23644,N_22672);
and U26944 (N_26944,N_21673,N_21862);
and U26945 (N_26945,N_21217,N_22062);
nand U26946 (N_26946,N_22519,N_22167);
xor U26947 (N_26947,N_22551,N_22197);
or U26948 (N_26948,N_21495,N_22524);
nor U26949 (N_26949,N_22345,N_22653);
nand U26950 (N_26950,N_22160,N_21320);
or U26951 (N_26951,N_22316,N_23017);
nand U26952 (N_26952,N_23548,N_21587);
and U26953 (N_26953,N_21721,N_21777);
xor U26954 (N_26954,N_21684,N_21527);
or U26955 (N_26955,N_23848,N_21140);
nand U26956 (N_26956,N_22325,N_22112);
xor U26957 (N_26957,N_21650,N_21238);
xor U26958 (N_26958,N_21436,N_23518);
and U26959 (N_26959,N_22561,N_22628);
or U26960 (N_26960,N_21294,N_21802);
xnor U26961 (N_26961,N_23351,N_21216);
or U26962 (N_26962,N_22792,N_21575);
nand U26963 (N_26963,N_23096,N_23705);
nand U26964 (N_26964,N_23986,N_22872);
or U26965 (N_26965,N_21997,N_23949);
nand U26966 (N_26966,N_22967,N_22700);
xor U26967 (N_26967,N_22018,N_23596);
nand U26968 (N_26968,N_22443,N_22823);
nor U26969 (N_26969,N_22977,N_22619);
nand U26970 (N_26970,N_23165,N_21768);
xor U26971 (N_26971,N_21984,N_21569);
xor U26972 (N_26972,N_23150,N_22083);
xnor U26973 (N_26973,N_21449,N_22007);
and U26974 (N_26974,N_22957,N_23106);
xnor U26975 (N_26975,N_23064,N_23763);
xnor U26976 (N_26976,N_23193,N_21278);
nand U26977 (N_26977,N_21631,N_21749);
nor U26978 (N_26978,N_22101,N_21752);
and U26979 (N_26979,N_23468,N_22577);
nor U26980 (N_26980,N_22804,N_21738);
and U26981 (N_26981,N_23797,N_23126);
nand U26982 (N_26982,N_23054,N_21829);
xor U26983 (N_26983,N_21407,N_21413);
and U26984 (N_26984,N_21310,N_21577);
and U26985 (N_26985,N_21199,N_22240);
nor U26986 (N_26986,N_21876,N_21283);
and U26987 (N_26987,N_23479,N_23452);
nand U26988 (N_26988,N_22647,N_23683);
nor U26989 (N_26989,N_21237,N_23388);
or U26990 (N_26990,N_21008,N_22070);
and U26991 (N_26991,N_21945,N_23200);
nand U26992 (N_26992,N_21851,N_23487);
nor U26993 (N_26993,N_22036,N_22479);
nor U26994 (N_26994,N_23763,N_21947);
or U26995 (N_26995,N_21728,N_22182);
nand U26996 (N_26996,N_23859,N_23825);
xnor U26997 (N_26997,N_21368,N_23488);
or U26998 (N_26998,N_22700,N_21993);
nand U26999 (N_26999,N_21214,N_23822);
xor U27000 (N_27000,N_25673,N_25612);
nand U27001 (N_27001,N_25309,N_24543);
and U27002 (N_27002,N_26106,N_26008);
xor U27003 (N_27003,N_24190,N_25846);
nand U27004 (N_27004,N_24551,N_26322);
and U27005 (N_27005,N_25529,N_26691);
xnor U27006 (N_27006,N_25955,N_26382);
nand U27007 (N_27007,N_25752,N_25352);
nand U27008 (N_27008,N_25844,N_26635);
nand U27009 (N_27009,N_25975,N_25656);
and U27010 (N_27010,N_25780,N_25029);
xnor U27011 (N_27011,N_24055,N_25927);
nor U27012 (N_27012,N_24455,N_25242);
or U27013 (N_27013,N_26113,N_25324);
nor U27014 (N_27014,N_25938,N_26619);
xnor U27015 (N_27015,N_24892,N_25197);
nor U27016 (N_27016,N_25199,N_25746);
nand U27017 (N_27017,N_26056,N_24705);
or U27018 (N_27018,N_26513,N_24809);
nor U27019 (N_27019,N_24471,N_26039);
or U27020 (N_27020,N_26125,N_25789);
or U27021 (N_27021,N_26249,N_26412);
and U27022 (N_27022,N_24421,N_25775);
nor U27023 (N_27023,N_25727,N_26343);
and U27024 (N_27024,N_26416,N_26243);
nor U27025 (N_27025,N_24383,N_26456);
nor U27026 (N_27026,N_26407,N_25383);
and U27027 (N_27027,N_26506,N_26897);
nor U27028 (N_27028,N_26973,N_26142);
nor U27029 (N_27029,N_25616,N_26172);
xor U27030 (N_27030,N_25390,N_25555);
nand U27031 (N_27031,N_26188,N_26858);
and U27032 (N_27032,N_26203,N_25883);
xnor U27033 (N_27033,N_25837,N_26624);
and U27034 (N_27034,N_24032,N_24107);
and U27035 (N_27035,N_25118,N_25804);
nor U27036 (N_27036,N_26392,N_24340);
xnor U27037 (N_27037,N_25295,N_25454);
or U27038 (N_27038,N_26176,N_26074);
nor U27039 (N_27039,N_25561,N_25298);
and U27040 (N_27040,N_25218,N_26457);
or U27041 (N_27041,N_25693,N_26841);
and U27042 (N_27042,N_24479,N_26484);
or U27043 (N_27043,N_24634,N_26028);
nand U27044 (N_27044,N_24270,N_25411);
or U27045 (N_27045,N_25822,N_24367);
or U27046 (N_27046,N_26238,N_24191);
nor U27047 (N_27047,N_26754,N_24748);
nor U27048 (N_27048,N_26546,N_25562);
nand U27049 (N_27049,N_26710,N_26356);
nand U27050 (N_27050,N_25914,N_24973);
xor U27051 (N_27051,N_26795,N_25901);
or U27052 (N_27052,N_25488,N_26094);
and U27053 (N_27053,N_25525,N_25668);
and U27054 (N_27054,N_25545,N_25340);
nor U27055 (N_27055,N_26913,N_24192);
and U27056 (N_27056,N_25297,N_24928);
xor U27057 (N_27057,N_24791,N_24038);
or U27058 (N_27058,N_25947,N_26507);
nor U27059 (N_27059,N_24310,N_24042);
and U27060 (N_27060,N_25660,N_25861);
xor U27061 (N_27061,N_24811,N_25318);
nand U27062 (N_27062,N_26420,N_24959);
and U27063 (N_27063,N_24929,N_25267);
and U27064 (N_27064,N_26267,N_25048);
or U27065 (N_27065,N_25217,N_24901);
nor U27066 (N_27066,N_24043,N_24004);
nor U27067 (N_27067,N_25294,N_26006);
or U27068 (N_27068,N_24537,N_24667);
or U27069 (N_27069,N_26571,N_24112);
nor U27070 (N_27070,N_24956,N_26399);
and U27071 (N_27071,N_24690,N_26823);
or U27072 (N_27072,N_26721,N_24681);
and U27073 (N_27073,N_26995,N_24234);
nor U27074 (N_27074,N_24179,N_25039);
nor U27075 (N_27075,N_24835,N_26562);
nand U27076 (N_27076,N_25253,N_26610);
nor U27077 (N_27077,N_25916,N_24418);
xor U27078 (N_27078,N_24309,N_25394);
xnor U27079 (N_27079,N_26859,N_24244);
xnor U27080 (N_27080,N_25892,N_24668);
nor U27081 (N_27081,N_25310,N_26538);
or U27082 (N_27082,N_25364,N_24064);
and U27083 (N_27083,N_25361,N_25317);
and U27084 (N_27084,N_24000,N_24049);
xor U27085 (N_27085,N_26964,N_26650);
and U27086 (N_27086,N_26334,N_25874);
nor U27087 (N_27087,N_26566,N_24328);
nand U27088 (N_27088,N_25675,N_24499);
nand U27089 (N_27089,N_24731,N_24530);
nor U27090 (N_27090,N_26477,N_26517);
or U27091 (N_27091,N_25836,N_26908);
nor U27092 (N_27092,N_26173,N_26625);
and U27093 (N_27093,N_24780,N_24905);
nand U27094 (N_27094,N_25401,N_26470);
xor U27095 (N_27095,N_24154,N_25589);
and U27096 (N_27096,N_25569,N_25246);
and U27097 (N_27097,N_25876,N_24075);
xor U27098 (N_27098,N_26946,N_25615);
nor U27099 (N_27099,N_25234,N_26579);
xor U27100 (N_27100,N_26344,N_24022);
nand U27101 (N_27101,N_26664,N_24862);
xnor U27102 (N_27102,N_25412,N_26421);
xnor U27103 (N_27103,N_26263,N_26910);
nand U27104 (N_27104,N_25858,N_25337);
and U27105 (N_27105,N_26554,N_26174);
xor U27106 (N_27106,N_26881,N_26530);
nor U27107 (N_27107,N_25802,N_24797);
or U27108 (N_27108,N_25951,N_24073);
nor U27109 (N_27109,N_25105,N_26775);
and U27110 (N_27110,N_26455,N_24206);
and U27111 (N_27111,N_24024,N_24060);
nand U27112 (N_27112,N_26527,N_24294);
xor U27113 (N_27113,N_26207,N_24239);
nand U27114 (N_27114,N_24723,N_26861);
xnor U27115 (N_27115,N_26069,N_24123);
and U27116 (N_27116,N_24896,N_25522);
or U27117 (N_27117,N_26269,N_24695);
or U27118 (N_27118,N_26866,N_26580);
and U27119 (N_27119,N_25015,N_24879);
or U27120 (N_27120,N_25765,N_24752);
xnor U27121 (N_27121,N_24981,N_24227);
and U27122 (N_27122,N_26864,N_26958);
nor U27123 (N_27123,N_26879,N_26501);
xnor U27124 (N_27124,N_25872,N_24618);
xnor U27125 (N_27125,N_25647,N_26091);
nor U27126 (N_27126,N_25950,N_25028);
nand U27127 (N_27127,N_25059,N_26418);
xnor U27128 (N_27128,N_26835,N_26242);
nand U27129 (N_27129,N_24156,N_25046);
nor U27130 (N_27130,N_24229,N_24617);
and U27131 (N_27131,N_26101,N_25308);
and U27132 (N_27132,N_26615,N_25447);
and U27133 (N_27133,N_26602,N_24846);
nor U27134 (N_27134,N_24373,N_25206);
and U27135 (N_27135,N_24980,N_25396);
or U27136 (N_27136,N_24619,N_24880);
nand U27137 (N_27137,N_25890,N_25508);
nand U27138 (N_27138,N_24703,N_25236);
nor U27139 (N_27139,N_26641,N_26902);
or U27140 (N_27140,N_25358,N_26651);
xor U27141 (N_27141,N_24574,N_25185);
and U27142 (N_27142,N_25651,N_25728);
nand U27143 (N_27143,N_24236,N_25828);
xnor U27144 (N_27144,N_26439,N_25176);
xor U27145 (N_27145,N_26260,N_26276);
nand U27146 (N_27146,N_26289,N_26849);
nor U27147 (N_27147,N_24364,N_25257);
and U27148 (N_27148,N_25993,N_24408);
and U27149 (N_27149,N_26525,N_25877);
or U27150 (N_27150,N_24856,N_24938);
nor U27151 (N_27151,N_26985,N_25605);
nand U27152 (N_27152,N_25027,N_26303);
xor U27153 (N_27153,N_24113,N_26743);
nand U27154 (N_27154,N_24608,N_26646);
and U27155 (N_27155,N_24825,N_25331);
or U27156 (N_27156,N_24068,N_24144);
or U27157 (N_27157,N_26131,N_24491);
nor U27158 (N_27158,N_24385,N_24838);
xor U27159 (N_27159,N_26895,N_26012);
and U27160 (N_27160,N_24553,N_24945);
nor U27161 (N_27161,N_26396,N_25426);
xor U27162 (N_27162,N_25229,N_26424);
nor U27163 (N_27163,N_25400,N_24867);
or U27164 (N_27164,N_25266,N_26603);
or U27165 (N_27165,N_26219,N_24097);
and U27166 (N_27166,N_26844,N_25868);
nand U27167 (N_27167,N_26768,N_25170);
nor U27168 (N_27168,N_26883,N_25944);
nand U27169 (N_27169,N_24369,N_25293);
and U27170 (N_27170,N_25946,N_25491);
and U27171 (N_27171,N_25187,N_26827);
xor U27172 (N_27172,N_24734,N_26676);
or U27173 (N_27173,N_25408,N_25722);
and U27174 (N_27174,N_25788,N_26792);
xor U27175 (N_27175,N_26857,N_25057);
or U27176 (N_27176,N_25597,N_25359);
nand U27177 (N_27177,N_24626,N_24743);
or U27178 (N_27178,N_26773,N_24869);
xor U27179 (N_27179,N_26612,N_26876);
nand U27180 (N_27180,N_24785,N_26248);
xnor U27181 (N_27181,N_24218,N_25035);
nand U27182 (N_27182,N_26962,N_24381);
or U27183 (N_27183,N_26842,N_26986);
and U27184 (N_27184,N_25280,N_25999);
nand U27185 (N_27185,N_26675,N_25891);
and U27186 (N_27186,N_26087,N_25754);
or U27187 (N_27187,N_26496,N_25099);
xnor U27188 (N_27188,N_25304,N_24061);
or U27189 (N_27189,N_26891,N_26965);
nand U27190 (N_27190,N_24217,N_24372);
nand U27191 (N_27191,N_26670,N_26159);
nand U27192 (N_27192,N_26297,N_25044);
nor U27193 (N_27193,N_25483,N_26605);
nand U27194 (N_27194,N_25150,N_26593);
nand U27195 (N_27195,N_26256,N_26787);
and U27196 (N_27196,N_24352,N_26863);
nor U27197 (N_27197,N_26317,N_25356);
or U27198 (N_27198,N_25879,N_26257);
and U27199 (N_27199,N_26930,N_24569);
nor U27200 (N_27200,N_24254,N_26555);
or U27201 (N_27201,N_25366,N_26002);
nand U27202 (N_27202,N_26824,N_24860);
xnor U27203 (N_27203,N_26868,N_26432);
nor U27204 (N_27204,N_25751,N_26552);
and U27205 (N_27205,N_26059,N_26954);
or U27206 (N_27206,N_26434,N_26960);
and U27207 (N_27207,N_25766,N_24761);
and U27208 (N_27208,N_25225,N_26089);
nor U27209 (N_27209,N_24787,N_25554);
nand U27210 (N_27210,N_24771,N_25959);
xor U27211 (N_27211,N_25496,N_26030);
xor U27212 (N_27212,N_26110,N_25908);
nor U27213 (N_27213,N_25943,N_26018);
nor U27214 (N_27214,N_24729,N_25537);
nand U27215 (N_27215,N_26678,N_25133);
xnor U27216 (N_27216,N_25138,N_26104);
xnor U27217 (N_27217,N_25051,N_25985);
and U27218 (N_27218,N_24323,N_25896);
xor U27219 (N_27219,N_26431,N_25988);
nand U27220 (N_27220,N_25781,N_25729);
nand U27221 (N_27221,N_24972,N_25523);
xnor U27222 (N_27222,N_25797,N_25041);
nor U27223 (N_27223,N_25388,N_24028);
or U27224 (N_27224,N_25047,N_24386);
nor U27225 (N_27225,N_24422,N_24268);
or U27226 (N_27226,N_25533,N_24519);
nand U27227 (N_27227,N_24442,N_26892);
or U27228 (N_27228,N_26004,N_26498);
xnor U27229 (N_27229,N_26674,N_24476);
nor U27230 (N_27230,N_25919,N_24498);
nor U27231 (N_27231,N_26482,N_25686);
or U27232 (N_27232,N_25012,N_24586);
nand U27233 (N_27233,N_25799,N_24711);
nor U27234 (N_27234,N_26323,N_26078);
and U27235 (N_27235,N_24348,N_24429);
nand U27236 (N_27236,N_26940,N_26193);
nand U27237 (N_27237,N_25974,N_25247);
or U27238 (N_27238,N_26802,N_26869);
and U27239 (N_27239,N_24092,N_24708);
xor U27240 (N_27240,N_26730,N_25205);
nand U27241 (N_27241,N_25121,N_25313);
nor U27242 (N_27242,N_24193,N_26911);
xor U27243 (N_27243,N_25184,N_25724);
xnor U27244 (N_27244,N_25092,N_26390);
and U27245 (N_27245,N_24046,N_26614);
xnor U27246 (N_27246,N_26592,N_25906);
and U27247 (N_27247,N_24987,N_26732);
nor U27248 (N_27248,N_26529,N_25903);
nand U27249 (N_27249,N_25747,N_26111);
xor U27250 (N_27250,N_24834,N_24589);
nand U27251 (N_27251,N_25220,N_25104);
nor U27252 (N_27252,N_26971,N_24641);
nand U27253 (N_27253,N_25885,N_25859);
nor U27254 (N_27254,N_26175,N_24267);
and U27255 (N_27255,N_25888,N_26847);
xor U27256 (N_27256,N_24549,N_26693);
nor U27257 (N_27257,N_24245,N_25543);
nor U27258 (N_27258,N_24450,N_26291);
nand U27259 (N_27259,N_24917,N_24189);
nand U27260 (N_27260,N_26274,N_25194);
or U27261 (N_27261,N_26575,N_25375);
and U27262 (N_27262,N_26015,N_26932);
xor U27263 (N_27263,N_24246,N_24152);
and U27264 (N_27264,N_26572,N_26262);
nand U27265 (N_27265,N_24011,N_24333);
and U27266 (N_27266,N_25466,N_25536);
and U27267 (N_27267,N_25532,N_25557);
or U27268 (N_27268,N_26411,N_24506);
xor U27269 (N_27269,N_25259,N_26444);
nand U27270 (N_27270,N_24793,N_25272);
and U27271 (N_27271,N_26545,N_26143);
or U27272 (N_27272,N_24345,N_24305);
nor U27273 (N_27273,N_26948,N_25648);
nor U27274 (N_27274,N_25886,N_26987);
and U27275 (N_27275,N_25434,N_26837);
or U27276 (N_27276,N_24117,N_24539);
nand U27277 (N_27277,N_24861,N_24565);
nor U27278 (N_27278,N_25431,N_24344);
nand U27279 (N_27279,N_25839,N_26682);
nor U27280 (N_27280,N_24767,N_25976);
xnor U27281 (N_27281,N_25702,N_24788);
and U27282 (N_27282,N_24240,N_25312);
nand U27283 (N_27283,N_26425,N_24993);
and U27284 (N_27284,N_25068,N_24492);
or U27285 (N_27285,N_24623,N_26618);
xnor U27286 (N_27286,N_25639,N_24392);
or U27287 (N_27287,N_24757,N_25725);
nor U27288 (N_27288,N_26372,N_24921);
or U27289 (N_27289,N_25827,N_25207);
nor U27290 (N_27290,N_26011,N_26123);
and U27291 (N_27291,N_24223,N_24394);
or U27292 (N_27292,N_25867,N_24276);
or U27293 (N_27293,N_26715,N_26244);
nor U27294 (N_27294,N_25601,N_26349);
xnor U27295 (N_27295,N_26124,N_24720);
nor U27296 (N_27296,N_25435,N_25215);
nand U27297 (N_27297,N_24495,N_26067);
and U27298 (N_27298,N_25924,N_25534);
nand U27299 (N_27299,N_24898,N_26966);
nor U27300 (N_27300,N_26254,N_25759);
xor U27301 (N_27301,N_24907,N_26413);
nor U27302 (N_27302,N_25241,N_24363);
and U27303 (N_27303,N_25347,N_25430);
nand U27304 (N_27304,N_25911,N_24315);
and U27305 (N_27305,N_26049,N_26326);
nor U27306 (N_27306,N_25991,N_24642);
or U27307 (N_27307,N_25037,N_24766);
and U27308 (N_27308,N_24978,N_24889);
xor U27309 (N_27309,N_26998,N_25657);
and U27310 (N_27310,N_26836,N_26443);
and U27311 (N_27311,N_25417,N_24427);
or U27312 (N_27312,N_25414,N_25492);
xnor U27313 (N_27313,N_25969,N_26989);
or U27314 (N_27314,N_24078,N_24090);
xor U27315 (N_27315,N_26728,N_26856);
and U27316 (N_27316,N_24451,N_26606);
nor U27317 (N_27317,N_25416,N_26268);
or U27318 (N_27318,N_24529,N_24319);
or U27319 (N_27319,N_24027,N_24709);
nand U27320 (N_27320,N_25973,N_25591);
nand U27321 (N_27321,N_25287,N_24604);
nand U27322 (N_27322,N_26955,N_26258);
xnor U27323 (N_27323,N_26312,N_25320);
or U27324 (N_27324,N_24958,N_25608);
nor U27325 (N_27325,N_25243,N_25026);
xor U27326 (N_27326,N_24253,N_26748);
xnor U27327 (N_27327,N_25147,N_24966);
and U27328 (N_27328,N_26817,N_25713);
nand U27329 (N_27329,N_24505,N_25278);
nor U27330 (N_27330,N_24955,N_25744);
nor U27331 (N_27331,N_25967,N_25820);
or U27332 (N_27332,N_24080,N_26947);
nand U27333 (N_27333,N_26819,N_25376);
and U27334 (N_27334,N_26638,N_25311);
and U27335 (N_27335,N_24969,N_25763);
xnor U27336 (N_27336,N_25263,N_26400);
and U27337 (N_27337,N_26631,N_26365);
or U27338 (N_27338,N_24868,N_25681);
and U27339 (N_27339,N_24658,N_26265);
and U27340 (N_27340,N_26634,N_24473);
xor U27341 (N_27341,N_26153,N_25101);
and U27342 (N_27342,N_26522,N_26843);
nand U27343 (N_27343,N_24178,N_25606);
nand U27344 (N_27344,N_24899,N_25449);
or U27345 (N_27345,N_24753,N_24388);
nand U27346 (N_27346,N_26723,N_24164);
and U27347 (N_27347,N_26611,N_26315);
nor U27348 (N_27348,N_26216,N_26133);
nor U27349 (N_27349,N_25004,N_24069);
xor U27350 (N_27350,N_26719,N_24976);
nor U27351 (N_27351,N_24754,N_24453);
nor U27352 (N_27352,N_26179,N_24226);
nor U27353 (N_27353,N_26832,N_25083);
xnor U27354 (N_27354,N_25638,N_26366);
xnor U27355 (N_27355,N_25108,N_24613);
or U27356 (N_27356,N_26384,N_25604);
and U27357 (N_27357,N_25032,N_26758);
nand U27358 (N_27358,N_25140,N_25952);
xor U27359 (N_27359,N_25462,N_26925);
xor U27360 (N_27360,N_25850,N_26241);
and U27361 (N_27361,N_24103,N_26387);
nor U27362 (N_27362,N_24630,N_25327);
nand U27363 (N_27363,N_26449,N_24895);
nand U27364 (N_27364,N_25678,N_24510);
nor U27365 (N_27365,N_26117,N_25010);
nand U27366 (N_27366,N_26929,N_24402);
nor U27367 (N_27367,N_24124,N_24607);
nor U27368 (N_27368,N_24298,N_26454);
nand U27369 (N_27369,N_25030,N_24412);
nor U27370 (N_27370,N_25459,N_26191);
or U27371 (N_27371,N_24170,N_24366);
or U27372 (N_27372,N_25995,N_25696);
and U27373 (N_27373,N_25233,N_26036);
xnor U27374 (N_27374,N_26846,N_25602);
nand U27375 (N_27375,N_24911,N_24849);
and U27376 (N_27376,N_24685,N_26669);
xor U27377 (N_27377,N_26829,N_25348);
or U27378 (N_27378,N_25553,N_26493);
and U27379 (N_27379,N_24303,N_24647);
nand U27380 (N_27380,N_25421,N_26550);
xnor U27381 (N_27381,N_26044,N_26630);
xor U27382 (N_27382,N_25189,N_26747);
nand U27383 (N_27383,N_26494,N_26724);
and U27384 (N_27384,N_24409,N_26043);
nand U27385 (N_27385,N_24930,N_26632);
xor U27386 (N_27386,N_25878,N_24198);
xnor U27387 (N_27387,N_26812,N_25962);
xor U27388 (N_27388,N_24926,N_25521);
and U27389 (N_27389,N_24775,N_26608);
xor U27390 (N_27390,N_26205,N_26616);
and U27391 (N_27391,N_24350,N_26027);
or U27392 (N_27392,N_24201,N_26272);
nand U27393 (N_27393,N_26488,N_26475);
xnor U27394 (N_27394,N_24670,N_26800);
nor U27395 (N_27395,N_26351,N_25214);
and U27396 (N_27396,N_24763,N_25934);
or U27397 (N_27397,N_24435,N_24019);
xor U27398 (N_27398,N_24238,N_25661);
nand U27399 (N_27399,N_25210,N_25931);
nor U27400 (N_27400,N_24745,N_26626);
nor U27401 (N_27401,N_24555,N_25464);
nor U27402 (N_27402,N_26275,N_24772);
or U27403 (N_27403,N_25814,N_24304);
xnor U27404 (N_27404,N_24095,N_24196);
nor U27405 (N_27405,N_24676,N_24398);
or U27406 (N_27406,N_24337,N_24516);
xor U27407 (N_27407,N_24532,N_25279);
and U27408 (N_27408,N_25631,N_25670);
and U27409 (N_27409,N_24378,N_24301);
nor U27410 (N_27410,N_25302,N_25831);
nand U27411 (N_27411,N_25600,N_25134);
and U27412 (N_27412,N_26548,N_25918);
xor U27413 (N_27413,N_25504,N_26686);
nor U27414 (N_27414,N_24354,N_24045);
and U27415 (N_27415,N_25418,N_24517);
and U27416 (N_27416,N_24628,N_25617);
or U27417 (N_27417,N_26515,N_24581);
or U27418 (N_27418,N_25107,N_26406);
nor U27419 (N_27419,N_26391,N_26290);
nor U27420 (N_27420,N_25611,N_24133);
and U27421 (N_27421,N_25900,N_24824);
xor U27422 (N_27422,N_25117,N_24329);
nand U27423 (N_27423,N_25330,N_26224);
and U27424 (N_27424,N_24052,N_26358);
xor U27425 (N_27425,N_26329,N_24806);
nor U27426 (N_27426,N_24454,N_24211);
and U27427 (N_27427,N_26689,N_25285);
and U27428 (N_27428,N_24284,N_25120);
or U27429 (N_27429,N_25904,N_24908);
nor U27430 (N_27430,N_26834,N_24759);
or U27431 (N_27431,N_24410,N_26361);
and U27432 (N_27432,N_24687,N_24698);
xnor U27433 (N_27433,N_25803,N_24233);
xnor U27434 (N_27434,N_24215,N_25568);
and U27435 (N_27435,N_26797,N_26588);
nor U27436 (N_27436,N_26814,N_24248);
and U27437 (N_27437,N_25873,N_24571);
xor U27438 (N_27438,N_26782,N_25080);
xnor U27439 (N_27439,N_25232,N_25477);
and U27440 (N_27440,N_25021,N_24612);
nor U27441 (N_27441,N_25110,N_26848);
nor U27442 (N_27442,N_26668,N_25219);
and U27443 (N_27443,N_24166,N_26983);
nor U27444 (N_27444,N_24620,N_25097);
nand U27445 (N_27445,N_24358,N_26453);
or U27446 (N_27446,N_25992,N_25392);
nor U27447 (N_27447,N_26389,N_24853);
xnor U27448 (N_27448,N_26707,N_25091);
or U27449 (N_27449,N_24674,N_25132);
nor U27450 (N_27450,N_24213,N_25453);
nor U27451 (N_27451,N_24437,N_24988);
and U27452 (N_27452,N_25957,N_25773);
nor U27453 (N_27453,N_24979,N_24464);
or U27454 (N_27454,N_25166,N_24768);
xnor U27455 (N_27455,N_24527,N_26574);
nor U27456 (N_27456,N_25432,N_24833);
or U27457 (N_27457,N_26316,N_24132);
or U27458 (N_27458,N_24953,N_26874);
or U27459 (N_27459,N_24736,N_25758);
or U27460 (N_27460,N_26048,N_26975);
xor U27461 (N_27461,N_24269,N_26499);
xor U27462 (N_27462,N_25982,N_25481);
nand U27463 (N_27463,N_24564,N_24325);
and U27464 (N_27464,N_25167,N_24286);
and U27465 (N_27465,N_26750,N_24405);
and U27466 (N_27466,N_26543,N_26705);
nand U27467 (N_27467,N_25405,N_24614);
xor U27468 (N_27468,N_26033,N_26127);
nor U27469 (N_27469,N_24995,N_25354);
nor U27470 (N_27470,N_26560,N_26502);
or U27471 (N_27471,N_24436,N_26234);
nor U27472 (N_27472,N_24082,N_24875);
and U27473 (N_27473,N_25755,N_24669);
nor U27474 (N_27474,N_24857,N_26557);
or U27475 (N_27475,N_26158,N_26704);
or U27476 (N_27476,N_24949,N_24120);
or U27477 (N_27477,N_26559,N_24523);
and U27478 (N_27478,N_26526,N_25960);
nor U27479 (N_27479,N_26586,N_24939);
nor U27480 (N_27480,N_25559,N_25177);
xor U27481 (N_27481,N_26516,N_26135);
nor U27482 (N_27482,N_24913,N_24327);
and U27483 (N_27483,N_24487,N_25123);
nand U27484 (N_27484,N_26473,N_26357);
and U27485 (N_27485,N_25428,N_25350);
nor U27486 (N_27486,N_25451,N_25694);
nand U27487 (N_27487,N_25077,N_26286);
and U27488 (N_27488,N_26239,N_25355);
or U27489 (N_27489,N_24462,N_25966);
nor U27490 (N_27490,N_26152,N_25855);
nand U27491 (N_27491,N_26833,N_25650);
nand U27492 (N_27492,N_25144,N_25475);
nand U27493 (N_27493,N_24118,N_25096);
and U27494 (N_27494,N_25192,N_24985);
nand U27495 (N_27495,N_26894,N_25701);
and U27496 (N_27496,N_25461,N_25753);
and U27497 (N_27497,N_24209,N_26259);
nand U27498 (N_27498,N_26500,N_25299);
xnor U27499 (N_27499,N_25180,N_25250);
xnor U27500 (N_27500,N_26565,N_26031);
nor U27501 (N_27501,N_24205,N_26569);
nor U27502 (N_27502,N_26957,N_26737);
nand U27503 (N_27503,N_24463,N_24362);
nor U27504 (N_27504,N_26505,N_26162);
and U27505 (N_27505,N_24430,N_25145);
nand U27506 (N_27506,N_24001,N_26665);
or U27507 (N_27507,N_26330,N_24468);
or U27508 (N_27508,N_24289,N_25685);
nor U27509 (N_27509,N_24514,N_26064);
nor U27510 (N_27510,N_24774,N_24792);
or U27511 (N_27511,N_26026,N_26582);
and U27512 (N_27512,N_24106,N_24314);
xnor U27513 (N_27513,N_25894,N_26130);
xnor U27514 (N_27514,N_26255,N_26717);
xor U27515 (N_27515,N_26383,N_24756);
nor U27516 (N_27516,N_24130,N_25023);
nand U27517 (N_27517,N_24762,N_25198);
nor U27518 (N_27518,N_24041,N_26250);
or U27519 (N_27519,N_24876,N_26001);
nor U27520 (N_27520,N_25905,N_24273);
nor U27521 (N_27521,N_26884,N_25663);
nor U27522 (N_27522,N_26972,N_25439);
nor U27523 (N_27523,N_24417,N_24025);
xnor U27524 (N_27524,N_25707,N_25811);
or U27525 (N_27525,N_25609,N_24906);
nor U27526 (N_27526,N_24307,N_26872);
xnor U27527 (N_27527,N_26215,N_25169);
nor U27528 (N_27528,N_24300,N_24382);
or U27529 (N_27529,N_25070,N_25996);
and U27530 (N_27530,N_26950,N_25619);
and U27531 (N_27531,N_24320,N_25446);
or U27532 (N_27532,N_24518,N_24677);
xnor U27533 (N_27533,N_26350,N_26165);
nand U27534 (N_27534,N_26054,N_26301);
nor U27535 (N_27535,N_26440,N_25863);
nand U27536 (N_27536,N_24472,N_26374);
and U27537 (N_27537,N_25706,N_24359);
xnor U27538 (N_27538,N_25457,N_24458);
nor U27539 (N_27539,N_24018,N_25761);
nand U27540 (N_27540,N_25128,N_26084);
nor U27541 (N_27541,N_24635,N_26898);
and U27542 (N_27542,N_26035,N_25816);
or U27543 (N_27543,N_25020,N_24143);
nand U27544 (N_27544,N_24904,N_24848);
nor U27545 (N_27545,N_26620,N_25042);
nor U27546 (N_27546,N_24016,N_26781);
and U27547 (N_27547,N_25472,N_25291);
or U27548 (N_27548,N_24513,N_25014);
or U27549 (N_27549,N_26659,N_24413);
and U27550 (N_27550,N_25588,N_24511);
or U27551 (N_27551,N_24807,N_24747);
and U27552 (N_27552,N_24950,N_24886);
xnor U27553 (N_27553,N_24679,N_24449);
nor U27554 (N_27554,N_25062,N_24675);
or U27555 (N_27555,N_25343,N_25898);
and U27556 (N_27556,N_24063,N_25164);
and U27557 (N_27557,N_24741,N_25641);
nand U27558 (N_27558,N_25520,N_26199);
or U27559 (N_27559,N_24556,N_25452);
nor U27560 (N_27560,N_25321,N_26694);
nand U27561 (N_27561,N_25902,N_25478);
and U27562 (N_27562,N_24989,N_26105);
or U27563 (N_27563,N_26144,N_24125);
nand U27564 (N_27564,N_25926,N_24440);
nor U27565 (N_27565,N_24704,N_26978);
xor U27566 (N_27566,N_26369,N_26777);
or U27567 (N_27567,N_25776,N_24952);
xnor U27568 (N_27568,N_24796,N_25018);
xor U27569 (N_27569,N_26007,N_26942);
and U27570 (N_27570,N_25281,N_26993);
or U27571 (N_27571,N_26311,N_25825);
xor U27572 (N_27572,N_26403,N_24007);
or U27573 (N_27573,N_26716,N_25049);
xor U27574 (N_27574,N_25531,N_25783);
or U27575 (N_27575,N_24694,N_26558);
or U27576 (N_27576,N_24802,N_26167);
nand U27577 (N_27577,N_25948,N_24331);
xnor U27578 (N_27578,N_24176,N_25190);
nor U27579 (N_27579,N_24087,N_24393);
and U27580 (N_27580,N_25270,N_24822);
or U27581 (N_27581,N_26486,N_25768);
or U27582 (N_27582,N_25642,N_26000);
xnor U27583 (N_27583,N_26821,N_26904);
or U27584 (N_27584,N_24592,N_24355);
and U27585 (N_27585,N_25530,N_24991);
and U27586 (N_27586,N_26916,N_24072);
nand U27587 (N_27587,N_26132,N_25201);
and U27588 (N_27588,N_24900,N_26109);
or U27589 (N_27589,N_25404,N_24026);
nor U27590 (N_27590,N_26685,N_25486);
or U27591 (N_27591,N_25407,N_26068);
nor U27592 (N_27592,N_24056,N_24466);
or U27593 (N_27593,N_24469,N_26483);
or U27594 (N_27594,N_26636,N_26663);
and U27595 (N_27595,N_25689,N_24817);
and U27596 (N_27596,N_24810,N_25627);
nand U27597 (N_27597,N_24021,N_25994);
xnor U27598 (N_27598,N_24291,N_26765);
nand U27599 (N_27599,N_26304,N_25316);
and U27600 (N_27600,N_25264,N_26447);
nor U27601 (N_27601,N_25239,N_24318);
nor U27602 (N_27602,N_25662,N_24664);
or U27603 (N_27603,N_25468,N_24660);
nor U27604 (N_27604,N_24122,N_26491);
xor U27605 (N_27605,N_24836,N_26660);
or U27606 (N_27606,N_24672,N_26598);
nor U27607 (N_27607,N_26564,N_24287);
and U27608 (N_27608,N_26789,N_26645);
nand U27609 (N_27609,N_26072,N_26367);
or U27610 (N_27610,N_26107,N_26979);
or U27611 (N_27611,N_26683,N_25249);
and U27612 (N_27612,N_25708,N_26838);
nor U27613 (N_27613,N_25618,N_26058);
and U27614 (N_27614,N_24962,N_25745);
nand U27615 (N_27615,N_25666,N_24292);
nand U27616 (N_27616,N_26283,N_25511);
xor U27617 (N_27617,N_24884,N_25260);
nand U27618 (N_27618,N_24415,N_25748);
nand U27619 (N_27619,N_24439,N_26793);
and U27620 (N_27620,N_25860,N_24459);
and U27621 (N_27621,N_25510,N_24339);
nand U27622 (N_27622,N_25547,N_25528);
or U27623 (N_27623,N_26353,N_26342);
or U27624 (N_27624,N_26233,N_26279);
nor U27625 (N_27625,N_26808,N_26534);
nor U27626 (N_27626,N_26873,N_25932);
and U27627 (N_27627,N_25305,N_26448);
nor U27628 (N_27628,N_24088,N_25289);
and U27629 (N_27629,N_24610,N_24841);
or U27630 (N_27630,N_24371,N_26034);
and U27631 (N_27631,N_26156,N_24582);
or U27632 (N_27632,N_26271,N_26761);
nand U27633 (N_27633,N_24065,N_25715);
xnor U27634 (N_27634,N_24081,N_25398);
nor U27635 (N_27635,N_25990,N_26200);
xor U27636 (N_27636,N_26753,N_25997);
nor U27637 (N_27637,N_26828,N_24560);
or U27638 (N_27638,N_24376,N_26146);
or U27639 (N_27639,N_26112,N_25186);
or U27640 (N_27640,N_26459,N_25275);
or U27641 (N_27641,N_24142,N_24591);
nand U27642 (N_27642,N_25319,N_24036);
nand U27643 (N_27643,N_25805,N_24770);
nor U27644 (N_27644,N_24139,N_24361);
xor U27645 (N_27645,N_26230,N_25777);
or U27646 (N_27646,N_26464,N_26292);
nand U27647 (N_27647,N_26968,N_24057);
and U27648 (N_27648,N_26512,N_25683);
nand U27649 (N_27649,N_25779,N_25550);
and U27650 (N_27650,N_24902,N_26338);
nor U27651 (N_27651,N_26760,N_25127);
or U27652 (N_27652,N_26914,N_24751);
xnor U27653 (N_27653,N_25500,N_25025);
or U27654 (N_27654,N_25565,N_26788);
and U27655 (N_27655,N_25502,N_24071);
xnor U27656 (N_27656,N_24540,N_24663);
nand U27657 (N_27657,N_24579,N_26170);
and U27658 (N_27658,N_25979,N_24724);
nor U27659 (N_27659,N_24483,N_25196);
nor U27660 (N_27660,N_24854,N_25181);
nor U27661 (N_27661,N_24659,N_25567);
or U27662 (N_27662,N_25684,N_25750);
nor U27663 (N_27663,N_24311,N_25594);
nand U27664 (N_27664,N_26264,N_25913);
nand U27665 (N_27665,N_25961,N_26196);
or U27666 (N_27666,N_26991,N_26887);
or U27667 (N_27667,N_26852,N_24850);
nor U27668 (N_27668,N_25235,N_26961);
nor U27669 (N_27669,N_25445,N_24525);
or U27670 (N_27670,N_25762,N_24404);
and U27671 (N_27671,N_25909,N_25625);
xor U27672 (N_27672,N_26769,N_24781);
and U27673 (N_27673,N_24477,N_26302);
nor U27674 (N_27674,N_24866,N_24522);
nand U27675 (N_27675,N_26161,N_25085);
or U27676 (N_27676,N_26734,N_24452);
nand U27677 (N_27677,N_26485,N_26013);
or U27678 (N_27678,N_25122,N_26941);
nor U27679 (N_27679,N_24353,N_26540);
xnor U27680 (N_27680,N_25437,N_24725);
nor U27681 (N_27681,N_24387,N_26436);
nand U27682 (N_27682,N_26115,N_24923);
xor U27683 (N_27683,N_25463,N_24322);
nand U27684 (N_27684,N_24086,N_24843);
xor U27685 (N_27685,N_24308,N_24534);
and U27686 (N_27686,N_25116,N_24666);
or U27687 (N_27687,N_26818,N_24277);
nand U27688 (N_27688,N_25503,N_24794);
nor U27689 (N_27689,N_25322,N_24374);
or U27690 (N_27690,N_24131,N_25810);
or U27691 (N_27691,N_24147,N_25283);
and U27692 (N_27692,N_25182,N_26981);
or U27693 (N_27693,N_24101,N_26820);
or U27694 (N_27694,N_24494,N_24249);
or U27695 (N_27695,N_25829,N_24338);
nand U27696 (N_27696,N_25143,N_24158);
and U27697 (N_27697,N_26251,N_25507);
nor U27698 (N_27698,N_24489,N_26997);
nor U27699 (N_27699,N_26921,N_25157);
nand U27700 (N_27700,N_24974,N_24598);
xor U27701 (N_27701,N_25254,N_24925);
nand U27702 (N_27702,N_26759,N_25323);
nand U27703 (N_27703,N_26318,N_26655);
or U27704 (N_27704,N_24157,N_26809);
nor U27705 (N_27705,N_25385,N_25734);
nor U27706 (N_27706,N_26282,N_24738);
or U27707 (N_27707,N_24365,N_25252);
xnor U27708 (N_27708,N_25476,N_24261);
nor U27709 (N_27709,N_26212,N_25692);
xor U27710 (N_27710,N_26394,N_26519);
nand U27711 (N_27711,N_26553,N_25887);
nor U27712 (N_27712,N_25209,N_26969);
xnor U27713 (N_27713,N_24058,N_25636);
or U27714 (N_27714,N_26229,N_26596);
xnor U27715 (N_27715,N_26801,N_25817);
and U27716 (N_27716,N_26232,N_26523);
or U27717 (N_27717,N_26549,N_25524);
nor U27718 (N_27718,N_24099,N_26147);
nand U27719 (N_27719,N_25968,N_26816);
xnor U27720 (N_27720,N_24710,N_24208);
or U27721 (N_27721,N_25493,N_25112);
xor U27722 (N_27722,N_25705,N_26798);
or U27723 (N_27723,N_26157,N_25422);
or U27724 (N_27724,N_26583,N_25490);
xnor U27725 (N_27725,N_24983,N_26647);
or U27726 (N_27726,N_26053,N_24758);
and U27727 (N_27727,N_24111,N_25301);
or U27728 (N_27728,N_26992,N_26749);
xnor U27729 (N_27729,N_25599,N_25942);
xor U27730 (N_27730,N_25163,N_25442);
nand U27731 (N_27731,N_26752,N_24247);
and U27732 (N_27732,N_24533,N_26168);
nor U27733 (N_27733,N_24638,N_24934);
xor U27734 (N_27734,N_26362,N_26755);
and U27735 (N_27735,N_25633,N_25223);
nor U27736 (N_27736,N_25749,N_26126);
nand U27737 (N_27737,N_25980,N_25760);
or U27738 (N_27738,N_24882,N_26308);
nand U27739 (N_27739,N_25494,N_26570);
xnor U27740 (N_27740,N_26469,N_24935);
nand U27741 (N_27741,N_24077,N_25251);
nor U27742 (N_27742,N_24181,N_24971);
or U27743 (N_27743,N_26936,N_25341);
and U27744 (N_27744,N_25596,N_25339);
nor U27745 (N_27745,N_25587,N_25643);
or U27746 (N_27746,N_25098,N_25470);
xnor U27747 (N_27747,N_26703,N_25130);
and U27748 (N_27748,N_24521,N_26221);
xnor U27749 (N_27749,N_25764,N_24400);
or U27750 (N_27750,N_24837,N_24031);
and U27751 (N_27751,N_25081,N_26671);
nor U27752 (N_27752,N_26584,N_24558);
nand U27753 (N_27753,N_24845,N_24151);
and U27754 (N_27754,N_25704,N_26096);
nand U27755 (N_27755,N_25495,N_25928);
and U27756 (N_27756,N_25815,N_26882);
nand U27757 (N_27757,N_25373,N_26364);
and U27758 (N_27758,N_26341,N_26273);
and U27759 (N_27759,N_25770,N_25677);
and U27760 (N_27760,N_25427,N_25929);
nor U27761 (N_27761,N_24783,N_25221);
nor U27762 (N_27762,N_24351,N_25832);
nand U27763 (N_27763,N_24411,N_24960);
nand U27764 (N_27764,N_24033,N_25469);
xnor U27765 (N_27765,N_24914,N_26590);
nand U27766 (N_27766,N_26017,N_25635);
xnor U27767 (N_27767,N_25935,N_24829);
nand U27768 (N_27768,N_26393,N_25579);
or U27769 (N_27769,N_26780,N_26514);
xor U27770 (N_27770,N_24174,N_25630);
and U27771 (N_27771,N_25771,N_26185);
xnor U27772 (N_27772,N_24927,N_24755);
or U27773 (N_27773,N_24335,N_24716);
xnor U27774 (N_27774,N_25620,N_24883);
nor U27775 (N_27775,N_26877,N_24448);
or U27776 (N_27776,N_25362,N_24357);
xor U27777 (N_27777,N_24403,N_24568);
and U27778 (N_27778,N_24282,N_25429);
or U27779 (N_27779,N_26120,N_26097);
or U27780 (N_27780,N_26414,N_24175);
nand U27781 (N_27781,N_25509,N_24688);
and U27782 (N_27782,N_24221,N_25972);
or U27783 (N_27783,N_24799,N_26458);
nor U27784 (N_27784,N_25054,N_25089);
nand U27785 (N_27785,N_26381,N_26662);
xnor U27786 (N_27786,N_24686,N_24546);
or U27787 (N_27787,N_26654,N_25440);
nor U27788 (N_27788,N_25655,N_24749);
xnor U27789 (N_27789,N_24079,N_25640);
nor U27790 (N_27790,N_25228,N_26071);
xor U27791 (N_27791,N_25971,N_26977);
and U27792 (N_27792,N_25512,N_24616);
xnor U27793 (N_27793,N_26567,N_24414);
and U27794 (N_27794,N_24800,N_26298);
nand U27795 (N_27795,N_26347,N_26294);
or U27796 (N_27796,N_25102,N_25721);
nand U27797 (N_27797,N_24002,N_25610);
nor U27798 (N_27798,N_26181,N_26083);
nand U27799 (N_27799,N_25807,N_24232);
nand U27800 (N_27800,N_26252,N_24813);
xnor U27801 (N_27801,N_25871,N_26184);
and U27802 (N_27802,N_26075,N_25148);
nor U27803 (N_27803,N_24632,N_24746);
xnor U27804 (N_27804,N_26644,N_24457);
or U27805 (N_27805,N_26319,N_26633);
nor U27806 (N_27806,N_25541,N_24645);
and U27807 (N_27807,N_25391,N_24346);
xor U27808 (N_27808,N_25989,N_26661);
nor U27809 (N_27809,N_24721,N_25153);
nor U27810 (N_27810,N_24484,N_24954);
xor U27811 (N_27811,N_26595,N_24203);
and U27812 (N_27812,N_26963,N_25146);
nor U27813 (N_27813,N_24020,N_26151);
and U27814 (N_27814,N_25699,N_24689);
nand U27815 (N_27815,N_26052,N_24153);
nor U27816 (N_27816,N_26093,N_24160);
and U27817 (N_27817,N_25227,N_26129);
and U27818 (N_27818,N_24627,N_24443);
xor U27819 (N_27819,N_25730,N_26024);
xnor U27820 (N_27820,N_25043,N_25303);
and U27821 (N_27821,N_25129,N_24067);
or U27822 (N_27822,N_26745,N_24187);
or U27823 (N_27823,N_24341,N_26673);
or U27824 (N_27824,N_24183,N_25821);
or U27825 (N_27825,N_26751,N_25843);
nand U27826 (N_27826,N_25598,N_24566);
nor U27827 (N_27827,N_26182,N_25344);
nand U27828 (N_27828,N_24732,N_25593);
nand U27829 (N_27829,N_25856,N_26463);
xnor U27830 (N_27830,N_24265,N_24076);
or U27831 (N_27831,N_25936,N_26321);
nand U27832 (N_27832,N_26442,N_26375);
or U27833 (N_27833,N_25329,N_24629);
and U27834 (N_27834,N_24920,N_24419);
and U27835 (N_27835,N_26122,N_24940);
and U27836 (N_27836,N_26460,N_24188);
and U27837 (N_27837,N_25109,N_26666);
nor U27838 (N_27838,N_25465,N_25794);
or U27839 (N_27839,N_24611,N_26649);
or U27840 (N_27840,N_26284,N_25716);
or U27841 (N_27841,N_26826,N_24595);
or U27842 (N_27842,N_25849,N_24219);
nor U27843 (N_27843,N_26076,N_24250);
or U27844 (N_27844,N_26430,N_26479);
and U27845 (N_27845,N_25142,N_26417);
nand U27846 (N_27846,N_26974,N_24275);
and U27847 (N_27847,N_25188,N_24136);
and U27848 (N_27848,N_26108,N_26497);
xor U27849 (N_27849,N_24281,N_24826);
xor U27850 (N_27850,N_24727,N_26187);
xor U27851 (N_27851,N_24128,N_25360);
nand U27852 (N_27852,N_25624,N_25515);
nand U27853 (N_27853,N_24587,N_26010);
and U27854 (N_27854,N_25769,N_24865);
nor U27855 (N_27855,N_26452,N_25086);
nor U27856 (N_27856,N_24808,N_26521);
or U27857 (N_27857,N_25482,N_25984);
and U27858 (N_27858,N_24737,N_25840);
nor U27859 (N_27859,N_24819,N_25718);
nor U27860 (N_27860,N_25288,N_25833);
xor U27861 (N_27861,N_25261,N_26733);
or U27862 (N_27862,N_25268,N_25058);
and U27863 (N_27863,N_24040,N_24601);
nand U27864 (N_27864,N_26306,N_26307);
or U27865 (N_27865,N_25024,N_24982);
or U27866 (N_27866,N_26907,N_26853);
nand U27867 (N_27867,N_25471,N_26851);
or U27868 (N_27868,N_26003,N_24470);
and U27869 (N_27869,N_25953,N_26735);
or U27870 (N_27870,N_26959,N_25152);
nor U27871 (N_27871,N_25379,N_24146);
nand U27872 (N_27872,N_25958,N_25274);
nand U27873 (N_27873,N_25248,N_25155);
and U27874 (N_27874,N_25306,N_26767);
nor U27875 (N_27875,N_26532,N_25586);
nand U27876 (N_27876,N_26335,N_24593);
and U27877 (N_27877,N_26220,N_24212);
or U27878 (N_27878,N_26277,N_24590);
and U27879 (N_27879,N_26040,N_25200);
xnor U27880 (N_27880,N_26601,N_24654);
xnor U27881 (N_27881,N_26180,N_26771);
nor U27882 (N_27882,N_25649,N_26285);
and U27883 (N_27883,N_24583,N_24655);
and U27884 (N_27884,N_24597,N_25862);
or U27885 (N_27885,N_26585,N_24047);
and U27886 (N_27886,N_25372,N_24726);
or U27887 (N_27887,N_25450,N_25881);
and U27888 (N_27888,N_24683,N_26726);
nand U27889 (N_27889,N_24885,N_24184);
or U27890 (N_27890,N_24515,N_26539);
or U27891 (N_27891,N_25017,N_25204);
nand U27892 (N_27892,N_25093,N_24909);
nand U27893 (N_27893,N_26831,N_25671);
and U27894 (N_27894,N_25033,N_24615);
nor U27895 (N_27895,N_26613,N_26287);
xnor U27896 (N_27896,N_26237,N_26537);
and U27897 (N_27897,N_24912,N_24573);
or U27898 (N_27898,N_25866,N_24456);
nand U27899 (N_27899,N_25497,N_24538);
xor U27900 (N_27900,N_26441,N_24119);
xor U27901 (N_27901,N_26472,N_25717);
nand U27902 (N_27902,N_25653,N_25371);
nand U27903 (N_27903,N_26918,N_25066);
nor U27904 (N_27904,N_24778,N_25369);
and U27905 (N_27905,N_24606,N_25577);
and U27906 (N_27906,N_26746,N_26652);
nand U27907 (N_27907,N_26092,N_25563);
nand U27908 (N_27908,N_25036,N_24633);
and U27909 (N_27909,N_26324,N_25540);
nor U27910 (N_27910,N_24013,N_25743);
nor U27911 (N_27911,N_24977,N_25193);
and U27912 (N_27912,N_25245,N_26401);
nand U27913 (N_27913,N_24501,N_26429);
or U27914 (N_27914,N_26348,N_26840);
nand U27915 (N_27915,N_24098,N_26041);
nand U27916 (N_27916,N_24624,N_24465);
or U27917 (N_27917,N_25050,N_24488);
xnor U27918 (N_27918,N_24924,N_25183);
xor U27919 (N_27919,N_25621,N_24048);
nor U27920 (N_27920,N_26388,N_25314);
nor U27921 (N_27921,N_26845,N_24951);
nor U27922 (N_27922,N_24173,N_24375);
xor U27923 (N_27923,N_25212,N_24576);
nand U27924 (N_27924,N_26806,N_24423);
nor U27925 (N_27925,N_24777,N_25741);
and U27926 (N_27926,N_24542,N_24126);
or U27927 (N_27927,N_26377,N_26967);
nand U27928 (N_27928,N_24652,N_25119);
or U27929 (N_27929,N_24008,N_26246);
and U27930 (N_27930,N_25680,N_26095);
nand U27931 (N_27931,N_24216,N_24091);
nand U27932 (N_27932,N_26169,N_24801);
and U27933 (N_27933,N_26510,N_25084);
and U27934 (N_27934,N_25224,N_26194);
nor U27935 (N_27935,N_26939,N_24750);
xnor U27936 (N_27936,N_24931,N_26197);
xor U27937 (N_27937,N_24544,N_26912);
xor U27938 (N_27938,N_24083,N_26687);
xnor U27939 (N_27939,N_26725,N_24863);
xnor U27940 (N_27940,N_25111,N_26055);
or U27941 (N_27941,N_25795,N_24278);
xnor U27942 (N_27942,N_24243,N_25165);
or U27943 (N_27943,N_24336,N_26467);
nor U27944 (N_27944,N_25527,N_24044);
nand U27945 (N_27945,N_24713,N_26223);
or U27946 (N_27946,N_24461,N_26427);
or U27947 (N_27947,N_25933,N_24948);
nand U27948 (N_27948,N_25087,N_24812);
nor U27949 (N_27949,N_25069,N_24177);
xnor U27950 (N_27950,N_25987,N_25880);
nand U27951 (N_27951,N_26581,N_24651);
xor U27952 (N_27952,N_25917,N_25216);
or U27953 (N_27953,N_25757,N_24992);
and U27954 (N_27954,N_24496,N_24640);
xor U27955 (N_27955,N_26415,N_25767);
xor U27956 (N_27956,N_24578,N_26934);
nand U27957 (N_27957,N_25742,N_24171);
or U27958 (N_27958,N_25920,N_24460);
or U27959 (N_27959,N_24968,N_26293);
nand U27960 (N_27960,N_25399,N_26145);
nor U27961 (N_27961,N_24194,N_26492);
or U27962 (N_27962,N_24650,N_26305);
xnor U27963 (N_27963,N_25941,N_24561);
nand U27964 (N_27964,N_24594,N_25443);
nand U27965 (N_27965,N_25402,N_25168);
or U27966 (N_27966,N_25970,N_24297);
nand U27967 (N_27967,N_24831,N_24163);
nor U27968 (N_27968,N_25045,N_25333);
and U27969 (N_27969,N_24888,N_25467);
and U27970 (N_27970,N_24535,N_25100);
xor U27971 (N_27971,N_26077,N_26079);
nand U27972 (N_27972,N_26166,N_24567);
or U27973 (N_27973,N_25056,N_24528);
and U27974 (N_27974,N_26825,N_25460);
nor U27975 (N_27975,N_26766,N_24182);
xnor U27976 (N_27976,N_25277,N_24399);
or U27977 (N_27977,N_25607,N_25103);
xor U27978 (N_27978,N_24200,N_25441);
and U27979 (N_27979,N_25672,N_26057);
xnor U27980 (N_27980,N_25230,N_25796);
nor U27981 (N_27981,N_26642,N_26450);
nand U27982 (N_27982,N_24631,N_26850);
and U27983 (N_27983,N_24148,N_25363);
nand U27984 (N_27984,N_25040,N_25202);
and U27985 (N_27985,N_25173,N_24438);
xnor U27986 (N_27986,N_24207,N_26927);
and U27987 (N_27987,N_25590,N_24881);
nand U27988 (N_27988,N_24998,N_26060);
nand U27989 (N_27989,N_24114,N_25517);
xnor U27990 (N_27990,N_25013,N_25079);
nand U27991 (N_27991,N_26438,N_26901);
xnor U27992 (N_27992,N_26280,N_26346);
nand U27993 (N_27993,N_24356,N_26171);
nor U27994 (N_27994,N_25409,N_25542);
nand U27995 (N_27995,N_26102,N_24214);
nor U27996 (N_27996,N_26042,N_24554);
nand U27997 (N_27997,N_24500,N_24444);
and U27998 (N_27998,N_26360,N_24548);
xor U27999 (N_27999,N_26478,N_24541);
and U28000 (N_28000,N_26370,N_25485);
xnor U28001 (N_28001,N_24859,N_25367);
nor U28002 (N_28002,N_26046,N_25149);
nor U28003 (N_28003,N_26628,N_24851);
nand U28004 (N_28004,N_26578,N_25580);
and U28005 (N_28005,N_24434,N_24512);
nand U28006 (N_28006,N_25981,N_24701);
nor U28007 (N_28007,N_25954,N_26922);
nor U28008 (N_28008,N_26890,N_26355);
nand U28009 (N_28009,N_24010,N_26712);
nor U28010 (N_28010,N_24682,N_24274);
nand U28011 (N_28011,N_24872,N_24066);
nand U28012 (N_28012,N_24782,N_25676);
nand U28013 (N_28013,N_24264,N_26536);
nor U28014 (N_28014,N_24858,N_25213);
nand U28015 (N_28015,N_25595,N_24486);
nor U28016 (N_28016,N_24054,N_24947);
nor U28017 (N_28017,N_24722,N_26148);
xnor U28018 (N_28018,N_24828,N_26062);
or U28019 (N_28019,N_24918,N_26803);
and U28020 (N_28020,N_24814,N_26422);
nand U28021 (N_28021,N_24266,N_25949);
and U28022 (N_28022,N_24696,N_25357);
or U28023 (N_28023,N_26813,N_26402);
nand U28024 (N_28024,N_26573,N_26698);
nand U28025 (N_28025,N_26688,N_26639);
nand U28026 (N_28026,N_25374,N_26038);
nor U28027 (N_28027,N_26903,N_24186);
nor U28028 (N_28028,N_25226,N_24823);
nor U28029 (N_28029,N_26378,N_26471);
xor U28030 (N_28030,N_25386,N_26480);
and U28031 (N_28031,N_24317,N_25945);
or U28032 (N_28032,N_26025,N_26711);
nor U28033 (N_28033,N_25790,N_25406);
xor U28034 (N_28034,N_26805,N_26032);
nor U28035 (N_28035,N_24441,N_26888);
nand U28036 (N_28036,N_25571,N_25682);
nor U28037 (N_28037,N_24684,N_26437);
and U28038 (N_28038,N_24271,N_25334);
nand U28039 (N_28039,N_26327,N_24015);
xor U28040 (N_28040,N_24504,N_24225);
and U28041 (N_28041,N_24552,N_26738);
or U28042 (N_28042,N_25284,N_25731);
or U28043 (N_28043,N_24636,N_26213);
xor U28044 (N_28044,N_26088,N_25458);
xnor U28045 (N_28045,N_24678,N_26050);
and U28046 (N_28046,N_25546,N_24199);
and U28047 (N_28047,N_26192,N_24657);
or U28048 (N_28048,N_25002,N_25195);
and U28049 (N_28049,N_24715,N_26935);
nor U28050 (N_28050,N_25256,N_25864);
nand U28051 (N_28051,N_24172,N_24493);
nand U28052 (N_28052,N_24110,N_25338);
nand U28053 (N_28053,N_26218,N_25582);
nand U28054 (N_28054,N_26086,N_25425);
or U28055 (N_28055,N_26937,N_24255);
and U28056 (N_28056,N_25688,N_25003);
or U28057 (N_28057,N_26770,N_24034);
nand U28058 (N_28058,N_24242,N_25793);
or U28059 (N_28059,N_25977,N_24467);
xnor U28060 (N_28060,N_25578,N_26518);
xnor U28061 (N_28061,N_25296,N_24997);
and U28062 (N_28062,N_26225,N_26830);
nor U28063 (N_28063,N_25151,N_25853);
xnor U28064 (N_28064,N_24967,N_24159);
or U28065 (N_28065,N_25778,N_24084);
xor U28066 (N_28066,N_25208,N_25570);
xnor U28067 (N_28067,N_25448,N_25346);
xor U28068 (N_28068,N_26713,N_25519);
or U28069 (N_28069,N_26541,N_26589);
or U28070 (N_28070,N_25179,N_25162);
nor U28071 (N_28071,N_26423,N_25551);
nand U28072 (N_28072,N_26511,N_24431);
and U28073 (N_28073,N_24490,N_26190);
and U28074 (N_28074,N_24379,N_24280);
nand U28075 (N_28075,N_24919,N_25548);
nor U28076 (N_28076,N_26599,N_25231);
nand U28077 (N_28077,N_24739,N_25711);
nor U28078 (N_28078,N_26600,N_25082);
xor U28079 (N_28079,N_24502,N_26217);
nor U28080 (N_28080,N_24827,N_24330);
xnor U28081 (N_28081,N_24603,N_25078);
xor U28082 (N_28082,N_24818,N_25124);
xor U28083 (N_28083,N_26296,N_24384);
xor U28084 (N_28084,N_26999,N_25126);
nor U28085 (N_28085,N_24145,N_26542);
xor U28086 (N_28086,N_24104,N_25576);
nand U28087 (N_28087,N_26186,N_26236);
nand U28088 (N_28088,N_26433,N_26933);
nor U28089 (N_28089,N_26658,N_24115);
or U28090 (N_28090,N_25703,N_24842);
nand U28091 (N_28091,N_25487,N_25965);
xnor U28092 (N_28092,N_26354,N_24984);
xnor U28093 (N_28093,N_24718,N_24005);
nand U28094 (N_28094,N_25738,N_25479);
and U28095 (N_28095,N_24296,N_24003);
nand U28096 (N_28096,N_26408,N_26435);
xnor U28097 (N_28097,N_24559,N_24150);
or U28098 (N_28098,N_26629,N_26461);
nor U28099 (N_28099,N_24116,N_26727);
nor U28100 (N_28100,N_26790,N_24481);
xnor U28101 (N_28101,N_25141,N_26149);
nor U28102 (N_28102,N_25172,N_24795);
xor U28103 (N_28103,N_25930,N_26697);
nor U28104 (N_28104,N_25063,N_25583);
nor U28105 (N_28105,N_25154,N_24893);
and U28106 (N_28106,N_26328,N_25792);
nor U28107 (N_28107,N_24702,N_26657);
or U28108 (N_28108,N_24508,N_25501);
nor U28109 (N_28109,N_26481,N_25016);
or U28110 (N_28110,N_24140,N_26214);
nor U28111 (N_28111,N_24263,N_24220);
nand U28112 (N_28112,N_24599,N_24562);
nor U28113 (N_28113,N_26862,N_26103);
nand U28114 (N_28114,N_26794,N_24138);
nand U28115 (N_28115,N_26373,N_26729);
or U28116 (N_28116,N_26783,N_26445);
xnor U28117 (N_28117,N_24990,N_24871);
nor U28118 (N_28118,N_26720,N_24299);
nand U28119 (N_28119,N_24070,N_25222);
nor U28120 (N_28120,N_26222,N_25106);
and U28121 (N_28121,N_26653,N_24584);
xnor U28122 (N_28122,N_25370,N_25161);
xnor U28123 (N_28123,N_24306,N_25895);
nor U28124 (N_28124,N_25823,N_26531);
xnor U28125 (N_28125,N_25574,N_26337);
nand U28126 (N_28126,N_26299,N_26568);
nor U28127 (N_28127,N_24230,N_24401);
and U28128 (N_28128,N_24798,N_24425);
and U28129 (N_28129,N_25368,N_25258);
or U28130 (N_28130,N_26762,N_25136);
xor U28131 (N_28131,N_24279,N_25211);
nand U28132 (N_28132,N_26063,N_25498);
or U28133 (N_28133,N_24520,N_25581);
and U28134 (N_28134,N_24326,N_26363);
nand U28135 (N_28135,N_24497,N_25269);
or U28136 (N_28136,N_26648,N_24149);
xnor U28137 (N_28137,N_26451,N_24742);
nand U28138 (N_28138,N_25654,N_24815);
xnor U28139 (N_28139,N_25413,N_24821);
or U28140 (N_28140,N_26051,N_25646);
xnor U28141 (N_28141,N_24023,N_24185);
and U28142 (N_28142,N_26178,N_25506);
or U28143 (N_28143,N_24693,N_26474);
nand U28144 (N_28144,N_24887,N_26426);
xor U28145 (N_28145,N_25473,N_25276);
and U28146 (N_28146,N_25326,N_24035);
nand U28147 (N_28147,N_26577,N_26875);
xnor U28148 (N_28148,N_26029,N_25645);
or U28149 (N_28149,N_24029,N_24580);
and U28150 (N_28150,N_25784,N_26352);
and U28151 (N_28151,N_26141,N_26270);
nand U28152 (N_28152,N_24673,N_25292);
or U28153 (N_28153,N_25921,N_26395);
nor U28154 (N_28154,N_26681,N_25697);
xnor U28155 (N_28155,N_26359,N_24765);
nor U28156 (N_28156,N_26982,N_25809);
nand U28157 (N_28157,N_26544,N_26886);
nor U28158 (N_28158,N_25573,N_25415);
and U28159 (N_28159,N_24963,N_26708);
nor U28160 (N_28160,N_26757,N_24816);
xor U28161 (N_28161,N_26547,N_26211);
or U28162 (N_28162,N_24349,N_26731);
and U28163 (N_28163,N_24017,N_26622);
nand U28164 (N_28164,N_25539,N_24210);
xor U28165 (N_28165,N_26462,N_26551);
and U28166 (N_28166,N_24121,N_25349);
xnor U28167 (N_28167,N_24832,N_26253);
and U28168 (N_28168,N_25072,N_25723);
or U28169 (N_28169,N_24874,N_25669);
xor U28170 (N_28170,N_24760,N_25572);
nor U28171 (N_28171,N_25786,N_26380);
nor U28172 (N_28172,N_24656,N_25782);
or U28173 (N_28173,N_24256,N_26509);
or U28174 (N_28174,N_24377,N_26928);
and U28175 (N_28175,N_25290,N_24946);
nand U28176 (N_28176,N_24432,N_26208);
or U28177 (N_28177,N_24482,N_25875);
nand U28178 (N_28178,N_26970,N_25191);
and U28179 (N_28179,N_24096,N_24779);
or U28180 (N_28180,N_25345,N_25552);
or U28181 (N_28181,N_25560,N_26684);
or U28182 (N_28182,N_24692,N_24714);
xor U28183 (N_28183,N_24910,N_24572);
xnor U28184 (N_28184,N_26504,N_26404);
and U28185 (N_28185,N_25830,N_24180);
nor U28186 (N_28186,N_26014,N_25806);
nor U28187 (N_28187,N_25740,N_25365);
or U28188 (N_28188,N_24053,N_25378);
nor U28189 (N_28189,N_25382,N_26915);
nor U28190 (N_28190,N_25912,N_26189);
nor U28191 (N_28191,N_24878,N_24890);
xnor U28192 (N_28192,N_24707,N_24740);
nand U28193 (N_28193,N_26885,N_25613);
and U28194 (N_28194,N_26202,N_26476);
or U28195 (N_28195,N_24407,N_25436);
xnor U28196 (N_28196,N_25489,N_24944);
xnor U28197 (N_28197,N_26022,N_26535);
or U28198 (N_28198,N_26150,N_26774);
nand U28199 (N_28199,N_26980,N_25818);
nand U28200 (N_28200,N_24545,N_24012);
xnor U28201 (N_28201,N_26736,N_25813);
or U28202 (N_28202,N_24855,N_25664);
or U28203 (N_28203,N_25005,N_25075);
nor U28204 (N_28204,N_26656,N_25691);
or U28205 (N_28205,N_26695,N_26855);
and U28206 (N_28206,N_24039,N_24202);
nor U28207 (N_28207,N_26085,N_26815);
and U28208 (N_28208,N_24109,N_24965);
nor U28209 (N_28209,N_26204,N_25137);
or U28210 (N_28210,N_25237,N_25238);
xor U28211 (N_28211,N_26870,N_26791);
xor U28212 (N_28212,N_25514,N_26714);
or U28213 (N_28213,N_24637,N_24733);
nor U28214 (N_28214,N_26066,N_26098);
and U28215 (N_28215,N_25732,N_24943);
xor U28216 (N_28216,N_25342,N_25756);
and U28217 (N_28217,N_26556,N_25518);
xnor U28218 (N_28218,N_25667,N_26637);
and U28219 (N_28219,N_24396,N_26776);
and U28220 (N_28220,N_25006,N_26090);
xnor U28221 (N_28221,N_26310,N_26081);
xor U28222 (N_28222,N_25065,N_26867);
or U28223 (N_28223,N_26976,N_24094);
and U28224 (N_28224,N_24847,N_26163);
nor U28225 (N_28225,N_25034,N_24428);
nand U28226 (N_28226,N_24609,N_24712);
nor U28227 (N_28227,N_26692,N_25998);
nor U28228 (N_28228,N_25526,N_24769);
or U28229 (N_28229,N_25160,N_26860);
xnor U28230 (N_28230,N_25687,N_25834);
nand U28231 (N_28231,N_26201,N_24332);
nand U28232 (N_28232,N_26245,N_26742);
xnor U28233 (N_28233,N_25847,N_25857);
nor U28234 (N_28234,N_25869,N_26368);
or U28235 (N_28235,N_24994,N_25038);
and U28236 (N_28236,N_26266,N_24550);
and U28237 (N_28237,N_24283,N_25848);
or U28238 (N_28238,N_26744,N_26508);
nor U28239 (N_28239,N_26865,N_25073);
nand U28240 (N_28240,N_26899,N_24204);
nor U28241 (N_28241,N_25739,N_25690);
xor U28242 (N_28242,N_26587,N_24155);
or U28243 (N_28243,N_24840,N_25852);
nand U28244 (N_28244,N_24621,N_26300);
and U28245 (N_28245,N_26627,N_25628);
nand U28246 (N_28246,N_25315,N_26994);
or U28247 (N_28247,N_26209,N_25698);
or U28248 (N_28248,N_25812,N_26495);
and U28249 (N_28249,N_25923,N_26118);
or U28250 (N_28250,N_24426,N_25964);
or U28251 (N_28251,N_24790,N_25865);
nor U28252 (N_28252,N_24380,N_26810);
nand U28253 (N_28253,N_26487,N_26807);
nor U28254 (N_28254,N_26871,N_26778);
nand U28255 (N_28255,N_26679,N_25353);
nor U28256 (N_28256,N_25456,N_26690);
nor U28257 (N_28257,N_25336,N_24108);
nand U28258 (N_28258,N_25939,N_25384);
xnor U28259 (N_28259,N_24602,N_25882);
xor U28260 (N_28260,N_24433,N_26137);
nor U28261 (N_28261,N_24916,N_25090);
nor U28262 (N_28262,N_25845,N_25785);
or U28263 (N_28263,N_25637,N_25710);
nor U28264 (N_28264,N_26138,N_25819);
nand U28265 (N_28265,N_26009,N_26528);
nor U28266 (N_28266,N_25244,N_25622);
and U28267 (N_28267,N_24258,N_24547);
nor U28268 (N_28268,N_25658,N_24162);
and U28269 (N_28269,N_25031,N_25135);
nor U28270 (N_28270,N_25899,N_24941);
or U28271 (N_28271,N_24447,N_24937);
nand U28272 (N_28272,N_25332,N_26134);
or U28273 (N_28273,N_25381,N_26121);
xor U28274 (N_28274,N_26739,N_25071);
xor U28275 (N_28275,N_25712,N_24915);
or U28276 (N_28276,N_24313,N_24285);
nand U28277 (N_28277,N_26839,N_26696);
and U28278 (N_28278,N_26164,N_24397);
nor U28279 (N_28279,N_24996,N_25735);
or U28280 (N_28280,N_26247,N_24773);
nand U28281 (N_28281,N_26953,N_24524);
xnor U28282 (N_28282,N_25064,N_26786);
xnor U28283 (N_28283,N_26905,N_25614);
nor U28284 (N_28284,N_25113,N_25907);
xnor U28285 (N_28285,N_24224,N_25171);
nor U28286 (N_28286,N_24416,N_24089);
and U28287 (N_28287,N_26339,N_25632);
and U28288 (N_28288,N_26938,N_26325);
and U28289 (N_28289,N_24252,N_24161);
xor U28290 (N_28290,N_24891,N_25986);
and U28291 (N_28291,N_26128,N_24334);
and U28292 (N_28292,N_25393,N_26667);
nand U28293 (N_28293,N_26709,N_24389);
or U28294 (N_28294,N_26295,N_24295);
nand U28295 (N_28295,N_24050,N_25131);
or U28296 (N_28296,N_24059,N_25841);
or U28297 (N_28297,N_24302,N_24744);
nor U28298 (N_28298,N_25910,N_25255);
nand U28299 (N_28299,N_25335,N_24764);
or U28300 (N_28300,N_26061,N_24730);
and U28301 (N_28301,N_25736,N_25851);
and U28302 (N_28302,N_26332,N_24009);
nor U28303 (N_28303,N_24316,N_24735);
nand U28304 (N_28304,N_26385,N_25139);
xor U28305 (N_28305,N_25420,N_26154);
xnor U28306 (N_28306,N_24942,N_25022);
nand U28307 (N_28307,N_25963,N_25055);
nand U28308 (N_28308,N_26718,N_24575);
or U28309 (N_28309,N_26533,N_26345);
xnor U28310 (N_28310,N_26990,N_26070);
nor U28311 (N_28311,N_25772,N_25455);
nand U28312 (N_28312,N_26195,N_24037);
or U28313 (N_28313,N_24127,N_26699);
and U28314 (N_28314,N_25592,N_26772);
nor U28315 (N_28315,N_26228,N_24728);
xnor U28316 (N_28316,N_25558,N_26945);
nor U28317 (N_28317,N_25240,N_26520);
nor U28318 (N_28318,N_24197,N_24605);
nand U28319 (N_28319,N_25328,N_26261);
nand U28320 (N_28320,N_25094,N_24557);
nand U28321 (N_28321,N_26398,N_25286);
xnor U28322 (N_28322,N_25019,N_26314);
xor U28323 (N_28323,N_26198,N_25053);
nand U28324 (N_28324,N_25265,N_24474);
or U28325 (N_28325,N_25659,N_26917);
or U28326 (N_28326,N_24360,N_25808);
or U28327 (N_28327,N_24420,N_24805);
nand U28328 (N_28328,N_25499,N_24137);
and U28329 (N_28329,N_25300,N_26386);
or U28330 (N_28330,N_26943,N_25505);
xnor U28331 (N_28331,N_25387,N_26466);
xor U28332 (N_28332,N_25726,N_26923);
nor U28333 (N_28333,N_24241,N_25444);
nor U28334 (N_28334,N_25800,N_25870);
xnor U28335 (N_28335,N_24424,N_25403);
xnor U28336 (N_28336,N_26524,N_25484);
xor U28337 (N_28337,N_25915,N_26226);
xnor U28338 (N_28338,N_26920,N_24665);
nor U28339 (N_28339,N_24646,N_24475);
xor U28340 (N_28340,N_25983,N_25854);
or U28341 (N_28341,N_25922,N_25007);
nor U28342 (N_28342,N_24235,N_25937);
nor U28343 (N_28343,N_24700,N_24932);
xnor U28344 (N_28344,N_24643,N_25203);
nand U28345 (N_28345,N_26563,N_25665);
nand U28346 (N_28346,N_24370,N_24933);
xnor U28347 (N_28347,N_26799,N_25842);
nor U28348 (N_28348,N_26896,N_26594);
nand U28349 (N_28349,N_24697,N_26490);
xor U28350 (N_28350,N_24321,N_24999);
nand U28351 (N_28351,N_26784,N_24894);
nor U28352 (N_28352,N_24343,N_25714);
and U28353 (N_28353,N_24970,N_26931);
nor U28354 (N_28354,N_26227,N_26591);
or U28355 (N_28355,N_26722,N_24784);
xor U28356 (N_28356,N_26082,N_24877);
and U28357 (N_28357,N_25088,N_24228);
nor U28358 (N_28358,N_24844,N_26376);
nor U28359 (N_28359,N_25838,N_26740);
nor U28360 (N_28360,N_25603,N_25544);
or U28361 (N_28361,N_26900,N_25516);
and U28362 (N_28362,N_24563,N_24526);
nor U28363 (N_28363,N_24165,N_26804);
nand U28364 (N_28364,N_25389,N_24719);
xnor U28365 (N_28365,N_25156,N_24648);
nand U28366 (N_28366,N_25674,N_24706);
nor U28367 (N_28367,N_26906,N_25273);
nand U28368 (N_28368,N_25397,N_25433);
nand U28369 (N_28369,N_25380,N_26037);
nor U28370 (N_28370,N_25623,N_26607);
nand U28371 (N_28371,N_25115,N_25001);
xor U28372 (N_28372,N_25791,N_25282);
xor U28373 (N_28373,N_26240,N_26988);
xnor U28374 (N_28374,N_25835,N_24480);
nor U28375 (N_28375,N_25513,N_24129);
or U28376 (N_28376,N_25095,N_25940);
and U28377 (N_28377,N_24536,N_24653);
nor U28378 (N_28378,N_24478,N_26672);
and U28379 (N_28379,N_24262,N_26309);
nand U28380 (N_28380,N_26741,N_26623);
nand U28381 (N_28381,N_24368,N_25733);
nor U28382 (N_28382,N_26854,N_25695);
nand U28383 (N_28383,N_26428,N_24406);
or U28384 (N_28384,N_24445,N_24312);
or U28385 (N_28385,N_26160,N_25824);
nand U28386 (N_28386,N_25000,N_25178);
or U28387 (N_28387,N_24342,N_26045);
or U28388 (N_28388,N_24644,N_24102);
or U28389 (N_28389,N_24093,N_25271);
or U28390 (N_28390,N_26597,N_25175);
and U28391 (N_28391,N_24585,N_26617);
and U28392 (N_28392,N_24717,N_25787);
nand U28393 (N_28393,N_25474,N_24135);
and U28394 (N_28394,N_25307,N_26333);
nor U28395 (N_28395,N_24957,N_26956);
nor U28396 (N_28396,N_24347,N_26183);
or U28397 (N_28397,N_25575,N_26926);
nor U28398 (N_28398,N_25438,N_26640);
nor U28399 (N_28399,N_25556,N_24507);
nor U28400 (N_28400,N_24839,N_24803);
and U28401 (N_28401,N_26281,N_24776);
xnor U28402 (N_28402,N_26114,N_26811);
nor U28403 (N_28403,N_24852,N_25564);
or U28404 (N_28404,N_26065,N_24290);
or U28405 (N_28405,N_24691,N_25629);
nor U28406 (N_28406,N_25125,N_24014);
xnor U28407 (N_28407,N_24820,N_26609);
or U28408 (N_28408,N_25011,N_24259);
nand U28409 (N_28409,N_26100,N_24671);
xor U28410 (N_28410,N_26763,N_26320);
and U28411 (N_28411,N_26278,N_24141);
or U28412 (N_28412,N_26136,N_26446);
xnor U28413 (N_28413,N_26468,N_26680);
nand U28414 (N_28414,N_25801,N_26576);
xnor U28415 (N_28415,N_26155,N_24870);
xor U28416 (N_28416,N_26023,N_25351);
and U28417 (N_28417,N_26073,N_24509);
or U28418 (N_28418,N_25419,N_26779);
or U28419 (N_28419,N_26288,N_26020);
and U28420 (N_28420,N_24570,N_26706);
nor U28421 (N_28421,N_26336,N_24168);
or U28422 (N_28422,N_24167,N_25074);
nand U28423 (N_28423,N_26643,N_25956);
nor U28424 (N_28424,N_24074,N_25480);
and U28425 (N_28425,N_25061,N_26331);
nand U28426 (N_28426,N_24830,N_24169);
nand U28427 (N_28427,N_25798,N_24030);
nor U28428 (N_28428,N_25737,N_25174);
or U28429 (N_28429,N_26419,N_24260);
nand U28430 (N_28430,N_24680,N_24195);
xor U28431 (N_28431,N_25709,N_26410);
nor U28432 (N_28432,N_26235,N_26621);
nand U28433 (N_28433,N_25549,N_24237);
nand U28434 (N_28434,N_25052,N_24964);
xnor U28435 (N_28435,N_26140,N_25159);
and U28436 (N_28436,N_26952,N_26701);
nand U28437 (N_28437,N_25700,N_24922);
nor U28438 (N_28438,N_25774,N_26021);
nor U28439 (N_28439,N_25325,N_25893);
xor U28440 (N_28440,N_24649,N_26177);
and U28441 (N_28441,N_24975,N_24395);
and U28442 (N_28442,N_25076,N_25008);
nand U28443 (N_28443,N_26785,N_25925);
or U28444 (N_28444,N_24873,N_26677);
xor U28445 (N_28445,N_24324,N_25395);
nand U28446 (N_28446,N_26313,N_25720);
nand U28447 (N_28447,N_26465,N_26099);
or U28448 (N_28448,N_24961,N_26822);
nand U28449 (N_28449,N_26080,N_24272);
xor U28450 (N_28450,N_26756,N_26016);
nand U28451 (N_28451,N_25884,N_24789);
nand U28452 (N_28452,N_25585,N_26880);
nor U28453 (N_28453,N_25009,N_26503);
nand U28454 (N_28454,N_24661,N_24625);
or U28455 (N_28455,N_24134,N_26889);
nand U28456 (N_28456,N_25634,N_24897);
and U28457 (N_28457,N_24662,N_26700);
nor U28458 (N_28458,N_25566,N_25114);
nor U28459 (N_28459,N_25826,N_25538);
and U28460 (N_28460,N_26909,N_24251);
xor U28461 (N_28461,N_24786,N_26116);
or U28462 (N_28462,N_26231,N_26561);
xor U28463 (N_28463,N_24105,N_26984);
nand U28464 (N_28464,N_24085,N_25424);
or U28465 (N_28465,N_25978,N_24596);
and U28466 (N_28466,N_26893,N_26139);
nand U28467 (N_28467,N_26206,N_24062);
and U28468 (N_28468,N_24100,N_26405);
or U28469 (N_28469,N_25262,N_24222);
nor U28470 (N_28470,N_24390,N_24503);
xnor U28471 (N_28471,N_26944,N_24986);
or U28472 (N_28472,N_26340,N_24864);
nand U28473 (N_28473,N_26379,N_24639);
and U28474 (N_28474,N_24006,N_24485);
xor U28475 (N_28475,N_26409,N_26796);
and U28476 (N_28476,N_25897,N_24804);
nor U28477 (N_28477,N_24293,N_25423);
nor U28478 (N_28478,N_26919,N_26764);
or U28479 (N_28479,N_25584,N_24446);
nand U28480 (N_28480,N_26604,N_24588);
and U28481 (N_28481,N_24622,N_24699);
xnor U28482 (N_28482,N_24257,N_25652);
nor U28483 (N_28483,N_26005,N_25060);
and U28484 (N_28484,N_24231,N_25158);
and U28485 (N_28485,N_26996,N_26924);
nor U28486 (N_28486,N_25067,N_24531);
nor U28487 (N_28487,N_25377,N_25410);
and U28488 (N_28488,N_26702,N_26489);
nor U28489 (N_28489,N_24051,N_26397);
nor U28490 (N_28490,N_24577,N_26951);
nand U28491 (N_28491,N_26371,N_24391);
xnor U28492 (N_28492,N_26047,N_25889);
or U28493 (N_28493,N_26119,N_26210);
or U28494 (N_28494,N_24936,N_25679);
or U28495 (N_28495,N_26949,N_25626);
nor U28496 (N_28496,N_24600,N_25535);
xor U28497 (N_28497,N_25719,N_26019);
and U28498 (N_28498,N_24903,N_26878);
xnor U28499 (N_28499,N_24288,N_25644);
or U28500 (N_28500,N_24985,N_25365);
and U28501 (N_28501,N_25663,N_26755);
and U28502 (N_28502,N_24502,N_24619);
or U28503 (N_28503,N_24907,N_25391);
and U28504 (N_28504,N_25947,N_25122);
and U28505 (N_28505,N_24709,N_26535);
nor U28506 (N_28506,N_24352,N_26334);
nand U28507 (N_28507,N_26340,N_26632);
xor U28508 (N_28508,N_25702,N_24337);
nor U28509 (N_28509,N_25392,N_26203);
or U28510 (N_28510,N_24078,N_24471);
or U28511 (N_28511,N_24894,N_24171);
xor U28512 (N_28512,N_25109,N_25930);
nand U28513 (N_28513,N_26154,N_25382);
xnor U28514 (N_28514,N_24024,N_26994);
or U28515 (N_28515,N_25884,N_25318);
nand U28516 (N_28516,N_24236,N_24578);
xor U28517 (N_28517,N_26737,N_26008);
nand U28518 (N_28518,N_25405,N_24248);
xor U28519 (N_28519,N_24954,N_26090);
and U28520 (N_28520,N_24023,N_26735);
or U28521 (N_28521,N_25685,N_25607);
nand U28522 (N_28522,N_25678,N_25369);
xor U28523 (N_28523,N_26209,N_25793);
or U28524 (N_28524,N_25560,N_25553);
nand U28525 (N_28525,N_25644,N_26045);
and U28526 (N_28526,N_25928,N_24782);
or U28527 (N_28527,N_24410,N_26323);
nor U28528 (N_28528,N_25093,N_26749);
xor U28529 (N_28529,N_25816,N_25227);
nor U28530 (N_28530,N_24285,N_24483);
nand U28531 (N_28531,N_26875,N_25240);
nor U28532 (N_28532,N_26327,N_24004);
nor U28533 (N_28533,N_25948,N_24790);
or U28534 (N_28534,N_25358,N_26296);
nand U28535 (N_28535,N_24622,N_25333);
xor U28536 (N_28536,N_24628,N_25136);
or U28537 (N_28537,N_25424,N_25491);
nor U28538 (N_28538,N_26079,N_26710);
or U28539 (N_28539,N_24843,N_24289);
nor U28540 (N_28540,N_25448,N_24725);
xnor U28541 (N_28541,N_26228,N_24850);
or U28542 (N_28542,N_24720,N_24933);
or U28543 (N_28543,N_24006,N_25000);
nor U28544 (N_28544,N_24432,N_25083);
xor U28545 (N_28545,N_24411,N_24823);
xor U28546 (N_28546,N_25055,N_26728);
and U28547 (N_28547,N_24885,N_24667);
xor U28548 (N_28548,N_25403,N_24003);
or U28549 (N_28549,N_26999,N_24523);
nor U28550 (N_28550,N_26915,N_25690);
nand U28551 (N_28551,N_26442,N_25652);
and U28552 (N_28552,N_26940,N_25925);
xnor U28553 (N_28553,N_24952,N_24478);
nand U28554 (N_28554,N_25593,N_24365);
nor U28555 (N_28555,N_24503,N_26254);
xor U28556 (N_28556,N_25633,N_24820);
or U28557 (N_28557,N_25977,N_25393);
or U28558 (N_28558,N_26143,N_24221);
nor U28559 (N_28559,N_24065,N_25833);
nand U28560 (N_28560,N_25159,N_24817);
nor U28561 (N_28561,N_25158,N_26472);
and U28562 (N_28562,N_25176,N_25072);
nand U28563 (N_28563,N_26038,N_24817);
and U28564 (N_28564,N_25545,N_25338);
and U28565 (N_28565,N_24428,N_26392);
and U28566 (N_28566,N_26868,N_26422);
and U28567 (N_28567,N_24614,N_26528);
nand U28568 (N_28568,N_25662,N_24127);
nor U28569 (N_28569,N_26145,N_26675);
or U28570 (N_28570,N_25796,N_26726);
and U28571 (N_28571,N_24515,N_24907);
nor U28572 (N_28572,N_24396,N_25317);
and U28573 (N_28573,N_26318,N_26067);
or U28574 (N_28574,N_26148,N_26152);
or U28575 (N_28575,N_26474,N_26197);
and U28576 (N_28576,N_26464,N_26498);
or U28577 (N_28577,N_26988,N_24768);
nor U28578 (N_28578,N_25361,N_25198);
or U28579 (N_28579,N_24734,N_26577);
or U28580 (N_28580,N_25744,N_26479);
and U28581 (N_28581,N_24622,N_26620);
nand U28582 (N_28582,N_26803,N_24908);
and U28583 (N_28583,N_25698,N_24222);
and U28584 (N_28584,N_26006,N_25580);
xnor U28585 (N_28585,N_25503,N_26123);
nor U28586 (N_28586,N_26186,N_25555);
xor U28587 (N_28587,N_24485,N_25971);
or U28588 (N_28588,N_25172,N_26247);
and U28589 (N_28589,N_26186,N_26478);
nand U28590 (N_28590,N_24873,N_26409);
or U28591 (N_28591,N_24504,N_24152);
or U28592 (N_28592,N_25177,N_25325);
and U28593 (N_28593,N_24122,N_24304);
and U28594 (N_28594,N_24362,N_26259);
xor U28595 (N_28595,N_24861,N_24451);
xnor U28596 (N_28596,N_26054,N_24913);
xnor U28597 (N_28597,N_26075,N_26542);
and U28598 (N_28598,N_24234,N_25172);
nor U28599 (N_28599,N_25765,N_26686);
xor U28600 (N_28600,N_26079,N_24894);
nor U28601 (N_28601,N_25177,N_26202);
nand U28602 (N_28602,N_24164,N_25004);
nor U28603 (N_28603,N_25363,N_26684);
xor U28604 (N_28604,N_26934,N_26767);
and U28605 (N_28605,N_26040,N_25939);
and U28606 (N_28606,N_24804,N_25979);
nor U28607 (N_28607,N_24522,N_25805);
xnor U28608 (N_28608,N_24808,N_25441);
and U28609 (N_28609,N_26598,N_24382);
nand U28610 (N_28610,N_26645,N_25831);
and U28611 (N_28611,N_25329,N_25585);
nor U28612 (N_28612,N_25874,N_24631);
nand U28613 (N_28613,N_26608,N_26446);
xnor U28614 (N_28614,N_24145,N_26097);
xor U28615 (N_28615,N_25765,N_24900);
nor U28616 (N_28616,N_26158,N_26853);
or U28617 (N_28617,N_26040,N_25546);
nand U28618 (N_28618,N_26313,N_25730);
nor U28619 (N_28619,N_26770,N_24568);
or U28620 (N_28620,N_26370,N_26349);
nor U28621 (N_28621,N_24610,N_26408);
nor U28622 (N_28622,N_26926,N_26499);
or U28623 (N_28623,N_26366,N_26698);
and U28624 (N_28624,N_25150,N_26278);
nand U28625 (N_28625,N_24489,N_26523);
and U28626 (N_28626,N_25697,N_25022);
and U28627 (N_28627,N_25867,N_25544);
xor U28628 (N_28628,N_24982,N_24607);
or U28629 (N_28629,N_24871,N_26794);
and U28630 (N_28630,N_25243,N_24371);
nand U28631 (N_28631,N_26806,N_24757);
nor U28632 (N_28632,N_25035,N_26763);
or U28633 (N_28633,N_26666,N_24022);
or U28634 (N_28634,N_25512,N_26624);
and U28635 (N_28635,N_24957,N_26011);
nor U28636 (N_28636,N_24472,N_25417);
and U28637 (N_28637,N_25512,N_24605);
xor U28638 (N_28638,N_26683,N_26088);
nand U28639 (N_28639,N_26761,N_25071);
or U28640 (N_28640,N_24893,N_25428);
nor U28641 (N_28641,N_24911,N_26866);
nand U28642 (N_28642,N_24922,N_24067);
nand U28643 (N_28643,N_26154,N_25845);
or U28644 (N_28644,N_26010,N_24196);
xnor U28645 (N_28645,N_26185,N_26768);
and U28646 (N_28646,N_26005,N_24266);
nor U28647 (N_28647,N_26594,N_25612);
or U28648 (N_28648,N_26118,N_26981);
nand U28649 (N_28649,N_25578,N_26590);
or U28650 (N_28650,N_25335,N_24585);
nor U28651 (N_28651,N_25863,N_26578);
nand U28652 (N_28652,N_26819,N_24712);
nor U28653 (N_28653,N_25996,N_24071);
or U28654 (N_28654,N_25667,N_26771);
nor U28655 (N_28655,N_25227,N_24346);
xnor U28656 (N_28656,N_26428,N_25397);
nor U28657 (N_28657,N_25617,N_26681);
or U28658 (N_28658,N_26523,N_24050);
nor U28659 (N_28659,N_24806,N_24083);
and U28660 (N_28660,N_24213,N_24025);
nor U28661 (N_28661,N_24178,N_24446);
or U28662 (N_28662,N_26049,N_24633);
nor U28663 (N_28663,N_26992,N_24471);
nor U28664 (N_28664,N_25664,N_24307);
or U28665 (N_28665,N_26965,N_24140);
or U28666 (N_28666,N_25051,N_24481);
nor U28667 (N_28667,N_26925,N_26068);
xnor U28668 (N_28668,N_24901,N_25509);
xor U28669 (N_28669,N_26456,N_24438);
or U28670 (N_28670,N_26584,N_24608);
or U28671 (N_28671,N_24420,N_24941);
nor U28672 (N_28672,N_25095,N_26541);
nand U28673 (N_28673,N_26077,N_25958);
nor U28674 (N_28674,N_25104,N_26413);
or U28675 (N_28675,N_25395,N_26268);
nor U28676 (N_28676,N_24845,N_25825);
nand U28677 (N_28677,N_25996,N_24062);
and U28678 (N_28678,N_26257,N_25192);
nor U28679 (N_28679,N_26815,N_25230);
and U28680 (N_28680,N_25297,N_26910);
nor U28681 (N_28681,N_26459,N_24708);
nand U28682 (N_28682,N_25747,N_25844);
xor U28683 (N_28683,N_24619,N_26132);
and U28684 (N_28684,N_26803,N_24692);
xor U28685 (N_28685,N_25614,N_26351);
nor U28686 (N_28686,N_26324,N_24696);
xnor U28687 (N_28687,N_26209,N_26863);
and U28688 (N_28688,N_25195,N_25600);
or U28689 (N_28689,N_25335,N_26426);
nand U28690 (N_28690,N_24430,N_26983);
nor U28691 (N_28691,N_25522,N_26685);
nor U28692 (N_28692,N_25471,N_24322);
or U28693 (N_28693,N_26249,N_24300);
and U28694 (N_28694,N_25229,N_25033);
xnor U28695 (N_28695,N_26191,N_24085);
xnor U28696 (N_28696,N_24748,N_24994);
xor U28697 (N_28697,N_24366,N_26866);
nor U28698 (N_28698,N_24480,N_25217);
and U28699 (N_28699,N_26226,N_26420);
and U28700 (N_28700,N_26127,N_26475);
nand U28701 (N_28701,N_24523,N_24452);
nor U28702 (N_28702,N_25958,N_26646);
and U28703 (N_28703,N_26113,N_26354);
xor U28704 (N_28704,N_26321,N_24777);
nor U28705 (N_28705,N_26611,N_24411);
or U28706 (N_28706,N_26850,N_26553);
or U28707 (N_28707,N_24727,N_26700);
and U28708 (N_28708,N_24636,N_26918);
nand U28709 (N_28709,N_26494,N_25872);
nor U28710 (N_28710,N_24056,N_24713);
or U28711 (N_28711,N_25114,N_25811);
nand U28712 (N_28712,N_24223,N_25621);
nand U28713 (N_28713,N_24175,N_25886);
xor U28714 (N_28714,N_24193,N_24443);
and U28715 (N_28715,N_25493,N_25679);
nand U28716 (N_28716,N_24613,N_26085);
nor U28717 (N_28717,N_26852,N_24186);
nand U28718 (N_28718,N_26407,N_26497);
xor U28719 (N_28719,N_26194,N_25177);
nor U28720 (N_28720,N_26358,N_25141);
xor U28721 (N_28721,N_24467,N_24028);
nor U28722 (N_28722,N_24591,N_26686);
nor U28723 (N_28723,N_26287,N_24565);
nor U28724 (N_28724,N_25878,N_26740);
xnor U28725 (N_28725,N_24497,N_26021);
nor U28726 (N_28726,N_24018,N_24308);
xnor U28727 (N_28727,N_25865,N_25712);
xor U28728 (N_28728,N_24226,N_24651);
xor U28729 (N_28729,N_24585,N_25249);
xnor U28730 (N_28730,N_24360,N_25620);
or U28731 (N_28731,N_25811,N_26181);
nand U28732 (N_28732,N_25466,N_26847);
nor U28733 (N_28733,N_24841,N_26270);
xnor U28734 (N_28734,N_25569,N_25128);
and U28735 (N_28735,N_24571,N_24906);
nor U28736 (N_28736,N_24073,N_24151);
nor U28737 (N_28737,N_26886,N_26030);
xnor U28738 (N_28738,N_26263,N_25066);
xor U28739 (N_28739,N_26763,N_25523);
xnor U28740 (N_28740,N_26951,N_24736);
nand U28741 (N_28741,N_26488,N_24698);
and U28742 (N_28742,N_25211,N_24540);
or U28743 (N_28743,N_25961,N_24603);
nor U28744 (N_28744,N_25808,N_25363);
or U28745 (N_28745,N_24579,N_26976);
nor U28746 (N_28746,N_24242,N_25309);
nor U28747 (N_28747,N_25218,N_26329);
xnor U28748 (N_28748,N_24993,N_24641);
xnor U28749 (N_28749,N_24420,N_26719);
nand U28750 (N_28750,N_24370,N_24970);
or U28751 (N_28751,N_26959,N_25612);
nand U28752 (N_28752,N_25987,N_25246);
and U28753 (N_28753,N_26748,N_24135);
or U28754 (N_28754,N_24001,N_25381);
nor U28755 (N_28755,N_25773,N_26758);
and U28756 (N_28756,N_26970,N_25887);
xnor U28757 (N_28757,N_26580,N_24735);
xnor U28758 (N_28758,N_26843,N_26970);
or U28759 (N_28759,N_25950,N_26004);
xnor U28760 (N_28760,N_25893,N_25524);
xor U28761 (N_28761,N_24667,N_24779);
and U28762 (N_28762,N_25492,N_26464);
xor U28763 (N_28763,N_24692,N_24495);
or U28764 (N_28764,N_25131,N_24805);
xnor U28765 (N_28765,N_24922,N_24258);
and U28766 (N_28766,N_25597,N_26228);
nor U28767 (N_28767,N_25165,N_24548);
or U28768 (N_28768,N_25260,N_25030);
nand U28769 (N_28769,N_24261,N_25229);
nor U28770 (N_28770,N_24839,N_25096);
nor U28771 (N_28771,N_25498,N_25493);
xor U28772 (N_28772,N_26007,N_25054);
xnor U28773 (N_28773,N_24166,N_26343);
and U28774 (N_28774,N_26648,N_25192);
nor U28775 (N_28775,N_26865,N_25383);
nor U28776 (N_28776,N_25123,N_24224);
or U28777 (N_28777,N_24454,N_26784);
xnor U28778 (N_28778,N_25103,N_25591);
nand U28779 (N_28779,N_25683,N_24896);
nor U28780 (N_28780,N_26752,N_25040);
nand U28781 (N_28781,N_26324,N_25377);
or U28782 (N_28782,N_25887,N_24763);
xor U28783 (N_28783,N_25793,N_26389);
xnor U28784 (N_28784,N_26518,N_24321);
nand U28785 (N_28785,N_26321,N_25312);
nor U28786 (N_28786,N_24299,N_24560);
nand U28787 (N_28787,N_24225,N_24633);
or U28788 (N_28788,N_25735,N_26166);
and U28789 (N_28789,N_25065,N_26525);
nand U28790 (N_28790,N_25796,N_24119);
nand U28791 (N_28791,N_26452,N_25091);
nand U28792 (N_28792,N_25737,N_25982);
or U28793 (N_28793,N_24933,N_25315);
or U28794 (N_28794,N_25815,N_24314);
nand U28795 (N_28795,N_25939,N_25133);
xor U28796 (N_28796,N_25628,N_26688);
or U28797 (N_28797,N_25557,N_25485);
or U28798 (N_28798,N_26874,N_24489);
or U28799 (N_28799,N_26122,N_25632);
xnor U28800 (N_28800,N_24458,N_25078);
nand U28801 (N_28801,N_26021,N_26142);
nand U28802 (N_28802,N_24811,N_25353);
xor U28803 (N_28803,N_24920,N_24868);
or U28804 (N_28804,N_24855,N_24472);
nor U28805 (N_28805,N_26486,N_25915);
xor U28806 (N_28806,N_26235,N_25171);
nand U28807 (N_28807,N_24179,N_26306);
xor U28808 (N_28808,N_24408,N_24160);
nor U28809 (N_28809,N_25013,N_26117);
nor U28810 (N_28810,N_25956,N_24809);
and U28811 (N_28811,N_26106,N_26701);
nand U28812 (N_28812,N_25106,N_26794);
nand U28813 (N_28813,N_24666,N_25942);
xnor U28814 (N_28814,N_26140,N_24182);
or U28815 (N_28815,N_24952,N_26103);
xor U28816 (N_28816,N_26443,N_25731);
nand U28817 (N_28817,N_24053,N_25581);
and U28818 (N_28818,N_26269,N_24050);
xnor U28819 (N_28819,N_26524,N_24467);
and U28820 (N_28820,N_24079,N_26783);
nor U28821 (N_28821,N_25737,N_24202);
nand U28822 (N_28822,N_24470,N_26604);
or U28823 (N_28823,N_26137,N_25860);
xor U28824 (N_28824,N_24157,N_24716);
nand U28825 (N_28825,N_26212,N_24375);
nor U28826 (N_28826,N_26850,N_26104);
nand U28827 (N_28827,N_26416,N_25451);
and U28828 (N_28828,N_26606,N_26670);
and U28829 (N_28829,N_24606,N_26833);
or U28830 (N_28830,N_25247,N_25042);
nor U28831 (N_28831,N_24690,N_26379);
nand U28832 (N_28832,N_25137,N_24195);
and U28833 (N_28833,N_25793,N_24844);
nand U28834 (N_28834,N_25090,N_24713);
or U28835 (N_28835,N_26029,N_24171);
nor U28836 (N_28836,N_25420,N_26267);
and U28837 (N_28837,N_24800,N_25384);
and U28838 (N_28838,N_24785,N_25934);
or U28839 (N_28839,N_26737,N_26929);
nand U28840 (N_28840,N_24510,N_24946);
or U28841 (N_28841,N_26732,N_24292);
xnor U28842 (N_28842,N_25414,N_26823);
nand U28843 (N_28843,N_26641,N_24527);
and U28844 (N_28844,N_26827,N_25968);
xor U28845 (N_28845,N_25555,N_26243);
nand U28846 (N_28846,N_26457,N_26594);
and U28847 (N_28847,N_25274,N_26008);
nor U28848 (N_28848,N_26178,N_24671);
nor U28849 (N_28849,N_24838,N_26194);
xor U28850 (N_28850,N_25921,N_24387);
and U28851 (N_28851,N_25116,N_26828);
nand U28852 (N_28852,N_24286,N_26911);
or U28853 (N_28853,N_25849,N_25777);
nor U28854 (N_28854,N_26515,N_25777);
and U28855 (N_28855,N_24949,N_25457);
nor U28856 (N_28856,N_25744,N_24231);
xnor U28857 (N_28857,N_24433,N_25054);
xnor U28858 (N_28858,N_25041,N_25936);
or U28859 (N_28859,N_25666,N_25904);
nor U28860 (N_28860,N_26409,N_24896);
nor U28861 (N_28861,N_26468,N_24668);
xor U28862 (N_28862,N_24969,N_25675);
or U28863 (N_28863,N_26041,N_25934);
or U28864 (N_28864,N_25201,N_24288);
xnor U28865 (N_28865,N_24719,N_24393);
xnor U28866 (N_28866,N_25470,N_26999);
xor U28867 (N_28867,N_26834,N_25481);
nor U28868 (N_28868,N_26405,N_24546);
nor U28869 (N_28869,N_24609,N_25461);
nand U28870 (N_28870,N_24361,N_24144);
or U28871 (N_28871,N_25030,N_25076);
xor U28872 (N_28872,N_24006,N_26565);
and U28873 (N_28873,N_25847,N_24450);
xnor U28874 (N_28874,N_25889,N_24956);
and U28875 (N_28875,N_24402,N_26807);
nand U28876 (N_28876,N_24223,N_24943);
or U28877 (N_28877,N_24967,N_24976);
and U28878 (N_28878,N_25410,N_26070);
and U28879 (N_28879,N_25301,N_26280);
xor U28880 (N_28880,N_26575,N_26823);
nand U28881 (N_28881,N_26198,N_24417);
or U28882 (N_28882,N_24525,N_26019);
and U28883 (N_28883,N_25349,N_25647);
and U28884 (N_28884,N_25188,N_24913);
xor U28885 (N_28885,N_24385,N_24331);
nand U28886 (N_28886,N_24433,N_24716);
nor U28887 (N_28887,N_26097,N_25077);
or U28888 (N_28888,N_24644,N_26178);
xor U28889 (N_28889,N_26752,N_26814);
xor U28890 (N_28890,N_25215,N_26665);
and U28891 (N_28891,N_26146,N_25038);
and U28892 (N_28892,N_25653,N_24633);
nor U28893 (N_28893,N_24046,N_24366);
nand U28894 (N_28894,N_24931,N_26343);
xnor U28895 (N_28895,N_24610,N_24067);
and U28896 (N_28896,N_26052,N_25909);
and U28897 (N_28897,N_26849,N_24775);
or U28898 (N_28898,N_24785,N_26259);
xor U28899 (N_28899,N_24315,N_24589);
nand U28900 (N_28900,N_26656,N_26086);
xnor U28901 (N_28901,N_26504,N_25227);
nand U28902 (N_28902,N_24266,N_24988);
xnor U28903 (N_28903,N_26281,N_25207);
xnor U28904 (N_28904,N_24744,N_24368);
or U28905 (N_28905,N_25521,N_25568);
or U28906 (N_28906,N_25436,N_26951);
nor U28907 (N_28907,N_24805,N_25491);
or U28908 (N_28908,N_24805,N_24825);
nor U28909 (N_28909,N_26125,N_25516);
nand U28910 (N_28910,N_26134,N_26900);
nand U28911 (N_28911,N_24383,N_24812);
nor U28912 (N_28912,N_25911,N_24369);
nor U28913 (N_28913,N_25347,N_25680);
nor U28914 (N_28914,N_25506,N_24125);
xor U28915 (N_28915,N_26253,N_24852);
or U28916 (N_28916,N_24446,N_26605);
and U28917 (N_28917,N_24141,N_25294);
nor U28918 (N_28918,N_26476,N_26484);
xnor U28919 (N_28919,N_25453,N_25889);
and U28920 (N_28920,N_24970,N_26623);
nor U28921 (N_28921,N_25852,N_25132);
nand U28922 (N_28922,N_25208,N_25475);
nor U28923 (N_28923,N_24723,N_26925);
or U28924 (N_28924,N_26132,N_24206);
nor U28925 (N_28925,N_25767,N_24890);
and U28926 (N_28926,N_26411,N_24323);
nor U28927 (N_28927,N_26540,N_25551);
or U28928 (N_28928,N_24094,N_26413);
and U28929 (N_28929,N_26084,N_25208);
xnor U28930 (N_28930,N_24214,N_25241);
xnor U28931 (N_28931,N_25782,N_24001);
nand U28932 (N_28932,N_24233,N_24066);
xor U28933 (N_28933,N_25123,N_24043);
xor U28934 (N_28934,N_25170,N_26059);
and U28935 (N_28935,N_24483,N_24856);
xnor U28936 (N_28936,N_26819,N_26064);
nand U28937 (N_28937,N_26431,N_25389);
and U28938 (N_28938,N_24787,N_24822);
or U28939 (N_28939,N_24639,N_26801);
nor U28940 (N_28940,N_24339,N_26838);
xnor U28941 (N_28941,N_24378,N_26055);
or U28942 (N_28942,N_26853,N_24579);
xnor U28943 (N_28943,N_24199,N_26792);
or U28944 (N_28944,N_26124,N_25692);
nand U28945 (N_28945,N_26331,N_25886);
nor U28946 (N_28946,N_26805,N_24017);
xnor U28947 (N_28947,N_25929,N_26985);
and U28948 (N_28948,N_24505,N_25735);
nor U28949 (N_28949,N_25977,N_26647);
nand U28950 (N_28950,N_25992,N_24540);
and U28951 (N_28951,N_25711,N_25287);
or U28952 (N_28952,N_25816,N_26826);
nand U28953 (N_28953,N_26899,N_24492);
nand U28954 (N_28954,N_26505,N_24580);
and U28955 (N_28955,N_25846,N_26483);
nand U28956 (N_28956,N_25993,N_26598);
and U28957 (N_28957,N_24375,N_25759);
or U28958 (N_28958,N_24425,N_24665);
nand U28959 (N_28959,N_24117,N_26574);
or U28960 (N_28960,N_24400,N_26700);
nor U28961 (N_28961,N_25474,N_26286);
nand U28962 (N_28962,N_24479,N_24091);
xor U28963 (N_28963,N_24247,N_24939);
xor U28964 (N_28964,N_25778,N_24548);
nand U28965 (N_28965,N_25988,N_26183);
nand U28966 (N_28966,N_25969,N_26285);
and U28967 (N_28967,N_24572,N_24806);
nor U28968 (N_28968,N_24624,N_25649);
nor U28969 (N_28969,N_25790,N_24777);
nor U28970 (N_28970,N_24132,N_24030);
nand U28971 (N_28971,N_26656,N_26915);
nor U28972 (N_28972,N_24191,N_24101);
or U28973 (N_28973,N_26516,N_26001);
and U28974 (N_28974,N_25441,N_25495);
nand U28975 (N_28975,N_26577,N_24719);
and U28976 (N_28976,N_25636,N_26637);
and U28977 (N_28977,N_26048,N_24884);
nand U28978 (N_28978,N_26999,N_26622);
nor U28979 (N_28979,N_25407,N_25374);
nand U28980 (N_28980,N_26791,N_26027);
nor U28981 (N_28981,N_26686,N_26032);
nor U28982 (N_28982,N_25479,N_25560);
or U28983 (N_28983,N_26307,N_25889);
nor U28984 (N_28984,N_24946,N_25278);
and U28985 (N_28985,N_24589,N_26499);
nor U28986 (N_28986,N_25239,N_26361);
nor U28987 (N_28987,N_24062,N_25749);
xor U28988 (N_28988,N_24626,N_24242);
and U28989 (N_28989,N_24894,N_25042);
nor U28990 (N_28990,N_24239,N_25631);
xor U28991 (N_28991,N_24258,N_26971);
nand U28992 (N_28992,N_26607,N_24222);
nand U28993 (N_28993,N_24636,N_26562);
and U28994 (N_28994,N_26988,N_24466);
nand U28995 (N_28995,N_24344,N_26422);
nor U28996 (N_28996,N_24244,N_24971);
or U28997 (N_28997,N_26388,N_26313);
nor U28998 (N_28998,N_24335,N_26466);
xor U28999 (N_28999,N_25773,N_26161);
nor U29000 (N_29000,N_25279,N_24294);
and U29001 (N_29001,N_26083,N_26429);
nor U29002 (N_29002,N_26736,N_26282);
xnor U29003 (N_29003,N_25870,N_26552);
or U29004 (N_29004,N_24241,N_26341);
or U29005 (N_29005,N_25344,N_24480);
nor U29006 (N_29006,N_24277,N_26576);
xnor U29007 (N_29007,N_26208,N_26983);
nand U29008 (N_29008,N_26781,N_26479);
or U29009 (N_29009,N_24323,N_25444);
nand U29010 (N_29010,N_24568,N_25860);
and U29011 (N_29011,N_25225,N_24927);
nand U29012 (N_29012,N_26968,N_26899);
or U29013 (N_29013,N_25713,N_24743);
and U29014 (N_29014,N_25821,N_24398);
xnor U29015 (N_29015,N_24285,N_24829);
nand U29016 (N_29016,N_24052,N_25020);
or U29017 (N_29017,N_25652,N_25641);
nand U29018 (N_29018,N_25363,N_25226);
or U29019 (N_29019,N_25646,N_24117);
and U29020 (N_29020,N_25314,N_26252);
nand U29021 (N_29021,N_26846,N_25755);
nand U29022 (N_29022,N_25030,N_24708);
and U29023 (N_29023,N_26878,N_24797);
and U29024 (N_29024,N_24918,N_26253);
or U29025 (N_29025,N_24098,N_26879);
or U29026 (N_29026,N_25154,N_24075);
and U29027 (N_29027,N_26429,N_25348);
or U29028 (N_29028,N_24415,N_25969);
nor U29029 (N_29029,N_24355,N_26061);
xnor U29030 (N_29030,N_25946,N_24572);
nor U29031 (N_29031,N_25945,N_25509);
or U29032 (N_29032,N_24631,N_24987);
and U29033 (N_29033,N_25081,N_26168);
or U29034 (N_29034,N_25623,N_26797);
nand U29035 (N_29035,N_25749,N_25609);
and U29036 (N_29036,N_25587,N_25733);
or U29037 (N_29037,N_26474,N_26228);
xnor U29038 (N_29038,N_24183,N_24915);
or U29039 (N_29039,N_25922,N_26497);
and U29040 (N_29040,N_25970,N_25476);
or U29041 (N_29041,N_25533,N_24033);
xor U29042 (N_29042,N_24123,N_24215);
xor U29043 (N_29043,N_26407,N_25501);
xor U29044 (N_29044,N_25238,N_24170);
nor U29045 (N_29045,N_25614,N_25512);
nor U29046 (N_29046,N_26511,N_26320);
and U29047 (N_29047,N_25093,N_26064);
nor U29048 (N_29048,N_25512,N_24103);
nor U29049 (N_29049,N_24657,N_26946);
xnor U29050 (N_29050,N_25437,N_24300);
nor U29051 (N_29051,N_24853,N_26723);
or U29052 (N_29052,N_25960,N_26761);
and U29053 (N_29053,N_26225,N_24430);
xor U29054 (N_29054,N_25905,N_26398);
and U29055 (N_29055,N_26210,N_24387);
and U29056 (N_29056,N_24040,N_26621);
nor U29057 (N_29057,N_25169,N_25040);
and U29058 (N_29058,N_24394,N_26337);
xnor U29059 (N_29059,N_26609,N_25884);
and U29060 (N_29060,N_26015,N_26877);
nand U29061 (N_29061,N_24178,N_25718);
xor U29062 (N_29062,N_26909,N_26549);
or U29063 (N_29063,N_25067,N_26014);
or U29064 (N_29064,N_25971,N_26875);
nor U29065 (N_29065,N_25369,N_24006);
nand U29066 (N_29066,N_26252,N_24793);
and U29067 (N_29067,N_24217,N_24485);
nor U29068 (N_29068,N_25090,N_26314);
nand U29069 (N_29069,N_24497,N_24496);
or U29070 (N_29070,N_25704,N_25920);
and U29071 (N_29071,N_26785,N_24900);
and U29072 (N_29072,N_24878,N_25482);
and U29073 (N_29073,N_24568,N_24077);
nor U29074 (N_29074,N_25931,N_26909);
xnor U29075 (N_29075,N_26181,N_24604);
xor U29076 (N_29076,N_24244,N_25979);
nor U29077 (N_29077,N_25227,N_25075);
or U29078 (N_29078,N_24203,N_25226);
nor U29079 (N_29079,N_24597,N_26801);
nand U29080 (N_29080,N_24178,N_26798);
xor U29081 (N_29081,N_24963,N_24016);
xnor U29082 (N_29082,N_25600,N_26765);
nor U29083 (N_29083,N_24917,N_26724);
or U29084 (N_29084,N_26398,N_25374);
nor U29085 (N_29085,N_26288,N_26707);
and U29086 (N_29086,N_26515,N_24797);
or U29087 (N_29087,N_25190,N_25666);
or U29088 (N_29088,N_25605,N_24031);
and U29089 (N_29089,N_25679,N_26690);
nand U29090 (N_29090,N_25026,N_26289);
and U29091 (N_29091,N_24359,N_24561);
and U29092 (N_29092,N_24355,N_25266);
and U29093 (N_29093,N_26496,N_24866);
xnor U29094 (N_29094,N_25839,N_26278);
xnor U29095 (N_29095,N_26219,N_25027);
nand U29096 (N_29096,N_25925,N_26164);
or U29097 (N_29097,N_25514,N_24467);
and U29098 (N_29098,N_24422,N_25611);
or U29099 (N_29099,N_25859,N_25819);
and U29100 (N_29100,N_24488,N_24912);
nor U29101 (N_29101,N_25469,N_26572);
nand U29102 (N_29102,N_24097,N_24831);
xor U29103 (N_29103,N_26598,N_24533);
xor U29104 (N_29104,N_25173,N_26502);
nand U29105 (N_29105,N_25139,N_26585);
nor U29106 (N_29106,N_24756,N_26608);
or U29107 (N_29107,N_24063,N_24722);
nor U29108 (N_29108,N_24349,N_24896);
and U29109 (N_29109,N_25665,N_25285);
or U29110 (N_29110,N_26523,N_24071);
nand U29111 (N_29111,N_25548,N_25653);
nor U29112 (N_29112,N_24725,N_25377);
or U29113 (N_29113,N_24194,N_24523);
nand U29114 (N_29114,N_26118,N_26650);
nand U29115 (N_29115,N_26775,N_25275);
nand U29116 (N_29116,N_24997,N_25497);
or U29117 (N_29117,N_26543,N_24878);
nand U29118 (N_29118,N_25851,N_26422);
and U29119 (N_29119,N_24468,N_25683);
xnor U29120 (N_29120,N_25803,N_25406);
and U29121 (N_29121,N_25927,N_25702);
and U29122 (N_29122,N_25577,N_24480);
xor U29123 (N_29123,N_26900,N_25417);
and U29124 (N_29124,N_24817,N_24430);
nand U29125 (N_29125,N_26858,N_24566);
and U29126 (N_29126,N_25352,N_24662);
nand U29127 (N_29127,N_24793,N_26616);
and U29128 (N_29128,N_25767,N_24553);
nor U29129 (N_29129,N_26865,N_24226);
and U29130 (N_29130,N_24090,N_25549);
xor U29131 (N_29131,N_24924,N_24873);
and U29132 (N_29132,N_24347,N_24279);
nor U29133 (N_29133,N_25633,N_25443);
xnor U29134 (N_29134,N_24736,N_24181);
or U29135 (N_29135,N_26870,N_26112);
xnor U29136 (N_29136,N_26366,N_24053);
or U29137 (N_29137,N_24697,N_26523);
and U29138 (N_29138,N_25045,N_25881);
nand U29139 (N_29139,N_25685,N_25151);
nand U29140 (N_29140,N_24861,N_25867);
nor U29141 (N_29141,N_25854,N_26217);
nor U29142 (N_29142,N_24807,N_25757);
or U29143 (N_29143,N_26826,N_24958);
nand U29144 (N_29144,N_26482,N_26107);
nor U29145 (N_29145,N_25947,N_24413);
xor U29146 (N_29146,N_25161,N_25036);
nand U29147 (N_29147,N_25191,N_24611);
nor U29148 (N_29148,N_24916,N_26764);
nand U29149 (N_29149,N_26345,N_26131);
or U29150 (N_29150,N_26902,N_24572);
and U29151 (N_29151,N_26732,N_26971);
nor U29152 (N_29152,N_24946,N_26487);
nand U29153 (N_29153,N_25910,N_24630);
nor U29154 (N_29154,N_24092,N_26286);
and U29155 (N_29155,N_25910,N_24510);
xnor U29156 (N_29156,N_24310,N_24522);
nor U29157 (N_29157,N_26010,N_26993);
or U29158 (N_29158,N_26394,N_25408);
nor U29159 (N_29159,N_25132,N_25868);
nand U29160 (N_29160,N_25447,N_24791);
nor U29161 (N_29161,N_25633,N_24363);
nand U29162 (N_29162,N_26363,N_25001);
or U29163 (N_29163,N_25633,N_26334);
or U29164 (N_29164,N_25902,N_26837);
xnor U29165 (N_29165,N_26084,N_26494);
or U29166 (N_29166,N_26365,N_24554);
nor U29167 (N_29167,N_25290,N_25943);
or U29168 (N_29168,N_25076,N_24432);
nor U29169 (N_29169,N_26334,N_26260);
xnor U29170 (N_29170,N_26445,N_25048);
nor U29171 (N_29171,N_24161,N_25505);
nor U29172 (N_29172,N_25716,N_25736);
or U29173 (N_29173,N_25835,N_24872);
nor U29174 (N_29174,N_25762,N_24038);
nor U29175 (N_29175,N_25670,N_25233);
or U29176 (N_29176,N_24377,N_26517);
and U29177 (N_29177,N_25154,N_26484);
and U29178 (N_29178,N_26171,N_25587);
or U29179 (N_29179,N_24764,N_26822);
nand U29180 (N_29180,N_24607,N_26719);
xnor U29181 (N_29181,N_24925,N_24857);
nand U29182 (N_29182,N_25867,N_26774);
nand U29183 (N_29183,N_25198,N_25954);
nor U29184 (N_29184,N_25653,N_25436);
xor U29185 (N_29185,N_25140,N_25195);
nor U29186 (N_29186,N_26801,N_26058);
xnor U29187 (N_29187,N_24995,N_24195);
nand U29188 (N_29188,N_26601,N_24818);
or U29189 (N_29189,N_25035,N_26153);
xnor U29190 (N_29190,N_25025,N_26320);
nand U29191 (N_29191,N_25787,N_25612);
or U29192 (N_29192,N_24847,N_26593);
and U29193 (N_29193,N_24976,N_26456);
and U29194 (N_29194,N_25526,N_24832);
nand U29195 (N_29195,N_24553,N_26051);
and U29196 (N_29196,N_26106,N_25911);
nor U29197 (N_29197,N_24448,N_25041);
nor U29198 (N_29198,N_26729,N_24481);
nand U29199 (N_29199,N_24374,N_24075);
and U29200 (N_29200,N_26910,N_24479);
xor U29201 (N_29201,N_26552,N_26700);
nand U29202 (N_29202,N_24448,N_24328);
or U29203 (N_29203,N_25882,N_25805);
or U29204 (N_29204,N_26349,N_26276);
or U29205 (N_29205,N_26901,N_24234);
nor U29206 (N_29206,N_24700,N_24412);
nand U29207 (N_29207,N_26590,N_24535);
or U29208 (N_29208,N_25553,N_24290);
nand U29209 (N_29209,N_26376,N_24641);
nor U29210 (N_29210,N_24249,N_25264);
nor U29211 (N_29211,N_26428,N_26388);
nand U29212 (N_29212,N_24948,N_25967);
or U29213 (N_29213,N_26125,N_25082);
and U29214 (N_29214,N_24550,N_25742);
or U29215 (N_29215,N_26269,N_26747);
or U29216 (N_29216,N_26648,N_25699);
xnor U29217 (N_29217,N_26381,N_24115);
or U29218 (N_29218,N_26234,N_24090);
xnor U29219 (N_29219,N_24621,N_25216);
nand U29220 (N_29220,N_25031,N_26806);
or U29221 (N_29221,N_26950,N_25568);
and U29222 (N_29222,N_24407,N_24418);
nor U29223 (N_29223,N_25987,N_25295);
nor U29224 (N_29224,N_24245,N_24894);
xor U29225 (N_29225,N_24467,N_24752);
nand U29226 (N_29226,N_24950,N_26991);
or U29227 (N_29227,N_25774,N_24496);
nor U29228 (N_29228,N_26280,N_24292);
nand U29229 (N_29229,N_26533,N_24917);
nand U29230 (N_29230,N_25112,N_25730);
nor U29231 (N_29231,N_25673,N_25472);
nand U29232 (N_29232,N_26491,N_25392);
and U29233 (N_29233,N_24259,N_24181);
and U29234 (N_29234,N_24637,N_25575);
nand U29235 (N_29235,N_25416,N_25730);
xor U29236 (N_29236,N_25974,N_24913);
xnor U29237 (N_29237,N_25890,N_24914);
or U29238 (N_29238,N_26235,N_26573);
nand U29239 (N_29239,N_24822,N_24457);
nand U29240 (N_29240,N_24575,N_25690);
nand U29241 (N_29241,N_24410,N_26497);
or U29242 (N_29242,N_24038,N_25559);
xor U29243 (N_29243,N_26236,N_25741);
nor U29244 (N_29244,N_24893,N_24151);
nor U29245 (N_29245,N_26171,N_25996);
and U29246 (N_29246,N_26354,N_25522);
nand U29247 (N_29247,N_25590,N_24660);
or U29248 (N_29248,N_25390,N_26184);
nand U29249 (N_29249,N_24034,N_26798);
or U29250 (N_29250,N_24786,N_26716);
and U29251 (N_29251,N_26404,N_25549);
or U29252 (N_29252,N_26094,N_26313);
nor U29253 (N_29253,N_25084,N_24163);
nand U29254 (N_29254,N_24251,N_26875);
and U29255 (N_29255,N_24772,N_24513);
or U29256 (N_29256,N_25906,N_26312);
and U29257 (N_29257,N_26240,N_24285);
nand U29258 (N_29258,N_24291,N_26615);
or U29259 (N_29259,N_24823,N_25520);
xor U29260 (N_29260,N_25112,N_25761);
or U29261 (N_29261,N_24905,N_26162);
and U29262 (N_29262,N_24105,N_24529);
and U29263 (N_29263,N_24174,N_24630);
or U29264 (N_29264,N_25897,N_26046);
nand U29265 (N_29265,N_24783,N_26449);
nor U29266 (N_29266,N_24669,N_24557);
nor U29267 (N_29267,N_25238,N_24519);
and U29268 (N_29268,N_24595,N_25974);
and U29269 (N_29269,N_25080,N_25663);
or U29270 (N_29270,N_24773,N_24996);
nand U29271 (N_29271,N_24981,N_24509);
nor U29272 (N_29272,N_24630,N_25201);
nor U29273 (N_29273,N_25766,N_26260);
or U29274 (N_29274,N_25732,N_25867);
nand U29275 (N_29275,N_24831,N_25704);
and U29276 (N_29276,N_25720,N_24713);
xnor U29277 (N_29277,N_26193,N_24212);
xnor U29278 (N_29278,N_24756,N_24278);
or U29279 (N_29279,N_24003,N_25338);
nor U29280 (N_29280,N_25723,N_25370);
nor U29281 (N_29281,N_24573,N_25962);
and U29282 (N_29282,N_25505,N_24952);
nand U29283 (N_29283,N_25080,N_24371);
and U29284 (N_29284,N_26114,N_25110);
nor U29285 (N_29285,N_25692,N_26665);
nand U29286 (N_29286,N_24953,N_24590);
nand U29287 (N_29287,N_26531,N_25317);
xor U29288 (N_29288,N_25317,N_26110);
nor U29289 (N_29289,N_24858,N_25918);
and U29290 (N_29290,N_25896,N_26920);
xor U29291 (N_29291,N_26832,N_25094);
nor U29292 (N_29292,N_26185,N_24897);
or U29293 (N_29293,N_25463,N_26387);
or U29294 (N_29294,N_24195,N_25452);
xnor U29295 (N_29295,N_24326,N_25280);
xor U29296 (N_29296,N_25945,N_26638);
nand U29297 (N_29297,N_24936,N_24301);
xnor U29298 (N_29298,N_24732,N_24230);
nor U29299 (N_29299,N_25434,N_26093);
nor U29300 (N_29300,N_25983,N_24300);
nor U29301 (N_29301,N_25666,N_26224);
nor U29302 (N_29302,N_26678,N_26654);
nor U29303 (N_29303,N_25211,N_25653);
or U29304 (N_29304,N_25085,N_26925);
nand U29305 (N_29305,N_26278,N_26479);
xnor U29306 (N_29306,N_26757,N_24966);
xor U29307 (N_29307,N_24076,N_24025);
nand U29308 (N_29308,N_25366,N_26698);
xnor U29309 (N_29309,N_26017,N_24403);
nor U29310 (N_29310,N_24802,N_25098);
or U29311 (N_29311,N_26036,N_25355);
nand U29312 (N_29312,N_24243,N_25412);
and U29313 (N_29313,N_24424,N_26858);
nand U29314 (N_29314,N_26828,N_26207);
nand U29315 (N_29315,N_25127,N_26908);
nor U29316 (N_29316,N_26785,N_26854);
or U29317 (N_29317,N_26888,N_24147);
nand U29318 (N_29318,N_25417,N_24763);
and U29319 (N_29319,N_25886,N_24153);
nand U29320 (N_29320,N_26347,N_25377);
and U29321 (N_29321,N_26270,N_24416);
nor U29322 (N_29322,N_24125,N_26335);
nor U29323 (N_29323,N_26745,N_24077);
xor U29324 (N_29324,N_26870,N_26286);
xnor U29325 (N_29325,N_25907,N_24703);
and U29326 (N_29326,N_24528,N_25549);
nand U29327 (N_29327,N_24249,N_26229);
xnor U29328 (N_29328,N_25220,N_24544);
or U29329 (N_29329,N_24428,N_25310);
nand U29330 (N_29330,N_26378,N_24398);
nor U29331 (N_29331,N_24246,N_26220);
or U29332 (N_29332,N_25923,N_26687);
and U29333 (N_29333,N_26904,N_25099);
nand U29334 (N_29334,N_26014,N_26948);
nand U29335 (N_29335,N_25165,N_26291);
xnor U29336 (N_29336,N_24468,N_25466);
and U29337 (N_29337,N_26245,N_25705);
and U29338 (N_29338,N_26712,N_26731);
nor U29339 (N_29339,N_24552,N_26560);
or U29340 (N_29340,N_25078,N_26611);
xor U29341 (N_29341,N_25261,N_25507);
nand U29342 (N_29342,N_24824,N_25011);
nor U29343 (N_29343,N_26615,N_26502);
and U29344 (N_29344,N_26743,N_26789);
or U29345 (N_29345,N_24759,N_25072);
or U29346 (N_29346,N_25082,N_24431);
nor U29347 (N_29347,N_24967,N_26014);
or U29348 (N_29348,N_24423,N_25543);
xnor U29349 (N_29349,N_26532,N_25200);
or U29350 (N_29350,N_24991,N_25755);
and U29351 (N_29351,N_26703,N_25603);
and U29352 (N_29352,N_24192,N_25222);
and U29353 (N_29353,N_25530,N_24757);
nor U29354 (N_29354,N_25441,N_26726);
or U29355 (N_29355,N_25059,N_24727);
nor U29356 (N_29356,N_24438,N_25267);
nand U29357 (N_29357,N_26200,N_26482);
nand U29358 (N_29358,N_25209,N_24639);
and U29359 (N_29359,N_26337,N_26597);
nor U29360 (N_29360,N_25125,N_25828);
nand U29361 (N_29361,N_26495,N_26629);
and U29362 (N_29362,N_26974,N_24074);
nor U29363 (N_29363,N_25608,N_24312);
xnor U29364 (N_29364,N_26846,N_24675);
or U29365 (N_29365,N_26759,N_26762);
nand U29366 (N_29366,N_24842,N_25499);
nor U29367 (N_29367,N_25061,N_24363);
nor U29368 (N_29368,N_24768,N_26353);
and U29369 (N_29369,N_24141,N_26055);
nor U29370 (N_29370,N_24520,N_26448);
and U29371 (N_29371,N_24902,N_24121);
nor U29372 (N_29372,N_25451,N_26843);
nand U29373 (N_29373,N_25163,N_24827);
xor U29374 (N_29374,N_25087,N_26059);
nor U29375 (N_29375,N_26314,N_25524);
nor U29376 (N_29376,N_26625,N_25363);
xor U29377 (N_29377,N_25947,N_25596);
and U29378 (N_29378,N_24445,N_25415);
or U29379 (N_29379,N_26911,N_25345);
xnor U29380 (N_29380,N_25310,N_24632);
or U29381 (N_29381,N_25692,N_24476);
nand U29382 (N_29382,N_24585,N_24346);
nor U29383 (N_29383,N_25174,N_26286);
nand U29384 (N_29384,N_25315,N_26705);
xnor U29385 (N_29385,N_25992,N_25385);
nand U29386 (N_29386,N_24241,N_24283);
nor U29387 (N_29387,N_25030,N_26951);
nand U29388 (N_29388,N_24512,N_24544);
nand U29389 (N_29389,N_26646,N_24628);
and U29390 (N_29390,N_24212,N_24629);
nor U29391 (N_29391,N_24750,N_26588);
xor U29392 (N_29392,N_26070,N_24591);
or U29393 (N_29393,N_24309,N_24367);
nand U29394 (N_29394,N_25652,N_25089);
nand U29395 (N_29395,N_25778,N_24666);
or U29396 (N_29396,N_26354,N_25757);
xor U29397 (N_29397,N_26702,N_24569);
or U29398 (N_29398,N_26006,N_26623);
nand U29399 (N_29399,N_26113,N_26468);
nand U29400 (N_29400,N_26932,N_24206);
nand U29401 (N_29401,N_25664,N_26789);
or U29402 (N_29402,N_25421,N_26963);
or U29403 (N_29403,N_26945,N_26572);
xor U29404 (N_29404,N_24871,N_25844);
nor U29405 (N_29405,N_24656,N_25504);
nor U29406 (N_29406,N_24474,N_24708);
and U29407 (N_29407,N_25192,N_26271);
nor U29408 (N_29408,N_26084,N_24692);
and U29409 (N_29409,N_26687,N_24161);
and U29410 (N_29410,N_26206,N_24308);
nor U29411 (N_29411,N_26325,N_24122);
or U29412 (N_29412,N_26764,N_25840);
nand U29413 (N_29413,N_25848,N_26578);
nand U29414 (N_29414,N_25221,N_26909);
xor U29415 (N_29415,N_26389,N_25640);
nand U29416 (N_29416,N_26131,N_24046);
xnor U29417 (N_29417,N_25132,N_26002);
nor U29418 (N_29418,N_26468,N_24157);
nand U29419 (N_29419,N_24809,N_24877);
or U29420 (N_29420,N_24621,N_26555);
xor U29421 (N_29421,N_25131,N_26728);
nor U29422 (N_29422,N_25573,N_26149);
or U29423 (N_29423,N_26672,N_24601);
xor U29424 (N_29424,N_26352,N_24118);
nand U29425 (N_29425,N_24969,N_24866);
or U29426 (N_29426,N_24947,N_26820);
nor U29427 (N_29427,N_24256,N_25598);
nor U29428 (N_29428,N_24377,N_25918);
nor U29429 (N_29429,N_26502,N_24659);
xor U29430 (N_29430,N_26956,N_25212);
or U29431 (N_29431,N_26157,N_25720);
nor U29432 (N_29432,N_26436,N_24251);
nand U29433 (N_29433,N_26871,N_26507);
xor U29434 (N_29434,N_24824,N_24921);
nor U29435 (N_29435,N_24854,N_26541);
nand U29436 (N_29436,N_24143,N_25667);
and U29437 (N_29437,N_25352,N_24504);
xnor U29438 (N_29438,N_24842,N_25914);
or U29439 (N_29439,N_25863,N_25111);
nor U29440 (N_29440,N_25037,N_26929);
xor U29441 (N_29441,N_26998,N_26731);
xnor U29442 (N_29442,N_26859,N_24617);
or U29443 (N_29443,N_24041,N_24159);
xor U29444 (N_29444,N_26410,N_25606);
xnor U29445 (N_29445,N_24768,N_24496);
xor U29446 (N_29446,N_24940,N_26480);
nor U29447 (N_29447,N_24468,N_25438);
and U29448 (N_29448,N_24596,N_24320);
and U29449 (N_29449,N_24342,N_26818);
and U29450 (N_29450,N_25941,N_26251);
and U29451 (N_29451,N_25960,N_24777);
nand U29452 (N_29452,N_26599,N_26864);
and U29453 (N_29453,N_26964,N_24795);
nand U29454 (N_29454,N_26765,N_25875);
or U29455 (N_29455,N_25992,N_24299);
or U29456 (N_29456,N_25941,N_24475);
and U29457 (N_29457,N_26513,N_24356);
nor U29458 (N_29458,N_26198,N_24867);
nand U29459 (N_29459,N_25833,N_26078);
xor U29460 (N_29460,N_25695,N_25705);
or U29461 (N_29461,N_24157,N_24669);
and U29462 (N_29462,N_25233,N_26445);
nor U29463 (N_29463,N_24882,N_25036);
nor U29464 (N_29464,N_25502,N_25847);
and U29465 (N_29465,N_24778,N_26691);
xnor U29466 (N_29466,N_26677,N_26423);
nor U29467 (N_29467,N_25942,N_26651);
and U29468 (N_29468,N_24033,N_24219);
and U29469 (N_29469,N_25505,N_25728);
nand U29470 (N_29470,N_25613,N_24998);
xor U29471 (N_29471,N_25918,N_25066);
nor U29472 (N_29472,N_25406,N_25925);
xor U29473 (N_29473,N_25004,N_25798);
or U29474 (N_29474,N_24624,N_26729);
xor U29475 (N_29475,N_24158,N_26585);
nand U29476 (N_29476,N_25903,N_24641);
xnor U29477 (N_29477,N_24826,N_25518);
nand U29478 (N_29478,N_24395,N_25735);
nand U29479 (N_29479,N_26683,N_26395);
and U29480 (N_29480,N_24423,N_24372);
nor U29481 (N_29481,N_26924,N_25734);
or U29482 (N_29482,N_24060,N_25749);
xor U29483 (N_29483,N_26590,N_26832);
or U29484 (N_29484,N_24523,N_26447);
xnor U29485 (N_29485,N_25978,N_24907);
nor U29486 (N_29486,N_26849,N_25715);
and U29487 (N_29487,N_25104,N_25994);
xnor U29488 (N_29488,N_24881,N_25010);
or U29489 (N_29489,N_24359,N_24266);
nand U29490 (N_29490,N_25409,N_26991);
and U29491 (N_29491,N_24714,N_25264);
xor U29492 (N_29492,N_26538,N_25317);
or U29493 (N_29493,N_24072,N_24504);
xnor U29494 (N_29494,N_25763,N_25480);
xor U29495 (N_29495,N_26600,N_25476);
nand U29496 (N_29496,N_24841,N_26261);
nor U29497 (N_29497,N_24535,N_25139);
and U29498 (N_29498,N_24637,N_26094);
xor U29499 (N_29499,N_25862,N_25421);
nand U29500 (N_29500,N_24961,N_26984);
or U29501 (N_29501,N_24319,N_26992);
nand U29502 (N_29502,N_26269,N_25103);
and U29503 (N_29503,N_25485,N_25871);
or U29504 (N_29504,N_25575,N_26759);
nand U29505 (N_29505,N_25668,N_25758);
nand U29506 (N_29506,N_24704,N_24565);
or U29507 (N_29507,N_26569,N_26735);
and U29508 (N_29508,N_24934,N_26703);
and U29509 (N_29509,N_25962,N_26795);
and U29510 (N_29510,N_24805,N_25709);
and U29511 (N_29511,N_26004,N_24190);
or U29512 (N_29512,N_25763,N_24789);
nor U29513 (N_29513,N_26883,N_25356);
nand U29514 (N_29514,N_26027,N_24202);
xnor U29515 (N_29515,N_26060,N_26951);
xor U29516 (N_29516,N_26142,N_26487);
xor U29517 (N_29517,N_26425,N_26818);
xnor U29518 (N_29518,N_25520,N_24702);
nand U29519 (N_29519,N_25776,N_25833);
nor U29520 (N_29520,N_24570,N_24664);
nor U29521 (N_29521,N_25314,N_26354);
xnor U29522 (N_29522,N_26199,N_26537);
nand U29523 (N_29523,N_25892,N_26036);
or U29524 (N_29524,N_24127,N_26950);
nand U29525 (N_29525,N_24292,N_26916);
nor U29526 (N_29526,N_25423,N_24775);
nand U29527 (N_29527,N_25786,N_24253);
nor U29528 (N_29528,N_25666,N_24322);
nand U29529 (N_29529,N_25576,N_24771);
nor U29530 (N_29530,N_25241,N_25031);
nand U29531 (N_29531,N_24925,N_26915);
xor U29532 (N_29532,N_24029,N_24636);
nor U29533 (N_29533,N_24136,N_24364);
or U29534 (N_29534,N_25465,N_25058);
xor U29535 (N_29535,N_24320,N_25454);
and U29536 (N_29536,N_25999,N_24086);
xor U29537 (N_29537,N_26003,N_24372);
xor U29538 (N_29538,N_26237,N_24300);
nor U29539 (N_29539,N_24337,N_25707);
or U29540 (N_29540,N_24289,N_24546);
nand U29541 (N_29541,N_26828,N_26745);
and U29542 (N_29542,N_26584,N_24265);
or U29543 (N_29543,N_25397,N_26386);
nor U29544 (N_29544,N_24998,N_26260);
xor U29545 (N_29545,N_26403,N_24044);
or U29546 (N_29546,N_24595,N_24794);
or U29547 (N_29547,N_26554,N_26759);
xor U29548 (N_29548,N_25844,N_26720);
nor U29549 (N_29549,N_25306,N_26753);
nor U29550 (N_29550,N_24212,N_25400);
and U29551 (N_29551,N_25263,N_26049);
or U29552 (N_29552,N_25488,N_25280);
or U29553 (N_29553,N_26118,N_26510);
xor U29554 (N_29554,N_24844,N_24365);
nand U29555 (N_29555,N_26918,N_25626);
or U29556 (N_29556,N_24245,N_24288);
and U29557 (N_29557,N_24700,N_24494);
nand U29558 (N_29558,N_24900,N_25549);
nand U29559 (N_29559,N_24435,N_25879);
and U29560 (N_29560,N_24040,N_25038);
nand U29561 (N_29561,N_26684,N_25461);
nor U29562 (N_29562,N_24050,N_26784);
and U29563 (N_29563,N_25178,N_26760);
or U29564 (N_29564,N_26100,N_25642);
nand U29565 (N_29565,N_26620,N_25003);
nand U29566 (N_29566,N_25925,N_24549);
xor U29567 (N_29567,N_25587,N_26478);
xnor U29568 (N_29568,N_25583,N_24378);
or U29569 (N_29569,N_26981,N_26812);
nor U29570 (N_29570,N_26880,N_25536);
xnor U29571 (N_29571,N_26631,N_26117);
and U29572 (N_29572,N_24220,N_24105);
nand U29573 (N_29573,N_25703,N_24402);
or U29574 (N_29574,N_25096,N_26198);
and U29575 (N_29575,N_26973,N_25786);
and U29576 (N_29576,N_24380,N_26106);
nand U29577 (N_29577,N_26338,N_25953);
and U29578 (N_29578,N_24585,N_25911);
or U29579 (N_29579,N_26567,N_26220);
nand U29580 (N_29580,N_25984,N_26088);
xnor U29581 (N_29581,N_25429,N_25892);
or U29582 (N_29582,N_26617,N_24456);
and U29583 (N_29583,N_24969,N_25392);
xor U29584 (N_29584,N_24865,N_25588);
xnor U29585 (N_29585,N_26690,N_25190);
nor U29586 (N_29586,N_24360,N_25197);
and U29587 (N_29587,N_25917,N_26303);
xor U29588 (N_29588,N_24560,N_24048);
nand U29589 (N_29589,N_26808,N_24895);
or U29590 (N_29590,N_25152,N_25842);
nor U29591 (N_29591,N_25256,N_26860);
and U29592 (N_29592,N_25441,N_25120);
xnor U29593 (N_29593,N_24641,N_26020);
or U29594 (N_29594,N_26174,N_24543);
nand U29595 (N_29595,N_26665,N_25954);
xor U29596 (N_29596,N_26386,N_26377);
and U29597 (N_29597,N_25771,N_24561);
xor U29598 (N_29598,N_25470,N_24444);
nor U29599 (N_29599,N_24998,N_26160);
and U29600 (N_29600,N_26992,N_24042);
nor U29601 (N_29601,N_24320,N_25317);
and U29602 (N_29602,N_24585,N_25186);
or U29603 (N_29603,N_24620,N_26134);
xnor U29604 (N_29604,N_26328,N_26696);
nand U29605 (N_29605,N_24262,N_24612);
nor U29606 (N_29606,N_26894,N_26424);
and U29607 (N_29607,N_26228,N_24925);
nor U29608 (N_29608,N_26789,N_25459);
or U29609 (N_29609,N_25346,N_26672);
xnor U29610 (N_29610,N_25694,N_26361);
xnor U29611 (N_29611,N_26309,N_24390);
nand U29612 (N_29612,N_26918,N_24975);
xor U29613 (N_29613,N_25973,N_25502);
xor U29614 (N_29614,N_25179,N_25440);
xnor U29615 (N_29615,N_26974,N_25385);
or U29616 (N_29616,N_25353,N_24986);
nand U29617 (N_29617,N_25820,N_24924);
and U29618 (N_29618,N_26992,N_24182);
or U29619 (N_29619,N_24903,N_26591);
and U29620 (N_29620,N_25177,N_25558);
xnor U29621 (N_29621,N_26318,N_26234);
nor U29622 (N_29622,N_26331,N_24950);
or U29623 (N_29623,N_26901,N_26894);
nand U29624 (N_29624,N_26949,N_25654);
or U29625 (N_29625,N_25495,N_26646);
xnor U29626 (N_29626,N_24292,N_24907);
and U29627 (N_29627,N_25314,N_24643);
or U29628 (N_29628,N_24421,N_24086);
nor U29629 (N_29629,N_26584,N_24117);
or U29630 (N_29630,N_26365,N_26937);
or U29631 (N_29631,N_25751,N_26477);
nand U29632 (N_29632,N_25343,N_24774);
and U29633 (N_29633,N_24341,N_24596);
or U29634 (N_29634,N_25370,N_24101);
nand U29635 (N_29635,N_24204,N_26725);
nor U29636 (N_29636,N_24997,N_26867);
and U29637 (N_29637,N_24582,N_26006);
nor U29638 (N_29638,N_24713,N_24997);
nor U29639 (N_29639,N_26241,N_26257);
nand U29640 (N_29640,N_24158,N_25638);
nor U29641 (N_29641,N_25522,N_24592);
and U29642 (N_29642,N_24211,N_26896);
and U29643 (N_29643,N_25874,N_25472);
nand U29644 (N_29644,N_26115,N_24952);
and U29645 (N_29645,N_25999,N_24483);
xnor U29646 (N_29646,N_25064,N_26948);
nor U29647 (N_29647,N_25079,N_25168);
nor U29648 (N_29648,N_25621,N_25830);
xor U29649 (N_29649,N_25312,N_24264);
xnor U29650 (N_29650,N_26567,N_25410);
nor U29651 (N_29651,N_24854,N_25407);
and U29652 (N_29652,N_25712,N_24672);
nand U29653 (N_29653,N_25506,N_26626);
xnor U29654 (N_29654,N_25674,N_24617);
nand U29655 (N_29655,N_24247,N_24330);
nand U29656 (N_29656,N_24561,N_24818);
nand U29657 (N_29657,N_25618,N_26354);
nand U29658 (N_29658,N_26643,N_26777);
xnor U29659 (N_29659,N_26980,N_26598);
nor U29660 (N_29660,N_25978,N_24521);
xnor U29661 (N_29661,N_24775,N_26445);
or U29662 (N_29662,N_26105,N_25369);
and U29663 (N_29663,N_25693,N_25299);
nor U29664 (N_29664,N_25605,N_24483);
xor U29665 (N_29665,N_24755,N_24011);
or U29666 (N_29666,N_24469,N_24201);
nor U29667 (N_29667,N_26599,N_24564);
and U29668 (N_29668,N_25695,N_24571);
nor U29669 (N_29669,N_26710,N_24881);
nor U29670 (N_29670,N_24684,N_24527);
and U29671 (N_29671,N_25659,N_24920);
and U29672 (N_29672,N_26983,N_25860);
and U29673 (N_29673,N_25865,N_25291);
and U29674 (N_29674,N_25954,N_24048);
xor U29675 (N_29675,N_24333,N_26637);
nor U29676 (N_29676,N_25572,N_24680);
xnor U29677 (N_29677,N_24626,N_24480);
nand U29678 (N_29678,N_26656,N_24533);
xor U29679 (N_29679,N_26944,N_26133);
nand U29680 (N_29680,N_26606,N_24579);
and U29681 (N_29681,N_24960,N_25528);
nand U29682 (N_29682,N_26612,N_25229);
nand U29683 (N_29683,N_26567,N_24080);
nand U29684 (N_29684,N_26081,N_24127);
nor U29685 (N_29685,N_26284,N_26652);
and U29686 (N_29686,N_26720,N_24030);
xnor U29687 (N_29687,N_24709,N_26199);
xor U29688 (N_29688,N_26368,N_25911);
or U29689 (N_29689,N_25404,N_24509);
and U29690 (N_29690,N_25289,N_26894);
nand U29691 (N_29691,N_24518,N_26726);
nor U29692 (N_29692,N_24896,N_24248);
xnor U29693 (N_29693,N_25903,N_24319);
nor U29694 (N_29694,N_24698,N_25032);
nor U29695 (N_29695,N_24324,N_26296);
xnor U29696 (N_29696,N_25077,N_24200);
or U29697 (N_29697,N_26103,N_25729);
or U29698 (N_29698,N_26095,N_24526);
nor U29699 (N_29699,N_24520,N_24045);
xnor U29700 (N_29700,N_25306,N_26792);
and U29701 (N_29701,N_26165,N_25844);
and U29702 (N_29702,N_26609,N_25836);
xor U29703 (N_29703,N_25712,N_25149);
nor U29704 (N_29704,N_25677,N_25562);
and U29705 (N_29705,N_26218,N_24680);
or U29706 (N_29706,N_26134,N_25621);
or U29707 (N_29707,N_25721,N_24864);
xor U29708 (N_29708,N_26005,N_26239);
and U29709 (N_29709,N_26587,N_24691);
and U29710 (N_29710,N_24339,N_24032);
and U29711 (N_29711,N_26818,N_24243);
nor U29712 (N_29712,N_25855,N_26150);
and U29713 (N_29713,N_26247,N_26019);
nand U29714 (N_29714,N_26888,N_24075);
or U29715 (N_29715,N_25560,N_24368);
xnor U29716 (N_29716,N_26840,N_25005);
or U29717 (N_29717,N_25320,N_26503);
or U29718 (N_29718,N_25321,N_25657);
nor U29719 (N_29719,N_24977,N_24012);
and U29720 (N_29720,N_26034,N_26945);
xor U29721 (N_29721,N_24819,N_25246);
nand U29722 (N_29722,N_25103,N_24426);
and U29723 (N_29723,N_24655,N_26346);
nor U29724 (N_29724,N_25877,N_24902);
and U29725 (N_29725,N_24017,N_26589);
and U29726 (N_29726,N_26803,N_25422);
nand U29727 (N_29727,N_26406,N_25973);
and U29728 (N_29728,N_26169,N_24916);
or U29729 (N_29729,N_26940,N_25769);
xor U29730 (N_29730,N_26286,N_24345);
or U29731 (N_29731,N_24788,N_24370);
or U29732 (N_29732,N_25353,N_25419);
nor U29733 (N_29733,N_26323,N_26659);
xnor U29734 (N_29734,N_24482,N_26861);
xnor U29735 (N_29735,N_26206,N_25464);
nand U29736 (N_29736,N_24734,N_24635);
nand U29737 (N_29737,N_26687,N_25842);
nand U29738 (N_29738,N_26180,N_24855);
xnor U29739 (N_29739,N_24204,N_24656);
and U29740 (N_29740,N_25159,N_24916);
xnor U29741 (N_29741,N_26079,N_26251);
nand U29742 (N_29742,N_24165,N_25026);
or U29743 (N_29743,N_24226,N_25286);
nor U29744 (N_29744,N_25749,N_26857);
nor U29745 (N_29745,N_24179,N_25752);
nand U29746 (N_29746,N_24824,N_25003);
nor U29747 (N_29747,N_24328,N_26882);
nor U29748 (N_29748,N_26750,N_25578);
or U29749 (N_29749,N_25694,N_26082);
or U29750 (N_29750,N_25963,N_24920);
or U29751 (N_29751,N_26961,N_26540);
xnor U29752 (N_29752,N_25679,N_24822);
nand U29753 (N_29753,N_24770,N_26669);
or U29754 (N_29754,N_25310,N_25128);
nand U29755 (N_29755,N_26985,N_25393);
or U29756 (N_29756,N_25839,N_25688);
or U29757 (N_29757,N_24153,N_24235);
or U29758 (N_29758,N_25146,N_24943);
or U29759 (N_29759,N_24141,N_26735);
xnor U29760 (N_29760,N_24680,N_25680);
and U29761 (N_29761,N_26222,N_24768);
nor U29762 (N_29762,N_26977,N_24169);
and U29763 (N_29763,N_25320,N_25814);
and U29764 (N_29764,N_25194,N_25477);
or U29765 (N_29765,N_26111,N_24905);
nand U29766 (N_29766,N_26623,N_26040);
xnor U29767 (N_29767,N_25250,N_24737);
and U29768 (N_29768,N_24005,N_25356);
nand U29769 (N_29769,N_24192,N_24128);
xor U29770 (N_29770,N_26140,N_25412);
nand U29771 (N_29771,N_26405,N_24994);
or U29772 (N_29772,N_24837,N_26202);
nor U29773 (N_29773,N_24671,N_25339);
nand U29774 (N_29774,N_24086,N_24029);
or U29775 (N_29775,N_26637,N_25387);
nor U29776 (N_29776,N_25568,N_24649);
xor U29777 (N_29777,N_25697,N_25916);
and U29778 (N_29778,N_25297,N_24262);
or U29779 (N_29779,N_26084,N_24235);
and U29780 (N_29780,N_26043,N_26694);
and U29781 (N_29781,N_26561,N_25456);
nand U29782 (N_29782,N_26086,N_26385);
or U29783 (N_29783,N_26019,N_26280);
nor U29784 (N_29784,N_25254,N_24736);
or U29785 (N_29785,N_25735,N_24338);
or U29786 (N_29786,N_25068,N_25292);
and U29787 (N_29787,N_25663,N_25158);
xor U29788 (N_29788,N_25554,N_24962);
or U29789 (N_29789,N_25707,N_24964);
or U29790 (N_29790,N_25334,N_25595);
nor U29791 (N_29791,N_26569,N_24408);
nand U29792 (N_29792,N_26055,N_26464);
nand U29793 (N_29793,N_24335,N_25580);
and U29794 (N_29794,N_26993,N_25241);
nand U29795 (N_29795,N_25496,N_24765);
or U29796 (N_29796,N_26828,N_25374);
or U29797 (N_29797,N_25822,N_25560);
or U29798 (N_29798,N_24642,N_24991);
xor U29799 (N_29799,N_26159,N_24824);
nor U29800 (N_29800,N_25963,N_26636);
and U29801 (N_29801,N_24937,N_24332);
nor U29802 (N_29802,N_24894,N_26017);
nor U29803 (N_29803,N_26997,N_24284);
xnor U29804 (N_29804,N_25289,N_26141);
nand U29805 (N_29805,N_25833,N_24636);
nor U29806 (N_29806,N_26978,N_26690);
nor U29807 (N_29807,N_26584,N_26415);
and U29808 (N_29808,N_26260,N_26874);
xor U29809 (N_29809,N_24153,N_25725);
nor U29810 (N_29810,N_26767,N_26904);
nor U29811 (N_29811,N_26112,N_26350);
xnor U29812 (N_29812,N_25853,N_25701);
xor U29813 (N_29813,N_25596,N_25494);
or U29814 (N_29814,N_25488,N_24603);
nor U29815 (N_29815,N_26451,N_25998);
or U29816 (N_29816,N_24448,N_25634);
and U29817 (N_29817,N_25767,N_25718);
xnor U29818 (N_29818,N_25178,N_26694);
nor U29819 (N_29819,N_24877,N_25061);
or U29820 (N_29820,N_24760,N_24607);
nor U29821 (N_29821,N_26045,N_24001);
or U29822 (N_29822,N_26037,N_24854);
nand U29823 (N_29823,N_25431,N_25885);
or U29824 (N_29824,N_25047,N_24673);
or U29825 (N_29825,N_24027,N_24871);
xnor U29826 (N_29826,N_24038,N_24134);
nand U29827 (N_29827,N_26702,N_24679);
and U29828 (N_29828,N_25079,N_25513);
nor U29829 (N_29829,N_24818,N_25545);
xor U29830 (N_29830,N_26188,N_26012);
nand U29831 (N_29831,N_24232,N_25654);
or U29832 (N_29832,N_25388,N_25408);
xnor U29833 (N_29833,N_24775,N_25078);
nand U29834 (N_29834,N_26968,N_25771);
nand U29835 (N_29835,N_25162,N_26783);
xnor U29836 (N_29836,N_24050,N_25087);
or U29837 (N_29837,N_24759,N_26362);
nor U29838 (N_29838,N_26759,N_26610);
nand U29839 (N_29839,N_25094,N_25021);
xnor U29840 (N_29840,N_26543,N_24028);
and U29841 (N_29841,N_26599,N_26441);
xor U29842 (N_29842,N_26372,N_24662);
nand U29843 (N_29843,N_25118,N_26702);
nand U29844 (N_29844,N_24041,N_26440);
nand U29845 (N_29845,N_24822,N_25451);
and U29846 (N_29846,N_24497,N_24674);
nor U29847 (N_29847,N_24407,N_26528);
nor U29848 (N_29848,N_24466,N_25532);
nand U29849 (N_29849,N_26178,N_26569);
and U29850 (N_29850,N_26110,N_24180);
or U29851 (N_29851,N_25419,N_26260);
xor U29852 (N_29852,N_26949,N_25486);
or U29853 (N_29853,N_25845,N_26683);
or U29854 (N_29854,N_24592,N_24291);
nand U29855 (N_29855,N_24188,N_26852);
xor U29856 (N_29856,N_26069,N_25645);
and U29857 (N_29857,N_25536,N_24951);
nor U29858 (N_29858,N_24845,N_24185);
xor U29859 (N_29859,N_25872,N_24776);
or U29860 (N_29860,N_25256,N_24274);
nor U29861 (N_29861,N_26085,N_26123);
nor U29862 (N_29862,N_24581,N_25337);
and U29863 (N_29863,N_24859,N_24056);
nor U29864 (N_29864,N_26419,N_26108);
xor U29865 (N_29865,N_26172,N_24383);
nor U29866 (N_29866,N_25160,N_25193);
xnor U29867 (N_29867,N_24496,N_24115);
and U29868 (N_29868,N_26827,N_26986);
or U29869 (N_29869,N_26831,N_25483);
nand U29870 (N_29870,N_24524,N_26671);
or U29871 (N_29871,N_25155,N_24596);
nand U29872 (N_29872,N_24535,N_26417);
and U29873 (N_29873,N_26028,N_24867);
nor U29874 (N_29874,N_26870,N_24848);
and U29875 (N_29875,N_24042,N_24220);
nor U29876 (N_29876,N_26369,N_24782);
xnor U29877 (N_29877,N_25077,N_25671);
nand U29878 (N_29878,N_24365,N_25321);
or U29879 (N_29879,N_26804,N_24230);
xnor U29880 (N_29880,N_25876,N_25084);
nor U29881 (N_29881,N_24598,N_25956);
and U29882 (N_29882,N_24879,N_26568);
and U29883 (N_29883,N_24234,N_25340);
xor U29884 (N_29884,N_26142,N_26928);
nor U29885 (N_29885,N_25727,N_24338);
nor U29886 (N_29886,N_26426,N_24849);
nand U29887 (N_29887,N_24631,N_24371);
nand U29888 (N_29888,N_24973,N_25328);
xor U29889 (N_29889,N_24747,N_25384);
nand U29890 (N_29890,N_26466,N_26168);
xor U29891 (N_29891,N_25869,N_26630);
nand U29892 (N_29892,N_26284,N_25392);
and U29893 (N_29893,N_25558,N_25343);
nor U29894 (N_29894,N_26577,N_24193);
nand U29895 (N_29895,N_25834,N_26677);
nor U29896 (N_29896,N_25172,N_24024);
xor U29897 (N_29897,N_24143,N_24943);
or U29898 (N_29898,N_25377,N_26794);
and U29899 (N_29899,N_26566,N_26561);
and U29900 (N_29900,N_24930,N_26674);
xnor U29901 (N_29901,N_24539,N_24524);
or U29902 (N_29902,N_26608,N_24443);
nor U29903 (N_29903,N_24309,N_26369);
nor U29904 (N_29904,N_24483,N_25077);
and U29905 (N_29905,N_24556,N_25900);
nand U29906 (N_29906,N_26115,N_24760);
nand U29907 (N_29907,N_25306,N_25614);
xnor U29908 (N_29908,N_24449,N_24361);
or U29909 (N_29909,N_26858,N_26516);
nor U29910 (N_29910,N_24007,N_24421);
and U29911 (N_29911,N_26739,N_26196);
xnor U29912 (N_29912,N_25081,N_24315);
nor U29913 (N_29913,N_26700,N_25541);
nor U29914 (N_29914,N_26195,N_26965);
xnor U29915 (N_29915,N_24756,N_24339);
or U29916 (N_29916,N_24090,N_25967);
xnor U29917 (N_29917,N_25897,N_25249);
or U29918 (N_29918,N_25586,N_25681);
xnor U29919 (N_29919,N_26918,N_25178);
and U29920 (N_29920,N_26694,N_26854);
nor U29921 (N_29921,N_26757,N_25714);
nand U29922 (N_29922,N_24048,N_26894);
nand U29923 (N_29923,N_24128,N_26159);
or U29924 (N_29924,N_25511,N_26171);
nand U29925 (N_29925,N_25694,N_26233);
nand U29926 (N_29926,N_24750,N_24690);
and U29927 (N_29927,N_26507,N_24326);
nor U29928 (N_29928,N_25112,N_25561);
xnor U29929 (N_29929,N_26745,N_26765);
xnor U29930 (N_29930,N_26848,N_24086);
nor U29931 (N_29931,N_25606,N_25930);
nor U29932 (N_29932,N_25699,N_26357);
xnor U29933 (N_29933,N_25689,N_24508);
nand U29934 (N_29934,N_26556,N_25730);
or U29935 (N_29935,N_24447,N_25536);
nor U29936 (N_29936,N_25165,N_24131);
nand U29937 (N_29937,N_25301,N_24886);
nor U29938 (N_29938,N_25892,N_25419);
and U29939 (N_29939,N_24696,N_26397);
or U29940 (N_29940,N_26462,N_25563);
and U29941 (N_29941,N_26965,N_25169);
nor U29942 (N_29942,N_24515,N_26100);
or U29943 (N_29943,N_24137,N_24287);
nor U29944 (N_29944,N_26554,N_26997);
xor U29945 (N_29945,N_24672,N_26307);
nor U29946 (N_29946,N_24206,N_24007);
nand U29947 (N_29947,N_25356,N_26656);
xor U29948 (N_29948,N_24619,N_25391);
nor U29949 (N_29949,N_24092,N_26217);
xnor U29950 (N_29950,N_25812,N_24859);
nor U29951 (N_29951,N_24106,N_24268);
or U29952 (N_29952,N_26974,N_25699);
nor U29953 (N_29953,N_25509,N_24839);
nor U29954 (N_29954,N_26956,N_26829);
nand U29955 (N_29955,N_25755,N_24072);
nand U29956 (N_29956,N_25394,N_25490);
or U29957 (N_29957,N_24149,N_24054);
and U29958 (N_29958,N_24895,N_25090);
xor U29959 (N_29959,N_25702,N_25097);
xnor U29960 (N_29960,N_25091,N_25688);
nand U29961 (N_29961,N_24151,N_26331);
nor U29962 (N_29962,N_25516,N_24862);
xor U29963 (N_29963,N_25345,N_25495);
nor U29964 (N_29964,N_24495,N_26304);
xor U29965 (N_29965,N_26847,N_25758);
and U29966 (N_29966,N_26739,N_25811);
and U29967 (N_29967,N_25984,N_26223);
nor U29968 (N_29968,N_24061,N_24265);
nand U29969 (N_29969,N_24004,N_25778);
nand U29970 (N_29970,N_26200,N_24360);
nor U29971 (N_29971,N_26836,N_25669);
nand U29972 (N_29972,N_25083,N_25390);
nand U29973 (N_29973,N_26617,N_26302);
or U29974 (N_29974,N_26107,N_24989);
nor U29975 (N_29975,N_24501,N_25446);
nand U29976 (N_29976,N_26507,N_24325);
nor U29977 (N_29977,N_26174,N_25232);
nand U29978 (N_29978,N_26732,N_25072);
nand U29979 (N_29979,N_26084,N_24352);
or U29980 (N_29980,N_26532,N_25019);
nand U29981 (N_29981,N_25063,N_26238);
or U29982 (N_29982,N_26421,N_25586);
nor U29983 (N_29983,N_26295,N_25420);
xnor U29984 (N_29984,N_26454,N_24973);
nand U29985 (N_29985,N_26350,N_25286);
xor U29986 (N_29986,N_26138,N_25567);
nand U29987 (N_29987,N_24701,N_26806);
nand U29988 (N_29988,N_26022,N_25874);
nand U29989 (N_29989,N_24621,N_26356);
nand U29990 (N_29990,N_25217,N_25205);
and U29991 (N_29991,N_24850,N_24374);
nor U29992 (N_29992,N_25768,N_25095);
and U29993 (N_29993,N_26443,N_25981);
nand U29994 (N_29994,N_26366,N_26904);
nand U29995 (N_29995,N_25728,N_26078);
xnor U29996 (N_29996,N_24930,N_26120);
xor U29997 (N_29997,N_24586,N_25651);
and U29998 (N_29998,N_25284,N_26466);
xnor U29999 (N_29999,N_24403,N_26153);
nor UO_0 (O_0,N_29110,N_28673);
and UO_1 (O_1,N_28222,N_29898);
xnor UO_2 (O_2,N_28899,N_27986);
nor UO_3 (O_3,N_27051,N_28060);
nor UO_4 (O_4,N_28982,N_27730);
and UO_5 (O_5,N_27486,N_29504);
nor UO_6 (O_6,N_29880,N_27722);
or UO_7 (O_7,N_29402,N_29695);
nand UO_8 (O_8,N_27893,N_29046);
nor UO_9 (O_9,N_29177,N_27620);
or UO_10 (O_10,N_28170,N_29420);
xor UO_11 (O_11,N_27152,N_27208);
nand UO_12 (O_12,N_29203,N_29915);
and UO_13 (O_13,N_27126,N_28489);
nand UO_14 (O_14,N_27200,N_27279);
nor UO_15 (O_15,N_27170,N_27876);
or UO_16 (O_16,N_29388,N_29316);
or UO_17 (O_17,N_29913,N_27927);
nor UO_18 (O_18,N_28200,N_27463);
nand UO_19 (O_19,N_27064,N_28439);
nand UO_20 (O_20,N_27540,N_29395);
xnor UO_21 (O_21,N_29999,N_27036);
and UO_22 (O_22,N_28594,N_27163);
nor UO_23 (O_23,N_27456,N_28580);
nand UO_24 (O_24,N_29277,N_28588);
nor UO_25 (O_25,N_28452,N_27910);
or UO_26 (O_26,N_28744,N_27470);
and UO_27 (O_27,N_29372,N_28967);
or UO_28 (O_28,N_28848,N_29176);
nor UO_29 (O_29,N_27849,N_28813);
nand UO_30 (O_30,N_28742,N_27076);
or UO_31 (O_31,N_28267,N_29934);
xnor UO_32 (O_32,N_29831,N_27184);
or UO_33 (O_33,N_29047,N_27260);
or UO_34 (O_34,N_29423,N_28649);
nand UO_35 (O_35,N_27637,N_27975);
xor UO_36 (O_36,N_29692,N_27443);
or UO_37 (O_37,N_28665,N_28701);
nor UO_38 (O_38,N_29171,N_27274);
nand UO_39 (O_39,N_27179,N_29376);
or UO_40 (O_40,N_28343,N_27324);
or UO_41 (O_41,N_27081,N_27994);
and UO_42 (O_42,N_29178,N_28781);
and UO_43 (O_43,N_28191,N_27901);
nor UO_44 (O_44,N_29845,N_29725);
nand UO_45 (O_45,N_27804,N_28412);
or UO_46 (O_46,N_27531,N_29606);
and UO_47 (O_47,N_27723,N_28745);
nor UO_48 (O_48,N_29299,N_28415);
nor UO_49 (O_49,N_28668,N_27213);
xor UO_50 (O_50,N_29335,N_27414);
nand UO_51 (O_51,N_28463,N_28532);
and UO_52 (O_52,N_27845,N_29525);
xnor UO_53 (O_53,N_29529,N_27916);
nor UO_54 (O_54,N_29200,N_29717);
and UO_55 (O_55,N_29647,N_27333);
or UO_56 (O_56,N_28359,N_28315);
and UO_57 (O_57,N_28661,N_28909);
or UO_58 (O_58,N_27570,N_28888);
nor UO_59 (O_59,N_29865,N_29422);
nand UO_60 (O_60,N_29764,N_29303);
nor UO_61 (O_61,N_28945,N_29440);
nor UO_62 (O_62,N_29615,N_28783);
or UO_63 (O_63,N_27968,N_29225);
nor UO_64 (O_64,N_29539,N_29071);
and UO_65 (O_65,N_27568,N_29685);
or UO_66 (O_66,N_29911,N_28239);
xnor UO_67 (O_67,N_29001,N_29494);
xnor UO_68 (O_68,N_28876,N_27834);
and UO_69 (O_69,N_27792,N_27817);
and UO_70 (O_70,N_27437,N_29327);
and UO_71 (O_71,N_28894,N_29951);
xnor UO_72 (O_72,N_28216,N_29584);
nor UO_73 (O_73,N_27614,N_27041);
or UO_74 (O_74,N_27821,N_29863);
xor UO_75 (O_75,N_28131,N_29321);
xor UO_76 (O_76,N_27546,N_27543);
nor UO_77 (O_77,N_27815,N_28006);
xor UO_78 (O_78,N_28423,N_29519);
nor UO_79 (O_79,N_27692,N_29229);
nor UO_80 (O_80,N_29445,N_27832);
nor UO_81 (O_81,N_29185,N_29527);
xor UO_82 (O_82,N_28393,N_27493);
nor UO_83 (O_83,N_28310,N_28160);
nand UO_84 (O_84,N_27079,N_27471);
xnor UO_85 (O_85,N_29884,N_29318);
nor UO_86 (O_86,N_28620,N_29645);
xor UO_87 (O_87,N_27572,N_28853);
xor UO_88 (O_88,N_27118,N_29594);
nor UO_89 (O_89,N_28571,N_29574);
nor UO_90 (O_90,N_27077,N_27226);
nand UO_91 (O_91,N_28126,N_28688);
and UO_92 (O_92,N_29389,N_27367);
or UO_93 (O_93,N_29595,N_29686);
nand UO_94 (O_94,N_27631,N_27703);
nand UO_95 (O_95,N_29187,N_28047);
or UO_96 (O_96,N_28923,N_27453);
and UO_97 (O_97,N_28291,N_28054);
xor UO_98 (O_98,N_27518,N_29380);
and UO_99 (O_99,N_27830,N_28318);
and UO_100 (O_100,N_28065,N_28406);
nor UO_101 (O_101,N_28019,N_27833);
xnor UO_102 (O_102,N_29867,N_28547);
nand UO_103 (O_103,N_29995,N_28007);
nand UO_104 (O_104,N_29705,N_29446);
nand UO_105 (O_105,N_28572,N_27672);
and UO_106 (O_106,N_29320,N_27828);
or UO_107 (O_107,N_29699,N_28248);
xor UO_108 (O_108,N_29065,N_27819);
xnor UO_109 (O_109,N_28598,N_27303);
xor UO_110 (O_110,N_27252,N_28378);
or UO_111 (O_111,N_28635,N_27446);
or UO_112 (O_112,N_27476,N_29363);
nand UO_113 (O_113,N_27482,N_29581);
or UO_114 (O_114,N_29561,N_28893);
nand UO_115 (O_115,N_29862,N_28785);
and UO_116 (O_116,N_28313,N_27108);
and UO_117 (O_117,N_28187,N_28186);
nor UO_118 (O_118,N_28583,N_29718);
nand UO_119 (O_119,N_28308,N_29608);
nor UO_120 (O_120,N_29554,N_29360);
nor UO_121 (O_121,N_28995,N_29112);
and UO_122 (O_122,N_27043,N_28787);
xor UO_123 (O_123,N_27773,N_28613);
or UO_124 (O_124,N_29752,N_28618);
and UO_125 (O_125,N_28137,N_28014);
and UO_126 (O_126,N_28907,N_27989);
nor UO_127 (O_127,N_27805,N_28684);
and UO_128 (O_128,N_27014,N_29450);
xor UO_129 (O_129,N_28669,N_28299);
xnor UO_130 (O_130,N_29710,N_27313);
nor UO_131 (O_131,N_27988,N_28775);
and UO_132 (O_132,N_29116,N_29905);
and UO_133 (O_133,N_27566,N_27537);
xor UO_134 (O_134,N_27534,N_28424);
xor UO_135 (O_135,N_29501,N_29691);
xnor UO_136 (O_136,N_28537,N_29459);
nand UO_137 (O_137,N_29713,N_29920);
and UO_138 (O_138,N_27510,N_29857);
or UO_139 (O_139,N_27438,N_29025);
xor UO_140 (O_140,N_27706,N_28244);
nor UO_141 (O_141,N_27924,N_29707);
and UO_142 (O_142,N_29728,N_27281);
and UO_143 (O_143,N_27030,N_29137);
or UO_144 (O_144,N_29205,N_29131);
or UO_145 (O_145,N_27061,N_29899);
xor UO_146 (O_146,N_29506,N_29179);
nand UO_147 (O_147,N_29281,N_29304);
xnor UO_148 (O_148,N_27465,N_28324);
or UO_149 (O_149,N_28402,N_28646);
xnor UO_150 (O_150,N_27445,N_27549);
nand UO_151 (O_151,N_27584,N_29997);
xnor UO_152 (O_152,N_29133,N_29503);
nand UO_153 (O_153,N_27981,N_28314);
xnor UO_154 (O_154,N_29596,N_28386);
xnor UO_155 (O_155,N_29130,N_29088);
and UO_156 (O_156,N_29773,N_27604);
and UO_157 (O_157,N_27195,N_28487);
nor UO_158 (O_158,N_28297,N_29429);
nand UO_159 (O_159,N_27073,N_27530);
xnor UO_160 (O_160,N_29268,N_27918);
nor UO_161 (O_161,N_27268,N_28912);
and UO_162 (O_162,N_28838,N_27746);
xnor UO_163 (O_163,N_29602,N_28431);
and UO_164 (O_164,N_29684,N_28334);
or UO_165 (O_165,N_29356,N_29151);
nor UO_166 (O_166,N_29086,N_28805);
and UO_167 (O_167,N_27411,N_29148);
xor UO_168 (O_168,N_28855,N_28056);
nand UO_169 (O_169,N_28215,N_27273);
xnor UO_170 (O_170,N_27002,N_27171);
or UO_171 (O_171,N_29127,N_29122);
nand UO_172 (O_172,N_28440,N_27348);
xor UO_173 (O_173,N_29374,N_27858);
xnor UO_174 (O_174,N_28005,N_29084);
and UO_175 (O_175,N_28260,N_29189);
xnor UO_176 (O_176,N_28333,N_28933);
or UO_177 (O_177,N_29157,N_28063);
xor UO_178 (O_178,N_27949,N_28189);
nand UO_179 (O_179,N_28540,N_29948);
or UO_180 (O_180,N_27814,N_27410);
xor UO_181 (O_181,N_27305,N_29550);
or UO_182 (O_182,N_28766,N_27952);
or UO_183 (O_183,N_29531,N_27272);
nor UO_184 (O_184,N_27104,N_29285);
nor UO_185 (O_185,N_29023,N_27478);
xnor UO_186 (O_186,N_29230,N_27287);
nand UO_187 (O_187,N_28573,N_28528);
and UO_188 (O_188,N_27444,N_27450);
or UO_189 (O_189,N_29985,N_29201);
and UO_190 (O_190,N_29246,N_28699);
and UO_191 (O_191,N_28714,N_28847);
xor UO_192 (O_192,N_29106,N_28416);
nor UO_193 (O_193,N_28003,N_27498);
or UO_194 (O_194,N_28103,N_27078);
or UO_195 (O_195,N_29342,N_28685);
or UO_196 (O_196,N_29368,N_27701);
or UO_197 (O_197,N_27965,N_28567);
nor UO_198 (O_198,N_27366,N_27027);
nand UO_199 (O_199,N_29290,N_27236);
and UO_200 (O_200,N_28413,N_28789);
and UO_201 (O_201,N_29099,N_29977);
nand UO_202 (O_202,N_27275,N_27033);
nand UO_203 (O_203,N_27539,N_29590);
nand UO_204 (O_204,N_27661,N_29734);
or UO_205 (O_205,N_27558,N_29015);
nand UO_206 (O_206,N_29297,N_29258);
nor UO_207 (O_207,N_27675,N_28767);
xor UO_208 (O_208,N_28071,N_28551);
xnor UO_209 (O_209,N_28691,N_29757);
nand UO_210 (O_210,N_27882,N_28041);
or UO_211 (O_211,N_28417,N_27159);
xor UO_212 (O_212,N_29377,N_27899);
and UO_213 (O_213,N_27325,N_29618);
and UO_214 (O_214,N_27824,N_28199);
and UO_215 (O_215,N_29500,N_28956);
nand UO_216 (O_216,N_28459,N_29700);
and UO_217 (O_217,N_27978,N_27392);
xor UO_218 (O_218,N_28905,N_29220);
xor UO_219 (O_219,N_29719,N_28761);
xnor UO_220 (O_220,N_28686,N_29243);
and UO_221 (O_221,N_27067,N_28364);
and UO_222 (O_222,N_29777,N_28279);
nor UO_223 (O_223,N_29944,N_28846);
and UO_224 (O_224,N_29996,N_29628);
nand UO_225 (O_225,N_28536,N_29149);
or UO_226 (O_226,N_29808,N_28389);
nor UO_227 (O_227,N_28960,N_28175);
and UO_228 (O_228,N_29776,N_28095);
xnor UO_229 (O_229,N_29090,N_29159);
or UO_230 (O_230,N_28645,N_27563);
xor UO_231 (O_231,N_29639,N_29624);
nor UO_232 (O_232,N_29903,N_27137);
or UO_233 (O_233,N_29658,N_29031);
nand UO_234 (O_234,N_28653,N_28827);
or UO_235 (O_235,N_29465,N_29016);
nor UO_236 (O_236,N_28350,N_28173);
and UO_237 (O_237,N_28721,N_27875);
and UO_238 (O_238,N_27435,N_29682);
or UO_239 (O_239,N_29330,N_29505);
nand UO_240 (O_240,N_29917,N_29732);
xor UO_241 (O_241,N_29417,N_29787);
or UO_242 (O_242,N_28149,N_28689);
nor UO_243 (O_243,N_27642,N_29011);
xnor UO_244 (O_244,N_28821,N_28422);
and UO_245 (O_245,N_29514,N_29952);
and UO_246 (O_246,N_29066,N_29902);
nand UO_247 (O_247,N_28471,N_29694);
or UO_248 (O_248,N_28290,N_29912);
nor UO_249 (O_249,N_29266,N_29984);
nor UO_250 (O_250,N_28480,N_29708);
xor UO_251 (O_251,N_28832,N_28032);
and UO_252 (O_252,N_28533,N_28446);
nand UO_253 (O_253,N_27726,N_29324);
or UO_254 (O_254,N_28400,N_27688);
or UO_255 (O_255,N_29562,N_27685);
nor UO_256 (O_256,N_29462,N_28401);
nand UO_257 (O_257,N_29154,N_28954);
nor UO_258 (O_258,N_28118,N_28702);
xnor UO_259 (O_259,N_27071,N_28205);
or UO_260 (O_260,N_29323,N_28811);
or UO_261 (O_261,N_27878,N_27094);
nor UO_262 (O_262,N_27113,N_29730);
xor UO_263 (O_263,N_27358,N_27283);
and UO_264 (O_264,N_28859,N_27863);
nor UO_265 (O_265,N_29126,N_29235);
and UO_266 (O_266,N_28079,N_29345);
and UO_267 (O_267,N_29021,N_29916);
nor UO_268 (O_268,N_27120,N_29383);
nand UO_269 (O_269,N_29488,N_28085);
xor UO_270 (O_270,N_29928,N_27255);
and UO_271 (O_271,N_29400,N_27948);
xnor UO_272 (O_272,N_27601,N_28615);
or UO_273 (O_273,N_28419,N_28771);
nor UO_274 (O_274,N_28106,N_29766);
nor UO_275 (O_275,N_27295,N_28915);
nor UO_276 (O_276,N_28100,N_28352);
and UO_277 (O_277,N_27095,N_27848);
or UO_278 (O_278,N_28753,N_27473);
nand UO_279 (O_279,N_27502,N_29314);
xnor UO_280 (O_280,N_29036,N_27810);
or UO_281 (O_281,N_29767,N_27117);
or UO_282 (O_282,N_27775,N_29118);
nand UO_283 (O_283,N_27785,N_27233);
xnor UO_284 (O_284,N_28347,N_27951);
or UO_285 (O_285,N_27322,N_28449);
nand UO_286 (O_286,N_28433,N_28479);
or UO_287 (O_287,N_28790,N_27182);
and UO_288 (O_288,N_27280,N_29536);
nor UO_289 (O_289,N_27732,N_29067);
or UO_290 (O_290,N_27559,N_28969);
and UO_291 (O_291,N_28942,N_29035);
nor UO_292 (O_292,N_27423,N_28751);
nor UO_293 (O_293,N_29929,N_27944);
nand UO_294 (O_294,N_28800,N_27700);
nand UO_295 (O_295,N_28822,N_28037);
nand UO_296 (O_296,N_28087,N_28955);
or UO_297 (O_297,N_27576,N_27603);
and UO_298 (O_298,N_27357,N_29978);
nand UO_299 (O_299,N_29901,N_27351);
and UO_300 (O_300,N_28365,N_29540);
and UO_301 (O_301,N_28834,N_28112);
or UO_302 (O_302,N_27447,N_28280);
nor UO_303 (O_303,N_27232,N_27044);
nand UO_304 (O_304,N_29315,N_27336);
or UO_305 (O_305,N_27711,N_28602);
and UO_306 (O_306,N_28704,N_27683);
nand UO_307 (O_307,N_29262,N_29742);
or UO_308 (O_308,N_27598,N_28801);
nor UO_309 (O_309,N_27632,N_27749);
or UO_310 (O_310,N_27579,N_28523);
nor UO_311 (O_311,N_28733,N_27135);
nor UO_312 (O_312,N_27408,N_27983);
or UO_313 (O_313,N_27271,N_27215);
or UO_314 (O_314,N_27887,N_28990);
xnor UO_315 (O_315,N_29816,N_27640);
and UO_316 (O_316,N_28937,N_29257);
or UO_317 (O_317,N_29336,N_29559);
xor UO_318 (O_318,N_29333,N_29308);
or UO_319 (O_319,N_29829,N_28287);
nor UO_320 (O_320,N_29869,N_27102);
nor UO_321 (O_321,N_28709,N_28303);
nor UO_322 (O_322,N_28376,N_27340);
nand UO_323 (O_323,N_29100,N_29399);
nand UO_324 (O_324,N_27448,N_29190);
xnor UO_325 (O_325,N_28329,N_29089);
or UO_326 (O_326,N_28717,N_29234);
or UO_327 (O_327,N_28803,N_28275);
or UO_328 (O_328,N_27254,N_28575);
nand UO_329 (O_329,N_27883,N_28695);
xnor UO_330 (O_330,N_29104,N_27143);
and UO_331 (O_331,N_29347,N_28251);
or UO_332 (O_332,N_28289,N_29723);
and UO_333 (O_333,N_29238,N_27263);
or UO_334 (O_334,N_28693,N_29761);
and UO_335 (O_335,N_29775,N_27580);
and UO_336 (O_336,N_29407,N_29976);
and UO_337 (O_337,N_28786,N_28232);
or UO_338 (O_338,N_27211,N_28099);
xnor UO_339 (O_339,N_29212,N_27713);
or UO_340 (O_340,N_28619,N_27057);
nor UO_341 (O_341,N_28256,N_28860);
or UO_342 (O_342,N_29936,N_29969);
xnor UO_343 (O_343,N_28578,N_29398);
nand UO_344 (O_344,N_29659,N_28158);
or UO_345 (O_345,N_27181,N_28243);
xnor UO_346 (O_346,N_29874,N_28074);
or UO_347 (O_347,N_28478,N_29836);
and UO_348 (O_348,N_28388,N_29250);
xnor UO_349 (O_349,N_27622,N_29599);
and UO_350 (O_350,N_27220,N_27925);
or UO_351 (O_351,N_27237,N_27926);
nand UO_352 (O_352,N_27240,N_29741);
and UO_353 (O_353,N_28913,N_27130);
xor UO_354 (O_354,N_27318,N_27866);
xnor UO_355 (O_355,N_27720,N_29312);
or UO_356 (O_356,N_28295,N_28760);
and UO_357 (O_357,N_29019,N_28869);
nand UO_358 (O_358,N_29319,N_27754);
and UO_359 (O_359,N_29340,N_28294);
xnor UO_360 (O_360,N_27147,N_27401);
or UO_361 (O_361,N_27393,N_29068);
nor UO_362 (O_362,N_28252,N_27072);
and UO_363 (O_363,N_27767,N_29875);
xor UO_364 (O_364,N_27452,N_27793);
nor UO_365 (O_365,N_27103,N_27600);
nand UO_366 (O_366,N_28096,N_28421);
xnor UO_367 (O_367,N_29577,N_27852);
xor UO_368 (O_368,N_28652,N_29772);
nand UO_369 (O_369,N_29676,N_29961);
xnor UO_370 (O_370,N_27124,N_29269);
and UO_371 (O_371,N_29150,N_27835);
xor UO_372 (O_372,N_29062,N_28762);
and UO_373 (O_373,N_29716,N_28698);
or UO_374 (O_374,N_27514,N_28824);
xnor UO_375 (O_375,N_27046,N_29560);
and UO_376 (O_376,N_28127,N_27122);
xor UO_377 (O_377,N_28513,N_29393);
xnor UO_378 (O_378,N_27455,N_27731);
and UO_379 (O_379,N_29800,N_28975);
or UO_380 (O_380,N_27363,N_27062);
and UO_381 (O_381,N_27947,N_29251);
and UO_382 (O_382,N_29231,N_28778);
or UO_383 (O_383,N_27180,N_29956);
xor UO_384 (O_384,N_28012,N_28468);
or UO_385 (O_385,N_27854,N_29334);
nand UO_386 (O_386,N_27157,N_28107);
xnor UO_387 (O_387,N_27856,N_28872);
xnor UO_388 (O_388,N_27187,N_28732);
nor UO_389 (O_389,N_29704,N_28076);
nor UO_390 (O_390,N_27302,N_27466);
xor UO_391 (O_391,N_29288,N_27016);
or UO_392 (O_392,N_29744,N_27290);
xnor UO_393 (O_393,N_29582,N_28504);
nand UO_394 (O_394,N_29102,N_27705);
xor UO_395 (O_395,N_27991,N_27651);
nor UO_396 (O_396,N_27140,N_29939);
and UO_397 (O_397,N_29910,N_28736);
and UO_398 (O_398,N_29515,N_27996);
or UO_399 (O_399,N_28181,N_29853);
xor UO_400 (O_400,N_28068,N_29381);
xor UO_401 (O_401,N_28934,N_27052);
nor UO_402 (O_402,N_29408,N_29292);
nand UO_403 (O_403,N_28238,N_29498);
nand UO_404 (O_404,N_27436,N_27574);
nand UO_405 (O_405,N_28283,N_27054);
nor UO_406 (O_406,N_29635,N_29240);
nand UO_407 (O_407,N_27299,N_28823);
nand UO_408 (O_408,N_29825,N_28162);
or UO_409 (O_409,N_29548,N_29897);
nand UO_410 (O_410,N_29282,N_28470);
nand UO_411 (O_411,N_29534,N_27578);
and UO_412 (O_412,N_27250,N_28520);
and UO_413 (O_413,N_29485,N_29932);
nand UO_414 (O_414,N_27507,N_29010);
nor UO_415 (O_415,N_28024,N_29632);
nor UO_416 (O_416,N_27868,N_27082);
or UO_417 (O_417,N_27591,N_29894);
nand UO_418 (O_418,N_28121,N_28209);
nor UO_419 (O_419,N_28984,N_29696);
or UO_420 (O_420,N_28552,N_28502);
nand UO_421 (O_421,N_29366,N_28368);
nor UO_422 (O_422,N_27379,N_27128);
or UO_423 (O_423,N_28515,N_29163);
nand UO_424 (O_424,N_28507,N_29747);
nor UO_425 (O_425,N_27904,N_27974);
and UO_426 (O_426,N_28179,N_27425);
nand UO_427 (O_427,N_28172,N_27842);
or UO_428 (O_428,N_27013,N_28151);
nand UO_429 (O_429,N_28219,N_27586);
and UO_430 (O_430,N_27555,N_29538);
xnor UO_431 (O_431,N_29702,N_28606);
nor UO_432 (O_432,N_28857,N_28569);
xor UO_433 (O_433,N_27429,N_28772);
nor UO_434 (O_434,N_28815,N_28554);
nor UO_435 (O_435,N_27010,N_28974);
and UO_436 (O_436,N_29522,N_27345);
or UO_437 (O_437,N_28875,N_28867);
xor UO_438 (O_438,N_27310,N_29057);
xnor UO_439 (O_439,N_29410,N_28946);
nor UO_440 (O_440,N_29173,N_27234);
nand UO_441 (O_441,N_29868,N_29332);
nor UO_442 (O_442,N_27323,N_29837);
xor UO_443 (O_443,N_28488,N_28462);
nand UO_444 (O_444,N_28730,N_29481);
or UO_445 (O_445,N_27206,N_29672);
or UO_446 (O_446,N_28426,N_27747);
nor UO_447 (O_447,N_29169,N_27554);
or UO_448 (O_448,N_27733,N_29338);
nand UO_449 (O_449,N_28769,N_28676);
or UO_450 (O_450,N_28548,N_28804);
nor UO_451 (O_451,N_29779,N_28999);
or UO_452 (O_452,N_28113,N_29247);
xor UO_453 (O_453,N_29495,N_29771);
and UO_454 (O_454,N_28675,N_28261);
nand UO_455 (O_455,N_29714,N_29499);
nor UO_456 (O_456,N_27488,N_28935);
xnor UO_457 (O_457,N_27116,N_27162);
or UO_458 (O_458,N_28114,N_29487);
nor UO_459 (O_459,N_29475,N_28941);
and UO_460 (O_460,N_28963,N_29824);
and UO_461 (O_461,N_27816,N_28657);
nor UO_462 (O_462,N_28779,N_27647);
and UO_463 (O_463,N_27442,N_27099);
nand UO_464 (O_464,N_28817,N_27468);
and UO_465 (O_465,N_27355,N_29115);
and UO_466 (O_466,N_29575,N_29186);
or UO_467 (O_467,N_27224,N_27018);
or UO_468 (O_468,N_29619,N_29386);
nand UO_469 (O_469,N_27803,N_28166);
or UO_470 (O_470,N_27686,N_27619);
nand UO_471 (O_471,N_27551,N_28921);
or UO_472 (O_472,N_27676,N_27156);
nor UO_473 (O_473,N_29098,N_29451);
and UO_474 (O_474,N_29063,N_27627);
nor UO_475 (O_475,N_28739,N_28278);
or UO_476 (O_476,N_28473,N_28146);
nor UO_477 (O_477,N_29017,N_27879);
nand UO_478 (O_478,N_29852,N_28756);
and UO_479 (O_479,N_28831,N_27249);
or UO_480 (O_480,N_27007,N_29878);
nand UO_481 (O_481,N_27541,N_28271);
nor UO_482 (O_482,N_29080,N_27296);
or UO_483 (O_483,N_27420,N_27898);
nand UO_484 (O_484,N_28370,N_27025);
nand UO_485 (O_485,N_28241,N_28616);
or UO_486 (O_486,N_27148,N_28784);
nor UO_487 (O_487,N_28381,N_29217);
and UO_488 (O_488,N_27219,N_27264);
nand UO_489 (O_489,N_27090,N_29027);
xor UO_490 (O_490,N_29192,N_28609);
xor UO_491 (O_491,N_29546,N_28020);
and UO_492 (O_492,N_28926,N_28067);
nand UO_493 (O_493,N_28247,N_27964);
nor UO_494 (O_494,N_27520,N_28595);
xor UO_495 (O_495,N_27214,N_27769);
xnor UO_496 (O_496,N_29795,N_28980);
or UO_497 (O_497,N_28994,N_28321);
and UO_498 (O_498,N_27630,N_28511);
nor UO_499 (O_499,N_27693,N_29828);
xnor UO_500 (O_500,N_29182,N_29507);
nand UO_501 (O_501,N_29101,N_29729);
xnor UO_502 (O_502,N_27350,N_27506);
nand UO_503 (O_503,N_28361,N_28622);
or UO_504 (O_504,N_27841,N_28929);
nand UO_505 (O_505,N_27519,N_29322);
nor UO_506 (O_506,N_29083,N_28327);
or UO_507 (O_507,N_27480,N_27462);
xor UO_508 (O_508,N_28670,N_28397);
or UO_509 (O_509,N_29135,N_29138);
nor UO_510 (O_510,N_28667,N_27158);
xnor UO_511 (O_511,N_29832,N_27075);
and UO_512 (O_512,N_28952,N_28549);
or UO_513 (O_513,N_29973,N_28841);
or UO_514 (O_514,N_28125,N_28447);
nand UO_515 (O_515,N_29896,N_29403);
nand UO_516 (O_516,N_29037,N_27458);
or UO_517 (O_517,N_27553,N_28094);
and UO_518 (O_518,N_28521,N_28161);
and UO_519 (O_519,N_28582,N_27781);
xor UO_520 (O_520,N_29387,N_27282);
or UO_521 (O_521,N_28558,N_27394);
xor UO_522 (O_522,N_27011,N_27297);
nand UO_523 (O_523,N_29195,N_28078);
and UO_524 (O_524,N_27101,N_27998);
xnor UO_525 (O_525,N_29349,N_27331);
nand UO_526 (O_526,N_29468,N_28363);
and UO_527 (O_527,N_28214,N_29419);
nand UO_528 (O_528,N_27963,N_29491);
and UO_529 (O_529,N_28040,N_27742);
nand UO_530 (O_530,N_27657,N_27021);
xnor UO_531 (O_531,N_27006,N_29311);
nand UO_532 (O_532,N_29341,N_28164);
and UO_533 (O_533,N_28908,N_29518);
xor UO_534 (O_534,N_28249,N_29156);
and UO_535 (O_535,N_28868,N_28776);
nor UO_536 (O_536,N_28202,N_29166);
or UO_537 (O_537,N_29052,N_29317);
xnor UO_538 (O_538,N_29447,N_28072);
nand UO_539 (O_539,N_27535,N_29449);
or UO_540 (O_540,N_29430,N_27877);
or UO_541 (O_541,N_28155,N_27190);
and UO_542 (O_542,N_27939,N_27851);
xnor UO_543 (O_543,N_27431,N_28375);
or UO_544 (O_544,N_27610,N_27068);
nand UO_545 (O_545,N_29044,N_28264);
nand UO_546 (O_546,N_28250,N_28633);
or UO_547 (O_547,N_29219,N_27903);
or UO_548 (O_548,N_27608,N_27381);
nand UO_549 (O_549,N_29081,N_29587);
and UO_550 (O_550,N_28976,N_27193);
and UO_551 (O_551,N_29191,N_28183);
nand UO_552 (O_552,N_29919,N_29687);
nor UO_553 (O_553,N_28798,N_28052);
xnor UO_554 (O_554,N_27396,N_27251);
nand UO_555 (O_555,N_29076,N_28639);
xnor UO_556 (O_556,N_27623,N_29993);
nand UO_557 (O_557,N_27716,N_27434);
and UO_558 (O_558,N_28996,N_27748);
nand UO_559 (O_559,N_27505,N_29746);
and UO_560 (O_560,N_28840,N_28140);
xor UO_561 (O_561,N_29987,N_29737);
nor UO_562 (O_562,N_29543,N_27384);
or UO_563 (O_563,N_28434,N_28658);
xnor UO_564 (O_564,N_27669,N_27426);
and UO_565 (O_565,N_27405,N_29401);
or UO_566 (O_566,N_29649,N_29535);
nor UO_567 (O_567,N_29119,N_29558);
nand UO_568 (O_568,N_29502,N_27550);
and UO_569 (O_569,N_29456,N_28262);
nor UO_570 (O_570,N_28895,N_29454);
xnor UO_571 (O_571,N_28038,N_27525);
and UO_572 (O_572,N_28405,N_29541);
nand UO_573 (O_573,N_27886,N_27844);
and UO_574 (O_574,N_27668,N_27865);
or UO_575 (O_575,N_29061,N_27421);
and UO_576 (O_576,N_27908,N_29041);
and UO_577 (O_577,N_29160,N_29841);
or UO_578 (O_578,N_29774,N_29123);
xor UO_579 (O_579,N_27618,N_29199);
and UO_580 (O_580,N_28025,N_27613);
nand UO_581 (O_581,N_27504,N_29000);
nand UO_582 (O_582,N_28965,N_28508);
nor UO_583 (O_583,N_28810,N_29600);
nand UO_584 (O_584,N_29680,N_28302);
nand UO_585 (O_585,N_28884,N_27461);
or UO_586 (O_586,N_28541,N_27795);
nand UO_587 (O_587,N_27406,N_29979);
nand UO_588 (O_588,N_28430,N_27929);
nor UO_589 (O_589,N_27689,N_27241);
xor UO_590 (O_590,N_28743,N_29593);
nand UO_591 (O_591,N_27422,N_28950);
or UO_592 (O_592,N_29981,N_29028);
nor UO_593 (O_593,N_28932,N_28044);
and UO_594 (O_594,N_27387,N_28027);
xor UO_595 (O_595,N_28971,N_28842);
xnor UO_596 (O_596,N_27378,N_28176);
nor UO_597 (O_597,N_29612,N_28768);
and UO_598 (O_598,N_28750,N_27413);
or UO_599 (O_599,N_29648,N_29034);
xnor UO_600 (O_600,N_28436,N_29768);
or UO_601 (O_601,N_29823,N_29556);
and UO_602 (O_602,N_28339,N_27380);
nand UO_603 (O_603,N_29733,N_29662);
nand UO_604 (O_604,N_28512,N_28224);
and UO_605 (O_605,N_28061,N_27796);
or UO_606 (O_606,N_28089,N_28726);
xor UO_607 (O_607,N_29866,N_27982);
nand UO_608 (O_608,N_29588,N_27097);
nor UO_609 (O_609,N_27125,N_27086);
xor UO_610 (O_610,N_29585,N_28298);
xnor UO_611 (O_611,N_29147,N_27564);
xnor UO_612 (O_612,N_27015,N_28009);
or UO_613 (O_613,N_28904,N_28396);
and UO_614 (O_614,N_28435,N_28408);
nand UO_615 (O_615,N_28097,N_27884);
and UO_616 (O_616,N_29143,N_29183);
and UO_617 (O_617,N_29992,N_28135);
and UO_618 (O_618,N_27093,N_29629);
nand UO_619 (O_619,N_28837,N_29844);
nand UO_620 (O_620,N_27459,N_28105);
xnor UO_621 (O_621,N_29809,N_27261);
and UO_622 (O_622,N_28188,N_27373);
nor UO_623 (O_623,N_28013,N_29232);
xor UO_624 (O_624,N_29617,N_27349);
and UO_625 (O_625,N_29598,N_29881);
nand UO_626 (O_626,N_29762,N_29671);
or UO_627 (O_627,N_27375,N_28498);
nor UO_628 (O_628,N_28174,N_29132);
and UO_629 (O_629,N_27867,N_28632);
nand UO_630 (O_630,N_29667,N_29925);
nor UO_631 (O_631,N_27751,N_27060);
xnor UO_632 (O_632,N_27503,N_27311);
nor UO_633 (O_633,N_27943,N_28124);
nor UO_634 (O_634,N_27416,N_28070);
xor UO_635 (O_635,N_29609,N_28634);
or UO_636 (O_636,N_27308,N_27037);
nor UO_637 (O_637,N_28242,N_28000);
xnor UO_638 (O_638,N_27958,N_29655);
nand UO_639 (O_639,N_29942,N_28590);
or UO_640 (O_640,N_27881,N_29117);
xnor UO_641 (O_641,N_29326,N_29657);
or UO_642 (O_642,N_27110,N_28168);
and UO_643 (O_643,N_27621,N_27146);
nand UO_644 (O_644,N_27872,N_27826);
xnor UO_645 (O_645,N_28650,N_29244);
nand UO_646 (O_646,N_27873,N_29167);
and UO_647 (O_647,N_28833,N_27780);
and UO_648 (O_648,N_29409,N_29074);
or UO_649 (O_649,N_28142,N_27155);
xor UO_650 (O_650,N_28208,N_27267);
or UO_651 (O_651,N_28050,N_28640);
nand UO_652 (O_652,N_27753,N_27529);
nand UO_653 (O_653,N_29623,N_29136);
nor UO_654 (O_654,N_29313,N_29876);
nand UO_655 (O_655,N_27892,N_27752);
and UO_656 (O_656,N_27307,N_28080);
or UO_657 (O_657,N_27650,N_27439);
nor UO_658 (O_658,N_29093,N_27049);
nand UO_659 (O_659,N_28203,N_29945);
nand UO_660 (O_660,N_28506,N_27698);
nor UO_661 (O_661,N_29339,N_28293);
or UO_662 (O_662,N_29208,N_27160);
and UO_663 (O_663,N_28420,N_27798);
or UO_664 (O_664,N_29770,N_28845);
xor UO_665 (O_665,N_28088,N_29847);
nor UO_666 (O_666,N_28226,N_29206);
xnor UO_667 (O_667,N_27999,N_28445);
or UO_668 (O_668,N_29164,N_28898);
nand UO_669 (O_669,N_27891,N_28972);
and UO_670 (O_670,N_28958,N_28342);
nor UO_671 (O_671,N_27808,N_28409);
and UO_672 (O_672,N_27801,N_28553);
nor UO_673 (O_673,N_28887,N_27244);
xnor UO_674 (O_674,N_27391,N_28077);
xnor UO_675 (O_675,N_28557,N_28662);
nand UO_676 (O_676,N_29210,N_27334);
and UO_677 (O_677,N_27167,N_28273);
nand UO_678 (O_678,N_29362,N_29471);
and UO_679 (O_679,N_28165,N_28782);
nand UO_680 (O_680,N_28390,N_29424);
nor UO_681 (O_681,N_27369,N_27327);
or UO_682 (O_682,N_27709,N_28951);
and UO_683 (O_683,N_27256,N_28542);
or UO_684 (O_684,N_27654,N_27496);
or UO_685 (O_685,N_29302,N_27909);
nand UO_686 (O_686,N_29477,N_27969);
xor UO_687 (O_687,N_28223,N_29394);
xor UO_688 (O_688,N_29390,N_27790);
xnor UO_689 (O_689,N_29275,N_29194);
or UO_690 (O_690,N_28902,N_27900);
or UO_691 (O_691,N_27000,N_29161);
or UO_692 (O_692,N_27149,N_28826);
nand UO_693 (O_693,N_29140,N_27825);
nor UO_694 (O_694,N_27836,N_28608);
xnor UO_695 (O_695,N_28889,N_28643);
and UO_696 (O_696,N_29972,N_28231);
nor UO_697 (O_697,N_28877,N_28254);
xnor UO_698 (O_698,N_27395,N_29797);
or UO_699 (O_699,N_28957,N_28051);
xnor UO_700 (O_700,N_27596,N_29975);
nor UO_701 (O_701,N_27389,N_27577);
or UO_702 (O_702,N_28073,N_29107);
and UO_703 (O_703,N_28429,N_27940);
nand UO_704 (O_704,N_27352,N_27972);
xnor UO_705 (O_705,N_27734,N_27533);
or UO_706 (O_706,N_28484,N_28555);
nand UO_707 (O_707,N_29361,N_27048);
nor UO_708 (O_708,N_28991,N_29273);
and UO_709 (O_709,N_27776,N_27398);
or UO_710 (O_710,N_29105,N_29872);
xor UO_711 (O_711,N_29470,N_29196);
and UO_712 (O_712,N_28611,N_27223);
nand UO_713 (O_713,N_29480,N_28539);
and UO_714 (O_714,N_28117,N_29964);
xor UO_715 (O_715,N_29427,N_28286);
nand UO_716 (O_716,N_27638,N_27133);
nand UO_717 (O_717,N_27499,N_29991);
nor UO_718 (O_718,N_27995,N_27739);
xor UO_719 (O_719,N_27597,N_27690);
and UO_720 (O_720,N_27207,N_27040);
nand UO_721 (O_721,N_28530,N_29885);
nand UO_722 (O_722,N_27727,N_29780);
or UO_723 (O_723,N_27174,N_29072);
nand UO_724 (O_724,N_28526,N_29329);
nand UO_725 (O_725,N_28922,N_27191);
nor UO_726 (O_726,N_29121,N_29020);
or UO_727 (O_727,N_28332,N_27797);
xnor UO_728 (O_728,N_29544,N_27977);
nor UO_729 (O_729,N_28659,N_29849);
nor UO_730 (O_730,N_28481,N_28637);
and UO_731 (O_731,N_28544,N_29895);
xnor UO_732 (O_732,N_29683,N_28167);
nand UO_733 (O_733,N_29656,N_28494);
nor UO_734 (O_734,N_28692,N_27293);
xnor UO_735 (O_735,N_27919,N_27616);
and UO_736 (O_736,N_28660,N_29375);
nand UO_737 (O_737,N_28773,N_29030);
nor UO_738 (O_738,N_28819,N_27508);
or UO_739 (O_739,N_28740,N_28258);
and UO_740 (O_740,N_28944,N_28055);
nand UO_741 (O_741,N_27756,N_27121);
nor UO_742 (O_742,N_28749,N_27356);
and UO_743 (O_743,N_28272,N_27528);
nand UO_744 (O_744,N_29763,N_27624);
and UO_745 (O_745,N_29564,N_27031);
nand UO_746 (O_746,N_27084,N_29605);
nor UO_747 (O_747,N_28818,N_28943);
xor UO_748 (O_748,N_29631,N_27585);
or UO_749 (O_749,N_29859,N_28683);
and UO_750 (O_750,N_27658,N_27778);
and UO_751 (O_751,N_27500,N_27284);
nand UO_752 (O_752,N_27001,N_27659);
nor UO_753 (O_753,N_27679,N_29069);
xnor UO_754 (O_754,N_27341,N_28198);
nand UO_755 (O_755,N_29239,N_29567);
and UO_756 (O_756,N_29698,N_29579);
nand UO_757 (O_757,N_29437,N_28522);
nand UO_758 (O_758,N_27083,N_29367);
or UO_759 (O_759,N_28719,N_28927);
nand UO_760 (O_760,N_28373,N_28372);
or UO_761 (O_761,N_29855,N_27818);
nand UO_762 (O_762,N_28201,N_29812);
xnor UO_763 (O_763,N_29358,N_29927);
and UO_764 (O_764,N_27230,N_29139);
nor UO_765 (O_765,N_29039,N_29727);
xnor UO_766 (O_766,N_27058,N_29788);
nand UO_767 (O_767,N_27681,N_29755);
and UO_768 (O_768,N_28228,N_28820);
or UO_769 (O_769,N_27984,N_27098);
or UO_770 (O_770,N_28792,N_27065);
xnor UO_771 (O_771,N_29611,N_27359);
nor UO_772 (O_772,N_27581,N_28312);
nand UO_773 (O_773,N_27243,N_29861);
or UO_774 (O_774,N_28138,N_28010);
nand UO_775 (O_775,N_28983,N_29738);
nor UO_776 (O_776,N_28410,N_28403);
nor UO_777 (O_777,N_28034,N_29412);
and UO_778 (O_778,N_29842,N_27802);
nand UO_779 (O_779,N_28492,N_28947);
or UO_780 (O_780,N_27885,N_28906);
nand UO_781 (O_781,N_29007,N_29675);
xnor UO_782 (O_782,N_27298,N_29509);
nand UO_783 (O_783,N_28197,N_29079);
and UO_784 (O_784,N_28033,N_29793);
or UO_785 (O_785,N_27204,N_27602);
nand UO_786 (O_786,N_28565,N_29254);
and UO_787 (O_787,N_28023,N_28655);
or UO_788 (O_788,N_27248,N_27329);
nor UO_789 (O_789,N_28259,N_28110);
nand UO_790 (O_790,N_27870,N_27860);
nand UO_791 (O_791,N_29938,N_27107);
nor UO_792 (O_792,N_27629,N_29963);
and UO_793 (O_793,N_29778,N_28900);
nor UO_794 (O_794,N_27164,N_28331);
and UO_795 (O_795,N_27491,N_27038);
xor UO_796 (O_796,N_27532,N_28236);
nand UO_797 (O_797,N_27105,N_27628);
nand UO_798 (O_798,N_29726,N_29309);
or UO_799 (O_799,N_27262,N_29745);
and UO_800 (O_800,N_28752,N_29889);
and UO_801 (O_801,N_27513,N_28677);
and UO_802 (O_802,N_28441,N_28850);
xor UO_803 (O_803,N_28281,N_28196);
and UO_804 (O_804,N_27145,N_29353);
or UO_805 (O_805,N_27209,N_27593);
or UO_806 (O_806,N_29789,N_27301);
and UO_807 (O_807,N_27912,N_28240);
nor UO_808 (O_808,N_28914,N_27561);
and UO_809 (O_809,N_27134,N_29530);
nand UO_810 (O_810,N_29786,N_29385);
xor UO_811 (O_811,N_29802,N_28337);
or UO_812 (O_812,N_29242,N_28008);
nand UO_813 (O_813,N_27289,N_27612);
nor UO_814 (O_814,N_27938,N_29630);
xor UO_815 (O_815,N_27292,N_28550);
nand UO_816 (O_816,N_28057,N_27512);
nor UO_817 (O_817,N_29267,N_27326);
nand UO_818 (O_818,N_27216,N_28593);
and UO_819 (O_819,N_29613,N_27740);
nand UO_820 (O_820,N_29357,N_27066);
or UO_821 (O_821,N_28453,N_29478);
nand UO_822 (O_822,N_27056,N_28374);
nand UO_823 (O_823,N_28369,N_29168);
nor UO_824 (O_824,N_27997,N_29960);
nor UO_825 (O_825,N_29124,N_28797);
xor UO_826 (O_826,N_27022,N_29472);
or UO_827 (O_827,N_29520,N_27625);
xnor UO_828 (O_828,N_27365,N_28729);
nand UO_829 (O_829,N_28036,N_28391);
xor UO_830 (O_830,N_28873,N_29949);
and UO_831 (O_831,N_27695,N_28938);
and UO_832 (O_832,N_29043,N_28614);
or UO_833 (O_833,N_27454,N_28039);
and UO_834 (O_834,N_27154,N_27059);
or UO_835 (O_835,N_27869,N_29392);
and UO_836 (O_836,N_29378,N_29642);
xor UO_837 (O_837,N_27360,N_29578);
and UO_838 (O_838,N_27966,N_28348);
or UO_839 (O_839,N_29382,N_28133);
nand UO_840 (O_840,N_28328,N_29965);
xor UO_841 (O_841,N_29643,N_28438);
or UO_842 (O_842,N_29153,N_29678);
and UO_843 (O_843,N_29265,N_27721);
nand UO_844 (O_844,N_27106,N_29970);
or UO_845 (O_845,N_29024,N_29109);
xnor UO_846 (O_846,N_28679,N_27590);
nor UO_847 (O_847,N_28132,N_28664);
xnor UO_848 (O_848,N_29352,N_27791);
xor UO_849 (O_849,N_28234,N_29059);
xnor UO_850 (O_850,N_29583,N_29523);
xor UO_851 (O_851,N_29009,N_28104);
nor UO_852 (O_852,N_29653,N_27542);
or UO_853 (O_853,N_27890,N_28081);
and UO_854 (O_854,N_29891,N_29483);
nand UO_855 (O_855,N_28882,N_29586);
or UO_856 (O_856,N_28973,N_29283);
and UO_857 (O_857,N_28472,N_28207);
nand UO_858 (O_858,N_27003,N_27376);
and UO_859 (O_859,N_29804,N_28586);
or UO_860 (O_860,N_27189,N_28152);
nor UO_861 (O_861,N_28414,N_27704);
nand UO_862 (O_862,N_29442,N_29223);
or UO_863 (O_863,N_27123,N_29679);
xor UO_864 (O_864,N_29888,N_27403);
nor UO_865 (O_865,N_29280,N_29426);
nor UO_866 (O_866,N_27492,N_28687);
xnor UO_867 (O_867,N_28754,N_28525);
and UO_868 (O_868,N_29563,N_28765);
and UO_869 (O_869,N_27678,N_27332);
and UO_870 (O_870,N_28128,N_29873);
nand UO_871 (O_871,N_29758,N_29094);
xnor UO_872 (O_872,N_27418,N_29073);
nor UO_873 (O_873,N_27605,N_27151);
or UO_874 (O_874,N_28581,N_27479);
nor UO_875 (O_875,N_27197,N_27484);
nand UO_876 (O_876,N_29301,N_27930);
and UO_877 (O_877,N_28903,N_29170);
or UO_878 (O_878,N_28589,N_28854);
nand UO_879 (O_879,N_29644,N_27132);
nor UO_880 (O_880,N_28496,N_27684);
or UO_881 (O_881,N_29397,N_29328);
xnor UO_882 (O_882,N_28418,N_27788);
xnor UO_883 (O_883,N_28048,N_28322);
xor UO_884 (O_884,N_29144,N_27897);
xnor UO_885 (O_885,N_27080,N_29572);
or UO_886 (O_886,N_28384,N_28710);
and UO_887 (O_887,N_27960,N_29005);
nor UO_888 (O_888,N_28119,N_27192);
xnor UO_889 (O_889,N_28828,N_28678);
nor UO_890 (O_890,N_29103,N_28723);
xnor UO_891 (O_891,N_29736,N_28284);
nand UO_892 (O_892,N_29940,N_27607);
and UO_893 (O_893,N_28856,N_27115);
nor UO_894 (O_894,N_27346,N_27840);
nand UO_895 (O_895,N_27758,N_28469);
nor UO_896 (O_896,N_27343,N_28362);
and UO_897 (O_897,N_29370,N_28092);
nor UO_898 (O_898,N_27633,N_29722);
and UO_899 (O_899,N_27269,N_29528);
or UO_900 (O_900,N_29822,N_28576);
nor UO_901 (O_901,N_29990,N_29819);
and UO_902 (O_902,N_28728,N_29620);
nand UO_903 (O_903,N_27092,N_29870);
nand UO_904 (O_904,N_29490,N_29049);
nor UO_905 (O_905,N_29850,N_27674);
nor UO_906 (O_906,N_29621,N_28849);
nand UO_907 (O_907,N_29078,N_29803);
or UO_908 (O_908,N_28451,N_28706);
or UO_909 (O_909,N_29337,N_29484);
and UO_910 (O_910,N_29815,N_28344);
nor UO_911 (O_911,N_28367,N_27111);
and UO_912 (O_912,N_28531,N_28538);
nor UO_913 (O_913,N_28371,N_27644);
nor UO_914 (O_914,N_28101,N_29614);
nand UO_915 (O_915,N_27074,N_28163);
xor UO_916 (O_916,N_29310,N_29557);
or UO_917 (O_917,N_28004,N_27666);
and UO_918 (O_918,N_27569,N_27501);
or UO_919 (O_919,N_28353,N_28134);
nor UO_920 (O_920,N_27242,N_29141);
nand UO_921 (O_921,N_29489,N_28747);
nor UO_922 (O_922,N_27599,N_29551);
xor UO_923 (O_923,N_28911,N_29511);
nor UO_924 (O_924,N_29048,N_27475);
nor UO_925 (O_925,N_27257,N_27979);
or UO_926 (O_926,N_27228,N_27489);
xnor UO_927 (O_927,N_27911,N_28460);
nor UO_928 (O_928,N_28204,N_27522);
nand UO_929 (O_929,N_27567,N_28809);
nor UO_930 (O_930,N_28064,N_28255);
nor UO_931 (O_931,N_27009,N_27687);
nor UO_932 (O_932,N_29967,N_28225);
or UO_933 (O_933,N_28734,N_28432);
and UO_934 (O_934,N_28961,N_29843);
xnor UO_935 (O_935,N_29467,N_29848);
and UO_936 (O_936,N_28604,N_28084);
and UO_937 (O_937,N_27970,N_27371);
and UO_938 (O_938,N_27635,N_27728);
nor UO_939 (O_939,N_27588,N_27670);
nor UO_940 (O_940,N_29790,N_27286);
and UO_941 (O_941,N_28722,N_28148);
and UO_942 (O_942,N_27494,N_28763);
nand UO_943 (O_943,N_29120,N_27440);
nor UO_944 (O_944,N_29271,N_28193);
nor UO_945 (O_945,N_29134,N_28150);
or UO_946 (O_946,N_27913,N_29184);
nand UO_947 (O_947,N_29425,N_29050);
or UO_948 (O_948,N_27178,N_28886);
xnor UO_949 (O_949,N_28159,N_28851);
nor UO_950 (O_950,N_27433,N_29709);
nand UO_951 (O_951,N_29464,N_28083);
nand UO_952 (O_952,N_27432,N_29756);
nand UO_953 (O_953,N_28865,N_27547);
xor UO_954 (O_954,N_27750,N_27645);
and UO_955 (O_955,N_28880,N_29592);
or UO_956 (O_956,N_27441,N_29346);
and UO_957 (O_957,N_27617,N_29209);
nor UO_958 (O_958,N_27464,N_27368);
and UO_959 (O_959,N_27417,N_28600);
xnor UO_960 (O_960,N_29458,N_28901);
xnor UO_961 (O_961,N_27481,N_28529);
nor UO_962 (O_962,N_27285,N_28011);
and UO_963 (O_963,N_27931,N_28724);
nand UO_964 (O_964,N_28448,N_29783);
or UO_965 (O_965,N_29261,N_29807);
and UO_966 (O_966,N_28596,N_28697);
and UO_967 (O_967,N_27655,N_28579);
xor UO_968 (O_968,N_28171,N_28497);
and UO_969 (O_969,N_29731,N_29834);
nand UO_970 (O_970,N_29966,N_28816);
or UO_971 (O_971,N_29415,N_28574);
nand UO_972 (O_972,N_28715,N_28195);
xnor UO_973 (O_973,N_27715,N_29055);
nand UO_974 (O_974,N_29950,N_28970);
nand UO_975 (O_975,N_27278,N_27495);
or UO_976 (O_976,N_27524,N_28916);
or UO_977 (O_977,N_27962,N_28392);
and UO_978 (O_978,N_29513,N_28794);
or UO_979 (O_979,N_29782,N_28210);
nand UO_980 (O_980,N_29715,N_28712);
nor UO_981 (O_981,N_28269,N_29827);
and UO_982 (O_982,N_29263,N_27229);
nand UO_983 (O_983,N_28534,N_29452);
nand UO_984 (O_984,N_28123,N_29222);
nand UO_985 (O_985,N_28311,N_28323);
and UO_986 (O_986,N_29674,N_28561);
and UO_987 (O_987,N_27194,N_28516);
xor UO_988 (O_988,N_28870,N_28940);
xnor UO_989 (O_989,N_28212,N_28120);
xor UO_990 (O_990,N_27407,N_29735);
nand UO_991 (O_991,N_27321,N_28979);
nor UO_992 (O_992,N_28184,N_28192);
or UO_993 (O_993,N_27270,N_29463);
nand UO_994 (O_994,N_29096,N_27100);
nand UO_995 (O_995,N_27987,N_28221);
and UO_996 (O_996,N_29014,N_29526);
xnor UO_997 (O_997,N_29721,N_27276);
nand UO_998 (O_998,N_29510,N_27609);
and UO_999 (O_999,N_29636,N_27888);
or UO_1000 (O_1000,N_27774,N_28185);
and UO_1001 (O_1001,N_28626,N_29369);
nand UO_1002 (O_1002,N_29759,N_28257);
nor UO_1003 (O_1003,N_29637,N_29053);
nand UO_1004 (O_1004,N_27088,N_28977);
nand UO_1005 (O_1005,N_27766,N_29054);
nand UO_1006 (O_1006,N_29989,N_27712);
xor UO_1007 (O_1007,N_27544,N_29221);
nor UO_1008 (O_1008,N_27218,N_27779);
and UO_1009 (O_1009,N_27527,N_27029);
nor UO_1010 (O_1010,N_28500,N_29641);
or UO_1011 (O_1011,N_29580,N_29032);
xor UO_1012 (O_1012,N_29724,N_29276);
or UO_1013 (O_1013,N_29278,N_29441);
nand UO_1014 (O_1014,N_29508,N_28491);
xnor UO_1015 (O_1015,N_27702,N_27880);
and UO_1016 (O_1016,N_27935,N_28317);
or UO_1017 (O_1017,N_29002,N_29835);
nor UO_1018 (O_1018,N_29542,N_29610);
nor UO_1019 (O_1019,N_28519,N_29175);
or UO_1020 (O_1020,N_28493,N_27364);
and UO_1021 (O_1021,N_28919,N_27521);
and UO_1022 (O_1022,N_27847,N_29298);
nand UO_1023 (O_1023,N_29207,N_29858);
or UO_1024 (O_1024,N_27724,N_27129);
xor UO_1025 (O_1025,N_29661,N_28285);
xor UO_1026 (O_1026,N_27469,N_28566);
or UO_1027 (O_1027,N_27217,N_28156);
or UO_1028 (O_1028,N_27172,N_29817);
nor UO_1029 (O_1029,N_28021,N_27587);
and UO_1030 (O_1030,N_27166,N_27717);
or UO_1031 (O_1031,N_27428,N_29688);
nor UO_1032 (O_1032,N_28737,N_28987);
and UO_1033 (O_1033,N_28154,N_28871);
and UO_1034 (O_1034,N_29248,N_28814);
or UO_1035 (O_1035,N_27238,N_29983);
and UO_1036 (O_1036,N_29255,N_27063);
xor UO_1037 (O_1037,N_27783,N_29474);
or UO_1038 (O_1038,N_29887,N_27399);
nor UO_1039 (O_1039,N_29604,N_28475);
nand UO_1040 (O_1040,N_28812,N_28319);
xor UO_1041 (O_1041,N_28464,N_27487);
or UO_1042 (O_1042,N_27859,N_29029);
and UO_1043 (O_1043,N_28377,N_29749);
or UO_1044 (O_1044,N_28220,N_28398);
or UO_1045 (O_1045,N_29750,N_28109);
and UO_1046 (O_1046,N_27789,N_29864);
or UO_1047 (O_1047,N_28379,N_29555);
nor UO_1048 (O_1048,N_28304,N_29396);
and UO_1049 (O_1049,N_28617,N_28265);
or UO_1050 (O_1050,N_27954,N_29260);
or UO_1051 (O_1051,N_28277,N_28458);
or UO_1052 (O_1052,N_28235,N_28336);
nand UO_1053 (O_1053,N_29466,N_27460);
xnor UO_1054 (O_1054,N_27594,N_28301);
and UO_1055 (O_1055,N_28647,N_28610);
xor UO_1056 (O_1056,N_27096,N_27227);
nand UO_1057 (O_1057,N_29533,N_27959);
and UO_1058 (O_1058,N_29058,N_27091);
or UO_1059 (O_1059,N_28546,N_28562);
or UO_1060 (O_1060,N_29359,N_29486);
and UO_1061 (O_1061,N_28108,N_29038);
xnor UO_1062 (O_1062,N_28612,N_29552);
nand UO_1063 (O_1063,N_29284,N_27552);
or UO_1064 (O_1064,N_29413,N_27412);
or UO_1065 (O_1065,N_27490,N_27032);
xnor UO_1066 (O_1066,N_28641,N_28425);
or UO_1067 (O_1067,N_28354,N_27634);
xnor UO_1068 (O_1068,N_29224,N_27198);
nand UO_1069 (O_1069,N_28383,N_27347);
nor UO_1070 (O_1070,N_29801,N_27765);
nor UO_1071 (O_1071,N_28862,N_27141);
xnor UO_1072 (O_1072,N_27827,N_28059);
or UO_1073 (O_1073,N_27812,N_28276);
nand UO_1074 (O_1074,N_29607,N_29754);
nand UO_1075 (O_1075,N_27708,N_27763);
nor UO_1076 (O_1076,N_28029,N_28793);
nor UO_1077 (O_1077,N_28233,N_27385);
nor UO_1078 (O_1078,N_27811,N_27934);
nand UO_1079 (O_1079,N_27053,N_29625);
and UO_1080 (O_1080,N_28360,N_27794);
nor UO_1081 (O_1081,N_27928,N_27755);
nand UO_1082 (O_1082,N_28157,N_28345);
xor UO_1083 (O_1083,N_27993,N_28320);
xnor UO_1084 (O_1084,N_27714,N_27853);
xnor UO_1085 (O_1085,N_28288,N_29924);
nand UO_1086 (O_1086,N_27258,N_29958);
xor UO_1087 (O_1087,N_28382,N_29022);
and UO_1088 (O_1088,N_27342,N_28351);
xor UO_1089 (O_1089,N_29091,N_28644);
nand UO_1090 (O_1090,N_27222,N_28879);
nor UO_1091 (O_1091,N_29406,N_29496);
and UO_1092 (O_1092,N_28229,N_29434);
or UO_1093 (O_1093,N_29909,N_28356);
nor UO_1094 (O_1094,N_27175,N_27646);
xor UO_1095 (O_1095,N_28989,N_28058);
or UO_1096 (O_1096,N_27070,N_28672);
or UO_1097 (O_1097,N_28514,N_27026);
nand UO_1098 (O_1098,N_29253,N_27665);
nor UO_1099 (O_1099,N_27335,N_28093);
nor UO_1100 (O_1100,N_28018,N_28237);
and UO_1101 (O_1101,N_27855,N_29051);
and UO_1102 (O_1102,N_29287,N_27536);
and UO_1103 (O_1103,N_28177,N_27304);
nor UO_1104 (O_1104,N_29971,N_28780);
nand UO_1105 (O_1105,N_28727,N_28585);
xnor UO_1106 (O_1106,N_28454,N_29270);
or UO_1107 (O_1107,N_29013,N_27139);
or UO_1108 (O_1108,N_28268,N_29565);
or UO_1109 (O_1109,N_27933,N_28263);
or UO_1110 (O_1110,N_27807,N_27344);
nor UO_1111 (O_1111,N_27677,N_29082);
or UO_1112 (O_1112,N_28925,N_27922);
and UO_1113 (O_1113,N_28731,N_27383);
nand UO_1114 (O_1114,N_28666,N_27699);
xor UO_1115 (O_1115,N_27697,N_29438);
and UO_1116 (O_1116,N_29634,N_27136);
and UO_1117 (O_1117,N_29660,N_27523);
and UO_1118 (O_1118,N_29211,N_29354);
nor UO_1119 (O_1119,N_29128,N_28490);
and UO_1120 (O_1120,N_28002,N_28428);
xor UO_1121 (O_1121,N_29720,N_29416);
or UO_1122 (O_1122,N_27300,N_28066);
nor UO_1123 (O_1123,N_27641,N_27291);
nand UO_1124 (O_1124,N_27316,N_28631);
nand UO_1125 (O_1125,N_29576,N_29988);
and UO_1126 (O_1126,N_28129,N_28136);
xnor UO_1127 (O_1127,N_27961,N_29213);
nand UO_1128 (O_1128,N_28930,N_27573);
nand UO_1129 (O_1129,N_27906,N_29300);
and UO_1130 (O_1130,N_28022,N_27761);
and UO_1131 (O_1131,N_27202,N_27509);
nand UO_1132 (O_1132,N_28495,N_28296);
nand UO_1133 (O_1133,N_28366,N_28651);
or UO_1134 (O_1134,N_29097,N_29982);
and UO_1135 (O_1135,N_28625,N_29204);
xnor UO_1136 (O_1136,N_29129,N_27680);
and UO_1137 (O_1137,N_29087,N_28629);
xor UO_1138 (O_1138,N_29070,N_28988);
xnor UO_1139 (O_1139,N_29931,N_29893);
nor UO_1140 (O_1140,N_29638,N_29348);
or UO_1141 (O_1141,N_28325,N_28510);
nor UO_1142 (O_1142,N_27902,N_28966);
and UO_1143 (O_1143,N_29233,N_29974);
and UO_1144 (O_1144,N_29791,N_29241);
or UO_1145 (O_1145,N_29492,N_28505);
nand UO_1146 (O_1146,N_27402,N_29545);
nor UO_1147 (O_1147,N_29085,N_29799);
or UO_1148 (O_1148,N_28046,N_28091);
and UO_1149 (O_1149,N_28407,N_28654);
nand UO_1150 (O_1150,N_28992,N_28796);
or UO_1151 (O_1151,N_27538,N_28962);
or UO_1152 (O_1152,N_27864,N_28671);
xor UO_1153 (O_1153,N_29517,N_29821);
and UO_1154 (O_1154,N_27427,N_29042);
nand UO_1155 (O_1155,N_27370,N_27643);
nand UO_1156 (O_1156,N_28305,N_29008);
nand UO_1157 (O_1157,N_27921,N_29740);
or UO_1158 (O_1158,N_27131,N_29296);
or UO_1159 (O_1159,N_28543,N_29673);
nand UO_1160 (O_1160,N_29214,N_28245);
nor UO_1161 (O_1161,N_27377,N_29669);
nor UO_1162 (O_1162,N_27735,N_27397);
xor UO_1163 (O_1163,N_28300,N_27639);
nor UO_1164 (O_1164,N_29493,N_27266);
and UO_1165 (O_1165,N_28274,N_27012);
and UO_1166 (O_1166,N_27203,N_29521);
or UO_1167 (O_1167,N_29953,N_27294);
xnor UO_1168 (O_1168,N_28049,N_27400);
nor UO_1169 (O_1169,N_29218,N_29664);
xor UO_1170 (O_1170,N_29549,N_29418);
nand UO_1171 (O_1171,N_27176,N_28450);
xnor UO_1172 (O_1172,N_29784,N_27306);
and UO_1173 (O_1173,N_27743,N_29411);
or UO_1174 (O_1174,N_27784,N_28597);
xor UO_1175 (O_1175,N_27517,N_29077);
xnor UO_1176 (O_1176,N_29180,N_28563);
or UO_1177 (O_1177,N_27338,N_29959);
nor UO_1178 (O_1178,N_29703,N_28711);
and UO_1179 (O_1179,N_29060,N_29236);
nor UO_1180 (O_1180,N_27451,N_29482);
xor UO_1181 (O_1181,N_27757,N_29457);
xor UO_1182 (O_1182,N_27737,N_28404);
nor UO_1183 (O_1183,N_27388,N_28335);
and UO_1184 (O_1184,N_27087,N_29935);
nor UO_1185 (O_1185,N_29569,N_29603);
nor UO_1186 (O_1186,N_29045,N_29202);
nand UO_1187 (O_1187,N_29379,N_29012);
xor UO_1188 (O_1188,N_28349,N_28564);
nor UO_1189 (O_1189,N_27953,N_28843);
xor UO_1190 (O_1190,N_29479,N_29461);
xnor UO_1191 (O_1191,N_29181,N_28122);
nor UO_1192 (O_1192,N_29839,N_28764);
xor UO_1193 (O_1193,N_29930,N_27069);
nand UO_1194 (O_1194,N_28062,N_27235);
nand UO_1195 (O_1195,N_29701,N_28716);
nor UO_1196 (O_1196,N_28357,N_29882);
nand UO_1197 (O_1197,N_27361,N_29331);
xnor UO_1198 (O_1198,N_29307,N_29677);
nor UO_1199 (O_1199,N_29162,N_29792);
nor UO_1200 (O_1200,N_29690,N_29125);
or UO_1201 (O_1201,N_27682,N_28031);
nand UO_1202 (O_1202,N_27004,N_29404);
nor UO_1203 (O_1203,N_28111,N_27595);
nor UO_1204 (O_1204,N_28456,N_28139);
xnor UO_1205 (O_1205,N_28774,N_28053);
xnor UO_1206 (O_1206,N_29226,N_28985);
xor UO_1207 (O_1207,N_29274,N_27457);
nand UO_1208 (O_1208,N_28830,N_27199);
and UO_1209 (O_1209,N_28881,N_28102);
or UO_1210 (O_1210,N_27315,N_28759);
nor UO_1211 (O_1211,N_27142,N_29198);
nor UO_1212 (O_1212,N_29769,N_27372);
and UO_1213 (O_1213,N_29516,N_28545);
nand UO_1214 (O_1214,N_27648,N_27127);
nand UO_1215 (O_1215,N_27330,N_29432);
and UO_1216 (O_1216,N_28266,N_29883);
and UO_1217 (O_1217,N_27950,N_27449);
and UO_1218 (O_1218,N_27915,N_28924);
nor UO_1219 (O_1219,N_27526,N_27386);
or UO_1220 (O_1220,N_28928,N_27477);
nor UO_1221 (O_1221,N_27839,N_27738);
or UO_1222 (O_1222,N_29796,N_28601);
nor UO_1223 (O_1223,N_28130,N_27545);
nor UO_1224 (O_1224,N_28455,N_27777);
or UO_1225 (O_1225,N_27247,N_27895);
xnor UO_1226 (O_1226,N_29670,N_27353);
nor UO_1227 (O_1227,N_27565,N_28852);
or UO_1228 (O_1228,N_29075,N_27894);
or UO_1229 (O_1229,N_27045,N_27221);
nor UO_1230 (O_1230,N_27606,N_27165);
nand UO_1231 (O_1231,N_28939,N_29568);
and UO_1232 (O_1232,N_28910,N_27516);
xor UO_1233 (O_1233,N_28028,N_28292);
nor UO_1234 (O_1234,N_27838,N_27560);
or UO_1235 (O_1235,N_29986,N_28892);
xnor UO_1236 (O_1236,N_27649,N_29165);
and UO_1237 (O_1237,N_29497,N_27799);
and UO_1238 (O_1238,N_28948,N_28457);
nand UO_1239 (O_1239,N_28738,N_27288);
xor UO_1240 (O_1240,N_29152,N_28682);
xnor UO_1241 (O_1241,N_28694,N_29364);
nor UO_1242 (O_1242,N_27729,N_28141);
nor UO_1243 (O_1243,N_28807,N_29892);
nand UO_1244 (O_1244,N_29092,N_29907);
and UO_1245 (O_1245,N_28998,N_28016);
xor UO_1246 (O_1246,N_28599,N_29431);
and UO_1247 (O_1247,N_27225,N_29350);
nor UO_1248 (O_1248,N_29926,N_28623);
nor UO_1249 (O_1249,N_28705,N_28964);
and UO_1250 (O_1250,N_28395,N_28517);
nand UO_1251 (O_1251,N_27515,N_27320);
or UO_1252 (O_1252,N_28444,N_29524);
nor UO_1253 (O_1253,N_28341,N_27404);
and UO_1254 (O_1254,N_29941,N_27626);
nor UO_1255 (O_1255,N_27034,N_29980);
or UO_1256 (O_1256,N_27153,N_29616);
xnor UO_1257 (O_1257,N_27161,N_27239);
and UO_1258 (O_1258,N_27557,N_27850);
xnor UO_1259 (O_1259,N_29111,N_28656);
nor UO_1260 (O_1260,N_29854,N_27089);
and UO_1261 (O_1261,N_28355,N_27782);
or UO_1262 (O_1262,N_27354,N_29840);
nand UO_1263 (O_1263,N_29306,N_28098);
nor UO_1264 (O_1264,N_28802,N_28795);
nand UO_1265 (O_1265,N_27656,N_29439);
nand UO_1266 (O_1266,N_28791,N_29146);
xor UO_1267 (O_1267,N_27212,N_28603);
xor UO_1268 (O_1268,N_29830,N_27231);
nor UO_1269 (O_1269,N_29227,N_29295);
nand UO_1270 (O_1270,N_27762,N_29904);
nor UO_1271 (O_1271,N_28217,N_27362);
nand UO_1272 (O_1272,N_28153,N_28936);
or UO_1273 (O_1273,N_29455,N_29751);
nand UO_1274 (O_1274,N_27589,N_27932);
and UO_1275 (O_1275,N_27183,N_28559);
nand UO_1276 (O_1276,N_29806,N_28863);
or UO_1277 (O_1277,N_28636,N_29933);
nand UO_1278 (O_1278,N_28568,N_27772);
nand UO_1279 (O_1279,N_28180,N_27673);
and UO_1280 (O_1280,N_27409,N_29197);
nand UO_1281 (O_1281,N_29706,N_27809);
nor UO_1282 (O_1282,N_27874,N_27985);
nor UO_1283 (O_1283,N_28949,N_28621);
nor UO_1284 (O_1284,N_27474,N_28486);
or UO_1285 (O_1285,N_29325,N_27188);
and UO_1286 (O_1286,N_29890,N_29900);
and UO_1287 (O_1287,N_28017,N_28777);
nor UO_1288 (O_1288,N_27664,N_28213);
xor UO_1289 (O_1289,N_29846,N_29279);
xor UO_1290 (O_1290,N_28147,N_27485);
and UO_1291 (O_1291,N_27871,N_29739);
nand UO_1292 (O_1292,N_27472,N_28835);
xor UO_1293 (O_1293,N_28144,N_27483);
xor UO_1294 (O_1294,N_29760,N_28839);
nor UO_1295 (O_1295,N_29108,N_29646);
and UO_1296 (O_1296,N_27337,N_27923);
nor UO_1297 (O_1297,N_29697,N_27694);
and UO_1298 (O_1298,N_27050,N_28015);
and UO_1299 (O_1299,N_28836,N_27907);
or UO_1300 (O_1300,N_29665,N_29294);
and UO_1301 (O_1301,N_29689,N_27138);
xnor UO_1302 (O_1302,N_29879,N_29877);
xnor UO_1303 (O_1303,N_28591,N_28427);
or UO_1304 (O_1304,N_27319,N_27945);
nand UO_1305 (O_1305,N_27941,N_27663);
nand UO_1306 (O_1306,N_28206,N_29272);
or UO_1307 (O_1307,N_28309,N_29851);
nand UO_1308 (O_1308,N_27759,N_28316);
and UO_1309 (O_1309,N_27831,N_27210);
and UO_1310 (O_1310,N_29650,N_28358);
nor UO_1311 (O_1311,N_27760,N_29838);
nor UO_1312 (O_1312,N_27020,N_28035);
nand UO_1313 (O_1313,N_29460,N_28858);
nand UO_1314 (O_1314,N_29908,N_27415);
and UO_1315 (O_1315,N_27511,N_29663);
xnor UO_1316 (O_1316,N_28953,N_29968);
nor UO_1317 (O_1317,N_27942,N_28917);
nand UO_1318 (O_1318,N_28499,N_28959);
or UO_1319 (O_1319,N_29444,N_29256);
nor UO_1320 (O_1320,N_29537,N_29946);
and UO_1321 (O_1321,N_27671,N_28253);
nand UO_1322 (O_1322,N_28890,N_28075);
or UO_1323 (O_1323,N_27719,N_27662);
or UO_1324 (O_1324,N_28680,N_28556);
nand UO_1325 (O_1325,N_27035,N_27861);
xnor UO_1326 (O_1326,N_29814,N_29289);
xnor UO_1327 (O_1327,N_28399,N_29622);
nor UO_1328 (O_1328,N_29937,N_29040);
nand UO_1329 (O_1329,N_28587,N_27023);
nand UO_1330 (O_1330,N_28788,N_28607);
nand UO_1331 (O_1331,N_27055,N_29573);
and UO_1332 (O_1332,N_27725,N_27768);
xor UO_1333 (O_1333,N_27309,N_27660);
and UO_1334 (O_1334,N_28748,N_28825);
nand UO_1335 (O_1335,N_28211,N_29343);
and UO_1336 (O_1336,N_29193,N_27980);
nor UO_1337 (O_1337,N_29469,N_29597);
and UO_1338 (O_1338,N_29633,N_29820);
nand UO_1339 (O_1339,N_28042,N_29532);
or UO_1340 (O_1340,N_27846,N_27956);
xor UO_1341 (O_1341,N_27205,N_29943);
xnor UO_1342 (O_1342,N_27317,N_28270);
xor UO_1343 (O_1343,N_28674,N_29033);
or UO_1344 (O_1344,N_29114,N_27973);
or UO_1345 (O_1345,N_28700,N_27497);
and UO_1346 (O_1346,N_28878,N_27259);
nand UO_1347 (O_1347,N_29259,N_29651);
and UO_1348 (O_1348,N_27047,N_29681);
xnor UO_1349 (O_1349,N_28896,N_28627);
and UO_1350 (O_1350,N_28227,N_27005);
xnor UO_1351 (O_1351,N_27169,N_28861);
or UO_1352 (O_1352,N_27314,N_29955);
xor UO_1353 (O_1353,N_27829,N_28527);
nor UO_1354 (O_1354,N_29344,N_28501);
or UO_1355 (O_1355,N_27736,N_28182);
nor UO_1356 (O_1356,N_27787,N_28808);
and UO_1357 (O_1357,N_29566,N_28628);
nor UO_1358 (O_1358,N_28026,N_27920);
and UO_1359 (O_1359,N_29145,N_28690);
nand UO_1360 (O_1360,N_27390,N_27889);
xnor UO_1361 (O_1361,N_29448,N_29906);
nand UO_1362 (O_1362,N_27837,N_29794);
and UO_1363 (O_1363,N_28758,N_27246);
xnor UO_1364 (O_1364,N_27823,N_28986);
or UO_1365 (O_1365,N_28770,N_28535);
xnor UO_1366 (O_1366,N_29962,N_27820);
xnor UO_1367 (O_1367,N_28330,N_27786);
nand UO_1368 (O_1368,N_29056,N_29652);
nor UO_1369 (O_1369,N_27937,N_29810);
xor UO_1370 (O_1370,N_27718,N_27024);
nor UO_1371 (O_1371,N_27575,N_29026);
or UO_1372 (O_1372,N_27571,N_28465);
xor UO_1373 (O_1373,N_27008,N_29818);
nand UO_1374 (O_1374,N_28638,N_29743);
or UO_1375 (O_1375,N_27967,N_27744);
nor UO_1376 (O_1376,N_29591,N_29693);
or UO_1377 (O_1377,N_29405,N_27424);
and UO_1378 (O_1378,N_29371,N_27976);
or UO_1379 (O_1379,N_29286,N_28194);
nand UO_1380 (O_1380,N_29384,N_29391);
xor UO_1381 (O_1381,N_27562,N_28741);
nand UO_1382 (O_1382,N_27245,N_28503);
nor UO_1383 (O_1383,N_28394,N_27382);
and UO_1384 (O_1384,N_28385,N_28560);
and UO_1385 (O_1385,N_29476,N_28997);
nand UO_1386 (O_1386,N_27467,N_29922);
and UO_1387 (O_1387,N_28735,N_29712);
xor UO_1388 (O_1388,N_27990,N_29813);
nor UO_1389 (O_1389,N_28642,N_29805);
nor UO_1390 (O_1390,N_27186,N_27277);
or UO_1391 (O_1391,N_28338,N_28461);
nor UO_1392 (O_1392,N_28897,N_29954);
and UO_1393 (O_1393,N_29095,N_28509);
and UO_1394 (O_1394,N_28190,N_27653);
nor UO_1395 (O_1395,N_27857,N_28624);
and UO_1396 (O_1396,N_27615,N_29293);
nand UO_1397 (O_1397,N_27253,N_27430);
xor UO_1398 (O_1398,N_29833,N_27109);
xor UO_1399 (O_1399,N_29601,N_28746);
nor UO_1400 (O_1400,N_29785,N_27896);
or UO_1401 (O_1401,N_29305,N_27905);
xor UO_1402 (O_1402,N_28681,N_29923);
nand UO_1403 (O_1403,N_27936,N_28725);
xor UO_1404 (O_1404,N_29436,N_28592);
or UO_1405 (O_1405,N_29453,N_29435);
and UO_1406 (O_1406,N_27017,N_28442);
and UO_1407 (O_1407,N_29264,N_28648);
or UO_1408 (O_1408,N_29640,N_28844);
and UO_1409 (O_1409,N_28978,N_29886);
xnor UO_1410 (O_1410,N_28030,N_29018);
and UO_1411 (O_1411,N_28340,N_28518);
nand UO_1412 (O_1412,N_28968,N_29355);
nor UO_1413 (O_1413,N_28466,N_27652);
and UO_1414 (O_1414,N_29798,N_28718);
or UO_1415 (O_1415,N_28920,N_27971);
xnor UO_1416 (O_1416,N_29158,N_28069);
nor UO_1417 (O_1417,N_27312,N_28306);
nand UO_1418 (O_1418,N_28806,N_28043);
nor UO_1419 (O_1419,N_29064,N_28437);
nor UO_1420 (O_1420,N_28485,N_27992);
nand UO_1421 (O_1421,N_27710,N_29245);
nand UO_1422 (O_1422,N_28829,N_29994);
xnor UO_1423 (O_1423,N_27042,N_29003);
nor UO_1424 (O_1424,N_29365,N_29113);
and UO_1425 (O_1425,N_29414,N_27955);
nand UO_1426 (O_1426,N_29373,N_28931);
nand UO_1427 (O_1427,N_29473,N_29433);
or UO_1428 (O_1428,N_28799,N_28630);
nor UO_1429 (O_1429,N_27707,N_27119);
xnor UO_1430 (O_1430,N_29428,N_28483);
or UO_1431 (O_1431,N_28346,N_28866);
or UO_1432 (O_1432,N_28482,N_28885);
nand UO_1433 (O_1433,N_28883,N_29753);
or UO_1434 (O_1434,N_27822,N_29668);
or UO_1435 (O_1435,N_29004,N_28891);
and UO_1436 (O_1436,N_28169,N_28476);
nand UO_1437 (O_1437,N_27177,N_29811);
or UO_1438 (O_1438,N_28874,N_29921);
or UO_1439 (O_1439,N_28143,N_27843);
nor UO_1440 (O_1440,N_29826,N_28713);
or UO_1441 (O_1441,N_28145,N_28326);
nand UO_1442 (O_1442,N_27265,N_29571);
nand UO_1443 (O_1443,N_28707,N_29553);
and UO_1444 (O_1444,N_28663,N_28918);
or UO_1445 (O_1445,N_29443,N_27770);
xnor UO_1446 (O_1446,N_28467,N_28474);
nor UO_1447 (O_1447,N_28993,N_28584);
and UO_1448 (O_1448,N_29174,N_28443);
or UO_1449 (O_1449,N_28178,N_27917);
nand UO_1450 (O_1450,N_29216,N_27168);
and UO_1451 (O_1451,N_29627,N_27800);
nor UO_1452 (O_1452,N_27374,N_29918);
xnor UO_1453 (O_1453,N_28001,N_27196);
or UO_1454 (O_1454,N_28282,N_27583);
nand UO_1455 (O_1455,N_27914,N_29871);
or UO_1456 (O_1456,N_27592,N_28045);
xnor UO_1457 (O_1457,N_27173,N_29188);
or UO_1458 (O_1458,N_27028,N_28524);
nand UO_1459 (O_1459,N_27636,N_28116);
nor UO_1460 (O_1460,N_27611,N_27548);
nand UO_1461 (O_1461,N_28387,N_28246);
or UO_1462 (O_1462,N_29547,N_29626);
or UO_1463 (O_1463,N_29765,N_27201);
xor UO_1464 (O_1464,N_28703,N_27339);
and UO_1465 (O_1465,N_29228,N_27144);
nand UO_1466 (O_1466,N_27039,N_28720);
and UO_1467 (O_1467,N_27150,N_28115);
nor UO_1468 (O_1468,N_28577,N_27691);
nand UO_1469 (O_1469,N_28380,N_29781);
or UO_1470 (O_1470,N_27019,N_27862);
nand UO_1471 (O_1471,N_28307,N_28757);
nand UO_1472 (O_1472,N_28864,N_29748);
and UO_1473 (O_1473,N_28411,N_29570);
xnor UO_1474 (O_1474,N_28696,N_27813);
nor UO_1475 (O_1475,N_29249,N_29998);
or UO_1476 (O_1476,N_27328,N_27957);
nand UO_1477 (O_1477,N_27419,N_29589);
nor UO_1478 (O_1478,N_27771,N_29172);
xor UO_1479 (O_1479,N_29666,N_29654);
nand UO_1480 (O_1480,N_27582,N_29252);
and UO_1481 (O_1481,N_27741,N_28477);
xor UO_1482 (O_1482,N_29711,N_29512);
xnor UO_1483 (O_1483,N_29947,N_28570);
or UO_1484 (O_1484,N_27667,N_28082);
xnor UO_1485 (O_1485,N_28981,N_29215);
xor UO_1486 (O_1486,N_27185,N_29006);
nand UO_1487 (O_1487,N_28605,N_29155);
xnor UO_1488 (O_1488,N_27764,N_28218);
xnor UO_1489 (O_1489,N_29914,N_27114);
and UO_1490 (O_1490,N_28755,N_27085);
nor UO_1491 (O_1491,N_29142,N_28708);
and UO_1492 (O_1492,N_29237,N_27696);
nand UO_1493 (O_1493,N_28090,N_27112);
nor UO_1494 (O_1494,N_27745,N_29856);
nor UO_1495 (O_1495,N_27946,N_29860);
xor UO_1496 (O_1496,N_28230,N_27806);
nand UO_1497 (O_1497,N_29421,N_29291);
and UO_1498 (O_1498,N_27556,N_28086);
xnor UO_1499 (O_1499,N_29957,N_29351);
or UO_1500 (O_1500,N_27010,N_27410);
or UO_1501 (O_1501,N_29125,N_29726);
xnor UO_1502 (O_1502,N_29679,N_28866);
nand UO_1503 (O_1503,N_29033,N_29886);
and UO_1504 (O_1504,N_27206,N_27824);
nor UO_1505 (O_1505,N_29016,N_27782);
or UO_1506 (O_1506,N_29475,N_27480);
nand UO_1507 (O_1507,N_29388,N_27570);
xor UO_1508 (O_1508,N_27127,N_29989);
xor UO_1509 (O_1509,N_29171,N_29989);
nor UO_1510 (O_1510,N_29601,N_29841);
and UO_1511 (O_1511,N_28529,N_27051);
nand UO_1512 (O_1512,N_28467,N_27180);
nor UO_1513 (O_1513,N_29400,N_29935);
nor UO_1514 (O_1514,N_28100,N_29836);
nor UO_1515 (O_1515,N_27852,N_27629);
nand UO_1516 (O_1516,N_28916,N_29142);
and UO_1517 (O_1517,N_27310,N_28748);
or UO_1518 (O_1518,N_29445,N_28677);
and UO_1519 (O_1519,N_29352,N_27063);
nor UO_1520 (O_1520,N_28447,N_29801);
nor UO_1521 (O_1521,N_27044,N_27806);
nor UO_1522 (O_1522,N_29406,N_27885);
nand UO_1523 (O_1523,N_27837,N_29258);
or UO_1524 (O_1524,N_27350,N_29313);
xnor UO_1525 (O_1525,N_29057,N_29231);
xor UO_1526 (O_1526,N_27960,N_28126);
and UO_1527 (O_1527,N_28720,N_28408);
and UO_1528 (O_1528,N_28153,N_29652);
nand UO_1529 (O_1529,N_28047,N_27885);
nand UO_1530 (O_1530,N_27286,N_29601);
and UO_1531 (O_1531,N_29583,N_29128);
and UO_1532 (O_1532,N_29256,N_27155);
or UO_1533 (O_1533,N_28616,N_27893);
nor UO_1534 (O_1534,N_29431,N_29651);
and UO_1535 (O_1535,N_29087,N_27226);
xnor UO_1536 (O_1536,N_29263,N_28120);
nand UO_1537 (O_1537,N_28342,N_29280);
nor UO_1538 (O_1538,N_28012,N_29620);
nor UO_1539 (O_1539,N_29265,N_29634);
or UO_1540 (O_1540,N_29043,N_28291);
xor UO_1541 (O_1541,N_27329,N_29992);
xor UO_1542 (O_1542,N_28910,N_27452);
nand UO_1543 (O_1543,N_29136,N_28400);
and UO_1544 (O_1544,N_28305,N_27859);
and UO_1545 (O_1545,N_29312,N_29529);
nand UO_1546 (O_1546,N_29336,N_29359);
nor UO_1547 (O_1547,N_29385,N_27016);
nand UO_1548 (O_1548,N_28007,N_27085);
and UO_1549 (O_1549,N_28382,N_27154);
nand UO_1550 (O_1550,N_28728,N_27528);
xor UO_1551 (O_1551,N_28523,N_27092);
nor UO_1552 (O_1552,N_28597,N_27893);
or UO_1553 (O_1553,N_27371,N_28948);
or UO_1554 (O_1554,N_28985,N_28228);
nand UO_1555 (O_1555,N_27085,N_27179);
xor UO_1556 (O_1556,N_28676,N_27457);
and UO_1557 (O_1557,N_28240,N_28111);
xnor UO_1558 (O_1558,N_29838,N_29742);
nor UO_1559 (O_1559,N_27728,N_29266);
xnor UO_1560 (O_1560,N_28679,N_28038);
nand UO_1561 (O_1561,N_27831,N_27713);
and UO_1562 (O_1562,N_28499,N_29305);
nand UO_1563 (O_1563,N_27213,N_28707);
xnor UO_1564 (O_1564,N_28365,N_28245);
xor UO_1565 (O_1565,N_29055,N_29350);
nor UO_1566 (O_1566,N_28796,N_27456);
and UO_1567 (O_1567,N_28898,N_29284);
nand UO_1568 (O_1568,N_28683,N_28105);
nor UO_1569 (O_1569,N_27462,N_28726);
xnor UO_1570 (O_1570,N_27870,N_27689);
and UO_1571 (O_1571,N_27722,N_27757);
nand UO_1572 (O_1572,N_27151,N_27640);
nand UO_1573 (O_1573,N_29814,N_27596);
or UO_1574 (O_1574,N_29323,N_29922);
xor UO_1575 (O_1575,N_27799,N_28811);
or UO_1576 (O_1576,N_28729,N_28345);
and UO_1577 (O_1577,N_27672,N_28001);
or UO_1578 (O_1578,N_29412,N_29876);
or UO_1579 (O_1579,N_29421,N_27977);
and UO_1580 (O_1580,N_29577,N_28418);
and UO_1581 (O_1581,N_27108,N_28185);
nand UO_1582 (O_1582,N_27248,N_29589);
xnor UO_1583 (O_1583,N_28726,N_29909);
nand UO_1584 (O_1584,N_27982,N_27046);
xnor UO_1585 (O_1585,N_27163,N_28023);
nand UO_1586 (O_1586,N_28239,N_29171);
xnor UO_1587 (O_1587,N_27396,N_29836);
and UO_1588 (O_1588,N_29556,N_28833);
nor UO_1589 (O_1589,N_28382,N_29891);
nand UO_1590 (O_1590,N_28850,N_27904);
nand UO_1591 (O_1591,N_29655,N_28246);
or UO_1592 (O_1592,N_29140,N_29793);
or UO_1593 (O_1593,N_27609,N_28566);
xor UO_1594 (O_1594,N_28799,N_29744);
nor UO_1595 (O_1595,N_28576,N_28534);
or UO_1596 (O_1596,N_28999,N_29540);
or UO_1597 (O_1597,N_29348,N_29928);
and UO_1598 (O_1598,N_29002,N_27380);
and UO_1599 (O_1599,N_27312,N_27249);
or UO_1600 (O_1600,N_27618,N_27362);
nand UO_1601 (O_1601,N_29148,N_28757);
xor UO_1602 (O_1602,N_28156,N_29573);
nor UO_1603 (O_1603,N_27805,N_28591);
nor UO_1604 (O_1604,N_29520,N_27004);
xor UO_1605 (O_1605,N_29858,N_27914);
nand UO_1606 (O_1606,N_29767,N_28646);
nor UO_1607 (O_1607,N_28193,N_28669);
and UO_1608 (O_1608,N_29774,N_27490);
and UO_1609 (O_1609,N_29761,N_27763);
nand UO_1610 (O_1610,N_28596,N_27205);
nand UO_1611 (O_1611,N_28075,N_27474);
nand UO_1612 (O_1612,N_29351,N_29699);
xor UO_1613 (O_1613,N_28697,N_28228);
nor UO_1614 (O_1614,N_27110,N_27037);
xnor UO_1615 (O_1615,N_28442,N_29414);
and UO_1616 (O_1616,N_29793,N_29338);
and UO_1617 (O_1617,N_27620,N_29524);
xnor UO_1618 (O_1618,N_28656,N_27093);
and UO_1619 (O_1619,N_29356,N_27255);
nand UO_1620 (O_1620,N_29759,N_28720);
and UO_1621 (O_1621,N_29782,N_29614);
and UO_1622 (O_1622,N_28513,N_28946);
nand UO_1623 (O_1623,N_27162,N_29544);
nand UO_1624 (O_1624,N_28055,N_29167);
or UO_1625 (O_1625,N_28028,N_29159);
and UO_1626 (O_1626,N_28795,N_27285);
xnor UO_1627 (O_1627,N_28731,N_27946);
xnor UO_1628 (O_1628,N_29341,N_27846);
nand UO_1629 (O_1629,N_28866,N_28331);
xor UO_1630 (O_1630,N_28777,N_29685);
nor UO_1631 (O_1631,N_28434,N_27348);
nand UO_1632 (O_1632,N_27396,N_29577);
or UO_1633 (O_1633,N_29047,N_29671);
nor UO_1634 (O_1634,N_28730,N_28031);
nor UO_1635 (O_1635,N_27303,N_27970);
xor UO_1636 (O_1636,N_27307,N_29174);
xnor UO_1637 (O_1637,N_28551,N_27345);
and UO_1638 (O_1638,N_27006,N_27143);
and UO_1639 (O_1639,N_29122,N_28710);
or UO_1640 (O_1640,N_28495,N_28840);
nor UO_1641 (O_1641,N_28775,N_29957);
and UO_1642 (O_1642,N_29599,N_28493);
xnor UO_1643 (O_1643,N_28945,N_27889);
nor UO_1644 (O_1644,N_29515,N_28570);
xnor UO_1645 (O_1645,N_27182,N_28727);
xnor UO_1646 (O_1646,N_27487,N_29116);
nor UO_1647 (O_1647,N_28969,N_28976);
xnor UO_1648 (O_1648,N_28162,N_28460);
or UO_1649 (O_1649,N_28981,N_29639);
xor UO_1650 (O_1650,N_28399,N_27418);
or UO_1651 (O_1651,N_28933,N_29866);
xor UO_1652 (O_1652,N_27683,N_27969);
nor UO_1653 (O_1653,N_27608,N_28358);
and UO_1654 (O_1654,N_28176,N_29209);
nand UO_1655 (O_1655,N_29112,N_29703);
nor UO_1656 (O_1656,N_28220,N_28631);
and UO_1657 (O_1657,N_27546,N_28253);
nor UO_1658 (O_1658,N_29801,N_28017);
xor UO_1659 (O_1659,N_29448,N_28346);
and UO_1660 (O_1660,N_28511,N_28204);
xnor UO_1661 (O_1661,N_28173,N_29236);
and UO_1662 (O_1662,N_29524,N_27621);
and UO_1663 (O_1663,N_28749,N_29746);
or UO_1664 (O_1664,N_29864,N_28424);
xor UO_1665 (O_1665,N_28917,N_27632);
xnor UO_1666 (O_1666,N_28664,N_29905);
nand UO_1667 (O_1667,N_27740,N_27634);
and UO_1668 (O_1668,N_27345,N_28821);
and UO_1669 (O_1669,N_27851,N_28465);
nand UO_1670 (O_1670,N_29623,N_27342);
and UO_1671 (O_1671,N_27314,N_27820);
xor UO_1672 (O_1672,N_28483,N_27436);
or UO_1673 (O_1673,N_28081,N_27336);
xnor UO_1674 (O_1674,N_27297,N_27561);
nand UO_1675 (O_1675,N_27050,N_29798);
nor UO_1676 (O_1676,N_29223,N_27098);
or UO_1677 (O_1677,N_29683,N_28236);
nor UO_1678 (O_1678,N_29831,N_29351);
and UO_1679 (O_1679,N_28702,N_27520);
xor UO_1680 (O_1680,N_27795,N_29427);
nand UO_1681 (O_1681,N_27537,N_29052);
nand UO_1682 (O_1682,N_28865,N_28531);
and UO_1683 (O_1683,N_27943,N_29797);
nor UO_1684 (O_1684,N_28161,N_27729);
nand UO_1685 (O_1685,N_29077,N_28638);
nor UO_1686 (O_1686,N_29714,N_28297);
nor UO_1687 (O_1687,N_28581,N_29351);
nand UO_1688 (O_1688,N_29533,N_28501);
or UO_1689 (O_1689,N_28076,N_29765);
nand UO_1690 (O_1690,N_27338,N_27122);
xor UO_1691 (O_1691,N_29654,N_29577);
or UO_1692 (O_1692,N_29258,N_28793);
nor UO_1693 (O_1693,N_29241,N_29895);
and UO_1694 (O_1694,N_29664,N_29792);
xor UO_1695 (O_1695,N_29441,N_29227);
or UO_1696 (O_1696,N_27431,N_27544);
nand UO_1697 (O_1697,N_27748,N_29764);
nand UO_1698 (O_1698,N_28435,N_28961);
nor UO_1699 (O_1699,N_28575,N_27022);
or UO_1700 (O_1700,N_27958,N_28711);
nand UO_1701 (O_1701,N_27866,N_28050);
and UO_1702 (O_1702,N_27247,N_28961);
or UO_1703 (O_1703,N_28461,N_29113);
nor UO_1704 (O_1704,N_28981,N_28448);
or UO_1705 (O_1705,N_29318,N_29356);
xnor UO_1706 (O_1706,N_29142,N_27328);
or UO_1707 (O_1707,N_27323,N_29008);
nand UO_1708 (O_1708,N_28825,N_27375);
xnor UO_1709 (O_1709,N_29666,N_28800);
nand UO_1710 (O_1710,N_28937,N_29579);
xor UO_1711 (O_1711,N_28762,N_28732);
or UO_1712 (O_1712,N_29994,N_29744);
and UO_1713 (O_1713,N_28256,N_29894);
or UO_1714 (O_1714,N_27487,N_29245);
and UO_1715 (O_1715,N_29867,N_28410);
or UO_1716 (O_1716,N_28603,N_29336);
nor UO_1717 (O_1717,N_28491,N_29481);
and UO_1718 (O_1718,N_29008,N_29557);
or UO_1719 (O_1719,N_28264,N_28602);
and UO_1720 (O_1720,N_27562,N_27561);
or UO_1721 (O_1721,N_29153,N_28379);
nand UO_1722 (O_1722,N_27125,N_27426);
or UO_1723 (O_1723,N_28636,N_27651);
xor UO_1724 (O_1724,N_29949,N_28093);
xor UO_1725 (O_1725,N_29434,N_27455);
xnor UO_1726 (O_1726,N_27091,N_27266);
and UO_1727 (O_1727,N_27921,N_27357);
or UO_1728 (O_1728,N_28874,N_27733);
nand UO_1729 (O_1729,N_27206,N_29942);
nand UO_1730 (O_1730,N_27120,N_27289);
and UO_1731 (O_1731,N_28340,N_28162);
and UO_1732 (O_1732,N_28496,N_29756);
and UO_1733 (O_1733,N_27793,N_28677);
nand UO_1734 (O_1734,N_29428,N_28507);
xnor UO_1735 (O_1735,N_29980,N_29191);
nor UO_1736 (O_1736,N_29178,N_28538);
xor UO_1737 (O_1737,N_27156,N_28645);
xor UO_1738 (O_1738,N_27924,N_29574);
or UO_1739 (O_1739,N_27083,N_27638);
nor UO_1740 (O_1740,N_27469,N_29486);
nand UO_1741 (O_1741,N_28711,N_29720);
nor UO_1742 (O_1742,N_28274,N_27449);
or UO_1743 (O_1743,N_28692,N_27354);
nor UO_1744 (O_1744,N_29635,N_29437);
nand UO_1745 (O_1745,N_27097,N_27281);
or UO_1746 (O_1746,N_28474,N_28759);
or UO_1747 (O_1747,N_29150,N_28980);
or UO_1748 (O_1748,N_28388,N_28689);
xor UO_1749 (O_1749,N_28434,N_28055);
nor UO_1750 (O_1750,N_29683,N_28584);
xor UO_1751 (O_1751,N_27658,N_27892);
and UO_1752 (O_1752,N_28596,N_27674);
nor UO_1753 (O_1753,N_29647,N_27148);
nand UO_1754 (O_1754,N_27340,N_29319);
or UO_1755 (O_1755,N_29621,N_27252);
and UO_1756 (O_1756,N_28529,N_29562);
nand UO_1757 (O_1757,N_27744,N_27366);
or UO_1758 (O_1758,N_27614,N_29615);
nor UO_1759 (O_1759,N_27683,N_27792);
nand UO_1760 (O_1760,N_29467,N_27071);
or UO_1761 (O_1761,N_27753,N_29103);
or UO_1762 (O_1762,N_29898,N_27055);
or UO_1763 (O_1763,N_27519,N_27238);
or UO_1764 (O_1764,N_28042,N_29305);
xor UO_1765 (O_1765,N_27554,N_28834);
xnor UO_1766 (O_1766,N_29228,N_27877);
or UO_1767 (O_1767,N_29129,N_29720);
nor UO_1768 (O_1768,N_29780,N_28932);
xor UO_1769 (O_1769,N_27055,N_28368);
xnor UO_1770 (O_1770,N_29623,N_27530);
or UO_1771 (O_1771,N_27049,N_29539);
or UO_1772 (O_1772,N_27264,N_29440);
or UO_1773 (O_1773,N_27360,N_27373);
nor UO_1774 (O_1774,N_29140,N_27727);
nand UO_1775 (O_1775,N_29355,N_28851);
or UO_1776 (O_1776,N_27764,N_28195);
and UO_1777 (O_1777,N_29030,N_27451);
nand UO_1778 (O_1778,N_29343,N_28676);
and UO_1779 (O_1779,N_29844,N_29930);
or UO_1780 (O_1780,N_28642,N_27959);
xnor UO_1781 (O_1781,N_27687,N_27593);
xnor UO_1782 (O_1782,N_29984,N_29620);
or UO_1783 (O_1783,N_27400,N_28462);
xnor UO_1784 (O_1784,N_27620,N_29079);
nand UO_1785 (O_1785,N_29041,N_27002);
nor UO_1786 (O_1786,N_27709,N_29766);
nand UO_1787 (O_1787,N_28086,N_27552);
nand UO_1788 (O_1788,N_29271,N_28662);
nand UO_1789 (O_1789,N_28519,N_27703);
nor UO_1790 (O_1790,N_28135,N_29125);
or UO_1791 (O_1791,N_28709,N_27178);
and UO_1792 (O_1792,N_29584,N_28017);
and UO_1793 (O_1793,N_28042,N_27132);
xor UO_1794 (O_1794,N_28411,N_29612);
nand UO_1795 (O_1795,N_29041,N_28115);
and UO_1796 (O_1796,N_28348,N_28096);
and UO_1797 (O_1797,N_29511,N_27746);
or UO_1798 (O_1798,N_27240,N_29586);
and UO_1799 (O_1799,N_28544,N_29850);
nand UO_1800 (O_1800,N_28698,N_28171);
nand UO_1801 (O_1801,N_28545,N_27062);
nor UO_1802 (O_1802,N_28029,N_28586);
or UO_1803 (O_1803,N_28692,N_29560);
nand UO_1804 (O_1804,N_29962,N_28755);
nand UO_1805 (O_1805,N_29123,N_28654);
nor UO_1806 (O_1806,N_28603,N_27561);
or UO_1807 (O_1807,N_29310,N_28661);
and UO_1808 (O_1808,N_29214,N_29464);
xnor UO_1809 (O_1809,N_27694,N_27948);
nand UO_1810 (O_1810,N_27693,N_28049);
nand UO_1811 (O_1811,N_29566,N_29891);
or UO_1812 (O_1812,N_27378,N_27477);
nor UO_1813 (O_1813,N_28631,N_28137);
or UO_1814 (O_1814,N_28383,N_27312);
xnor UO_1815 (O_1815,N_28660,N_29354);
and UO_1816 (O_1816,N_29758,N_28764);
xor UO_1817 (O_1817,N_27728,N_27302);
nor UO_1818 (O_1818,N_28687,N_29021);
xnor UO_1819 (O_1819,N_29105,N_28233);
or UO_1820 (O_1820,N_29668,N_27148);
xor UO_1821 (O_1821,N_27466,N_29871);
and UO_1822 (O_1822,N_29520,N_28267);
or UO_1823 (O_1823,N_27889,N_29277);
nor UO_1824 (O_1824,N_28375,N_28684);
xor UO_1825 (O_1825,N_28987,N_27444);
xnor UO_1826 (O_1826,N_29021,N_28869);
nor UO_1827 (O_1827,N_27323,N_28455);
or UO_1828 (O_1828,N_27583,N_29181);
nand UO_1829 (O_1829,N_28756,N_29955);
and UO_1830 (O_1830,N_28837,N_28695);
and UO_1831 (O_1831,N_28105,N_28578);
nand UO_1832 (O_1832,N_27399,N_27899);
nor UO_1833 (O_1833,N_28866,N_29532);
xor UO_1834 (O_1834,N_28419,N_29054);
and UO_1835 (O_1835,N_27647,N_29174);
nand UO_1836 (O_1836,N_27916,N_27703);
xor UO_1837 (O_1837,N_27971,N_27981);
nand UO_1838 (O_1838,N_27936,N_28940);
and UO_1839 (O_1839,N_27512,N_27268);
and UO_1840 (O_1840,N_28831,N_28527);
and UO_1841 (O_1841,N_28893,N_28575);
or UO_1842 (O_1842,N_28152,N_28164);
and UO_1843 (O_1843,N_28471,N_27731);
nor UO_1844 (O_1844,N_27341,N_29176);
or UO_1845 (O_1845,N_27565,N_28275);
xor UO_1846 (O_1846,N_27139,N_29268);
nand UO_1847 (O_1847,N_29010,N_29800);
nor UO_1848 (O_1848,N_28201,N_27673);
nor UO_1849 (O_1849,N_28127,N_27969);
nand UO_1850 (O_1850,N_27741,N_29193);
or UO_1851 (O_1851,N_27282,N_28495);
xor UO_1852 (O_1852,N_29494,N_28715);
nand UO_1853 (O_1853,N_27344,N_29201);
nand UO_1854 (O_1854,N_29918,N_29743);
nand UO_1855 (O_1855,N_28610,N_29750);
or UO_1856 (O_1856,N_27417,N_28791);
nor UO_1857 (O_1857,N_29021,N_27228);
or UO_1858 (O_1858,N_29782,N_27456);
nor UO_1859 (O_1859,N_27516,N_29449);
nand UO_1860 (O_1860,N_28122,N_28225);
or UO_1861 (O_1861,N_28736,N_28982);
and UO_1862 (O_1862,N_29148,N_27933);
nor UO_1863 (O_1863,N_29959,N_28900);
nor UO_1864 (O_1864,N_28997,N_29102);
nand UO_1865 (O_1865,N_29608,N_29126);
and UO_1866 (O_1866,N_29911,N_28765);
xor UO_1867 (O_1867,N_28141,N_29277);
nand UO_1868 (O_1868,N_28356,N_28824);
nand UO_1869 (O_1869,N_28497,N_28060);
nor UO_1870 (O_1870,N_27578,N_27027);
and UO_1871 (O_1871,N_29412,N_27398);
xnor UO_1872 (O_1872,N_28038,N_28542);
and UO_1873 (O_1873,N_27986,N_27103);
or UO_1874 (O_1874,N_29740,N_28501);
nand UO_1875 (O_1875,N_28482,N_27368);
or UO_1876 (O_1876,N_29091,N_27165);
and UO_1877 (O_1877,N_29408,N_27055);
and UO_1878 (O_1878,N_27723,N_28965);
xor UO_1879 (O_1879,N_29589,N_29854);
xor UO_1880 (O_1880,N_29960,N_29681);
xnor UO_1881 (O_1881,N_27216,N_27441);
nand UO_1882 (O_1882,N_29842,N_29158);
xnor UO_1883 (O_1883,N_29811,N_27504);
nor UO_1884 (O_1884,N_28931,N_29367);
and UO_1885 (O_1885,N_29649,N_28285);
and UO_1886 (O_1886,N_27180,N_29177);
nand UO_1887 (O_1887,N_27692,N_29196);
nand UO_1888 (O_1888,N_27249,N_29006);
xor UO_1889 (O_1889,N_29081,N_27520);
or UO_1890 (O_1890,N_28398,N_29990);
nand UO_1891 (O_1891,N_29460,N_29079);
nand UO_1892 (O_1892,N_27543,N_28016);
nand UO_1893 (O_1893,N_28798,N_27728);
or UO_1894 (O_1894,N_29417,N_29700);
and UO_1895 (O_1895,N_28162,N_28268);
nor UO_1896 (O_1896,N_28194,N_28456);
xnor UO_1897 (O_1897,N_27426,N_29410);
nand UO_1898 (O_1898,N_28019,N_28385);
or UO_1899 (O_1899,N_29866,N_27781);
xnor UO_1900 (O_1900,N_28380,N_29854);
xor UO_1901 (O_1901,N_27917,N_29682);
nor UO_1902 (O_1902,N_29928,N_28826);
nor UO_1903 (O_1903,N_27592,N_29838);
nand UO_1904 (O_1904,N_27599,N_29685);
nor UO_1905 (O_1905,N_29805,N_27015);
nor UO_1906 (O_1906,N_28058,N_27516);
nor UO_1907 (O_1907,N_28563,N_28494);
xor UO_1908 (O_1908,N_27411,N_28242);
or UO_1909 (O_1909,N_28131,N_29737);
and UO_1910 (O_1910,N_28596,N_27536);
nor UO_1911 (O_1911,N_27457,N_28331);
and UO_1912 (O_1912,N_28865,N_27916);
nand UO_1913 (O_1913,N_28963,N_27887);
or UO_1914 (O_1914,N_29932,N_28072);
and UO_1915 (O_1915,N_27369,N_29916);
nor UO_1916 (O_1916,N_28355,N_28302);
nand UO_1917 (O_1917,N_28944,N_28820);
or UO_1918 (O_1918,N_27037,N_29463);
or UO_1919 (O_1919,N_29011,N_28411);
and UO_1920 (O_1920,N_29402,N_29051);
nor UO_1921 (O_1921,N_29891,N_29939);
and UO_1922 (O_1922,N_29734,N_28050);
xor UO_1923 (O_1923,N_28979,N_28532);
or UO_1924 (O_1924,N_29345,N_27576);
or UO_1925 (O_1925,N_27457,N_28564);
nor UO_1926 (O_1926,N_28106,N_28452);
nand UO_1927 (O_1927,N_28915,N_29490);
nand UO_1928 (O_1928,N_29590,N_28513);
xnor UO_1929 (O_1929,N_28255,N_28745);
nand UO_1930 (O_1930,N_28092,N_27825);
nand UO_1931 (O_1931,N_27774,N_29258);
xor UO_1932 (O_1932,N_29646,N_27740);
or UO_1933 (O_1933,N_27741,N_28629);
xnor UO_1934 (O_1934,N_28575,N_27097);
xor UO_1935 (O_1935,N_28811,N_29119);
nor UO_1936 (O_1936,N_27557,N_28844);
xor UO_1937 (O_1937,N_29905,N_28343);
or UO_1938 (O_1938,N_27208,N_29082);
xnor UO_1939 (O_1939,N_27184,N_29113);
nor UO_1940 (O_1940,N_27967,N_29156);
or UO_1941 (O_1941,N_27063,N_29698);
and UO_1942 (O_1942,N_28627,N_29190);
xor UO_1943 (O_1943,N_29079,N_29525);
nand UO_1944 (O_1944,N_29647,N_27924);
nand UO_1945 (O_1945,N_29426,N_29494);
xor UO_1946 (O_1946,N_27885,N_27579);
xor UO_1947 (O_1947,N_27819,N_27052);
nand UO_1948 (O_1948,N_29172,N_29906);
and UO_1949 (O_1949,N_27042,N_27431);
nor UO_1950 (O_1950,N_29325,N_27045);
xnor UO_1951 (O_1951,N_27620,N_28682);
nor UO_1952 (O_1952,N_28428,N_27299);
and UO_1953 (O_1953,N_28679,N_29350);
xor UO_1954 (O_1954,N_28399,N_29249);
or UO_1955 (O_1955,N_29318,N_27235);
xor UO_1956 (O_1956,N_29244,N_27502);
xor UO_1957 (O_1957,N_29893,N_28136);
nand UO_1958 (O_1958,N_29844,N_29476);
nor UO_1959 (O_1959,N_27899,N_28243);
nor UO_1960 (O_1960,N_29332,N_27779);
nor UO_1961 (O_1961,N_28767,N_29721);
or UO_1962 (O_1962,N_27671,N_28271);
nand UO_1963 (O_1963,N_28738,N_27773);
xor UO_1964 (O_1964,N_29474,N_28124);
xnor UO_1965 (O_1965,N_29060,N_29328);
and UO_1966 (O_1966,N_29524,N_28917);
xnor UO_1967 (O_1967,N_27648,N_28374);
xnor UO_1968 (O_1968,N_27953,N_27913);
nor UO_1969 (O_1969,N_28115,N_27074);
nand UO_1970 (O_1970,N_29723,N_27521);
and UO_1971 (O_1971,N_27229,N_29306);
and UO_1972 (O_1972,N_29668,N_29252);
and UO_1973 (O_1973,N_29030,N_27563);
or UO_1974 (O_1974,N_27307,N_28056);
or UO_1975 (O_1975,N_28235,N_29423);
xor UO_1976 (O_1976,N_28350,N_29585);
or UO_1977 (O_1977,N_28220,N_27693);
or UO_1978 (O_1978,N_29665,N_28060);
or UO_1979 (O_1979,N_29199,N_28510);
and UO_1980 (O_1980,N_29118,N_28616);
or UO_1981 (O_1981,N_28162,N_28980);
nand UO_1982 (O_1982,N_29929,N_28155);
and UO_1983 (O_1983,N_27228,N_28437);
nand UO_1984 (O_1984,N_28050,N_27271);
nand UO_1985 (O_1985,N_28095,N_29911);
or UO_1986 (O_1986,N_29692,N_28456);
and UO_1987 (O_1987,N_27921,N_27654);
and UO_1988 (O_1988,N_27415,N_28199);
and UO_1989 (O_1989,N_29494,N_28275);
and UO_1990 (O_1990,N_27622,N_29361);
nor UO_1991 (O_1991,N_29072,N_27460);
or UO_1992 (O_1992,N_27087,N_27154);
and UO_1993 (O_1993,N_27648,N_28368);
nor UO_1994 (O_1994,N_28228,N_27365);
and UO_1995 (O_1995,N_27090,N_29926);
nor UO_1996 (O_1996,N_29027,N_28837);
or UO_1997 (O_1997,N_27687,N_27626);
nor UO_1998 (O_1998,N_27166,N_27501);
nand UO_1999 (O_1999,N_27056,N_29723);
nand UO_2000 (O_2000,N_27758,N_29078);
nand UO_2001 (O_2001,N_29861,N_27016);
xor UO_2002 (O_2002,N_29628,N_29072);
or UO_2003 (O_2003,N_28246,N_27798);
nand UO_2004 (O_2004,N_28172,N_28130);
xor UO_2005 (O_2005,N_29118,N_27371);
and UO_2006 (O_2006,N_27592,N_28576);
or UO_2007 (O_2007,N_29649,N_28656);
and UO_2008 (O_2008,N_28671,N_28362);
and UO_2009 (O_2009,N_28263,N_29458);
xnor UO_2010 (O_2010,N_27800,N_28099);
nor UO_2011 (O_2011,N_29105,N_27607);
xnor UO_2012 (O_2012,N_28253,N_27286);
nor UO_2013 (O_2013,N_28334,N_28007);
nand UO_2014 (O_2014,N_29540,N_29863);
or UO_2015 (O_2015,N_28641,N_27738);
and UO_2016 (O_2016,N_28364,N_29586);
nand UO_2017 (O_2017,N_29898,N_27320);
nand UO_2018 (O_2018,N_29793,N_27882);
nand UO_2019 (O_2019,N_28838,N_29914);
xnor UO_2020 (O_2020,N_29903,N_29303);
nor UO_2021 (O_2021,N_27556,N_28064);
and UO_2022 (O_2022,N_28196,N_28861);
or UO_2023 (O_2023,N_28151,N_27172);
nand UO_2024 (O_2024,N_27248,N_28937);
or UO_2025 (O_2025,N_28269,N_29833);
or UO_2026 (O_2026,N_29876,N_28643);
or UO_2027 (O_2027,N_29868,N_29841);
xor UO_2028 (O_2028,N_27560,N_29096);
and UO_2029 (O_2029,N_28994,N_29404);
nor UO_2030 (O_2030,N_29603,N_27651);
xor UO_2031 (O_2031,N_28631,N_29159);
nand UO_2032 (O_2032,N_27498,N_27711);
nand UO_2033 (O_2033,N_29209,N_29396);
or UO_2034 (O_2034,N_29817,N_28763);
nand UO_2035 (O_2035,N_29886,N_28951);
nor UO_2036 (O_2036,N_28028,N_29125);
or UO_2037 (O_2037,N_29241,N_27083);
and UO_2038 (O_2038,N_29708,N_29133);
and UO_2039 (O_2039,N_28462,N_27807);
xor UO_2040 (O_2040,N_29807,N_29954);
xor UO_2041 (O_2041,N_28929,N_29377);
nand UO_2042 (O_2042,N_28044,N_27598);
and UO_2043 (O_2043,N_28142,N_28171);
nand UO_2044 (O_2044,N_29140,N_29031);
nand UO_2045 (O_2045,N_28661,N_28341);
xor UO_2046 (O_2046,N_29707,N_29862);
nor UO_2047 (O_2047,N_29447,N_29695);
xnor UO_2048 (O_2048,N_28309,N_28565);
or UO_2049 (O_2049,N_29610,N_27206);
nor UO_2050 (O_2050,N_28379,N_29328);
nand UO_2051 (O_2051,N_28554,N_28887);
nand UO_2052 (O_2052,N_28313,N_28235);
or UO_2053 (O_2053,N_27092,N_29339);
or UO_2054 (O_2054,N_27924,N_29526);
nand UO_2055 (O_2055,N_28764,N_29866);
nand UO_2056 (O_2056,N_29752,N_27072);
and UO_2057 (O_2057,N_29894,N_27704);
and UO_2058 (O_2058,N_27509,N_28603);
xor UO_2059 (O_2059,N_28965,N_29635);
nor UO_2060 (O_2060,N_27146,N_28427);
xnor UO_2061 (O_2061,N_28088,N_27166);
nor UO_2062 (O_2062,N_28521,N_29571);
nor UO_2063 (O_2063,N_28819,N_27835);
nand UO_2064 (O_2064,N_27710,N_27085);
nand UO_2065 (O_2065,N_27353,N_27369);
nand UO_2066 (O_2066,N_27959,N_28715);
nand UO_2067 (O_2067,N_27628,N_29353);
nor UO_2068 (O_2068,N_28482,N_28767);
nor UO_2069 (O_2069,N_28182,N_28669);
nand UO_2070 (O_2070,N_27753,N_29590);
nand UO_2071 (O_2071,N_29191,N_29671);
or UO_2072 (O_2072,N_28340,N_29100);
xor UO_2073 (O_2073,N_28854,N_28014);
nor UO_2074 (O_2074,N_27895,N_28351);
or UO_2075 (O_2075,N_27291,N_29607);
and UO_2076 (O_2076,N_28584,N_27100);
nand UO_2077 (O_2077,N_28021,N_28221);
nor UO_2078 (O_2078,N_28205,N_28193);
and UO_2079 (O_2079,N_29423,N_27532);
nor UO_2080 (O_2080,N_28945,N_27334);
xor UO_2081 (O_2081,N_27313,N_29228);
xnor UO_2082 (O_2082,N_28964,N_29905);
nand UO_2083 (O_2083,N_29255,N_27458);
xor UO_2084 (O_2084,N_29467,N_29552);
nand UO_2085 (O_2085,N_27893,N_29428);
nand UO_2086 (O_2086,N_27924,N_29864);
nor UO_2087 (O_2087,N_27683,N_27546);
xor UO_2088 (O_2088,N_29793,N_29274);
xnor UO_2089 (O_2089,N_28647,N_27020);
nor UO_2090 (O_2090,N_28830,N_27836);
xor UO_2091 (O_2091,N_27049,N_29956);
and UO_2092 (O_2092,N_28434,N_27292);
nor UO_2093 (O_2093,N_28149,N_28571);
and UO_2094 (O_2094,N_28586,N_29292);
or UO_2095 (O_2095,N_27714,N_29278);
nand UO_2096 (O_2096,N_27897,N_29479);
or UO_2097 (O_2097,N_27620,N_28571);
or UO_2098 (O_2098,N_28033,N_28260);
xnor UO_2099 (O_2099,N_28227,N_29515);
and UO_2100 (O_2100,N_27840,N_27030);
and UO_2101 (O_2101,N_27777,N_28734);
and UO_2102 (O_2102,N_29305,N_27368);
or UO_2103 (O_2103,N_27968,N_27565);
xor UO_2104 (O_2104,N_27456,N_29137);
nor UO_2105 (O_2105,N_29459,N_29345);
nor UO_2106 (O_2106,N_28836,N_27738);
and UO_2107 (O_2107,N_28772,N_28876);
nor UO_2108 (O_2108,N_29541,N_29559);
or UO_2109 (O_2109,N_28303,N_27803);
nand UO_2110 (O_2110,N_29148,N_27828);
and UO_2111 (O_2111,N_29222,N_29664);
nor UO_2112 (O_2112,N_27822,N_29684);
xor UO_2113 (O_2113,N_29181,N_28660);
nand UO_2114 (O_2114,N_27767,N_29066);
xor UO_2115 (O_2115,N_27784,N_27881);
and UO_2116 (O_2116,N_28694,N_28448);
xnor UO_2117 (O_2117,N_27535,N_29128);
nor UO_2118 (O_2118,N_28243,N_28802);
or UO_2119 (O_2119,N_29689,N_28025);
or UO_2120 (O_2120,N_29199,N_27425);
nor UO_2121 (O_2121,N_28458,N_28435);
or UO_2122 (O_2122,N_29239,N_27407);
and UO_2123 (O_2123,N_27544,N_27578);
or UO_2124 (O_2124,N_28562,N_28479);
and UO_2125 (O_2125,N_28628,N_28874);
xor UO_2126 (O_2126,N_29516,N_29136);
and UO_2127 (O_2127,N_28195,N_29638);
nand UO_2128 (O_2128,N_29376,N_29791);
and UO_2129 (O_2129,N_27033,N_28939);
nand UO_2130 (O_2130,N_28248,N_27089);
xor UO_2131 (O_2131,N_27303,N_27917);
xnor UO_2132 (O_2132,N_27916,N_29280);
or UO_2133 (O_2133,N_27823,N_27982);
nor UO_2134 (O_2134,N_28887,N_27059);
nor UO_2135 (O_2135,N_28302,N_28601);
nor UO_2136 (O_2136,N_28762,N_27200);
and UO_2137 (O_2137,N_27363,N_29620);
and UO_2138 (O_2138,N_28383,N_29097);
and UO_2139 (O_2139,N_29456,N_28329);
and UO_2140 (O_2140,N_29205,N_28348);
and UO_2141 (O_2141,N_27890,N_28189);
or UO_2142 (O_2142,N_27522,N_28592);
or UO_2143 (O_2143,N_27878,N_28365);
and UO_2144 (O_2144,N_27561,N_29537);
nand UO_2145 (O_2145,N_29259,N_27894);
and UO_2146 (O_2146,N_29820,N_29777);
nand UO_2147 (O_2147,N_29736,N_28542);
xor UO_2148 (O_2148,N_28784,N_27705);
or UO_2149 (O_2149,N_29178,N_27804);
or UO_2150 (O_2150,N_28390,N_29252);
and UO_2151 (O_2151,N_29426,N_27494);
nor UO_2152 (O_2152,N_28560,N_27160);
and UO_2153 (O_2153,N_28935,N_27658);
or UO_2154 (O_2154,N_28106,N_28176);
xor UO_2155 (O_2155,N_28651,N_27576);
or UO_2156 (O_2156,N_27514,N_27110);
nor UO_2157 (O_2157,N_29933,N_29320);
xnor UO_2158 (O_2158,N_29284,N_28042);
and UO_2159 (O_2159,N_27465,N_27543);
xor UO_2160 (O_2160,N_28073,N_28893);
and UO_2161 (O_2161,N_29458,N_28228);
or UO_2162 (O_2162,N_28371,N_28348);
or UO_2163 (O_2163,N_27087,N_27185);
nand UO_2164 (O_2164,N_28286,N_29556);
nand UO_2165 (O_2165,N_29362,N_27288);
nand UO_2166 (O_2166,N_28099,N_29399);
and UO_2167 (O_2167,N_28122,N_27326);
and UO_2168 (O_2168,N_27182,N_29712);
nand UO_2169 (O_2169,N_29919,N_29400);
nor UO_2170 (O_2170,N_28316,N_29283);
or UO_2171 (O_2171,N_27840,N_29481);
xor UO_2172 (O_2172,N_29377,N_27179);
or UO_2173 (O_2173,N_28597,N_29179);
nand UO_2174 (O_2174,N_29469,N_28945);
or UO_2175 (O_2175,N_27126,N_28675);
and UO_2176 (O_2176,N_27425,N_27876);
and UO_2177 (O_2177,N_27896,N_27331);
nand UO_2178 (O_2178,N_27091,N_27694);
and UO_2179 (O_2179,N_29722,N_29097);
xnor UO_2180 (O_2180,N_27984,N_27702);
nor UO_2181 (O_2181,N_27707,N_29860);
xor UO_2182 (O_2182,N_28369,N_28998);
or UO_2183 (O_2183,N_28692,N_27381);
nand UO_2184 (O_2184,N_28439,N_29881);
or UO_2185 (O_2185,N_29777,N_27489);
nor UO_2186 (O_2186,N_27976,N_28950);
and UO_2187 (O_2187,N_27331,N_29933);
and UO_2188 (O_2188,N_27870,N_29937);
nor UO_2189 (O_2189,N_29978,N_28461);
and UO_2190 (O_2190,N_28216,N_28255);
nor UO_2191 (O_2191,N_29116,N_28795);
or UO_2192 (O_2192,N_27725,N_27035);
or UO_2193 (O_2193,N_28412,N_29627);
nor UO_2194 (O_2194,N_27279,N_27981);
nand UO_2195 (O_2195,N_29761,N_28300);
nor UO_2196 (O_2196,N_29435,N_28236);
nand UO_2197 (O_2197,N_28335,N_28494);
nand UO_2198 (O_2198,N_28082,N_28800);
nand UO_2199 (O_2199,N_27188,N_29394);
and UO_2200 (O_2200,N_29756,N_29068);
or UO_2201 (O_2201,N_28138,N_27931);
or UO_2202 (O_2202,N_29730,N_27807);
and UO_2203 (O_2203,N_29301,N_28131);
or UO_2204 (O_2204,N_28583,N_29803);
and UO_2205 (O_2205,N_28928,N_27911);
xnor UO_2206 (O_2206,N_29699,N_27119);
xor UO_2207 (O_2207,N_29201,N_29343);
nand UO_2208 (O_2208,N_27876,N_27524);
nor UO_2209 (O_2209,N_27621,N_27048);
nor UO_2210 (O_2210,N_27529,N_27840);
nand UO_2211 (O_2211,N_27843,N_28903);
or UO_2212 (O_2212,N_27195,N_28527);
xor UO_2213 (O_2213,N_27208,N_29207);
and UO_2214 (O_2214,N_28552,N_28176);
and UO_2215 (O_2215,N_29656,N_29079);
xor UO_2216 (O_2216,N_28423,N_28957);
xor UO_2217 (O_2217,N_28264,N_29117);
xor UO_2218 (O_2218,N_28519,N_28035);
nand UO_2219 (O_2219,N_29395,N_27580);
or UO_2220 (O_2220,N_29834,N_29269);
and UO_2221 (O_2221,N_29174,N_29754);
or UO_2222 (O_2222,N_28584,N_28947);
and UO_2223 (O_2223,N_29578,N_28153);
nand UO_2224 (O_2224,N_27168,N_29525);
xnor UO_2225 (O_2225,N_29823,N_27271);
xnor UO_2226 (O_2226,N_27797,N_28933);
and UO_2227 (O_2227,N_28025,N_27324);
or UO_2228 (O_2228,N_29350,N_28382);
nor UO_2229 (O_2229,N_27368,N_29927);
xnor UO_2230 (O_2230,N_27893,N_27181);
or UO_2231 (O_2231,N_28009,N_27517);
xnor UO_2232 (O_2232,N_28403,N_29282);
or UO_2233 (O_2233,N_29206,N_28767);
and UO_2234 (O_2234,N_29101,N_29567);
or UO_2235 (O_2235,N_27344,N_28622);
or UO_2236 (O_2236,N_28093,N_29277);
xnor UO_2237 (O_2237,N_28389,N_27771);
or UO_2238 (O_2238,N_28350,N_29879);
and UO_2239 (O_2239,N_28360,N_28922);
nand UO_2240 (O_2240,N_29614,N_29628);
nand UO_2241 (O_2241,N_28907,N_28792);
and UO_2242 (O_2242,N_28888,N_29172);
xnor UO_2243 (O_2243,N_29290,N_28883);
xor UO_2244 (O_2244,N_29979,N_28159);
and UO_2245 (O_2245,N_28803,N_28259);
or UO_2246 (O_2246,N_28628,N_29070);
and UO_2247 (O_2247,N_29597,N_28062);
and UO_2248 (O_2248,N_28811,N_27327);
xnor UO_2249 (O_2249,N_27989,N_27082);
xnor UO_2250 (O_2250,N_27803,N_29334);
or UO_2251 (O_2251,N_28257,N_29649);
and UO_2252 (O_2252,N_28698,N_27852);
nand UO_2253 (O_2253,N_27305,N_27282);
and UO_2254 (O_2254,N_28540,N_29524);
nor UO_2255 (O_2255,N_27911,N_29263);
or UO_2256 (O_2256,N_28833,N_27880);
and UO_2257 (O_2257,N_28075,N_28595);
xor UO_2258 (O_2258,N_29728,N_29875);
xnor UO_2259 (O_2259,N_29316,N_27725);
xor UO_2260 (O_2260,N_27607,N_28355);
and UO_2261 (O_2261,N_28626,N_27654);
or UO_2262 (O_2262,N_27637,N_27107);
xor UO_2263 (O_2263,N_29018,N_27573);
xor UO_2264 (O_2264,N_28077,N_29039);
xor UO_2265 (O_2265,N_28891,N_28134);
xnor UO_2266 (O_2266,N_27474,N_27102);
and UO_2267 (O_2267,N_29774,N_27297);
xnor UO_2268 (O_2268,N_27841,N_29154);
and UO_2269 (O_2269,N_29556,N_29229);
nor UO_2270 (O_2270,N_27000,N_27181);
or UO_2271 (O_2271,N_28648,N_27427);
or UO_2272 (O_2272,N_27732,N_28710);
nor UO_2273 (O_2273,N_27512,N_28502);
nand UO_2274 (O_2274,N_29687,N_28236);
or UO_2275 (O_2275,N_28932,N_28270);
and UO_2276 (O_2276,N_28065,N_29805);
nand UO_2277 (O_2277,N_28480,N_29859);
nor UO_2278 (O_2278,N_29465,N_27395);
xor UO_2279 (O_2279,N_29359,N_29745);
nand UO_2280 (O_2280,N_29875,N_28990);
and UO_2281 (O_2281,N_27048,N_27602);
and UO_2282 (O_2282,N_28438,N_28321);
nand UO_2283 (O_2283,N_28554,N_28422);
or UO_2284 (O_2284,N_29556,N_29476);
nand UO_2285 (O_2285,N_28885,N_28435);
xor UO_2286 (O_2286,N_29849,N_27830);
xor UO_2287 (O_2287,N_27586,N_28867);
xnor UO_2288 (O_2288,N_28065,N_29054);
or UO_2289 (O_2289,N_27656,N_27645);
or UO_2290 (O_2290,N_27478,N_27199);
nor UO_2291 (O_2291,N_29863,N_29542);
xor UO_2292 (O_2292,N_28039,N_28763);
xor UO_2293 (O_2293,N_28299,N_28864);
nor UO_2294 (O_2294,N_27884,N_29664);
or UO_2295 (O_2295,N_29305,N_27489);
xor UO_2296 (O_2296,N_27932,N_28340);
nand UO_2297 (O_2297,N_27397,N_28236);
and UO_2298 (O_2298,N_27247,N_29204);
and UO_2299 (O_2299,N_29292,N_28778);
nor UO_2300 (O_2300,N_29943,N_27746);
nand UO_2301 (O_2301,N_27513,N_29672);
xnor UO_2302 (O_2302,N_28337,N_27555);
xnor UO_2303 (O_2303,N_28330,N_28924);
xor UO_2304 (O_2304,N_28422,N_27151);
nand UO_2305 (O_2305,N_28987,N_28625);
xnor UO_2306 (O_2306,N_29548,N_28226);
nand UO_2307 (O_2307,N_29263,N_29575);
or UO_2308 (O_2308,N_29121,N_28950);
xor UO_2309 (O_2309,N_28789,N_29536);
or UO_2310 (O_2310,N_29564,N_29137);
nand UO_2311 (O_2311,N_28335,N_28888);
or UO_2312 (O_2312,N_27883,N_27150);
nor UO_2313 (O_2313,N_27344,N_29687);
and UO_2314 (O_2314,N_27262,N_27379);
xor UO_2315 (O_2315,N_28113,N_28231);
or UO_2316 (O_2316,N_27548,N_27782);
or UO_2317 (O_2317,N_27206,N_27322);
xor UO_2318 (O_2318,N_29212,N_28244);
and UO_2319 (O_2319,N_29819,N_29061);
nor UO_2320 (O_2320,N_29796,N_29177);
or UO_2321 (O_2321,N_27662,N_28351);
and UO_2322 (O_2322,N_28150,N_28645);
nor UO_2323 (O_2323,N_27248,N_28288);
nand UO_2324 (O_2324,N_27064,N_27988);
xnor UO_2325 (O_2325,N_28374,N_29355);
and UO_2326 (O_2326,N_29025,N_28441);
nor UO_2327 (O_2327,N_29482,N_27627);
xnor UO_2328 (O_2328,N_29555,N_29857);
xor UO_2329 (O_2329,N_28670,N_29774);
and UO_2330 (O_2330,N_28063,N_27215);
nor UO_2331 (O_2331,N_27233,N_28294);
xnor UO_2332 (O_2332,N_27230,N_28264);
nand UO_2333 (O_2333,N_28272,N_29496);
nand UO_2334 (O_2334,N_29335,N_27304);
or UO_2335 (O_2335,N_27766,N_28644);
nor UO_2336 (O_2336,N_29682,N_27319);
nand UO_2337 (O_2337,N_29797,N_29230);
or UO_2338 (O_2338,N_29913,N_27766);
nor UO_2339 (O_2339,N_27496,N_29811);
xor UO_2340 (O_2340,N_29469,N_27967);
nand UO_2341 (O_2341,N_29688,N_29774);
xnor UO_2342 (O_2342,N_28229,N_28038);
and UO_2343 (O_2343,N_29972,N_29947);
nor UO_2344 (O_2344,N_28305,N_28961);
nor UO_2345 (O_2345,N_29603,N_28296);
nand UO_2346 (O_2346,N_28631,N_28074);
xor UO_2347 (O_2347,N_29835,N_29893);
and UO_2348 (O_2348,N_27763,N_29129);
nand UO_2349 (O_2349,N_29049,N_28113);
and UO_2350 (O_2350,N_27754,N_27106);
or UO_2351 (O_2351,N_27170,N_28950);
nor UO_2352 (O_2352,N_27647,N_27142);
xor UO_2353 (O_2353,N_28638,N_28518);
nor UO_2354 (O_2354,N_29963,N_28480);
xor UO_2355 (O_2355,N_27900,N_28416);
nand UO_2356 (O_2356,N_27774,N_27430);
and UO_2357 (O_2357,N_27849,N_27353);
nor UO_2358 (O_2358,N_27867,N_28822);
nor UO_2359 (O_2359,N_29527,N_28752);
nor UO_2360 (O_2360,N_27723,N_28220);
nand UO_2361 (O_2361,N_29693,N_29405);
xnor UO_2362 (O_2362,N_29058,N_27807);
xnor UO_2363 (O_2363,N_29498,N_29475);
and UO_2364 (O_2364,N_27723,N_29393);
or UO_2365 (O_2365,N_28906,N_28055);
nand UO_2366 (O_2366,N_29699,N_28894);
nor UO_2367 (O_2367,N_27482,N_29935);
or UO_2368 (O_2368,N_29744,N_29588);
and UO_2369 (O_2369,N_28960,N_28029);
and UO_2370 (O_2370,N_29468,N_27009);
or UO_2371 (O_2371,N_28436,N_27560);
or UO_2372 (O_2372,N_29961,N_28525);
or UO_2373 (O_2373,N_27158,N_29928);
xnor UO_2374 (O_2374,N_27336,N_28225);
nor UO_2375 (O_2375,N_29397,N_28473);
or UO_2376 (O_2376,N_29190,N_28020);
nand UO_2377 (O_2377,N_29004,N_28694);
or UO_2378 (O_2378,N_29718,N_28052);
nor UO_2379 (O_2379,N_27301,N_28664);
nor UO_2380 (O_2380,N_27957,N_28007);
and UO_2381 (O_2381,N_29588,N_27711);
xor UO_2382 (O_2382,N_28450,N_28437);
nor UO_2383 (O_2383,N_29184,N_29999);
and UO_2384 (O_2384,N_28570,N_28128);
or UO_2385 (O_2385,N_28276,N_29372);
and UO_2386 (O_2386,N_27912,N_29125);
nor UO_2387 (O_2387,N_28306,N_29613);
nor UO_2388 (O_2388,N_27168,N_27851);
and UO_2389 (O_2389,N_28257,N_29048);
nor UO_2390 (O_2390,N_27829,N_27399);
nor UO_2391 (O_2391,N_27126,N_28427);
or UO_2392 (O_2392,N_27748,N_28744);
nand UO_2393 (O_2393,N_29902,N_29924);
or UO_2394 (O_2394,N_29268,N_28197);
nand UO_2395 (O_2395,N_27336,N_27978);
nand UO_2396 (O_2396,N_27382,N_27129);
xor UO_2397 (O_2397,N_29756,N_27325);
and UO_2398 (O_2398,N_28490,N_29375);
or UO_2399 (O_2399,N_27432,N_27961);
and UO_2400 (O_2400,N_29096,N_28422);
nand UO_2401 (O_2401,N_28459,N_28853);
xor UO_2402 (O_2402,N_27505,N_29259);
nand UO_2403 (O_2403,N_29689,N_28788);
or UO_2404 (O_2404,N_28438,N_28606);
or UO_2405 (O_2405,N_29015,N_28099);
xor UO_2406 (O_2406,N_28579,N_27468);
nand UO_2407 (O_2407,N_29596,N_27760);
xor UO_2408 (O_2408,N_28388,N_27668);
and UO_2409 (O_2409,N_29220,N_29790);
xor UO_2410 (O_2410,N_29820,N_29773);
xor UO_2411 (O_2411,N_28370,N_28834);
nor UO_2412 (O_2412,N_27298,N_28991);
nor UO_2413 (O_2413,N_29683,N_27532);
nand UO_2414 (O_2414,N_27954,N_28961);
and UO_2415 (O_2415,N_27737,N_29261);
nand UO_2416 (O_2416,N_29181,N_29830);
xnor UO_2417 (O_2417,N_29872,N_27598);
or UO_2418 (O_2418,N_29381,N_29452);
nand UO_2419 (O_2419,N_28961,N_29814);
nor UO_2420 (O_2420,N_29616,N_29738);
or UO_2421 (O_2421,N_28770,N_28489);
nand UO_2422 (O_2422,N_28194,N_28452);
nor UO_2423 (O_2423,N_28312,N_27232);
or UO_2424 (O_2424,N_28844,N_28380);
or UO_2425 (O_2425,N_29334,N_27746);
and UO_2426 (O_2426,N_28059,N_27782);
nor UO_2427 (O_2427,N_28737,N_29138);
xnor UO_2428 (O_2428,N_29992,N_28972);
nand UO_2429 (O_2429,N_28231,N_27951);
nand UO_2430 (O_2430,N_28664,N_29583);
nand UO_2431 (O_2431,N_27435,N_28352);
xnor UO_2432 (O_2432,N_28876,N_29642);
and UO_2433 (O_2433,N_29878,N_28933);
nand UO_2434 (O_2434,N_28577,N_27235);
and UO_2435 (O_2435,N_27783,N_27892);
or UO_2436 (O_2436,N_27712,N_28778);
xor UO_2437 (O_2437,N_29876,N_27548);
or UO_2438 (O_2438,N_28528,N_28033);
and UO_2439 (O_2439,N_27789,N_27187);
or UO_2440 (O_2440,N_28184,N_28151);
and UO_2441 (O_2441,N_27786,N_28986);
xor UO_2442 (O_2442,N_28255,N_29392);
xor UO_2443 (O_2443,N_28419,N_28678);
nand UO_2444 (O_2444,N_28071,N_27335);
and UO_2445 (O_2445,N_27764,N_28033);
xor UO_2446 (O_2446,N_27247,N_28347);
nor UO_2447 (O_2447,N_29626,N_29603);
nand UO_2448 (O_2448,N_27850,N_29259);
and UO_2449 (O_2449,N_27332,N_29385);
xnor UO_2450 (O_2450,N_28396,N_28865);
or UO_2451 (O_2451,N_27785,N_29241);
nand UO_2452 (O_2452,N_28559,N_28552);
or UO_2453 (O_2453,N_28742,N_28135);
nor UO_2454 (O_2454,N_28594,N_29046);
or UO_2455 (O_2455,N_29650,N_27077);
or UO_2456 (O_2456,N_28330,N_27696);
nor UO_2457 (O_2457,N_29185,N_28611);
nor UO_2458 (O_2458,N_27078,N_29054);
and UO_2459 (O_2459,N_29703,N_27529);
or UO_2460 (O_2460,N_29168,N_27532);
nor UO_2461 (O_2461,N_29944,N_29323);
nor UO_2462 (O_2462,N_29421,N_28295);
or UO_2463 (O_2463,N_27736,N_27699);
nand UO_2464 (O_2464,N_27893,N_28347);
or UO_2465 (O_2465,N_27543,N_27686);
or UO_2466 (O_2466,N_29673,N_29593);
xnor UO_2467 (O_2467,N_28799,N_28383);
nor UO_2468 (O_2468,N_29417,N_27925);
xnor UO_2469 (O_2469,N_27482,N_27258);
nand UO_2470 (O_2470,N_29361,N_29305);
nor UO_2471 (O_2471,N_27776,N_28121);
nand UO_2472 (O_2472,N_28249,N_29374);
and UO_2473 (O_2473,N_27446,N_29307);
nand UO_2474 (O_2474,N_28080,N_28340);
and UO_2475 (O_2475,N_29353,N_27712);
or UO_2476 (O_2476,N_29120,N_27845);
or UO_2477 (O_2477,N_29704,N_28239);
nand UO_2478 (O_2478,N_28679,N_29434);
or UO_2479 (O_2479,N_28761,N_27759);
or UO_2480 (O_2480,N_29091,N_29653);
xnor UO_2481 (O_2481,N_27801,N_28411);
or UO_2482 (O_2482,N_27658,N_27583);
nand UO_2483 (O_2483,N_27468,N_27999);
nand UO_2484 (O_2484,N_28095,N_28949);
and UO_2485 (O_2485,N_29036,N_27878);
or UO_2486 (O_2486,N_27500,N_28241);
or UO_2487 (O_2487,N_27136,N_27940);
nand UO_2488 (O_2488,N_29784,N_28842);
and UO_2489 (O_2489,N_28033,N_27833);
nand UO_2490 (O_2490,N_29324,N_28136);
xor UO_2491 (O_2491,N_28600,N_27529);
or UO_2492 (O_2492,N_28651,N_28215);
xor UO_2493 (O_2493,N_28501,N_29942);
nor UO_2494 (O_2494,N_27133,N_27368);
xor UO_2495 (O_2495,N_27767,N_27712);
xor UO_2496 (O_2496,N_28096,N_29392);
or UO_2497 (O_2497,N_28946,N_28699);
xor UO_2498 (O_2498,N_29295,N_27609);
or UO_2499 (O_2499,N_27478,N_29203);
nor UO_2500 (O_2500,N_27447,N_29031);
nor UO_2501 (O_2501,N_29522,N_28763);
and UO_2502 (O_2502,N_28087,N_27971);
or UO_2503 (O_2503,N_29457,N_28406);
xor UO_2504 (O_2504,N_29360,N_27517);
xor UO_2505 (O_2505,N_29520,N_29786);
or UO_2506 (O_2506,N_28987,N_29688);
xor UO_2507 (O_2507,N_27825,N_28995);
nor UO_2508 (O_2508,N_27154,N_27524);
and UO_2509 (O_2509,N_29604,N_29610);
and UO_2510 (O_2510,N_29452,N_29387);
nand UO_2511 (O_2511,N_28730,N_29219);
nor UO_2512 (O_2512,N_27027,N_29637);
nand UO_2513 (O_2513,N_28978,N_27243);
nor UO_2514 (O_2514,N_28051,N_27642);
nor UO_2515 (O_2515,N_27593,N_28410);
and UO_2516 (O_2516,N_29766,N_27538);
nor UO_2517 (O_2517,N_27422,N_29134);
and UO_2518 (O_2518,N_27195,N_28008);
xnor UO_2519 (O_2519,N_28755,N_27723);
xor UO_2520 (O_2520,N_29972,N_27050);
xor UO_2521 (O_2521,N_28745,N_27329);
nand UO_2522 (O_2522,N_27092,N_29943);
xnor UO_2523 (O_2523,N_27725,N_28460);
nand UO_2524 (O_2524,N_29956,N_28565);
xor UO_2525 (O_2525,N_28395,N_27911);
or UO_2526 (O_2526,N_27099,N_27375);
nand UO_2527 (O_2527,N_27975,N_27395);
and UO_2528 (O_2528,N_27692,N_28331);
xor UO_2529 (O_2529,N_28195,N_28660);
xor UO_2530 (O_2530,N_27695,N_28206);
and UO_2531 (O_2531,N_28802,N_29473);
nor UO_2532 (O_2532,N_29923,N_29681);
xor UO_2533 (O_2533,N_29541,N_28220);
nand UO_2534 (O_2534,N_27264,N_27654);
nand UO_2535 (O_2535,N_27492,N_27472);
xnor UO_2536 (O_2536,N_28411,N_29168);
xnor UO_2537 (O_2537,N_28304,N_27186);
nor UO_2538 (O_2538,N_29476,N_27860);
and UO_2539 (O_2539,N_28741,N_28529);
and UO_2540 (O_2540,N_28108,N_27556);
nand UO_2541 (O_2541,N_27080,N_27823);
nor UO_2542 (O_2542,N_27958,N_27787);
nand UO_2543 (O_2543,N_29991,N_27273);
or UO_2544 (O_2544,N_28574,N_29197);
xor UO_2545 (O_2545,N_28677,N_29950);
or UO_2546 (O_2546,N_27325,N_27017);
and UO_2547 (O_2547,N_28849,N_29965);
xor UO_2548 (O_2548,N_27373,N_28931);
or UO_2549 (O_2549,N_29723,N_29740);
xor UO_2550 (O_2550,N_27540,N_29324);
xnor UO_2551 (O_2551,N_29677,N_27233);
nor UO_2552 (O_2552,N_28984,N_27748);
or UO_2553 (O_2553,N_27094,N_29480);
or UO_2554 (O_2554,N_28706,N_27624);
nor UO_2555 (O_2555,N_29569,N_28670);
nand UO_2556 (O_2556,N_28539,N_29885);
or UO_2557 (O_2557,N_29165,N_27327);
and UO_2558 (O_2558,N_29425,N_29114);
and UO_2559 (O_2559,N_27360,N_29179);
or UO_2560 (O_2560,N_27013,N_27869);
and UO_2561 (O_2561,N_27285,N_29548);
nand UO_2562 (O_2562,N_28860,N_29675);
or UO_2563 (O_2563,N_27380,N_28248);
nor UO_2564 (O_2564,N_29687,N_28957);
nor UO_2565 (O_2565,N_27005,N_28956);
nor UO_2566 (O_2566,N_28171,N_28293);
nor UO_2567 (O_2567,N_29826,N_29641);
and UO_2568 (O_2568,N_29853,N_28879);
nand UO_2569 (O_2569,N_28979,N_28104);
or UO_2570 (O_2570,N_27976,N_29396);
nor UO_2571 (O_2571,N_29513,N_28646);
xnor UO_2572 (O_2572,N_29568,N_27474);
nor UO_2573 (O_2573,N_28216,N_29977);
xor UO_2574 (O_2574,N_28713,N_29167);
nand UO_2575 (O_2575,N_29196,N_29246);
nand UO_2576 (O_2576,N_27945,N_29364);
xnor UO_2577 (O_2577,N_27169,N_29118);
nand UO_2578 (O_2578,N_29553,N_28829);
nand UO_2579 (O_2579,N_29926,N_29663);
xor UO_2580 (O_2580,N_27016,N_28018);
or UO_2581 (O_2581,N_28663,N_28214);
xnor UO_2582 (O_2582,N_28460,N_28790);
nand UO_2583 (O_2583,N_29904,N_28506);
nand UO_2584 (O_2584,N_29268,N_28529);
xor UO_2585 (O_2585,N_28219,N_29102);
nor UO_2586 (O_2586,N_27090,N_29907);
nand UO_2587 (O_2587,N_28602,N_27392);
and UO_2588 (O_2588,N_28460,N_28515);
xor UO_2589 (O_2589,N_29232,N_27506);
xor UO_2590 (O_2590,N_29847,N_28665);
xor UO_2591 (O_2591,N_29251,N_27068);
nor UO_2592 (O_2592,N_27258,N_29741);
or UO_2593 (O_2593,N_27678,N_27460);
or UO_2594 (O_2594,N_29673,N_27958);
nand UO_2595 (O_2595,N_29792,N_29111);
or UO_2596 (O_2596,N_29938,N_29615);
nand UO_2597 (O_2597,N_27650,N_29105);
and UO_2598 (O_2598,N_27460,N_29291);
or UO_2599 (O_2599,N_28960,N_27373);
or UO_2600 (O_2600,N_28946,N_27343);
or UO_2601 (O_2601,N_27326,N_28562);
nand UO_2602 (O_2602,N_28041,N_28096);
nand UO_2603 (O_2603,N_29215,N_28455);
nor UO_2604 (O_2604,N_28876,N_29071);
or UO_2605 (O_2605,N_27599,N_27780);
and UO_2606 (O_2606,N_27010,N_28991);
and UO_2607 (O_2607,N_29762,N_28330);
xor UO_2608 (O_2608,N_27265,N_28410);
xor UO_2609 (O_2609,N_28273,N_27261);
or UO_2610 (O_2610,N_27349,N_29714);
nand UO_2611 (O_2611,N_29614,N_28534);
and UO_2612 (O_2612,N_28808,N_29181);
or UO_2613 (O_2613,N_27294,N_28226);
or UO_2614 (O_2614,N_28785,N_27207);
or UO_2615 (O_2615,N_29278,N_27082);
xor UO_2616 (O_2616,N_28298,N_28899);
and UO_2617 (O_2617,N_28168,N_27031);
and UO_2618 (O_2618,N_29353,N_29542);
or UO_2619 (O_2619,N_29502,N_28239);
nand UO_2620 (O_2620,N_27315,N_27763);
and UO_2621 (O_2621,N_29841,N_27382);
xor UO_2622 (O_2622,N_28211,N_27554);
xor UO_2623 (O_2623,N_28604,N_28838);
and UO_2624 (O_2624,N_27436,N_28157);
nand UO_2625 (O_2625,N_29820,N_29408);
nand UO_2626 (O_2626,N_29326,N_27677);
or UO_2627 (O_2627,N_29521,N_27990);
nor UO_2628 (O_2628,N_29677,N_27150);
xor UO_2629 (O_2629,N_29731,N_28542);
nor UO_2630 (O_2630,N_28090,N_29872);
xor UO_2631 (O_2631,N_28107,N_29492);
or UO_2632 (O_2632,N_29145,N_27781);
or UO_2633 (O_2633,N_27079,N_28297);
and UO_2634 (O_2634,N_29040,N_29922);
and UO_2635 (O_2635,N_28391,N_29413);
xor UO_2636 (O_2636,N_29037,N_28225);
nand UO_2637 (O_2637,N_29147,N_29983);
nand UO_2638 (O_2638,N_28123,N_29449);
or UO_2639 (O_2639,N_27699,N_29363);
nor UO_2640 (O_2640,N_28081,N_29225);
or UO_2641 (O_2641,N_27416,N_28465);
and UO_2642 (O_2642,N_29577,N_29251);
nand UO_2643 (O_2643,N_29625,N_28705);
xor UO_2644 (O_2644,N_28318,N_28803);
nand UO_2645 (O_2645,N_29051,N_28662);
nand UO_2646 (O_2646,N_27155,N_27224);
and UO_2647 (O_2647,N_29399,N_29608);
and UO_2648 (O_2648,N_28308,N_29894);
nor UO_2649 (O_2649,N_27170,N_27873);
xnor UO_2650 (O_2650,N_27293,N_29859);
nand UO_2651 (O_2651,N_27625,N_28726);
nand UO_2652 (O_2652,N_27468,N_29812);
and UO_2653 (O_2653,N_29056,N_29708);
nand UO_2654 (O_2654,N_28523,N_27609);
and UO_2655 (O_2655,N_27823,N_27311);
or UO_2656 (O_2656,N_29310,N_29221);
nand UO_2657 (O_2657,N_29420,N_27627);
xor UO_2658 (O_2658,N_27419,N_28654);
nor UO_2659 (O_2659,N_27438,N_29226);
or UO_2660 (O_2660,N_28617,N_29231);
nor UO_2661 (O_2661,N_27703,N_28523);
xor UO_2662 (O_2662,N_27936,N_29139);
nand UO_2663 (O_2663,N_27644,N_29587);
xor UO_2664 (O_2664,N_29950,N_29402);
and UO_2665 (O_2665,N_27130,N_29012);
nand UO_2666 (O_2666,N_29358,N_27838);
xnor UO_2667 (O_2667,N_28787,N_29150);
and UO_2668 (O_2668,N_27690,N_28989);
nor UO_2669 (O_2669,N_27253,N_29809);
nand UO_2670 (O_2670,N_29799,N_29885);
and UO_2671 (O_2671,N_27027,N_27316);
xnor UO_2672 (O_2672,N_28187,N_29031);
nor UO_2673 (O_2673,N_28450,N_27471);
nand UO_2674 (O_2674,N_28872,N_29560);
or UO_2675 (O_2675,N_27218,N_27348);
and UO_2676 (O_2676,N_28252,N_27919);
and UO_2677 (O_2677,N_27200,N_27966);
nand UO_2678 (O_2678,N_28630,N_27741);
nor UO_2679 (O_2679,N_27477,N_28445);
nand UO_2680 (O_2680,N_28934,N_29939);
and UO_2681 (O_2681,N_29641,N_29689);
and UO_2682 (O_2682,N_29760,N_27229);
nand UO_2683 (O_2683,N_28034,N_28573);
and UO_2684 (O_2684,N_29568,N_28648);
xor UO_2685 (O_2685,N_28431,N_28929);
and UO_2686 (O_2686,N_29210,N_27356);
and UO_2687 (O_2687,N_27692,N_28442);
nand UO_2688 (O_2688,N_27778,N_28906);
and UO_2689 (O_2689,N_29830,N_27354);
and UO_2690 (O_2690,N_27755,N_29473);
and UO_2691 (O_2691,N_27204,N_28410);
nand UO_2692 (O_2692,N_27588,N_28014);
xor UO_2693 (O_2693,N_28776,N_28238);
nand UO_2694 (O_2694,N_29576,N_27276);
or UO_2695 (O_2695,N_28237,N_27442);
nand UO_2696 (O_2696,N_29252,N_29886);
and UO_2697 (O_2697,N_27938,N_29892);
nand UO_2698 (O_2698,N_29118,N_29070);
xor UO_2699 (O_2699,N_28533,N_29756);
or UO_2700 (O_2700,N_28817,N_28960);
nor UO_2701 (O_2701,N_29990,N_28846);
or UO_2702 (O_2702,N_28317,N_27924);
xnor UO_2703 (O_2703,N_28128,N_29637);
or UO_2704 (O_2704,N_28423,N_27495);
and UO_2705 (O_2705,N_28874,N_28476);
or UO_2706 (O_2706,N_27257,N_29751);
or UO_2707 (O_2707,N_28989,N_29087);
or UO_2708 (O_2708,N_29071,N_28058);
nand UO_2709 (O_2709,N_28168,N_27038);
nor UO_2710 (O_2710,N_29301,N_27460);
nor UO_2711 (O_2711,N_28582,N_28812);
nand UO_2712 (O_2712,N_27186,N_29934);
nand UO_2713 (O_2713,N_27996,N_27346);
and UO_2714 (O_2714,N_28542,N_29741);
xnor UO_2715 (O_2715,N_27324,N_29094);
nand UO_2716 (O_2716,N_29133,N_29172);
nor UO_2717 (O_2717,N_27268,N_29542);
and UO_2718 (O_2718,N_29389,N_28641);
or UO_2719 (O_2719,N_28475,N_28236);
and UO_2720 (O_2720,N_27659,N_28964);
nand UO_2721 (O_2721,N_28398,N_29742);
nand UO_2722 (O_2722,N_28899,N_28675);
nor UO_2723 (O_2723,N_27457,N_29122);
nand UO_2724 (O_2724,N_29508,N_27270);
or UO_2725 (O_2725,N_29036,N_27333);
nor UO_2726 (O_2726,N_28155,N_29832);
or UO_2727 (O_2727,N_28643,N_28289);
nand UO_2728 (O_2728,N_27067,N_27178);
or UO_2729 (O_2729,N_28797,N_29253);
nor UO_2730 (O_2730,N_29260,N_27894);
nor UO_2731 (O_2731,N_29154,N_28659);
xor UO_2732 (O_2732,N_27340,N_27994);
nand UO_2733 (O_2733,N_27516,N_29292);
and UO_2734 (O_2734,N_29838,N_28898);
nor UO_2735 (O_2735,N_29799,N_27484);
and UO_2736 (O_2736,N_27570,N_27766);
xor UO_2737 (O_2737,N_28561,N_27483);
nand UO_2738 (O_2738,N_28266,N_29871);
xor UO_2739 (O_2739,N_27005,N_29078);
or UO_2740 (O_2740,N_27310,N_29524);
nand UO_2741 (O_2741,N_29589,N_27488);
or UO_2742 (O_2742,N_28055,N_27540);
and UO_2743 (O_2743,N_27600,N_28213);
nor UO_2744 (O_2744,N_29667,N_27076);
nand UO_2745 (O_2745,N_27354,N_29407);
or UO_2746 (O_2746,N_29537,N_29355);
xor UO_2747 (O_2747,N_27855,N_29853);
nand UO_2748 (O_2748,N_28613,N_27185);
or UO_2749 (O_2749,N_27112,N_27741);
or UO_2750 (O_2750,N_28553,N_27293);
xor UO_2751 (O_2751,N_28126,N_27090);
nand UO_2752 (O_2752,N_29019,N_29747);
nor UO_2753 (O_2753,N_29848,N_27790);
and UO_2754 (O_2754,N_29446,N_29776);
xnor UO_2755 (O_2755,N_27456,N_28497);
nand UO_2756 (O_2756,N_29640,N_27020);
or UO_2757 (O_2757,N_29443,N_29888);
nand UO_2758 (O_2758,N_28554,N_27434);
xor UO_2759 (O_2759,N_28433,N_29372);
nor UO_2760 (O_2760,N_28575,N_27386);
nand UO_2761 (O_2761,N_28186,N_29036);
nor UO_2762 (O_2762,N_29323,N_29463);
and UO_2763 (O_2763,N_27003,N_27290);
nand UO_2764 (O_2764,N_29384,N_27932);
xor UO_2765 (O_2765,N_27625,N_28991);
nor UO_2766 (O_2766,N_27670,N_28381);
or UO_2767 (O_2767,N_28536,N_29391);
nor UO_2768 (O_2768,N_27049,N_27844);
xor UO_2769 (O_2769,N_28958,N_28113);
nor UO_2770 (O_2770,N_28913,N_29115);
xor UO_2771 (O_2771,N_28600,N_29872);
or UO_2772 (O_2772,N_28172,N_29856);
xnor UO_2773 (O_2773,N_28495,N_28293);
xor UO_2774 (O_2774,N_28312,N_28753);
or UO_2775 (O_2775,N_28477,N_29552);
and UO_2776 (O_2776,N_29971,N_29529);
and UO_2777 (O_2777,N_29297,N_29674);
xor UO_2778 (O_2778,N_27329,N_29982);
xor UO_2779 (O_2779,N_27386,N_28414);
nor UO_2780 (O_2780,N_27504,N_28368);
xnor UO_2781 (O_2781,N_29753,N_28846);
nand UO_2782 (O_2782,N_27346,N_29489);
nor UO_2783 (O_2783,N_28167,N_27068);
xnor UO_2784 (O_2784,N_27076,N_27349);
xor UO_2785 (O_2785,N_27177,N_27620);
or UO_2786 (O_2786,N_27084,N_29553);
nor UO_2787 (O_2787,N_27113,N_27771);
xnor UO_2788 (O_2788,N_29744,N_28682);
or UO_2789 (O_2789,N_29824,N_27735);
and UO_2790 (O_2790,N_28673,N_28577);
nand UO_2791 (O_2791,N_29496,N_28631);
nand UO_2792 (O_2792,N_28969,N_27100);
nand UO_2793 (O_2793,N_29469,N_29942);
nand UO_2794 (O_2794,N_28764,N_27752);
nand UO_2795 (O_2795,N_29386,N_28274);
or UO_2796 (O_2796,N_27832,N_28653);
nand UO_2797 (O_2797,N_29503,N_28413);
nor UO_2798 (O_2798,N_29515,N_27229);
and UO_2799 (O_2799,N_27503,N_27361);
nor UO_2800 (O_2800,N_29337,N_27780);
nand UO_2801 (O_2801,N_29458,N_28845);
xor UO_2802 (O_2802,N_27639,N_27876);
or UO_2803 (O_2803,N_27416,N_28020);
nand UO_2804 (O_2804,N_29820,N_27839);
nand UO_2805 (O_2805,N_27486,N_27465);
xnor UO_2806 (O_2806,N_29363,N_27818);
or UO_2807 (O_2807,N_27726,N_28467);
xnor UO_2808 (O_2808,N_29163,N_28919);
xor UO_2809 (O_2809,N_27919,N_28582);
nor UO_2810 (O_2810,N_27486,N_28118);
nor UO_2811 (O_2811,N_28108,N_27168);
xor UO_2812 (O_2812,N_28130,N_29129);
nor UO_2813 (O_2813,N_27082,N_28185);
nand UO_2814 (O_2814,N_29740,N_27002);
xnor UO_2815 (O_2815,N_29415,N_27618);
nor UO_2816 (O_2816,N_27373,N_27020);
nand UO_2817 (O_2817,N_29794,N_28876);
nor UO_2818 (O_2818,N_29208,N_28894);
nand UO_2819 (O_2819,N_29862,N_28363);
nand UO_2820 (O_2820,N_28746,N_29835);
and UO_2821 (O_2821,N_29366,N_27872);
or UO_2822 (O_2822,N_29858,N_29212);
and UO_2823 (O_2823,N_29197,N_29847);
xnor UO_2824 (O_2824,N_27653,N_27419);
nor UO_2825 (O_2825,N_28001,N_28703);
and UO_2826 (O_2826,N_29825,N_27203);
or UO_2827 (O_2827,N_27588,N_28638);
xnor UO_2828 (O_2828,N_29771,N_27506);
or UO_2829 (O_2829,N_27302,N_27295);
and UO_2830 (O_2830,N_27805,N_28993);
and UO_2831 (O_2831,N_27145,N_29500);
xor UO_2832 (O_2832,N_27782,N_29527);
nand UO_2833 (O_2833,N_29333,N_27953);
nand UO_2834 (O_2834,N_29578,N_27572);
xnor UO_2835 (O_2835,N_29580,N_28941);
xnor UO_2836 (O_2836,N_29792,N_28055);
and UO_2837 (O_2837,N_28953,N_29974);
nand UO_2838 (O_2838,N_29725,N_27100);
or UO_2839 (O_2839,N_27469,N_29017);
xnor UO_2840 (O_2840,N_29671,N_27278);
xor UO_2841 (O_2841,N_29792,N_29820);
and UO_2842 (O_2842,N_29597,N_28277);
nor UO_2843 (O_2843,N_29933,N_29281);
or UO_2844 (O_2844,N_29440,N_28581);
or UO_2845 (O_2845,N_27084,N_28893);
or UO_2846 (O_2846,N_28580,N_29281);
nor UO_2847 (O_2847,N_27676,N_27762);
and UO_2848 (O_2848,N_27117,N_29389);
or UO_2849 (O_2849,N_28364,N_28032);
nand UO_2850 (O_2850,N_29244,N_29522);
or UO_2851 (O_2851,N_29864,N_27621);
xnor UO_2852 (O_2852,N_28422,N_29894);
and UO_2853 (O_2853,N_27617,N_27867);
nor UO_2854 (O_2854,N_27176,N_28613);
or UO_2855 (O_2855,N_28120,N_27423);
or UO_2856 (O_2856,N_28031,N_28879);
or UO_2857 (O_2857,N_29683,N_27339);
xnor UO_2858 (O_2858,N_28823,N_27550);
or UO_2859 (O_2859,N_29768,N_27377);
xor UO_2860 (O_2860,N_29386,N_29600);
xor UO_2861 (O_2861,N_29343,N_27912);
or UO_2862 (O_2862,N_29805,N_27571);
xor UO_2863 (O_2863,N_27009,N_28983);
xor UO_2864 (O_2864,N_28871,N_28734);
xor UO_2865 (O_2865,N_27505,N_29438);
nand UO_2866 (O_2866,N_27142,N_29527);
nand UO_2867 (O_2867,N_27871,N_27751);
nor UO_2868 (O_2868,N_27548,N_29633);
xor UO_2869 (O_2869,N_28645,N_28695);
nand UO_2870 (O_2870,N_28184,N_28878);
xnor UO_2871 (O_2871,N_27509,N_29457);
xnor UO_2872 (O_2872,N_27757,N_28909);
and UO_2873 (O_2873,N_28530,N_29429);
nor UO_2874 (O_2874,N_27285,N_28873);
nor UO_2875 (O_2875,N_29023,N_27010);
or UO_2876 (O_2876,N_28876,N_28873);
nor UO_2877 (O_2877,N_29883,N_28430);
and UO_2878 (O_2878,N_29885,N_29154);
or UO_2879 (O_2879,N_27500,N_28671);
nor UO_2880 (O_2880,N_27038,N_28222);
nor UO_2881 (O_2881,N_28627,N_27156);
xor UO_2882 (O_2882,N_27817,N_28414);
xor UO_2883 (O_2883,N_27217,N_28339);
and UO_2884 (O_2884,N_28419,N_28578);
and UO_2885 (O_2885,N_28899,N_29934);
xnor UO_2886 (O_2886,N_27199,N_27543);
nand UO_2887 (O_2887,N_27786,N_28542);
nand UO_2888 (O_2888,N_28836,N_29503);
or UO_2889 (O_2889,N_27763,N_29821);
xnor UO_2890 (O_2890,N_28199,N_28880);
and UO_2891 (O_2891,N_29090,N_28487);
and UO_2892 (O_2892,N_29168,N_27960);
xnor UO_2893 (O_2893,N_28125,N_28184);
and UO_2894 (O_2894,N_27746,N_27809);
or UO_2895 (O_2895,N_29282,N_28973);
and UO_2896 (O_2896,N_29425,N_28649);
and UO_2897 (O_2897,N_28193,N_28351);
and UO_2898 (O_2898,N_29964,N_28872);
or UO_2899 (O_2899,N_27141,N_28675);
or UO_2900 (O_2900,N_29335,N_29343);
nor UO_2901 (O_2901,N_28487,N_28618);
and UO_2902 (O_2902,N_29611,N_27027);
nand UO_2903 (O_2903,N_27964,N_27705);
xnor UO_2904 (O_2904,N_29848,N_29230);
and UO_2905 (O_2905,N_28250,N_28984);
and UO_2906 (O_2906,N_28731,N_29694);
nand UO_2907 (O_2907,N_27014,N_27120);
and UO_2908 (O_2908,N_27707,N_27298);
or UO_2909 (O_2909,N_29352,N_27939);
nand UO_2910 (O_2910,N_28250,N_29319);
or UO_2911 (O_2911,N_29248,N_28368);
nand UO_2912 (O_2912,N_27452,N_28882);
xor UO_2913 (O_2913,N_29095,N_29880);
or UO_2914 (O_2914,N_28686,N_29975);
nand UO_2915 (O_2915,N_28715,N_27900);
and UO_2916 (O_2916,N_28292,N_27107);
nand UO_2917 (O_2917,N_28681,N_28095);
nor UO_2918 (O_2918,N_29250,N_29821);
nor UO_2919 (O_2919,N_29275,N_29931);
nor UO_2920 (O_2920,N_27655,N_27046);
nor UO_2921 (O_2921,N_27195,N_28525);
or UO_2922 (O_2922,N_29629,N_27311);
or UO_2923 (O_2923,N_27576,N_27157);
or UO_2924 (O_2924,N_28987,N_28508);
nor UO_2925 (O_2925,N_28498,N_28658);
nand UO_2926 (O_2926,N_27464,N_29500);
nand UO_2927 (O_2927,N_28656,N_27390);
nand UO_2928 (O_2928,N_27201,N_28588);
and UO_2929 (O_2929,N_27131,N_29326);
or UO_2930 (O_2930,N_27838,N_27286);
or UO_2931 (O_2931,N_28628,N_29419);
or UO_2932 (O_2932,N_29984,N_28498);
and UO_2933 (O_2933,N_29172,N_27418);
nand UO_2934 (O_2934,N_27871,N_27864);
nand UO_2935 (O_2935,N_28493,N_28532);
and UO_2936 (O_2936,N_29069,N_27993);
or UO_2937 (O_2937,N_29953,N_27387);
or UO_2938 (O_2938,N_28294,N_28971);
xor UO_2939 (O_2939,N_29541,N_27948);
and UO_2940 (O_2940,N_27870,N_29449);
and UO_2941 (O_2941,N_29001,N_29947);
nor UO_2942 (O_2942,N_27406,N_27254);
nor UO_2943 (O_2943,N_27701,N_27591);
xnor UO_2944 (O_2944,N_27555,N_27955);
nand UO_2945 (O_2945,N_29254,N_28668);
xnor UO_2946 (O_2946,N_29102,N_27172);
nand UO_2947 (O_2947,N_27101,N_29474);
nand UO_2948 (O_2948,N_28254,N_27684);
xor UO_2949 (O_2949,N_27323,N_27521);
nor UO_2950 (O_2950,N_27944,N_29645);
nor UO_2951 (O_2951,N_29673,N_28065);
xor UO_2952 (O_2952,N_28665,N_27262);
nand UO_2953 (O_2953,N_27748,N_28036);
nand UO_2954 (O_2954,N_29698,N_28393);
and UO_2955 (O_2955,N_27266,N_28486);
and UO_2956 (O_2956,N_28101,N_27671);
and UO_2957 (O_2957,N_29700,N_28392);
xor UO_2958 (O_2958,N_28766,N_27092);
or UO_2959 (O_2959,N_28893,N_27122);
xnor UO_2960 (O_2960,N_29033,N_29115);
xnor UO_2961 (O_2961,N_28876,N_28601);
nor UO_2962 (O_2962,N_28074,N_27667);
nand UO_2963 (O_2963,N_27804,N_27741);
nor UO_2964 (O_2964,N_28848,N_27444);
or UO_2965 (O_2965,N_28732,N_28408);
nor UO_2966 (O_2966,N_27269,N_27452);
and UO_2967 (O_2967,N_28428,N_28326);
nor UO_2968 (O_2968,N_29292,N_28267);
nand UO_2969 (O_2969,N_28161,N_29021);
xnor UO_2970 (O_2970,N_28008,N_27363);
or UO_2971 (O_2971,N_28681,N_28078);
nor UO_2972 (O_2972,N_29865,N_29108);
xnor UO_2973 (O_2973,N_27946,N_29661);
nand UO_2974 (O_2974,N_29494,N_28863);
or UO_2975 (O_2975,N_28472,N_29492);
or UO_2976 (O_2976,N_27662,N_28858);
nor UO_2977 (O_2977,N_28016,N_27862);
nor UO_2978 (O_2978,N_29648,N_29517);
nor UO_2979 (O_2979,N_28168,N_28890);
or UO_2980 (O_2980,N_27234,N_28461);
or UO_2981 (O_2981,N_29186,N_27869);
xor UO_2982 (O_2982,N_28483,N_29005);
nor UO_2983 (O_2983,N_27329,N_29663);
nor UO_2984 (O_2984,N_27851,N_27486);
or UO_2985 (O_2985,N_28800,N_27887);
xor UO_2986 (O_2986,N_28179,N_29406);
or UO_2987 (O_2987,N_27018,N_27078);
and UO_2988 (O_2988,N_29899,N_27383);
and UO_2989 (O_2989,N_29331,N_28887);
and UO_2990 (O_2990,N_27947,N_27979);
xor UO_2991 (O_2991,N_27672,N_29888);
xor UO_2992 (O_2992,N_27362,N_27132);
nor UO_2993 (O_2993,N_29243,N_29090);
nand UO_2994 (O_2994,N_29532,N_28395);
nand UO_2995 (O_2995,N_29031,N_27432);
nand UO_2996 (O_2996,N_29404,N_28686);
xor UO_2997 (O_2997,N_28804,N_29301);
or UO_2998 (O_2998,N_29880,N_28104);
nor UO_2999 (O_2999,N_28678,N_29346);
or UO_3000 (O_3000,N_28051,N_27081);
nor UO_3001 (O_3001,N_29551,N_27292);
nor UO_3002 (O_3002,N_29576,N_28024);
nor UO_3003 (O_3003,N_29574,N_29247);
or UO_3004 (O_3004,N_29056,N_29919);
or UO_3005 (O_3005,N_27378,N_28346);
nor UO_3006 (O_3006,N_29616,N_28992);
nor UO_3007 (O_3007,N_27846,N_28789);
nor UO_3008 (O_3008,N_27810,N_28794);
nand UO_3009 (O_3009,N_29937,N_27346);
xnor UO_3010 (O_3010,N_27859,N_29238);
xor UO_3011 (O_3011,N_27717,N_28782);
and UO_3012 (O_3012,N_27088,N_27347);
and UO_3013 (O_3013,N_28808,N_28995);
nand UO_3014 (O_3014,N_28842,N_28438);
nand UO_3015 (O_3015,N_27605,N_27483);
xnor UO_3016 (O_3016,N_27042,N_27937);
or UO_3017 (O_3017,N_29568,N_28474);
nand UO_3018 (O_3018,N_29898,N_29195);
and UO_3019 (O_3019,N_28447,N_27052);
nand UO_3020 (O_3020,N_29174,N_27037);
or UO_3021 (O_3021,N_27072,N_27183);
nor UO_3022 (O_3022,N_27832,N_29958);
or UO_3023 (O_3023,N_27197,N_27575);
nand UO_3024 (O_3024,N_27949,N_27526);
nand UO_3025 (O_3025,N_27008,N_28025);
xor UO_3026 (O_3026,N_27123,N_27951);
and UO_3027 (O_3027,N_28611,N_28785);
and UO_3028 (O_3028,N_28987,N_27838);
nand UO_3029 (O_3029,N_29320,N_28354);
or UO_3030 (O_3030,N_28289,N_29518);
xor UO_3031 (O_3031,N_27895,N_28462);
or UO_3032 (O_3032,N_27620,N_28518);
or UO_3033 (O_3033,N_28027,N_27110);
nand UO_3034 (O_3034,N_29794,N_27447);
nand UO_3035 (O_3035,N_28190,N_29332);
nand UO_3036 (O_3036,N_27831,N_27287);
or UO_3037 (O_3037,N_28770,N_29742);
nand UO_3038 (O_3038,N_29100,N_27294);
xnor UO_3039 (O_3039,N_29204,N_28329);
nor UO_3040 (O_3040,N_27285,N_28696);
or UO_3041 (O_3041,N_29609,N_28312);
nor UO_3042 (O_3042,N_27239,N_27768);
nor UO_3043 (O_3043,N_27793,N_29070);
nor UO_3044 (O_3044,N_27040,N_28552);
nand UO_3045 (O_3045,N_29220,N_28233);
and UO_3046 (O_3046,N_29960,N_28109);
nor UO_3047 (O_3047,N_28928,N_27697);
and UO_3048 (O_3048,N_29589,N_28590);
nor UO_3049 (O_3049,N_28280,N_28349);
and UO_3050 (O_3050,N_27496,N_27167);
or UO_3051 (O_3051,N_28176,N_27938);
xnor UO_3052 (O_3052,N_28600,N_27065);
nor UO_3053 (O_3053,N_29589,N_27647);
xnor UO_3054 (O_3054,N_28733,N_28414);
nor UO_3055 (O_3055,N_28486,N_29093);
nand UO_3056 (O_3056,N_28716,N_28072);
nand UO_3057 (O_3057,N_28878,N_27453);
nand UO_3058 (O_3058,N_28572,N_28774);
nor UO_3059 (O_3059,N_27055,N_27858);
nand UO_3060 (O_3060,N_27785,N_29069);
or UO_3061 (O_3061,N_28356,N_27527);
xnor UO_3062 (O_3062,N_29732,N_29527);
and UO_3063 (O_3063,N_27103,N_27445);
or UO_3064 (O_3064,N_29415,N_29815);
nor UO_3065 (O_3065,N_28175,N_27128);
or UO_3066 (O_3066,N_27585,N_28015);
nand UO_3067 (O_3067,N_29616,N_27064);
nor UO_3068 (O_3068,N_27900,N_28319);
nor UO_3069 (O_3069,N_28264,N_27729);
xnor UO_3070 (O_3070,N_28621,N_27795);
or UO_3071 (O_3071,N_29032,N_27357);
nor UO_3072 (O_3072,N_27285,N_27895);
xor UO_3073 (O_3073,N_28662,N_29399);
or UO_3074 (O_3074,N_28786,N_29375);
nor UO_3075 (O_3075,N_28917,N_29667);
xor UO_3076 (O_3076,N_27749,N_27235);
xor UO_3077 (O_3077,N_28665,N_29082);
and UO_3078 (O_3078,N_29691,N_29622);
nor UO_3079 (O_3079,N_27057,N_28595);
nor UO_3080 (O_3080,N_28514,N_27704);
and UO_3081 (O_3081,N_29086,N_27337);
xnor UO_3082 (O_3082,N_29763,N_29432);
or UO_3083 (O_3083,N_28915,N_28104);
nand UO_3084 (O_3084,N_29859,N_28265);
nand UO_3085 (O_3085,N_28593,N_28476);
or UO_3086 (O_3086,N_29529,N_28214);
nand UO_3087 (O_3087,N_28845,N_28563);
and UO_3088 (O_3088,N_29102,N_27442);
xnor UO_3089 (O_3089,N_27808,N_29189);
xnor UO_3090 (O_3090,N_27904,N_28373);
nor UO_3091 (O_3091,N_29788,N_29401);
or UO_3092 (O_3092,N_29404,N_28886);
and UO_3093 (O_3093,N_29714,N_27892);
nor UO_3094 (O_3094,N_27875,N_28274);
or UO_3095 (O_3095,N_29817,N_29455);
and UO_3096 (O_3096,N_27096,N_29904);
or UO_3097 (O_3097,N_27414,N_27693);
or UO_3098 (O_3098,N_27391,N_27861);
or UO_3099 (O_3099,N_29345,N_29548);
nor UO_3100 (O_3100,N_28072,N_29668);
or UO_3101 (O_3101,N_29413,N_29653);
and UO_3102 (O_3102,N_28074,N_29148);
nor UO_3103 (O_3103,N_29833,N_27068);
xor UO_3104 (O_3104,N_29163,N_28743);
xor UO_3105 (O_3105,N_29842,N_29549);
xor UO_3106 (O_3106,N_27973,N_29087);
nand UO_3107 (O_3107,N_29566,N_28556);
and UO_3108 (O_3108,N_29130,N_28528);
xnor UO_3109 (O_3109,N_28131,N_29190);
and UO_3110 (O_3110,N_29292,N_29947);
xor UO_3111 (O_3111,N_27352,N_29090);
and UO_3112 (O_3112,N_29801,N_28030);
and UO_3113 (O_3113,N_28733,N_28428);
xnor UO_3114 (O_3114,N_28785,N_28557);
xor UO_3115 (O_3115,N_29784,N_29348);
nor UO_3116 (O_3116,N_27106,N_28602);
nor UO_3117 (O_3117,N_29833,N_28970);
nand UO_3118 (O_3118,N_27458,N_29957);
and UO_3119 (O_3119,N_27293,N_29596);
or UO_3120 (O_3120,N_28800,N_29821);
or UO_3121 (O_3121,N_27897,N_29341);
nor UO_3122 (O_3122,N_28246,N_29489);
nand UO_3123 (O_3123,N_29574,N_27155);
and UO_3124 (O_3124,N_29867,N_28302);
nand UO_3125 (O_3125,N_28880,N_27124);
or UO_3126 (O_3126,N_28651,N_28120);
nand UO_3127 (O_3127,N_29291,N_29870);
and UO_3128 (O_3128,N_28999,N_29295);
and UO_3129 (O_3129,N_29998,N_27561);
or UO_3130 (O_3130,N_27075,N_29050);
nand UO_3131 (O_3131,N_29552,N_29936);
nand UO_3132 (O_3132,N_29768,N_29621);
xnor UO_3133 (O_3133,N_28231,N_28402);
and UO_3134 (O_3134,N_29619,N_28946);
nand UO_3135 (O_3135,N_28739,N_29456);
nor UO_3136 (O_3136,N_29524,N_28344);
xor UO_3137 (O_3137,N_27120,N_28059);
and UO_3138 (O_3138,N_29501,N_27497);
or UO_3139 (O_3139,N_29095,N_27882);
and UO_3140 (O_3140,N_27500,N_28119);
xnor UO_3141 (O_3141,N_29234,N_28157);
or UO_3142 (O_3142,N_29309,N_28580);
nand UO_3143 (O_3143,N_28660,N_27377);
and UO_3144 (O_3144,N_27430,N_28629);
xor UO_3145 (O_3145,N_29383,N_29841);
nor UO_3146 (O_3146,N_28832,N_28488);
nand UO_3147 (O_3147,N_29081,N_28275);
nor UO_3148 (O_3148,N_28835,N_29527);
or UO_3149 (O_3149,N_28286,N_28467);
and UO_3150 (O_3150,N_29755,N_29766);
and UO_3151 (O_3151,N_28914,N_28799);
nand UO_3152 (O_3152,N_29509,N_28984);
or UO_3153 (O_3153,N_29485,N_27996);
xor UO_3154 (O_3154,N_28280,N_28037);
or UO_3155 (O_3155,N_29372,N_29604);
xnor UO_3156 (O_3156,N_28467,N_29869);
nor UO_3157 (O_3157,N_29094,N_28905);
xnor UO_3158 (O_3158,N_28950,N_27400);
nand UO_3159 (O_3159,N_29201,N_29683);
nand UO_3160 (O_3160,N_28009,N_27756);
xnor UO_3161 (O_3161,N_28061,N_27468);
nand UO_3162 (O_3162,N_28674,N_27291);
and UO_3163 (O_3163,N_27135,N_29147);
and UO_3164 (O_3164,N_29841,N_27209);
xor UO_3165 (O_3165,N_28790,N_29310);
nand UO_3166 (O_3166,N_27250,N_28084);
or UO_3167 (O_3167,N_28773,N_29032);
nand UO_3168 (O_3168,N_28875,N_27990);
nand UO_3169 (O_3169,N_29876,N_29260);
xnor UO_3170 (O_3170,N_29282,N_29221);
or UO_3171 (O_3171,N_29672,N_29863);
or UO_3172 (O_3172,N_28772,N_29448);
xor UO_3173 (O_3173,N_28296,N_28577);
nand UO_3174 (O_3174,N_28567,N_27707);
nor UO_3175 (O_3175,N_27871,N_27888);
or UO_3176 (O_3176,N_29009,N_28712);
nor UO_3177 (O_3177,N_28843,N_27156);
xnor UO_3178 (O_3178,N_27934,N_27974);
nor UO_3179 (O_3179,N_28377,N_28865);
nor UO_3180 (O_3180,N_28180,N_28317);
nor UO_3181 (O_3181,N_28048,N_28959);
nand UO_3182 (O_3182,N_27293,N_29418);
or UO_3183 (O_3183,N_28788,N_28690);
or UO_3184 (O_3184,N_29043,N_28984);
or UO_3185 (O_3185,N_27571,N_29792);
nor UO_3186 (O_3186,N_28497,N_29986);
nand UO_3187 (O_3187,N_29226,N_29965);
nor UO_3188 (O_3188,N_27270,N_27783);
nand UO_3189 (O_3189,N_27175,N_29654);
or UO_3190 (O_3190,N_29017,N_28777);
and UO_3191 (O_3191,N_28381,N_29818);
nor UO_3192 (O_3192,N_29730,N_27049);
nor UO_3193 (O_3193,N_27534,N_28907);
xor UO_3194 (O_3194,N_27163,N_29788);
and UO_3195 (O_3195,N_29318,N_29446);
nor UO_3196 (O_3196,N_29872,N_27225);
xor UO_3197 (O_3197,N_29658,N_28097);
and UO_3198 (O_3198,N_28158,N_27434);
and UO_3199 (O_3199,N_28415,N_28540);
nand UO_3200 (O_3200,N_27522,N_27649);
nand UO_3201 (O_3201,N_28661,N_29024);
xnor UO_3202 (O_3202,N_27335,N_27394);
and UO_3203 (O_3203,N_27320,N_27856);
and UO_3204 (O_3204,N_27106,N_29675);
or UO_3205 (O_3205,N_27826,N_29550);
or UO_3206 (O_3206,N_29799,N_29268);
nor UO_3207 (O_3207,N_27887,N_29992);
or UO_3208 (O_3208,N_28809,N_29283);
or UO_3209 (O_3209,N_27554,N_28463);
and UO_3210 (O_3210,N_27408,N_27351);
xor UO_3211 (O_3211,N_29100,N_28912);
nor UO_3212 (O_3212,N_28133,N_27365);
nand UO_3213 (O_3213,N_28446,N_28033);
nor UO_3214 (O_3214,N_27817,N_29318);
nor UO_3215 (O_3215,N_27559,N_27767);
nand UO_3216 (O_3216,N_27868,N_28097);
nor UO_3217 (O_3217,N_28934,N_27806);
and UO_3218 (O_3218,N_27699,N_27274);
xor UO_3219 (O_3219,N_27608,N_29514);
xor UO_3220 (O_3220,N_27816,N_29815);
or UO_3221 (O_3221,N_29544,N_29459);
nor UO_3222 (O_3222,N_29947,N_29417);
nor UO_3223 (O_3223,N_28332,N_29462);
or UO_3224 (O_3224,N_28906,N_29479);
xnor UO_3225 (O_3225,N_27865,N_27913);
xnor UO_3226 (O_3226,N_28451,N_28923);
and UO_3227 (O_3227,N_28726,N_27472);
and UO_3228 (O_3228,N_29517,N_27311);
or UO_3229 (O_3229,N_29639,N_27993);
or UO_3230 (O_3230,N_29709,N_29762);
nor UO_3231 (O_3231,N_29634,N_28412);
nand UO_3232 (O_3232,N_27012,N_29660);
xor UO_3233 (O_3233,N_27055,N_29061);
and UO_3234 (O_3234,N_29048,N_29437);
nor UO_3235 (O_3235,N_27730,N_27599);
nand UO_3236 (O_3236,N_29733,N_27604);
and UO_3237 (O_3237,N_27725,N_27547);
nor UO_3238 (O_3238,N_27742,N_27002);
xor UO_3239 (O_3239,N_27381,N_29154);
xor UO_3240 (O_3240,N_27575,N_27825);
and UO_3241 (O_3241,N_29652,N_27771);
nor UO_3242 (O_3242,N_29925,N_28969);
or UO_3243 (O_3243,N_28401,N_27777);
nand UO_3244 (O_3244,N_28414,N_28152);
nand UO_3245 (O_3245,N_29714,N_28912);
or UO_3246 (O_3246,N_29194,N_27645);
xor UO_3247 (O_3247,N_28939,N_29061);
nor UO_3248 (O_3248,N_27074,N_29501);
xnor UO_3249 (O_3249,N_27740,N_27285);
nor UO_3250 (O_3250,N_29997,N_28012);
and UO_3251 (O_3251,N_29314,N_28664);
xor UO_3252 (O_3252,N_28555,N_28870);
nor UO_3253 (O_3253,N_29829,N_28052);
or UO_3254 (O_3254,N_28062,N_27068);
nor UO_3255 (O_3255,N_27925,N_27450);
nand UO_3256 (O_3256,N_27170,N_29299);
nor UO_3257 (O_3257,N_28315,N_28705);
and UO_3258 (O_3258,N_28040,N_28264);
and UO_3259 (O_3259,N_28889,N_29263);
xor UO_3260 (O_3260,N_29879,N_28564);
nor UO_3261 (O_3261,N_27632,N_27451);
nand UO_3262 (O_3262,N_29444,N_27501);
or UO_3263 (O_3263,N_28572,N_28760);
nor UO_3264 (O_3264,N_29999,N_27300);
or UO_3265 (O_3265,N_27585,N_27505);
nor UO_3266 (O_3266,N_29071,N_29902);
and UO_3267 (O_3267,N_28798,N_29277);
xor UO_3268 (O_3268,N_28132,N_28790);
nand UO_3269 (O_3269,N_28949,N_29430);
nor UO_3270 (O_3270,N_29103,N_27934);
nand UO_3271 (O_3271,N_29513,N_27287);
xor UO_3272 (O_3272,N_29373,N_29940);
nand UO_3273 (O_3273,N_28089,N_27942);
nor UO_3274 (O_3274,N_27507,N_29878);
or UO_3275 (O_3275,N_29213,N_29964);
and UO_3276 (O_3276,N_29191,N_27416);
nor UO_3277 (O_3277,N_29443,N_29977);
or UO_3278 (O_3278,N_29789,N_27227);
or UO_3279 (O_3279,N_29235,N_27111);
nand UO_3280 (O_3280,N_27626,N_27029);
or UO_3281 (O_3281,N_27665,N_28774);
or UO_3282 (O_3282,N_28233,N_28253);
or UO_3283 (O_3283,N_29724,N_29700);
xnor UO_3284 (O_3284,N_28451,N_29505);
xnor UO_3285 (O_3285,N_29634,N_27006);
or UO_3286 (O_3286,N_29285,N_29179);
nand UO_3287 (O_3287,N_27000,N_29473);
nor UO_3288 (O_3288,N_28707,N_28642);
nand UO_3289 (O_3289,N_28110,N_27064);
xnor UO_3290 (O_3290,N_28754,N_27897);
or UO_3291 (O_3291,N_28230,N_28956);
nand UO_3292 (O_3292,N_28379,N_28954);
and UO_3293 (O_3293,N_27940,N_29393);
nand UO_3294 (O_3294,N_29372,N_27598);
or UO_3295 (O_3295,N_27242,N_29804);
nand UO_3296 (O_3296,N_28580,N_27762);
and UO_3297 (O_3297,N_28963,N_27928);
nand UO_3298 (O_3298,N_27318,N_27325);
nand UO_3299 (O_3299,N_27899,N_29180);
or UO_3300 (O_3300,N_27867,N_28071);
nor UO_3301 (O_3301,N_27357,N_28581);
xor UO_3302 (O_3302,N_29037,N_28643);
nand UO_3303 (O_3303,N_28642,N_28893);
nor UO_3304 (O_3304,N_28929,N_28643);
or UO_3305 (O_3305,N_28994,N_27933);
xor UO_3306 (O_3306,N_27137,N_28190);
nor UO_3307 (O_3307,N_27412,N_29934);
nor UO_3308 (O_3308,N_29100,N_28377);
or UO_3309 (O_3309,N_28221,N_27679);
or UO_3310 (O_3310,N_28644,N_28421);
xor UO_3311 (O_3311,N_29060,N_28240);
and UO_3312 (O_3312,N_29568,N_29589);
xnor UO_3313 (O_3313,N_27570,N_28637);
or UO_3314 (O_3314,N_29027,N_28036);
nor UO_3315 (O_3315,N_29239,N_28054);
or UO_3316 (O_3316,N_29712,N_27264);
and UO_3317 (O_3317,N_27528,N_28235);
xor UO_3318 (O_3318,N_28365,N_27170);
or UO_3319 (O_3319,N_29391,N_28302);
xor UO_3320 (O_3320,N_27345,N_28450);
or UO_3321 (O_3321,N_27512,N_29615);
or UO_3322 (O_3322,N_28858,N_28626);
xor UO_3323 (O_3323,N_27215,N_27889);
and UO_3324 (O_3324,N_27322,N_27523);
xor UO_3325 (O_3325,N_29246,N_27701);
xor UO_3326 (O_3326,N_27936,N_29739);
or UO_3327 (O_3327,N_27714,N_29258);
and UO_3328 (O_3328,N_28889,N_27597);
and UO_3329 (O_3329,N_27879,N_28317);
or UO_3330 (O_3330,N_29428,N_28283);
nand UO_3331 (O_3331,N_28045,N_29921);
xnor UO_3332 (O_3332,N_27751,N_28989);
or UO_3333 (O_3333,N_29036,N_29896);
xor UO_3334 (O_3334,N_29998,N_27624);
or UO_3335 (O_3335,N_29507,N_28639);
and UO_3336 (O_3336,N_27910,N_29910);
nand UO_3337 (O_3337,N_27877,N_27684);
and UO_3338 (O_3338,N_29248,N_29339);
or UO_3339 (O_3339,N_27820,N_27378);
and UO_3340 (O_3340,N_27084,N_27419);
xor UO_3341 (O_3341,N_29045,N_28540);
or UO_3342 (O_3342,N_29769,N_27196);
nor UO_3343 (O_3343,N_29453,N_27786);
and UO_3344 (O_3344,N_29889,N_29178);
and UO_3345 (O_3345,N_27544,N_27434);
xnor UO_3346 (O_3346,N_29615,N_28557);
and UO_3347 (O_3347,N_28804,N_28304);
nand UO_3348 (O_3348,N_28421,N_27383);
and UO_3349 (O_3349,N_28550,N_27125);
nor UO_3350 (O_3350,N_27684,N_29942);
xor UO_3351 (O_3351,N_29773,N_27172);
or UO_3352 (O_3352,N_29567,N_27587);
nor UO_3353 (O_3353,N_28233,N_27616);
or UO_3354 (O_3354,N_28926,N_27190);
xnor UO_3355 (O_3355,N_29166,N_29889);
nand UO_3356 (O_3356,N_29001,N_27116);
or UO_3357 (O_3357,N_27634,N_29179);
or UO_3358 (O_3358,N_28055,N_28629);
nor UO_3359 (O_3359,N_28053,N_29596);
nor UO_3360 (O_3360,N_28437,N_28402);
xor UO_3361 (O_3361,N_27920,N_28711);
and UO_3362 (O_3362,N_28812,N_29545);
xnor UO_3363 (O_3363,N_27795,N_29130);
and UO_3364 (O_3364,N_28065,N_29580);
or UO_3365 (O_3365,N_28888,N_27740);
xor UO_3366 (O_3366,N_27263,N_27411);
nor UO_3367 (O_3367,N_27966,N_29477);
nor UO_3368 (O_3368,N_27674,N_27960);
or UO_3369 (O_3369,N_28957,N_29709);
xor UO_3370 (O_3370,N_29887,N_29637);
nand UO_3371 (O_3371,N_27540,N_27431);
nor UO_3372 (O_3372,N_29586,N_28826);
xnor UO_3373 (O_3373,N_29328,N_27693);
nor UO_3374 (O_3374,N_28560,N_28092);
and UO_3375 (O_3375,N_28965,N_27595);
nor UO_3376 (O_3376,N_29138,N_29427);
xnor UO_3377 (O_3377,N_29133,N_27763);
and UO_3378 (O_3378,N_27773,N_29609);
and UO_3379 (O_3379,N_29362,N_28190);
or UO_3380 (O_3380,N_28757,N_29442);
nor UO_3381 (O_3381,N_29826,N_29288);
nand UO_3382 (O_3382,N_28126,N_28504);
or UO_3383 (O_3383,N_29132,N_29707);
nand UO_3384 (O_3384,N_29368,N_27554);
or UO_3385 (O_3385,N_27430,N_27199);
or UO_3386 (O_3386,N_29298,N_28620);
and UO_3387 (O_3387,N_29179,N_29660);
and UO_3388 (O_3388,N_27210,N_29666);
nand UO_3389 (O_3389,N_28712,N_28423);
xor UO_3390 (O_3390,N_27672,N_28562);
nor UO_3391 (O_3391,N_27477,N_28040);
or UO_3392 (O_3392,N_28936,N_27419);
nand UO_3393 (O_3393,N_28071,N_28113);
xnor UO_3394 (O_3394,N_27787,N_27813);
and UO_3395 (O_3395,N_27399,N_28994);
nor UO_3396 (O_3396,N_29504,N_29618);
or UO_3397 (O_3397,N_27261,N_29756);
xnor UO_3398 (O_3398,N_27500,N_28884);
or UO_3399 (O_3399,N_28579,N_29166);
xor UO_3400 (O_3400,N_29790,N_27010);
nand UO_3401 (O_3401,N_27902,N_27346);
or UO_3402 (O_3402,N_29392,N_27770);
nand UO_3403 (O_3403,N_28092,N_29450);
and UO_3404 (O_3404,N_27836,N_29423);
nor UO_3405 (O_3405,N_27193,N_28479);
xor UO_3406 (O_3406,N_28128,N_28726);
and UO_3407 (O_3407,N_29274,N_29130);
nand UO_3408 (O_3408,N_27569,N_27329);
and UO_3409 (O_3409,N_29102,N_27296);
xnor UO_3410 (O_3410,N_29189,N_28424);
and UO_3411 (O_3411,N_29843,N_29473);
xor UO_3412 (O_3412,N_27389,N_28504);
nand UO_3413 (O_3413,N_29497,N_29838);
nand UO_3414 (O_3414,N_28055,N_29352);
and UO_3415 (O_3415,N_28019,N_28002);
nor UO_3416 (O_3416,N_27352,N_29352);
or UO_3417 (O_3417,N_27880,N_27084);
xnor UO_3418 (O_3418,N_27844,N_29349);
and UO_3419 (O_3419,N_27373,N_28150);
nand UO_3420 (O_3420,N_28000,N_28700);
nor UO_3421 (O_3421,N_27620,N_29179);
xor UO_3422 (O_3422,N_28222,N_27929);
nor UO_3423 (O_3423,N_27478,N_28159);
and UO_3424 (O_3424,N_29647,N_28060);
or UO_3425 (O_3425,N_27637,N_27383);
nor UO_3426 (O_3426,N_28610,N_29126);
nand UO_3427 (O_3427,N_27066,N_29511);
or UO_3428 (O_3428,N_27868,N_29222);
nand UO_3429 (O_3429,N_27509,N_28550);
nor UO_3430 (O_3430,N_27845,N_29936);
or UO_3431 (O_3431,N_27950,N_28837);
nor UO_3432 (O_3432,N_28357,N_29203);
and UO_3433 (O_3433,N_29742,N_29840);
nor UO_3434 (O_3434,N_29240,N_28706);
nand UO_3435 (O_3435,N_27397,N_27858);
or UO_3436 (O_3436,N_29315,N_29388);
xor UO_3437 (O_3437,N_28690,N_27102);
and UO_3438 (O_3438,N_29575,N_28599);
or UO_3439 (O_3439,N_27948,N_29512);
nor UO_3440 (O_3440,N_28217,N_27876);
nand UO_3441 (O_3441,N_29389,N_29830);
nand UO_3442 (O_3442,N_27108,N_28913);
nor UO_3443 (O_3443,N_27136,N_27559);
nor UO_3444 (O_3444,N_29176,N_28079);
nor UO_3445 (O_3445,N_28456,N_27132);
and UO_3446 (O_3446,N_29340,N_28730);
or UO_3447 (O_3447,N_29598,N_29832);
and UO_3448 (O_3448,N_28824,N_29586);
xnor UO_3449 (O_3449,N_29954,N_27474);
or UO_3450 (O_3450,N_27400,N_28285);
or UO_3451 (O_3451,N_29105,N_27361);
and UO_3452 (O_3452,N_28527,N_27893);
or UO_3453 (O_3453,N_29004,N_29109);
and UO_3454 (O_3454,N_28992,N_29906);
xnor UO_3455 (O_3455,N_27206,N_28194);
nand UO_3456 (O_3456,N_29652,N_29332);
or UO_3457 (O_3457,N_28656,N_29167);
xnor UO_3458 (O_3458,N_27262,N_29405);
nor UO_3459 (O_3459,N_29967,N_28780);
xnor UO_3460 (O_3460,N_28423,N_28024);
and UO_3461 (O_3461,N_27810,N_29008);
nor UO_3462 (O_3462,N_28019,N_28387);
and UO_3463 (O_3463,N_29587,N_28136);
or UO_3464 (O_3464,N_29418,N_28709);
or UO_3465 (O_3465,N_28087,N_27724);
or UO_3466 (O_3466,N_27884,N_28091);
xor UO_3467 (O_3467,N_27819,N_29914);
or UO_3468 (O_3468,N_29079,N_27856);
xor UO_3469 (O_3469,N_29956,N_28567);
nand UO_3470 (O_3470,N_28094,N_27348);
nand UO_3471 (O_3471,N_27609,N_27387);
or UO_3472 (O_3472,N_27955,N_27447);
nor UO_3473 (O_3473,N_28827,N_28531);
or UO_3474 (O_3474,N_29786,N_29279);
or UO_3475 (O_3475,N_27967,N_28259);
and UO_3476 (O_3476,N_29395,N_27835);
or UO_3477 (O_3477,N_29899,N_29020);
or UO_3478 (O_3478,N_29489,N_27810);
or UO_3479 (O_3479,N_28502,N_27513);
xor UO_3480 (O_3480,N_27585,N_27164);
nand UO_3481 (O_3481,N_27882,N_28632);
nor UO_3482 (O_3482,N_28669,N_28192);
xor UO_3483 (O_3483,N_29405,N_29030);
xnor UO_3484 (O_3484,N_29185,N_28051);
and UO_3485 (O_3485,N_27989,N_27190);
nand UO_3486 (O_3486,N_27461,N_28710);
and UO_3487 (O_3487,N_28721,N_27988);
and UO_3488 (O_3488,N_29708,N_29944);
and UO_3489 (O_3489,N_29779,N_28917);
or UO_3490 (O_3490,N_29304,N_28346);
and UO_3491 (O_3491,N_28905,N_28679);
nand UO_3492 (O_3492,N_29086,N_27845);
nor UO_3493 (O_3493,N_29607,N_29358);
nand UO_3494 (O_3494,N_27180,N_27500);
xnor UO_3495 (O_3495,N_29835,N_28681);
nand UO_3496 (O_3496,N_29004,N_29488);
xor UO_3497 (O_3497,N_29259,N_29535);
or UO_3498 (O_3498,N_29100,N_29671);
nor UO_3499 (O_3499,N_29709,N_28325);
endmodule