module basic_1000_10000_1500_20_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_868,In_761);
nor U1 (N_1,In_720,In_407);
nor U2 (N_2,In_713,In_65);
and U3 (N_3,In_875,In_665);
and U4 (N_4,In_397,In_624);
or U5 (N_5,In_616,In_18);
and U6 (N_6,In_648,In_615);
nand U7 (N_7,In_306,In_183);
nand U8 (N_8,In_205,In_423);
nand U9 (N_9,In_735,In_412);
or U10 (N_10,In_509,In_745);
nand U11 (N_11,In_706,In_20);
nand U12 (N_12,In_179,In_145);
and U13 (N_13,In_526,In_627);
nor U14 (N_14,In_344,In_670);
xor U15 (N_15,In_845,In_703);
nand U16 (N_16,In_912,In_592);
or U17 (N_17,In_81,In_346);
nor U18 (N_18,In_569,In_501);
and U19 (N_19,In_52,In_667);
nand U20 (N_20,In_785,In_202);
or U21 (N_21,In_764,In_176);
nand U22 (N_22,In_589,In_927);
nand U23 (N_23,In_477,In_654);
xor U24 (N_24,In_203,In_106);
nand U25 (N_25,In_283,In_859);
or U26 (N_26,In_227,In_951);
or U27 (N_27,In_623,In_947);
or U28 (N_28,In_548,In_19);
nor U29 (N_29,In_312,In_528);
nand U30 (N_30,In_893,In_175);
or U31 (N_31,In_308,In_460);
nand U32 (N_32,In_197,In_401);
or U33 (N_33,In_562,In_843);
nor U34 (N_34,In_290,In_726);
nand U35 (N_35,In_151,In_545);
and U36 (N_36,In_574,In_37);
and U37 (N_37,In_585,In_730);
nand U38 (N_38,In_458,In_400);
and U39 (N_39,In_136,In_661);
nand U40 (N_40,In_11,In_842);
or U41 (N_41,In_653,In_551);
and U42 (N_42,In_534,In_473);
nor U43 (N_43,In_610,In_274);
nand U44 (N_44,In_536,In_650);
and U45 (N_45,In_13,In_882);
xor U46 (N_46,In_802,In_728);
or U47 (N_47,In_261,In_838);
nor U48 (N_48,In_755,In_158);
and U49 (N_49,In_216,In_945);
nand U50 (N_50,In_191,In_823);
and U51 (N_51,In_722,In_935);
nor U52 (N_52,In_385,In_455);
or U53 (N_53,In_603,In_443);
or U54 (N_54,In_502,In_770);
nor U55 (N_55,In_300,In_877);
or U56 (N_56,In_192,In_212);
or U57 (N_57,In_114,In_673);
or U58 (N_58,In_375,In_517);
and U59 (N_59,In_839,In_527);
and U60 (N_60,In_532,In_871);
xor U61 (N_61,In_257,In_841);
and U62 (N_62,In_479,In_824);
nor U63 (N_63,In_121,In_91);
nand U64 (N_64,In_892,In_101);
nor U65 (N_65,In_90,In_22);
nand U66 (N_66,In_729,In_278);
or U67 (N_67,In_644,In_478);
nor U68 (N_68,In_487,In_629);
and U69 (N_69,In_438,In_668);
nor U70 (N_70,In_325,In_93);
or U71 (N_71,In_831,In_821);
nor U72 (N_72,In_529,In_565);
nand U73 (N_73,In_320,In_125);
or U74 (N_74,In_324,In_889);
and U75 (N_75,In_789,In_386);
nor U76 (N_76,In_638,In_17);
or U77 (N_77,In_832,In_498);
xnor U78 (N_78,In_905,In_470);
nand U79 (N_79,In_659,In_351);
nor U80 (N_80,In_568,In_512);
xor U81 (N_81,In_966,In_816);
xnor U82 (N_82,In_981,In_97);
or U83 (N_83,In_712,In_960);
and U84 (N_84,In_830,In_639);
xor U85 (N_85,In_812,In_642);
xnor U86 (N_86,In_88,In_856);
and U87 (N_87,In_747,In_281);
xnor U88 (N_88,In_983,In_384);
and U89 (N_89,In_356,In_500);
xor U90 (N_90,In_339,In_316);
and U91 (N_91,In_511,In_263);
nor U92 (N_92,In_128,In_298);
nand U93 (N_93,In_404,In_335);
or U94 (N_94,In_361,In_465);
or U95 (N_95,In_62,In_881);
nand U96 (N_96,In_430,In_996);
and U97 (N_97,In_612,In_457);
and U98 (N_98,In_631,In_736);
nand U99 (N_99,In_973,In_759);
or U100 (N_100,In_277,In_583);
xor U101 (N_101,In_119,In_146);
or U102 (N_102,In_558,In_166);
nand U103 (N_103,In_944,In_280);
xor U104 (N_104,In_756,In_535);
or U105 (N_105,In_15,In_766);
nand U106 (N_106,In_855,In_906);
nor U107 (N_107,In_452,In_161);
xor U108 (N_108,In_488,In_7);
or U109 (N_109,In_476,In_835);
nand U110 (N_110,In_322,In_311);
and U111 (N_111,In_826,In_507);
or U112 (N_112,In_890,In_991);
nor U113 (N_113,In_422,In_787);
xnor U114 (N_114,In_597,In_79);
or U115 (N_115,In_964,In_228);
nand U116 (N_116,In_891,In_1);
xnor U117 (N_117,In_825,In_464);
nand U118 (N_118,In_916,In_71);
or U119 (N_119,In_879,In_520);
and U120 (N_120,In_207,In_348);
nand U121 (N_121,In_750,In_997);
and U122 (N_122,In_137,In_472);
nor U123 (N_123,In_662,In_995);
nor U124 (N_124,In_931,In_525);
or U125 (N_125,In_748,In_87);
nand U126 (N_126,In_604,In_186);
xor U127 (N_127,In_625,In_499);
xor U128 (N_128,In_353,In_505);
nand U129 (N_129,In_854,In_572);
nor U130 (N_130,In_14,In_714);
xnor U131 (N_131,In_840,In_275);
nor U132 (N_132,In_682,In_948);
and U133 (N_133,In_704,In_561);
and U134 (N_134,In_211,In_968);
nor U135 (N_135,In_518,In_67);
and U136 (N_136,In_230,In_664);
or U137 (N_137,In_705,In_560);
nand U138 (N_138,In_873,In_396);
nand U139 (N_139,In_439,In_799);
nor U140 (N_140,In_446,In_986);
nand U141 (N_141,In_245,In_220);
or U142 (N_142,In_533,In_129);
or U143 (N_143,In_888,In_683);
xor U144 (N_144,In_946,In_955);
nor U145 (N_145,In_285,In_672);
nor U146 (N_146,In_926,In_651);
or U147 (N_147,In_780,In_21);
or U148 (N_148,In_159,In_177);
xnor U149 (N_149,In_406,In_915);
nor U150 (N_150,In_174,In_163);
or U151 (N_151,In_656,In_433);
and U152 (N_152,In_982,In_643);
nand U153 (N_153,In_420,In_934);
and U154 (N_154,In_149,In_963);
nor U155 (N_155,In_115,In_236);
or U156 (N_156,In_221,In_550);
or U157 (N_157,In_646,In_626);
nor U158 (N_158,In_850,In_640);
nor U159 (N_159,In_35,In_696);
nand U160 (N_160,In_33,In_674);
nor U161 (N_161,In_874,In_413);
or U162 (N_162,In_314,In_655);
nor U163 (N_163,In_942,In_330);
nor U164 (N_164,In_414,In_504);
and U165 (N_165,In_0,In_147);
and U166 (N_166,In_742,In_408);
and U167 (N_167,In_741,In_29);
nor U168 (N_168,In_961,In_164);
xnor U169 (N_169,In_169,In_899);
xor U170 (N_170,In_43,In_798);
nand U171 (N_171,In_480,In_497);
nor U172 (N_172,In_819,In_27);
and U173 (N_173,In_448,In_171);
xor U174 (N_174,In_48,In_666);
or U175 (N_175,In_219,In_657);
or U176 (N_176,In_194,In_286);
nand U177 (N_177,In_304,In_295);
and U178 (N_178,In_943,In_249);
and U179 (N_179,In_204,In_54);
nand U180 (N_180,In_309,In_813);
nand U181 (N_181,In_381,In_415);
nand U182 (N_182,In_250,In_669);
and U183 (N_183,In_323,In_617);
nand U184 (N_184,In_940,In_690);
nor U185 (N_185,In_282,In_393);
and U186 (N_186,In_793,In_224);
xnor U187 (N_187,In_738,In_395);
nor U188 (N_188,In_897,In_849);
nand U189 (N_189,In_894,In_442);
or U190 (N_190,In_768,In_707);
nor U191 (N_191,In_40,In_630);
and U192 (N_192,In_301,In_969);
and U193 (N_193,In_709,In_26);
nor U194 (N_194,In_794,In_688);
or U195 (N_195,In_242,In_89);
nand U196 (N_196,In_447,In_291);
nor U197 (N_197,In_368,In_345);
and U198 (N_198,In_698,In_701);
nor U199 (N_199,In_758,In_797);
and U200 (N_200,In_977,In_483);
nor U201 (N_201,In_811,In_59);
and U202 (N_202,In_270,In_784);
nand U203 (N_203,In_687,In_924);
nor U204 (N_204,In_240,In_421);
or U205 (N_205,In_697,In_681);
or U206 (N_206,In_123,In_699);
or U207 (N_207,In_466,In_660);
nand U208 (N_208,In_181,In_974);
nand U209 (N_209,In_402,In_84);
nand U210 (N_210,In_72,In_857);
nor U211 (N_211,In_636,In_445);
nor U212 (N_212,In_392,In_744);
and U213 (N_213,In_201,In_844);
and U214 (N_214,In_391,In_142);
and U215 (N_215,In_573,In_998);
and U216 (N_216,In_922,In_544);
nor U217 (N_217,In_635,In_833);
xnor U218 (N_218,In_156,In_69);
or U219 (N_219,In_941,In_410);
xor U220 (N_220,In_4,In_96);
and U221 (N_221,In_462,In_32);
and U222 (N_222,In_206,In_241);
nand U223 (N_223,In_820,In_321);
or U224 (N_224,In_564,In_231);
and U225 (N_225,In_73,In_437);
nand U226 (N_226,In_634,In_185);
nor U227 (N_227,In_853,In_307);
or U228 (N_228,In_710,In_343);
and U229 (N_229,In_394,In_131);
nor U230 (N_230,In_78,In_364);
nand U231 (N_231,In_515,In_866);
nand U232 (N_232,In_992,In_288);
and U233 (N_233,In_967,In_782);
nand U234 (N_234,In_456,In_210);
or U235 (N_235,In_869,In_349);
nor U236 (N_236,In_148,In_590);
nand U237 (N_237,In_426,In_723);
nor U238 (N_238,In_47,In_378);
nand U239 (N_239,In_896,In_676);
nand U240 (N_240,In_70,In_383);
nor U241 (N_241,In_104,In_938);
and U242 (N_242,In_804,In_584);
or U243 (N_243,In_399,In_276);
or U244 (N_244,In_6,In_555);
or U245 (N_245,In_130,In_632);
and U246 (N_246,In_746,In_503);
nand U247 (N_247,In_792,In_195);
and U248 (N_248,In_182,In_302);
nor U249 (N_249,In_918,In_593);
or U250 (N_250,In_783,In_108);
and U251 (N_251,In_379,In_39);
nor U252 (N_252,In_222,In_523);
nor U253 (N_253,In_340,In_425);
nand U254 (N_254,In_920,In_834);
and U255 (N_255,In_154,In_494);
nor U256 (N_256,In_461,In_82);
xnor U257 (N_257,In_75,In_567);
nand U258 (N_258,In_299,In_692);
nand U259 (N_259,In_482,In_815);
and U260 (N_260,In_170,In_923);
nor U261 (N_261,In_61,In_605);
and U262 (N_262,In_189,In_8);
xor U263 (N_263,In_398,In_700);
nand U264 (N_264,In_214,In_980);
nand U265 (N_265,In_264,In_380);
and U266 (N_266,In_272,In_847);
nor U267 (N_267,In_64,In_571);
nand U268 (N_268,In_577,In_901);
or U269 (N_269,In_602,In_733);
xnor U270 (N_270,In_454,In_489);
or U271 (N_271,In_435,In_342);
xnor U272 (N_272,In_2,In_484);
and U273 (N_273,In_576,In_658);
nand U274 (N_274,In_885,In_779);
or U275 (N_275,In_196,In_256);
and U276 (N_276,In_972,In_260);
and U277 (N_277,In_107,In_124);
nand U278 (N_278,In_332,In_519);
nor U279 (N_279,In_814,In_416);
nand U280 (N_280,In_717,In_836);
nor U281 (N_281,In_248,In_424);
nand U282 (N_282,In_749,In_810);
nand U283 (N_283,In_950,In_118);
and U284 (N_284,In_773,In_94);
xor U285 (N_285,In_979,In_315);
xnor U286 (N_286,In_587,In_247);
xnor U287 (N_287,In_258,In_864);
or U288 (N_288,In_215,In_600);
and U289 (N_289,In_134,In_575);
nor U290 (N_290,In_828,In_771);
and U291 (N_291,In_769,In_872);
nand U292 (N_292,In_50,In_900);
nor U293 (N_293,In_530,In_903);
and U294 (N_294,In_796,In_588);
and U295 (N_295,In_287,In_296);
and U296 (N_296,In_144,In_234);
xor U297 (N_297,In_988,In_428);
nor U298 (N_298,In_790,In_895);
xor U299 (N_299,In_334,In_508);
nor U300 (N_300,In_77,In_370);
nor U301 (N_301,In_141,In_579);
nand U302 (N_302,In_607,In_318);
or U303 (N_303,In_693,In_357);
and U304 (N_304,In_139,In_837);
or U305 (N_305,In_753,In_727);
nand U306 (N_306,In_358,In_41);
xor U307 (N_307,In_559,In_510);
nand U308 (N_308,In_239,In_266);
and U309 (N_309,In_861,In_450);
and U310 (N_310,In_279,In_209);
or U311 (N_311,In_172,In_788);
and U312 (N_312,In_369,In_902);
nor U313 (N_313,In_157,In_193);
and U314 (N_314,In_493,In_12);
nor U315 (N_315,In_467,In_725);
or U316 (N_316,In_611,In_880);
or U317 (N_317,In_786,In_829);
and U318 (N_318,In_313,In_990);
nor U319 (N_319,In_858,In_552);
and U320 (N_320,In_341,In_907);
or U321 (N_321,In_362,In_613);
or U322 (N_322,In_127,In_959);
and U323 (N_323,In_965,In_262);
or U324 (N_324,In_9,In_677);
xnor U325 (N_325,In_791,In_485);
nand U326 (N_326,In_367,In_949);
nand U327 (N_327,In_539,In_373);
nor U328 (N_328,In_16,In_122);
or U329 (N_329,In_958,In_580);
or U330 (N_330,In_956,In_419);
and U331 (N_331,In_776,In_388);
or U332 (N_332,In_876,In_581);
nand U333 (N_333,In_486,In_925);
or U334 (N_334,In_138,In_178);
nor U335 (N_335,In_652,In_740);
nor U336 (N_336,In_628,In_360);
nor U337 (N_337,In_173,In_721);
nand U338 (N_338,In_549,In_521);
xor U339 (N_339,In_524,In_95);
and U340 (N_340,In_781,In_724);
nor U341 (N_341,In_463,In_795);
nand U342 (N_342,In_80,In_808);
nor U343 (N_343,In_333,In_354);
and U344 (N_344,In_711,In_116);
xnor U345 (N_345,In_737,In_431);
nand U346 (N_346,In_365,In_265);
nand U347 (N_347,In_451,In_53);
or U348 (N_348,In_105,In_716);
nor U349 (N_349,In_774,In_363);
nand U350 (N_350,In_932,In_684);
nor U351 (N_351,In_994,In_474);
nor U352 (N_352,In_675,In_98);
nor U353 (N_353,In_468,In_514);
or U354 (N_354,In_165,In_42);
and U355 (N_355,In_685,In_237);
nor U356 (N_356,In_952,In_188);
or U357 (N_357,In_387,In_731);
and U358 (N_358,In_911,In_689);
nand U359 (N_359,In_347,In_389);
nor U360 (N_360,In_595,In_34);
nor U361 (N_361,In_51,In_453);
nand U362 (N_362,In_976,In_133);
nand U363 (N_363,In_200,In_752);
and U364 (N_364,In_112,In_310);
nor U365 (N_365,In_691,In_110);
nand U366 (N_366,In_546,In_678);
and U367 (N_367,In_235,In_49);
or U368 (N_368,In_327,In_143);
or U369 (N_369,In_3,In_765);
xnor U370 (N_370,In_23,In_594);
and U371 (N_371,In_60,In_553);
xor U372 (N_372,In_975,In_338);
or U373 (N_373,In_762,In_68);
nand U374 (N_374,In_556,In_601);
nand U375 (N_375,In_801,In_718);
and U376 (N_376,In_516,In_686);
nor U377 (N_377,In_582,In_459);
or U378 (N_378,In_427,In_243);
and U379 (N_379,In_74,In_86);
and U380 (N_380,In_140,In_492);
and U381 (N_381,In_83,In_754);
and U382 (N_382,In_294,In_971);
and U383 (N_383,In_827,In_647);
or U384 (N_384,In_403,In_641);
nand U385 (N_385,In_229,In_253);
nor U386 (N_386,In_168,In_541);
or U387 (N_387,In_329,In_45);
nor U388 (N_388,In_807,In_355);
nand U389 (N_389,In_56,In_619);
and U390 (N_390,In_190,In_44);
xor U391 (N_391,In_566,In_28);
nand U392 (N_392,In_25,In_293);
and U393 (N_393,In_198,In_429);
or U394 (N_394,In_244,In_36);
nand U395 (N_395,In_444,In_591);
and U396 (N_396,In_117,In_30);
or U397 (N_397,In_390,In_822);
nor U398 (N_398,In_38,In_702);
nand U399 (N_399,In_962,In_153);
or U400 (N_400,In_852,In_184);
nand U401 (N_401,In_273,In_618);
nor U402 (N_402,In_621,In_411);
nand U403 (N_403,In_109,In_238);
and U404 (N_404,In_268,In_679);
nor U405 (N_405,In_103,In_366);
and U406 (N_406,In_908,In_939);
xor U407 (N_407,In_863,In_805);
or U408 (N_408,In_649,In_531);
or U409 (N_409,In_606,In_24);
nor U410 (N_410,In_132,In_405);
nor U411 (N_411,In_297,In_883);
and U412 (N_412,In_162,In_490);
nand U413 (N_413,In_851,In_155);
and U414 (N_414,In_150,In_371);
and U415 (N_415,In_374,In_862);
nor U416 (N_416,In_85,In_884);
nor U417 (N_417,In_160,In_919);
nand U418 (N_418,In_914,In_817);
xnor U419 (N_419,In_58,In_126);
or U420 (N_420,In_475,In_251);
or U421 (N_421,In_233,In_985);
and U422 (N_422,In_609,In_92);
or U423 (N_423,In_775,In_31);
and U424 (N_424,In_680,In_436);
nor U425 (N_425,In_694,In_933);
nand U426 (N_426,In_496,In_100);
and U427 (N_427,In_246,In_557);
nand U428 (N_428,In_542,In_372);
nand U429 (N_429,In_999,In_989);
nand U430 (N_430,In_865,In_987);
nor U431 (N_431,In_481,In_937);
and U432 (N_432,In_113,In_695);
nand U433 (N_433,In_860,In_586);
nand U434 (N_434,In_441,In_870);
nand U435 (N_435,In_596,In_254);
nor U436 (N_436,In_760,In_887);
or U437 (N_437,In_570,In_910);
nand U438 (N_438,In_953,In_434);
or U439 (N_439,In_538,In_440);
nand U440 (N_440,In_331,In_547);
nor U441 (N_441,In_223,In_622);
nor U442 (N_442,In_317,In_232);
nand U443 (N_443,In_929,In_167);
or U444 (N_444,In_377,In_663);
or U445 (N_445,In_800,In_867);
and U446 (N_446,In_732,In_135);
nand U447 (N_447,In_715,In_671);
xnor U448 (N_448,In_614,In_848);
and U449 (N_449,In_708,In_772);
or U450 (N_450,In_252,In_225);
nor U451 (N_451,In_751,In_55);
and U452 (N_452,In_554,In_289);
nand U453 (N_453,In_350,In_213);
nand U454 (N_454,In_99,In_102);
or U455 (N_455,In_954,In_120);
nand U456 (N_456,In_846,In_767);
nand U457 (N_457,In_936,In_984);
or U458 (N_458,In_226,In_305);
and U459 (N_459,In_199,In_319);
xnor U460 (N_460,In_66,In_763);
nand U461 (N_461,In_208,In_292);
nand U462 (N_462,In_540,In_719);
nand U463 (N_463,In_608,In_777);
nand U464 (N_464,In_495,In_598);
nand U465 (N_465,In_620,In_469);
nand U466 (N_466,In_5,In_111);
nor U467 (N_467,In_382,In_303);
nand U468 (N_468,In_326,In_284);
nand U469 (N_469,In_417,In_46);
nor U470 (N_470,In_970,In_917);
and U471 (N_471,In_957,In_76);
and U472 (N_472,In_337,In_376);
nand U473 (N_473,In_359,In_409);
nand U474 (N_474,In_187,In_757);
or U475 (N_475,In_734,In_449);
or U476 (N_476,In_743,In_637);
and U477 (N_477,In_57,In_898);
or U478 (N_478,In_328,In_10);
nor U479 (N_479,In_904,In_152);
nor U480 (N_480,In_803,In_259);
nand U481 (N_481,In_739,In_336);
nor U482 (N_482,In_217,In_645);
xor U483 (N_483,In_930,In_255);
nor U484 (N_484,In_513,In_352);
and U485 (N_485,In_809,In_886);
and U486 (N_486,In_563,In_471);
or U487 (N_487,In_537,In_269);
nor U488 (N_488,In_778,In_432);
nor U489 (N_489,In_818,In_806);
xnor U490 (N_490,In_578,In_928);
or U491 (N_491,In_63,In_491);
xor U492 (N_492,In_506,In_978);
nor U493 (N_493,In_913,In_418);
and U494 (N_494,In_921,In_633);
nand U495 (N_495,In_878,In_267);
or U496 (N_496,In_522,In_993);
and U497 (N_497,In_271,In_218);
or U498 (N_498,In_599,In_543);
nor U499 (N_499,In_909,In_180);
and U500 (N_500,N_423,N_478);
or U501 (N_501,N_468,N_305);
nor U502 (N_502,N_157,N_449);
nand U503 (N_503,N_160,N_16);
or U504 (N_504,N_336,N_315);
nor U505 (N_505,N_233,N_13);
or U506 (N_506,N_284,N_314);
nor U507 (N_507,N_412,N_117);
and U508 (N_508,N_403,N_129);
or U509 (N_509,N_292,N_354);
and U510 (N_510,N_474,N_248);
xor U511 (N_511,N_279,N_422);
and U512 (N_512,N_113,N_216);
nand U513 (N_513,N_49,N_177);
and U514 (N_514,N_408,N_80);
or U515 (N_515,N_323,N_304);
and U516 (N_516,N_492,N_41);
nand U517 (N_517,N_320,N_379);
and U518 (N_518,N_184,N_458);
nor U519 (N_519,N_392,N_463);
xor U520 (N_520,N_446,N_209);
and U521 (N_521,N_33,N_81);
or U522 (N_522,N_60,N_466);
or U523 (N_523,N_413,N_208);
xor U524 (N_524,N_149,N_175);
or U525 (N_525,N_491,N_411);
xnor U526 (N_526,N_477,N_64);
and U527 (N_527,N_190,N_223);
nand U528 (N_528,N_493,N_438);
nor U529 (N_529,N_356,N_144);
nand U530 (N_530,N_455,N_38);
nand U531 (N_531,N_229,N_419);
and U532 (N_532,N_50,N_476);
nand U533 (N_533,N_258,N_274);
nand U534 (N_534,N_178,N_402);
and U535 (N_535,N_350,N_147);
or U536 (N_536,N_361,N_399);
and U537 (N_537,N_340,N_467);
or U538 (N_538,N_374,N_104);
nand U539 (N_539,N_161,N_246);
nor U540 (N_540,N_83,N_70);
or U541 (N_541,N_73,N_368);
and U542 (N_542,N_202,N_439);
or U543 (N_543,N_205,N_136);
and U544 (N_544,N_69,N_337);
or U545 (N_545,N_7,N_153);
nand U546 (N_546,N_25,N_358);
or U547 (N_547,N_196,N_357);
xor U548 (N_548,N_471,N_486);
nor U549 (N_549,N_297,N_420);
and U550 (N_550,N_164,N_311);
nand U551 (N_551,N_362,N_261);
nor U552 (N_552,N_448,N_231);
nor U553 (N_553,N_172,N_227);
and U554 (N_554,N_300,N_111);
nand U555 (N_555,N_228,N_351);
nor U556 (N_556,N_260,N_85);
or U557 (N_557,N_367,N_391);
and U558 (N_558,N_298,N_319);
or U559 (N_559,N_405,N_398);
nand U560 (N_560,N_397,N_309);
xor U561 (N_561,N_123,N_152);
nand U562 (N_562,N_185,N_285);
or U563 (N_563,N_487,N_109);
and U564 (N_564,N_95,N_203);
nor U565 (N_565,N_499,N_393);
and U566 (N_566,N_410,N_162);
and U567 (N_567,N_414,N_77);
nor U568 (N_568,N_212,N_101);
or U569 (N_569,N_465,N_89);
or U570 (N_570,N_127,N_37);
and U571 (N_571,N_306,N_135);
nor U572 (N_572,N_363,N_90);
nor U573 (N_573,N_473,N_295);
nand U574 (N_574,N_289,N_40);
nand U575 (N_575,N_333,N_121);
and U576 (N_576,N_443,N_469);
or U577 (N_577,N_51,N_247);
or U578 (N_578,N_325,N_384);
or U579 (N_579,N_226,N_28);
nor U580 (N_580,N_23,N_22);
and U581 (N_581,N_61,N_94);
and U582 (N_582,N_74,N_235);
nand U583 (N_583,N_97,N_312);
or U584 (N_584,N_34,N_338);
or U585 (N_585,N_479,N_360);
and U586 (N_586,N_276,N_441);
and U587 (N_587,N_106,N_232);
and U588 (N_588,N_19,N_26);
nand U589 (N_589,N_382,N_220);
nand U590 (N_590,N_464,N_238);
nand U591 (N_591,N_454,N_133);
and U592 (N_592,N_343,N_400);
and U593 (N_593,N_240,N_380);
or U594 (N_594,N_253,N_364);
and U595 (N_595,N_217,N_264);
nand U596 (N_596,N_198,N_98);
nor U597 (N_597,N_425,N_259);
xnor U598 (N_598,N_461,N_294);
nor U599 (N_599,N_495,N_15);
nor U600 (N_600,N_163,N_275);
nand U601 (N_601,N_225,N_291);
nand U602 (N_602,N_79,N_176);
and U603 (N_603,N_436,N_430);
nand U604 (N_604,N_122,N_293);
or U605 (N_605,N_245,N_349);
nand U606 (N_606,N_450,N_283);
nand U607 (N_607,N_145,N_103);
or U608 (N_608,N_317,N_99);
and U609 (N_609,N_58,N_386);
and U610 (N_610,N_407,N_183);
nor U611 (N_611,N_4,N_273);
xor U612 (N_612,N_472,N_262);
xnor U613 (N_613,N_329,N_255);
nor U614 (N_614,N_480,N_36);
nor U615 (N_615,N_130,N_482);
nand U616 (N_616,N_3,N_222);
or U617 (N_617,N_270,N_44);
or U618 (N_618,N_307,N_140);
or U619 (N_619,N_353,N_385);
xor U620 (N_620,N_490,N_375);
nand U621 (N_621,N_236,N_324);
or U622 (N_622,N_148,N_431);
nor U623 (N_623,N_271,N_32);
nand U624 (N_624,N_201,N_53);
nand U625 (N_625,N_366,N_137);
nor U626 (N_626,N_288,N_224);
nor U627 (N_627,N_207,N_125);
nand U628 (N_628,N_251,N_498);
nand U629 (N_629,N_330,N_310);
nor U630 (N_630,N_138,N_378);
nand U631 (N_631,N_266,N_355);
nand U632 (N_632,N_100,N_383);
and U633 (N_633,N_475,N_45);
nor U634 (N_634,N_29,N_387);
nor U635 (N_635,N_359,N_118);
nor U636 (N_636,N_352,N_54);
xnor U637 (N_637,N_20,N_332);
and U638 (N_638,N_277,N_115);
xnor U639 (N_639,N_286,N_17);
and U640 (N_640,N_327,N_415);
or U641 (N_641,N_179,N_56);
nor U642 (N_642,N_457,N_0);
xnor U643 (N_643,N_280,N_93);
nand U644 (N_644,N_9,N_8);
or U645 (N_645,N_460,N_150);
or U646 (N_646,N_5,N_67);
and U647 (N_647,N_341,N_86);
xnor U648 (N_648,N_348,N_142);
nand U649 (N_649,N_421,N_165);
and U650 (N_650,N_126,N_156);
nor U651 (N_651,N_427,N_59);
nor U652 (N_652,N_265,N_344);
nor U653 (N_653,N_401,N_11);
or U654 (N_654,N_120,N_43);
or U655 (N_655,N_47,N_418);
nor U656 (N_656,N_210,N_470);
or U657 (N_657,N_92,N_24);
and U658 (N_658,N_267,N_462);
nand U659 (N_659,N_192,N_167);
and U660 (N_660,N_76,N_447);
nand U661 (N_661,N_437,N_257);
or U662 (N_662,N_417,N_256);
xnor U663 (N_663,N_376,N_114);
and U664 (N_664,N_62,N_128);
and U665 (N_665,N_347,N_365);
or U666 (N_666,N_272,N_42);
nand U667 (N_667,N_200,N_102);
nand U668 (N_668,N_303,N_459);
xor U669 (N_669,N_389,N_174);
nand U670 (N_670,N_373,N_84);
and U671 (N_671,N_134,N_155);
and U672 (N_672,N_52,N_322);
and U673 (N_673,N_146,N_10);
or U674 (N_674,N_132,N_72);
or U675 (N_675,N_452,N_456);
and U676 (N_676,N_445,N_75);
nand U677 (N_677,N_369,N_168);
nand U678 (N_678,N_263,N_57);
or U679 (N_679,N_296,N_377);
and U680 (N_680,N_108,N_416);
nand U681 (N_681,N_234,N_21);
and U682 (N_682,N_440,N_370);
or U683 (N_683,N_318,N_381);
nand U684 (N_684,N_287,N_88);
and U685 (N_685,N_206,N_2);
and U686 (N_686,N_182,N_71);
and U687 (N_687,N_301,N_124);
nor U688 (N_688,N_268,N_131);
nand U689 (N_689,N_313,N_91);
nand U690 (N_690,N_243,N_494);
xnor U691 (N_691,N_12,N_55);
and U692 (N_692,N_335,N_302);
xnor U693 (N_693,N_46,N_171);
and U694 (N_694,N_31,N_143);
and U695 (N_695,N_424,N_194);
nor U696 (N_696,N_199,N_432);
or U697 (N_697,N_316,N_321);
or U698 (N_698,N_434,N_87);
or U699 (N_699,N_189,N_269);
nor U700 (N_700,N_394,N_483);
nand U701 (N_701,N_371,N_435);
nand U702 (N_702,N_6,N_396);
nand U703 (N_703,N_187,N_186);
xor U704 (N_704,N_404,N_308);
nand U705 (N_705,N_488,N_242);
and U706 (N_706,N_105,N_453);
nor U707 (N_707,N_154,N_82);
nand U708 (N_708,N_169,N_345);
and U709 (N_709,N_429,N_489);
nand U710 (N_710,N_299,N_188);
nor U711 (N_711,N_484,N_214);
xor U712 (N_712,N_342,N_249);
and U713 (N_713,N_78,N_1);
xnor U714 (N_714,N_444,N_426);
nor U715 (N_715,N_215,N_372);
or U716 (N_716,N_252,N_442);
or U717 (N_717,N_66,N_406);
nand U718 (N_718,N_290,N_151);
nor U719 (N_719,N_433,N_218);
nor U720 (N_720,N_241,N_139);
nor U721 (N_721,N_219,N_388);
nor U722 (N_722,N_409,N_346);
and U723 (N_723,N_254,N_244);
nand U724 (N_724,N_96,N_497);
nand U725 (N_725,N_428,N_339);
and U726 (N_726,N_110,N_221);
xnor U727 (N_727,N_166,N_112);
or U728 (N_728,N_68,N_119);
nand U729 (N_729,N_281,N_278);
xnor U730 (N_730,N_18,N_230);
and U731 (N_731,N_197,N_213);
nor U732 (N_732,N_237,N_282);
or U733 (N_733,N_395,N_239);
or U734 (N_734,N_141,N_331);
nand U735 (N_735,N_65,N_211);
nor U736 (N_736,N_250,N_158);
or U737 (N_737,N_173,N_107);
or U738 (N_738,N_170,N_451);
and U739 (N_739,N_496,N_48);
or U740 (N_740,N_30,N_334);
nand U741 (N_741,N_195,N_481);
nand U742 (N_742,N_390,N_180);
and U743 (N_743,N_181,N_116);
nand U744 (N_744,N_204,N_485);
and U745 (N_745,N_191,N_193);
nor U746 (N_746,N_159,N_14);
nand U747 (N_747,N_63,N_328);
or U748 (N_748,N_35,N_39);
or U749 (N_749,N_27,N_326);
nand U750 (N_750,N_93,N_333);
nor U751 (N_751,N_321,N_453);
nor U752 (N_752,N_374,N_199);
nand U753 (N_753,N_85,N_96);
or U754 (N_754,N_473,N_335);
nor U755 (N_755,N_256,N_479);
and U756 (N_756,N_319,N_242);
nor U757 (N_757,N_139,N_88);
nor U758 (N_758,N_461,N_168);
and U759 (N_759,N_249,N_384);
xnor U760 (N_760,N_279,N_133);
or U761 (N_761,N_171,N_427);
nor U762 (N_762,N_274,N_243);
nand U763 (N_763,N_163,N_231);
and U764 (N_764,N_176,N_69);
nor U765 (N_765,N_275,N_247);
and U766 (N_766,N_467,N_61);
nor U767 (N_767,N_495,N_304);
nor U768 (N_768,N_409,N_242);
nand U769 (N_769,N_16,N_0);
and U770 (N_770,N_174,N_454);
nand U771 (N_771,N_9,N_240);
or U772 (N_772,N_220,N_99);
nor U773 (N_773,N_324,N_34);
nand U774 (N_774,N_272,N_126);
nand U775 (N_775,N_195,N_356);
xnor U776 (N_776,N_349,N_236);
and U777 (N_777,N_149,N_55);
and U778 (N_778,N_442,N_432);
or U779 (N_779,N_306,N_181);
or U780 (N_780,N_121,N_356);
nand U781 (N_781,N_327,N_438);
and U782 (N_782,N_10,N_251);
and U783 (N_783,N_90,N_441);
nand U784 (N_784,N_53,N_416);
nand U785 (N_785,N_68,N_35);
nor U786 (N_786,N_194,N_452);
or U787 (N_787,N_58,N_271);
nor U788 (N_788,N_59,N_349);
and U789 (N_789,N_486,N_319);
nand U790 (N_790,N_316,N_404);
nand U791 (N_791,N_146,N_450);
or U792 (N_792,N_370,N_242);
nand U793 (N_793,N_265,N_129);
and U794 (N_794,N_187,N_273);
or U795 (N_795,N_67,N_118);
and U796 (N_796,N_290,N_431);
nand U797 (N_797,N_250,N_226);
nor U798 (N_798,N_160,N_383);
or U799 (N_799,N_290,N_93);
nand U800 (N_800,N_400,N_102);
nand U801 (N_801,N_126,N_111);
or U802 (N_802,N_71,N_117);
nor U803 (N_803,N_77,N_36);
or U804 (N_804,N_240,N_43);
nor U805 (N_805,N_3,N_383);
nand U806 (N_806,N_153,N_76);
or U807 (N_807,N_9,N_88);
and U808 (N_808,N_22,N_292);
or U809 (N_809,N_377,N_303);
nand U810 (N_810,N_489,N_147);
nor U811 (N_811,N_178,N_204);
xnor U812 (N_812,N_129,N_335);
nor U813 (N_813,N_195,N_332);
nand U814 (N_814,N_227,N_166);
nand U815 (N_815,N_40,N_338);
and U816 (N_816,N_131,N_403);
or U817 (N_817,N_310,N_15);
and U818 (N_818,N_390,N_267);
nor U819 (N_819,N_119,N_19);
nor U820 (N_820,N_258,N_380);
and U821 (N_821,N_147,N_129);
nor U822 (N_822,N_421,N_368);
and U823 (N_823,N_23,N_455);
and U824 (N_824,N_34,N_258);
or U825 (N_825,N_355,N_325);
or U826 (N_826,N_259,N_236);
and U827 (N_827,N_255,N_49);
and U828 (N_828,N_336,N_498);
nor U829 (N_829,N_228,N_381);
and U830 (N_830,N_242,N_5);
or U831 (N_831,N_440,N_412);
nand U832 (N_832,N_48,N_495);
and U833 (N_833,N_112,N_62);
and U834 (N_834,N_366,N_304);
or U835 (N_835,N_213,N_200);
and U836 (N_836,N_212,N_388);
and U837 (N_837,N_11,N_8);
and U838 (N_838,N_179,N_153);
and U839 (N_839,N_164,N_68);
nor U840 (N_840,N_35,N_310);
or U841 (N_841,N_26,N_9);
or U842 (N_842,N_224,N_130);
or U843 (N_843,N_87,N_34);
nand U844 (N_844,N_437,N_194);
nor U845 (N_845,N_105,N_273);
and U846 (N_846,N_379,N_20);
nand U847 (N_847,N_213,N_354);
nand U848 (N_848,N_28,N_181);
or U849 (N_849,N_12,N_414);
and U850 (N_850,N_132,N_242);
nor U851 (N_851,N_18,N_29);
or U852 (N_852,N_218,N_283);
or U853 (N_853,N_57,N_157);
nand U854 (N_854,N_179,N_110);
or U855 (N_855,N_254,N_119);
xnor U856 (N_856,N_490,N_199);
nand U857 (N_857,N_427,N_299);
nor U858 (N_858,N_490,N_494);
xnor U859 (N_859,N_0,N_237);
nand U860 (N_860,N_308,N_321);
and U861 (N_861,N_1,N_20);
nor U862 (N_862,N_70,N_380);
or U863 (N_863,N_100,N_84);
and U864 (N_864,N_165,N_416);
nand U865 (N_865,N_251,N_317);
or U866 (N_866,N_405,N_24);
and U867 (N_867,N_449,N_11);
and U868 (N_868,N_115,N_341);
nand U869 (N_869,N_252,N_430);
nor U870 (N_870,N_418,N_243);
nand U871 (N_871,N_34,N_39);
nor U872 (N_872,N_445,N_167);
nor U873 (N_873,N_44,N_488);
nand U874 (N_874,N_392,N_140);
nand U875 (N_875,N_202,N_64);
and U876 (N_876,N_318,N_332);
nor U877 (N_877,N_268,N_285);
and U878 (N_878,N_163,N_467);
and U879 (N_879,N_383,N_435);
nor U880 (N_880,N_277,N_195);
and U881 (N_881,N_296,N_174);
xnor U882 (N_882,N_113,N_217);
xnor U883 (N_883,N_397,N_112);
nand U884 (N_884,N_178,N_440);
nor U885 (N_885,N_151,N_234);
and U886 (N_886,N_286,N_125);
or U887 (N_887,N_158,N_144);
or U888 (N_888,N_275,N_452);
nor U889 (N_889,N_74,N_420);
nand U890 (N_890,N_37,N_30);
or U891 (N_891,N_139,N_314);
nor U892 (N_892,N_202,N_218);
xnor U893 (N_893,N_135,N_16);
xnor U894 (N_894,N_299,N_418);
and U895 (N_895,N_248,N_445);
or U896 (N_896,N_242,N_244);
nor U897 (N_897,N_416,N_102);
and U898 (N_898,N_154,N_131);
nor U899 (N_899,N_20,N_344);
nor U900 (N_900,N_157,N_485);
or U901 (N_901,N_78,N_348);
nor U902 (N_902,N_444,N_280);
nand U903 (N_903,N_193,N_479);
nor U904 (N_904,N_103,N_414);
or U905 (N_905,N_484,N_252);
and U906 (N_906,N_163,N_115);
nand U907 (N_907,N_18,N_434);
nand U908 (N_908,N_364,N_341);
and U909 (N_909,N_480,N_97);
and U910 (N_910,N_21,N_244);
nand U911 (N_911,N_452,N_351);
and U912 (N_912,N_426,N_132);
and U913 (N_913,N_180,N_283);
or U914 (N_914,N_354,N_430);
nand U915 (N_915,N_379,N_70);
nor U916 (N_916,N_85,N_161);
nand U917 (N_917,N_453,N_12);
or U918 (N_918,N_157,N_201);
or U919 (N_919,N_73,N_441);
or U920 (N_920,N_83,N_119);
nor U921 (N_921,N_342,N_234);
nor U922 (N_922,N_222,N_221);
or U923 (N_923,N_233,N_417);
or U924 (N_924,N_417,N_356);
xor U925 (N_925,N_132,N_262);
xor U926 (N_926,N_206,N_381);
nand U927 (N_927,N_59,N_153);
or U928 (N_928,N_356,N_214);
xnor U929 (N_929,N_389,N_108);
nor U930 (N_930,N_203,N_363);
or U931 (N_931,N_238,N_355);
or U932 (N_932,N_203,N_327);
nor U933 (N_933,N_5,N_11);
nand U934 (N_934,N_244,N_366);
or U935 (N_935,N_335,N_191);
nor U936 (N_936,N_249,N_312);
or U937 (N_937,N_266,N_427);
nor U938 (N_938,N_450,N_163);
nor U939 (N_939,N_433,N_87);
or U940 (N_940,N_458,N_319);
xnor U941 (N_941,N_306,N_114);
nand U942 (N_942,N_139,N_433);
nand U943 (N_943,N_214,N_154);
nand U944 (N_944,N_193,N_294);
or U945 (N_945,N_61,N_188);
and U946 (N_946,N_86,N_410);
xor U947 (N_947,N_133,N_61);
nand U948 (N_948,N_14,N_488);
and U949 (N_949,N_491,N_354);
and U950 (N_950,N_466,N_480);
nand U951 (N_951,N_225,N_299);
nor U952 (N_952,N_425,N_467);
xor U953 (N_953,N_411,N_378);
or U954 (N_954,N_377,N_17);
and U955 (N_955,N_390,N_86);
nand U956 (N_956,N_255,N_455);
nor U957 (N_957,N_434,N_93);
xor U958 (N_958,N_283,N_253);
or U959 (N_959,N_262,N_6);
or U960 (N_960,N_52,N_116);
nand U961 (N_961,N_403,N_328);
or U962 (N_962,N_440,N_240);
nor U963 (N_963,N_390,N_170);
and U964 (N_964,N_32,N_482);
and U965 (N_965,N_472,N_481);
or U966 (N_966,N_240,N_366);
and U967 (N_967,N_30,N_304);
or U968 (N_968,N_164,N_18);
nor U969 (N_969,N_314,N_81);
nor U970 (N_970,N_6,N_383);
or U971 (N_971,N_346,N_153);
xnor U972 (N_972,N_310,N_411);
and U973 (N_973,N_76,N_41);
and U974 (N_974,N_358,N_362);
nor U975 (N_975,N_1,N_286);
nor U976 (N_976,N_51,N_457);
nor U977 (N_977,N_253,N_122);
or U978 (N_978,N_261,N_379);
or U979 (N_979,N_47,N_185);
and U980 (N_980,N_430,N_472);
or U981 (N_981,N_411,N_443);
or U982 (N_982,N_63,N_422);
and U983 (N_983,N_219,N_5);
or U984 (N_984,N_343,N_476);
nor U985 (N_985,N_228,N_388);
nand U986 (N_986,N_156,N_89);
nand U987 (N_987,N_30,N_106);
nor U988 (N_988,N_23,N_176);
and U989 (N_989,N_64,N_361);
nand U990 (N_990,N_347,N_0);
or U991 (N_991,N_132,N_447);
and U992 (N_992,N_279,N_115);
or U993 (N_993,N_239,N_418);
nor U994 (N_994,N_324,N_97);
nand U995 (N_995,N_26,N_64);
or U996 (N_996,N_41,N_107);
nand U997 (N_997,N_117,N_96);
nor U998 (N_998,N_290,N_355);
and U999 (N_999,N_299,N_346);
nor U1000 (N_1000,N_819,N_566);
or U1001 (N_1001,N_848,N_772);
nand U1002 (N_1002,N_913,N_778);
and U1003 (N_1003,N_962,N_990);
and U1004 (N_1004,N_641,N_558);
nor U1005 (N_1005,N_878,N_787);
nand U1006 (N_1006,N_568,N_512);
and U1007 (N_1007,N_768,N_657);
or U1008 (N_1008,N_955,N_751);
nand U1009 (N_1009,N_977,N_814);
nor U1010 (N_1010,N_711,N_674);
nand U1011 (N_1011,N_600,N_598);
nor U1012 (N_1012,N_765,N_840);
nor U1013 (N_1013,N_827,N_922);
or U1014 (N_1014,N_527,N_627);
and U1015 (N_1015,N_638,N_549);
and U1016 (N_1016,N_694,N_681);
nand U1017 (N_1017,N_935,N_672);
xnor U1018 (N_1018,N_570,N_868);
nor U1019 (N_1019,N_552,N_893);
nor U1020 (N_1020,N_637,N_693);
nor U1021 (N_1021,N_924,N_669);
or U1022 (N_1022,N_722,N_979);
nand U1023 (N_1023,N_963,N_666);
or U1024 (N_1024,N_735,N_635);
nand U1025 (N_1025,N_952,N_554);
nor U1026 (N_1026,N_648,N_582);
nand U1027 (N_1027,N_896,N_576);
and U1028 (N_1028,N_695,N_523);
nor U1029 (N_1029,N_914,N_659);
or U1030 (N_1030,N_832,N_781);
and U1031 (N_1031,N_916,N_795);
nand U1032 (N_1032,N_583,N_629);
and U1033 (N_1033,N_730,N_759);
nor U1034 (N_1034,N_926,N_894);
nand U1035 (N_1035,N_531,N_766);
nand U1036 (N_1036,N_650,N_737);
or U1037 (N_1037,N_544,N_941);
xor U1038 (N_1038,N_587,N_954);
or U1039 (N_1039,N_520,N_621);
and U1040 (N_1040,N_615,N_713);
nand U1041 (N_1041,N_969,N_515);
nor U1042 (N_1042,N_890,N_804);
nand U1043 (N_1043,N_876,N_692);
or U1044 (N_1044,N_510,N_930);
and U1045 (N_1045,N_812,N_987);
xnor U1046 (N_1046,N_902,N_647);
nand U1047 (N_1047,N_503,N_780);
nor U1048 (N_1048,N_502,N_771);
or U1049 (N_1049,N_945,N_741);
nand U1050 (N_1050,N_698,N_517);
nand U1051 (N_1051,N_589,N_970);
nor U1052 (N_1052,N_511,N_709);
xnor U1053 (N_1053,N_883,N_733);
nor U1054 (N_1054,N_664,N_519);
nand U1055 (N_1055,N_953,N_701);
nand U1056 (N_1056,N_911,N_616);
and U1057 (N_1057,N_724,N_938);
or U1058 (N_1058,N_572,N_636);
or U1059 (N_1059,N_707,N_948);
xnor U1060 (N_1060,N_994,N_907);
nand U1061 (N_1061,N_956,N_612);
and U1062 (N_1062,N_861,N_599);
or U1063 (N_1063,N_833,N_667);
nand U1064 (N_1064,N_550,N_915);
or U1065 (N_1065,N_507,N_811);
nor U1066 (N_1066,N_597,N_988);
nand U1067 (N_1067,N_663,N_533);
nor U1068 (N_1068,N_508,N_714);
nand U1069 (N_1069,N_783,N_619);
or U1070 (N_1070,N_665,N_605);
and U1071 (N_1071,N_891,N_775);
nor U1072 (N_1072,N_660,N_836);
or U1073 (N_1073,N_633,N_983);
and U1074 (N_1074,N_539,N_606);
or U1075 (N_1075,N_720,N_951);
xor U1076 (N_1076,N_909,N_847);
and U1077 (N_1077,N_851,N_679);
and U1078 (N_1078,N_610,N_688);
nand U1079 (N_1079,N_573,N_949);
and U1080 (N_1080,N_680,N_564);
or U1081 (N_1081,N_622,N_927);
nand U1082 (N_1082,N_726,N_823);
or U1083 (N_1083,N_542,N_586);
or U1084 (N_1084,N_653,N_806);
or U1085 (N_1085,N_906,N_541);
or U1086 (N_1086,N_846,N_585);
nor U1087 (N_1087,N_630,N_905);
nand U1088 (N_1088,N_860,N_658);
or U1089 (N_1089,N_690,N_543);
nor U1090 (N_1090,N_723,N_639);
nor U1091 (N_1091,N_750,N_699);
nor U1092 (N_1092,N_535,N_863);
xor U1093 (N_1093,N_700,N_525);
and U1094 (N_1094,N_997,N_964);
xnor U1095 (N_1095,N_829,N_559);
and U1096 (N_1096,N_545,N_529);
nor U1097 (N_1097,N_798,N_601);
nand U1098 (N_1098,N_763,N_591);
and U1099 (N_1099,N_547,N_801);
nand U1100 (N_1100,N_805,N_675);
and U1101 (N_1101,N_684,N_626);
and U1102 (N_1102,N_501,N_875);
nand U1103 (N_1103,N_901,N_655);
and U1104 (N_1104,N_555,N_925);
or U1105 (N_1105,N_685,N_966);
and U1106 (N_1106,N_516,N_959);
xnor U1107 (N_1107,N_882,N_934);
nor U1108 (N_1108,N_683,N_594);
nor U1109 (N_1109,N_944,N_769);
and U1110 (N_1110,N_537,N_993);
or U1111 (N_1111,N_967,N_816);
nor U1112 (N_1112,N_887,N_578);
nor U1113 (N_1113,N_652,N_841);
and U1114 (N_1114,N_785,N_719);
or U1115 (N_1115,N_509,N_611);
nor U1116 (N_1116,N_839,N_689);
nand U1117 (N_1117,N_718,N_886);
or U1118 (N_1118,N_736,N_852);
and U1119 (N_1119,N_725,N_802);
xnor U1120 (N_1120,N_739,N_968);
nor U1121 (N_1121,N_603,N_928);
nor U1122 (N_1122,N_796,N_978);
nand U1123 (N_1123,N_793,N_834);
xnor U1124 (N_1124,N_831,N_874);
xor U1125 (N_1125,N_577,N_628);
nand U1126 (N_1126,N_943,N_682);
nand U1127 (N_1127,N_844,N_623);
nor U1128 (N_1128,N_872,N_818);
and U1129 (N_1129,N_743,N_538);
and U1130 (N_1130,N_734,N_620);
nand U1131 (N_1131,N_937,N_995);
xor U1132 (N_1132,N_705,N_703);
nor U1133 (N_1133,N_820,N_590);
nor U1134 (N_1134,N_624,N_755);
nand U1135 (N_1135,N_656,N_506);
nor U1136 (N_1136,N_923,N_644);
or U1137 (N_1137,N_731,N_563);
nor U1138 (N_1138,N_965,N_897);
nand U1139 (N_1139,N_746,N_727);
nand U1140 (N_1140,N_918,N_634);
nor U1141 (N_1141,N_807,N_957);
and U1142 (N_1142,N_546,N_526);
nor U1143 (N_1143,N_551,N_826);
or U1144 (N_1144,N_919,N_649);
or U1145 (N_1145,N_614,N_929);
or U1146 (N_1146,N_946,N_985);
and U1147 (N_1147,N_640,N_867);
nand U1148 (N_1148,N_749,N_940);
nand U1149 (N_1149,N_879,N_857);
or U1150 (N_1150,N_608,N_686);
nor U1151 (N_1151,N_961,N_996);
and U1152 (N_1152,N_976,N_855);
xor U1153 (N_1153,N_671,N_910);
nand U1154 (N_1154,N_975,N_715);
xor U1155 (N_1155,N_898,N_732);
nor U1156 (N_1156,N_782,N_748);
and U1157 (N_1157,N_895,N_654);
xor U1158 (N_1158,N_813,N_553);
nor U1159 (N_1159,N_838,N_609);
and U1160 (N_1160,N_604,N_788);
and U1161 (N_1161,N_595,N_702);
and U1162 (N_1162,N_642,N_825);
nor U1163 (N_1163,N_862,N_899);
nor U1164 (N_1164,N_856,N_774);
or U1165 (N_1165,N_842,N_903);
xor U1166 (N_1166,N_858,N_822);
nor U1167 (N_1167,N_540,N_973);
or U1168 (N_1168,N_728,N_933);
nand U1169 (N_1169,N_931,N_617);
nand U1170 (N_1170,N_631,N_687);
nor U1171 (N_1171,N_513,N_888);
or U1172 (N_1172,N_999,N_797);
and U1173 (N_1173,N_565,N_932);
or U1174 (N_1174,N_752,N_784);
or U1175 (N_1175,N_984,N_754);
nor U1176 (N_1176,N_717,N_625);
and U1177 (N_1177,N_921,N_668);
and U1178 (N_1178,N_974,N_697);
or U1179 (N_1179,N_849,N_579);
and U1180 (N_1180,N_505,N_528);
and U1181 (N_1181,N_602,N_869);
or U1182 (N_1182,N_767,N_691);
and U1183 (N_1183,N_518,N_696);
or U1184 (N_1184,N_871,N_661);
nor U1185 (N_1185,N_991,N_588);
xor U1186 (N_1186,N_950,N_877);
nand U1187 (N_1187,N_794,N_662);
nand U1188 (N_1188,N_845,N_676);
nand U1189 (N_1189,N_721,N_574);
or U1190 (N_1190,N_920,N_981);
or U1191 (N_1191,N_980,N_792);
or U1192 (N_1192,N_947,N_740);
or U1193 (N_1193,N_908,N_837);
or U1194 (N_1194,N_651,N_738);
nand U1195 (N_1195,N_853,N_548);
xor U1196 (N_1196,N_828,N_971);
nor U1197 (N_1197,N_799,N_557);
and U1198 (N_1198,N_561,N_912);
or U1199 (N_1199,N_810,N_989);
xnor U1200 (N_1200,N_998,N_534);
and U1201 (N_1201,N_881,N_884);
nor U1202 (N_1202,N_560,N_524);
nand U1203 (N_1203,N_789,N_607);
and U1204 (N_1204,N_581,N_569);
nand U1205 (N_1205,N_786,N_815);
nor U1206 (N_1206,N_678,N_972);
nand U1207 (N_1207,N_567,N_673);
nand U1208 (N_1208,N_632,N_514);
nor U1209 (N_1209,N_821,N_892);
nor U1210 (N_1210,N_521,N_936);
and U1211 (N_1211,N_764,N_939);
and U1212 (N_1212,N_779,N_777);
xnor U1213 (N_1213,N_530,N_817);
nor U1214 (N_1214,N_536,N_592);
or U1215 (N_1215,N_580,N_873);
or U1216 (N_1216,N_889,N_942);
nand U1217 (N_1217,N_790,N_850);
or U1218 (N_1218,N_646,N_865);
nor U1219 (N_1219,N_716,N_992);
nor U1220 (N_1220,N_762,N_562);
nand U1221 (N_1221,N_960,N_917);
nand U1222 (N_1222,N_677,N_500);
and U1223 (N_1223,N_835,N_770);
nand U1224 (N_1224,N_747,N_613);
xor U1225 (N_1225,N_532,N_824);
or U1226 (N_1226,N_885,N_758);
xor U1227 (N_1227,N_596,N_756);
or U1228 (N_1228,N_800,N_670);
nor U1229 (N_1229,N_556,N_859);
or U1230 (N_1230,N_986,N_982);
nor U1231 (N_1231,N_843,N_504);
and U1232 (N_1232,N_584,N_729);
xnor U1233 (N_1233,N_803,N_904);
nand U1234 (N_1234,N_593,N_643);
or U1235 (N_1235,N_900,N_773);
or U1236 (N_1236,N_864,N_830);
or U1237 (N_1237,N_706,N_809);
nor U1238 (N_1238,N_708,N_880);
nand U1239 (N_1239,N_757,N_571);
and U1240 (N_1240,N_870,N_791);
nor U1241 (N_1241,N_753,N_776);
and U1242 (N_1242,N_704,N_761);
nor U1243 (N_1243,N_712,N_854);
or U1244 (N_1244,N_808,N_866);
and U1245 (N_1245,N_618,N_958);
nor U1246 (N_1246,N_710,N_742);
and U1247 (N_1247,N_744,N_760);
and U1248 (N_1248,N_745,N_522);
nand U1249 (N_1249,N_645,N_575);
nor U1250 (N_1250,N_531,N_632);
nor U1251 (N_1251,N_997,N_527);
or U1252 (N_1252,N_540,N_534);
and U1253 (N_1253,N_529,N_838);
nand U1254 (N_1254,N_994,N_791);
nor U1255 (N_1255,N_885,N_674);
or U1256 (N_1256,N_877,N_506);
and U1257 (N_1257,N_912,N_768);
nor U1258 (N_1258,N_646,N_583);
and U1259 (N_1259,N_811,N_999);
or U1260 (N_1260,N_892,N_768);
nor U1261 (N_1261,N_691,N_971);
and U1262 (N_1262,N_526,N_631);
xnor U1263 (N_1263,N_955,N_770);
xnor U1264 (N_1264,N_873,N_625);
nor U1265 (N_1265,N_829,N_976);
and U1266 (N_1266,N_960,N_579);
nor U1267 (N_1267,N_803,N_980);
nand U1268 (N_1268,N_699,N_909);
or U1269 (N_1269,N_563,N_878);
or U1270 (N_1270,N_526,N_977);
xnor U1271 (N_1271,N_952,N_849);
nor U1272 (N_1272,N_664,N_654);
or U1273 (N_1273,N_796,N_649);
and U1274 (N_1274,N_893,N_701);
xor U1275 (N_1275,N_594,N_913);
nor U1276 (N_1276,N_714,N_904);
nor U1277 (N_1277,N_964,N_788);
nand U1278 (N_1278,N_780,N_671);
nor U1279 (N_1279,N_983,N_645);
or U1280 (N_1280,N_648,N_501);
nor U1281 (N_1281,N_831,N_807);
nor U1282 (N_1282,N_621,N_787);
xnor U1283 (N_1283,N_934,N_549);
or U1284 (N_1284,N_501,N_816);
and U1285 (N_1285,N_918,N_962);
or U1286 (N_1286,N_944,N_791);
nand U1287 (N_1287,N_975,N_723);
xor U1288 (N_1288,N_937,N_985);
or U1289 (N_1289,N_976,N_765);
nor U1290 (N_1290,N_770,N_890);
nor U1291 (N_1291,N_566,N_512);
and U1292 (N_1292,N_668,N_713);
and U1293 (N_1293,N_598,N_913);
nor U1294 (N_1294,N_534,N_719);
and U1295 (N_1295,N_872,N_739);
xor U1296 (N_1296,N_929,N_688);
nor U1297 (N_1297,N_676,N_593);
xor U1298 (N_1298,N_686,N_700);
or U1299 (N_1299,N_512,N_805);
and U1300 (N_1300,N_743,N_841);
and U1301 (N_1301,N_679,N_841);
and U1302 (N_1302,N_724,N_992);
xnor U1303 (N_1303,N_928,N_909);
and U1304 (N_1304,N_856,N_736);
or U1305 (N_1305,N_811,N_711);
xnor U1306 (N_1306,N_743,N_725);
nand U1307 (N_1307,N_561,N_865);
and U1308 (N_1308,N_667,N_636);
and U1309 (N_1309,N_889,N_687);
nor U1310 (N_1310,N_614,N_696);
or U1311 (N_1311,N_583,N_922);
or U1312 (N_1312,N_926,N_648);
nor U1313 (N_1313,N_824,N_997);
and U1314 (N_1314,N_957,N_603);
nor U1315 (N_1315,N_726,N_693);
nor U1316 (N_1316,N_670,N_501);
and U1317 (N_1317,N_730,N_940);
and U1318 (N_1318,N_968,N_605);
or U1319 (N_1319,N_779,N_818);
nand U1320 (N_1320,N_910,N_545);
or U1321 (N_1321,N_611,N_918);
nor U1322 (N_1322,N_952,N_828);
xnor U1323 (N_1323,N_962,N_868);
and U1324 (N_1324,N_564,N_787);
or U1325 (N_1325,N_809,N_872);
xnor U1326 (N_1326,N_541,N_663);
nand U1327 (N_1327,N_958,N_577);
nor U1328 (N_1328,N_927,N_941);
xor U1329 (N_1329,N_953,N_755);
nor U1330 (N_1330,N_573,N_607);
nand U1331 (N_1331,N_825,N_668);
and U1332 (N_1332,N_783,N_757);
or U1333 (N_1333,N_651,N_785);
nand U1334 (N_1334,N_810,N_770);
xnor U1335 (N_1335,N_600,N_656);
nand U1336 (N_1336,N_681,N_637);
nand U1337 (N_1337,N_876,N_693);
nand U1338 (N_1338,N_541,N_877);
nand U1339 (N_1339,N_698,N_910);
xnor U1340 (N_1340,N_951,N_873);
nor U1341 (N_1341,N_860,N_874);
or U1342 (N_1342,N_635,N_757);
xor U1343 (N_1343,N_531,N_783);
or U1344 (N_1344,N_534,N_907);
xor U1345 (N_1345,N_888,N_534);
nand U1346 (N_1346,N_532,N_874);
nor U1347 (N_1347,N_771,N_969);
nand U1348 (N_1348,N_748,N_966);
or U1349 (N_1349,N_548,N_762);
nor U1350 (N_1350,N_557,N_623);
or U1351 (N_1351,N_676,N_541);
nor U1352 (N_1352,N_746,N_545);
nor U1353 (N_1353,N_872,N_979);
nand U1354 (N_1354,N_915,N_624);
nand U1355 (N_1355,N_937,N_669);
nand U1356 (N_1356,N_535,N_699);
or U1357 (N_1357,N_638,N_546);
nand U1358 (N_1358,N_904,N_812);
or U1359 (N_1359,N_608,N_658);
xnor U1360 (N_1360,N_849,N_707);
nor U1361 (N_1361,N_718,N_588);
xnor U1362 (N_1362,N_671,N_836);
nand U1363 (N_1363,N_891,N_849);
xor U1364 (N_1364,N_544,N_530);
nand U1365 (N_1365,N_640,N_723);
xor U1366 (N_1366,N_731,N_674);
nand U1367 (N_1367,N_567,N_589);
or U1368 (N_1368,N_787,N_701);
xor U1369 (N_1369,N_799,N_578);
and U1370 (N_1370,N_927,N_964);
nand U1371 (N_1371,N_764,N_727);
and U1372 (N_1372,N_618,N_664);
or U1373 (N_1373,N_900,N_537);
nor U1374 (N_1374,N_987,N_552);
xor U1375 (N_1375,N_636,N_558);
nor U1376 (N_1376,N_709,N_792);
or U1377 (N_1377,N_964,N_822);
nand U1378 (N_1378,N_526,N_691);
and U1379 (N_1379,N_615,N_544);
nor U1380 (N_1380,N_565,N_550);
nand U1381 (N_1381,N_612,N_506);
nand U1382 (N_1382,N_835,N_924);
nand U1383 (N_1383,N_597,N_865);
or U1384 (N_1384,N_874,N_788);
xor U1385 (N_1385,N_682,N_973);
and U1386 (N_1386,N_750,N_603);
nand U1387 (N_1387,N_743,N_520);
or U1388 (N_1388,N_880,N_747);
nor U1389 (N_1389,N_701,N_890);
nand U1390 (N_1390,N_971,N_587);
and U1391 (N_1391,N_876,N_892);
and U1392 (N_1392,N_645,N_745);
nand U1393 (N_1393,N_863,N_918);
nand U1394 (N_1394,N_961,N_815);
nand U1395 (N_1395,N_536,N_542);
or U1396 (N_1396,N_907,N_666);
and U1397 (N_1397,N_960,N_510);
xnor U1398 (N_1398,N_504,N_951);
nand U1399 (N_1399,N_583,N_918);
nor U1400 (N_1400,N_632,N_913);
and U1401 (N_1401,N_872,N_747);
and U1402 (N_1402,N_842,N_835);
nand U1403 (N_1403,N_603,N_921);
nor U1404 (N_1404,N_557,N_814);
nor U1405 (N_1405,N_821,N_660);
and U1406 (N_1406,N_899,N_932);
or U1407 (N_1407,N_757,N_986);
nand U1408 (N_1408,N_615,N_611);
or U1409 (N_1409,N_757,N_514);
nor U1410 (N_1410,N_521,N_623);
and U1411 (N_1411,N_631,N_903);
and U1412 (N_1412,N_926,N_804);
and U1413 (N_1413,N_820,N_706);
nor U1414 (N_1414,N_851,N_526);
or U1415 (N_1415,N_921,N_679);
and U1416 (N_1416,N_552,N_755);
or U1417 (N_1417,N_729,N_792);
and U1418 (N_1418,N_651,N_735);
or U1419 (N_1419,N_697,N_648);
nor U1420 (N_1420,N_806,N_613);
nand U1421 (N_1421,N_771,N_978);
and U1422 (N_1422,N_877,N_882);
and U1423 (N_1423,N_872,N_532);
and U1424 (N_1424,N_706,N_691);
xnor U1425 (N_1425,N_834,N_812);
nand U1426 (N_1426,N_502,N_559);
and U1427 (N_1427,N_767,N_905);
nor U1428 (N_1428,N_939,N_530);
nand U1429 (N_1429,N_745,N_500);
nor U1430 (N_1430,N_581,N_918);
or U1431 (N_1431,N_679,N_842);
nor U1432 (N_1432,N_771,N_812);
nor U1433 (N_1433,N_903,N_509);
or U1434 (N_1434,N_796,N_793);
or U1435 (N_1435,N_518,N_516);
nand U1436 (N_1436,N_923,N_509);
or U1437 (N_1437,N_737,N_591);
and U1438 (N_1438,N_611,N_947);
nand U1439 (N_1439,N_532,N_559);
nand U1440 (N_1440,N_951,N_866);
and U1441 (N_1441,N_825,N_838);
and U1442 (N_1442,N_817,N_948);
nor U1443 (N_1443,N_925,N_563);
and U1444 (N_1444,N_665,N_586);
xor U1445 (N_1445,N_960,N_534);
nor U1446 (N_1446,N_741,N_593);
and U1447 (N_1447,N_783,N_550);
nor U1448 (N_1448,N_922,N_669);
or U1449 (N_1449,N_550,N_559);
and U1450 (N_1450,N_738,N_843);
and U1451 (N_1451,N_996,N_850);
or U1452 (N_1452,N_546,N_763);
or U1453 (N_1453,N_686,N_643);
nand U1454 (N_1454,N_577,N_736);
nor U1455 (N_1455,N_661,N_912);
and U1456 (N_1456,N_700,N_658);
nor U1457 (N_1457,N_511,N_967);
and U1458 (N_1458,N_590,N_892);
and U1459 (N_1459,N_769,N_510);
nor U1460 (N_1460,N_933,N_602);
nand U1461 (N_1461,N_782,N_764);
and U1462 (N_1462,N_724,N_990);
nand U1463 (N_1463,N_597,N_932);
or U1464 (N_1464,N_549,N_561);
xor U1465 (N_1465,N_953,N_835);
nor U1466 (N_1466,N_757,N_561);
nand U1467 (N_1467,N_847,N_609);
nand U1468 (N_1468,N_956,N_570);
or U1469 (N_1469,N_761,N_826);
and U1470 (N_1470,N_759,N_746);
and U1471 (N_1471,N_776,N_586);
xnor U1472 (N_1472,N_967,N_602);
and U1473 (N_1473,N_823,N_977);
nor U1474 (N_1474,N_923,N_651);
and U1475 (N_1475,N_567,N_746);
nor U1476 (N_1476,N_512,N_630);
nand U1477 (N_1477,N_605,N_800);
nor U1478 (N_1478,N_749,N_854);
nand U1479 (N_1479,N_856,N_661);
and U1480 (N_1480,N_557,N_524);
or U1481 (N_1481,N_520,N_598);
nand U1482 (N_1482,N_554,N_620);
and U1483 (N_1483,N_904,N_520);
nand U1484 (N_1484,N_506,N_644);
xor U1485 (N_1485,N_997,N_899);
nand U1486 (N_1486,N_807,N_703);
nand U1487 (N_1487,N_869,N_793);
and U1488 (N_1488,N_593,N_852);
or U1489 (N_1489,N_732,N_666);
and U1490 (N_1490,N_812,N_906);
or U1491 (N_1491,N_580,N_912);
and U1492 (N_1492,N_636,N_686);
and U1493 (N_1493,N_838,N_577);
and U1494 (N_1494,N_879,N_516);
or U1495 (N_1495,N_786,N_880);
xor U1496 (N_1496,N_796,N_788);
and U1497 (N_1497,N_687,N_812);
xnor U1498 (N_1498,N_717,N_769);
nor U1499 (N_1499,N_846,N_929);
or U1500 (N_1500,N_1295,N_1433);
nand U1501 (N_1501,N_1184,N_1408);
or U1502 (N_1502,N_1284,N_1423);
xnor U1503 (N_1503,N_1390,N_1254);
nor U1504 (N_1504,N_1221,N_1490);
or U1505 (N_1505,N_1217,N_1045);
nand U1506 (N_1506,N_1151,N_1074);
nand U1507 (N_1507,N_1168,N_1439);
or U1508 (N_1508,N_1305,N_1145);
nor U1509 (N_1509,N_1071,N_1154);
nand U1510 (N_1510,N_1068,N_1326);
and U1511 (N_1511,N_1426,N_1443);
nand U1512 (N_1512,N_1107,N_1122);
nor U1513 (N_1513,N_1409,N_1070);
nand U1514 (N_1514,N_1213,N_1281);
nor U1515 (N_1515,N_1231,N_1170);
nor U1516 (N_1516,N_1033,N_1123);
nor U1517 (N_1517,N_1324,N_1258);
xor U1518 (N_1518,N_1310,N_1178);
nand U1519 (N_1519,N_1169,N_1113);
and U1520 (N_1520,N_1028,N_1016);
or U1521 (N_1521,N_1472,N_1455);
or U1522 (N_1522,N_1108,N_1207);
nand U1523 (N_1523,N_1470,N_1088);
nor U1524 (N_1524,N_1488,N_1351);
nand U1525 (N_1525,N_1196,N_1462);
and U1526 (N_1526,N_1046,N_1319);
or U1527 (N_1527,N_1369,N_1388);
xor U1528 (N_1528,N_1224,N_1066);
xnor U1529 (N_1529,N_1360,N_1456);
or U1530 (N_1530,N_1348,N_1322);
nor U1531 (N_1531,N_1138,N_1427);
or U1532 (N_1532,N_1367,N_1252);
or U1533 (N_1533,N_1392,N_1090);
nor U1534 (N_1534,N_1054,N_1289);
and U1535 (N_1535,N_1299,N_1243);
and U1536 (N_1536,N_1082,N_1361);
nor U1537 (N_1537,N_1079,N_1304);
or U1538 (N_1538,N_1211,N_1004);
nor U1539 (N_1539,N_1349,N_1106);
or U1540 (N_1540,N_1134,N_1487);
xnor U1541 (N_1541,N_1063,N_1478);
or U1542 (N_1542,N_1204,N_1333);
xnor U1543 (N_1543,N_1429,N_1334);
and U1544 (N_1544,N_1386,N_1461);
or U1545 (N_1545,N_1125,N_1194);
xor U1546 (N_1546,N_1497,N_1047);
nor U1547 (N_1547,N_1007,N_1263);
or U1548 (N_1548,N_1378,N_1411);
nand U1549 (N_1549,N_1142,N_1301);
and U1550 (N_1550,N_1491,N_1446);
nor U1551 (N_1551,N_1286,N_1437);
or U1552 (N_1552,N_1012,N_1255);
or U1553 (N_1553,N_1019,N_1037);
xnor U1554 (N_1554,N_1148,N_1379);
nand U1555 (N_1555,N_1308,N_1156);
nand U1556 (N_1556,N_1459,N_1280);
nand U1557 (N_1557,N_1475,N_1331);
and U1558 (N_1558,N_1215,N_1352);
nor U1559 (N_1559,N_1273,N_1303);
and U1560 (N_1560,N_1422,N_1397);
xor U1561 (N_1561,N_1223,N_1257);
nand U1562 (N_1562,N_1401,N_1393);
or U1563 (N_1563,N_1230,N_1098);
and U1564 (N_1564,N_1262,N_1483);
or U1565 (N_1565,N_1067,N_1233);
nand U1566 (N_1566,N_1136,N_1132);
xnor U1567 (N_1567,N_1005,N_1155);
xnor U1568 (N_1568,N_1271,N_1009);
nor U1569 (N_1569,N_1244,N_1050);
nand U1570 (N_1570,N_1342,N_1246);
and U1571 (N_1571,N_1405,N_1064);
and U1572 (N_1572,N_1476,N_1293);
or U1573 (N_1573,N_1116,N_1274);
and U1574 (N_1574,N_1278,N_1372);
or U1575 (N_1575,N_1279,N_1402);
nor U1576 (N_1576,N_1094,N_1053);
nand U1577 (N_1577,N_1248,N_1103);
xor U1578 (N_1578,N_1292,N_1216);
and U1579 (N_1579,N_1049,N_1335);
nand U1580 (N_1580,N_1118,N_1022);
nor U1581 (N_1581,N_1198,N_1256);
nor U1582 (N_1582,N_1031,N_1466);
or U1583 (N_1583,N_1359,N_1077);
xnor U1584 (N_1584,N_1201,N_1172);
or U1585 (N_1585,N_1241,N_1374);
xnor U1586 (N_1586,N_1365,N_1384);
nand U1587 (N_1587,N_1339,N_1415);
nand U1588 (N_1588,N_1327,N_1385);
and U1589 (N_1589,N_1057,N_1364);
nor U1590 (N_1590,N_1105,N_1065);
nand U1591 (N_1591,N_1418,N_1164);
nand U1592 (N_1592,N_1381,N_1101);
nand U1593 (N_1593,N_1208,N_1355);
xnor U1594 (N_1594,N_1190,N_1083);
and U1595 (N_1595,N_1290,N_1084);
and U1596 (N_1596,N_1356,N_1314);
nand U1597 (N_1597,N_1311,N_1424);
xor U1598 (N_1598,N_1159,N_1078);
and U1599 (N_1599,N_1363,N_1099);
xor U1600 (N_1600,N_1102,N_1186);
nor U1601 (N_1601,N_1225,N_1160);
or U1602 (N_1602,N_1336,N_1171);
nand U1603 (N_1603,N_1344,N_1181);
nor U1604 (N_1604,N_1110,N_1152);
and U1605 (N_1605,N_1269,N_1484);
xor U1606 (N_1606,N_1234,N_1357);
or U1607 (N_1607,N_1307,N_1329);
or U1608 (N_1608,N_1345,N_1353);
nor U1609 (N_1609,N_1312,N_1195);
nor U1610 (N_1610,N_1149,N_1463);
xor U1611 (N_1611,N_1300,N_1062);
xnor U1612 (N_1612,N_1250,N_1283);
or U1613 (N_1613,N_1377,N_1193);
nand U1614 (N_1614,N_1086,N_1052);
nand U1615 (N_1615,N_1093,N_1180);
and U1616 (N_1616,N_1051,N_1163);
or U1617 (N_1617,N_1058,N_1153);
nand U1618 (N_1618,N_1400,N_1089);
nand U1619 (N_1619,N_1282,N_1436);
xnor U1620 (N_1620,N_1261,N_1450);
or U1621 (N_1621,N_1404,N_1027);
or U1622 (N_1622,N_1492,N_1496);
nor U1623 (N_1623,N_1120,N_1318);
and U1624 (N_1624,N_1410,N_1147);
or U1625 (N_1625,N_1416,N_1200);
nor U1626 (N_1626,N_1294,N_1471);
or U1627 (N_1627,N_1214,N_1115);
nor U1628 (N_1628,N_1347,N_1477);
or U1629 (N_1629,N_1238,N_1036);
xor U1630 (N_1630,N_1040,N_1112);
or U1631 (N_1631,N_1444,N_1001);
xnor U1632 (N_1632,N_1270,N_1288);
or U1633 (N_1633,N_1212,N_1403);
or U1634 (N_1634,N_1197,N_1267);
or U1635 (N_1635,N_1398,N_1265);
and U1636 (N_1636,N_1209,N_1465);
nor U1637 (N_1637,N_1218,N_1240);
xnor U1638 (N_1638,N_1239,N_1157);
and U1639 (N_1639,N_1126,N_1144);
nand U1640 (N_1640,N_1018,N_1495);
nor U1641 (N_1641,N_1006,N_1291);
or U1642 (N_1642,N_1366,N_1253);
and U1643 (N_1643,N_1296,N_1306);
nand U1644 (N_1644,N_1260,N_1313);
nand U1645 (N_1645,N_1371,N_1407);
xnor U1646 (N_1646,N_1376,N_1457);
nand U1647 (N_1647,N_1061,N_1259);
nor U1648 (N_1648,N_1245,N_1297);
and U1649 (N_1649,N_1174,N_1232);
nor U1650 (N_1650,N_1375,N_1023);
or U1651 (N_1651,N_1119,N_1150);
or U1652 (N_1652,N_1428,N_1185);
or U1653 (N_1653,N_1383,N_1141);
and U1654 (N_1654,N_1468,N_1104);
and U1655 (N_1655,N_1075,N_1338);
and U1656 (N_1656,N_1458,N_1453);
nor U1657 (N_1657,N_1073,N_1048);
and U1658 (N_1658,N_1128,N_1412);
and U1659 (N_1659,N_1399,N_1341);
and U1660 (N_1660,N_1220,N_1467);
nand U1661 (N_1661,N_1285,N_1121);
or U1662 (N_1662,N_1140,N_1362);
xor U1663 (N_1663,N_1124,N_1277);
or U1664 (N_1664,N_1056,N_1139);
xor U1665 (N_1665,N_1029,N_1039);
xnor U1666 (N_1666,N_1162,N_1100);
xor U1667 (N_1667,N_1229,N_1095);
xnor U1668 (N_1668,N_1130,N_1041);
or U1669 (N_1669,N_1191,N_1432);
nand U1670 (N_1670,N_1451,N_1203);
or U1671 (N_1671,N_1494,N_1275);
or U1672 (N_1672,N_1091,N_1069);
nand U1673 (N_1673,N_1021,N_1438);
nand U1674 (N_1674,N_1222,N_1354);
or U1675 (N_1675,N_1435,N_1413);
nor U1676 (N_1676,N_1445,N_1043);
nand U1677 (N_1677,N_1146,N_1396);
nor U1678 (N_1678,N_1205,N_1109);
nor U1679 (N_1679,N_1481,N_1264);
nor U1680 (N_1680,N_1173,N_1228);
and U1681 (N_1681,N_1420,N_1325);
nand U1682 (N_1682,N_1251,N_1340);
nor U1683 (N_1683,N_1485,N_1008);
and U1684 (N_1684,N_1454,N_1202);
or U1685 (N_1685,N_1013,N_1449);
and U1686 (N_1686,N_1085,N_1489);
or U1687 (N_1687,N_1117,N_1072);
and U1688 (N_1688,N_1431,N_1176);
nor U1689 (N_1689,N_1421,N_1323);
and U1690 (N_1690,N_1235,N_1189);
nor U1691 (N_1691,N_1135,N_1441);
xor U1692 (N_1692,N_1442,N_1080);
or U1693 (N_1693,N_1486,N_1425);
nand U1694 (N_1694,N_1014,N_1317);
nor U1695 (N_1695,N_1346,N_1414);
nand U1696 (N_1696,N_1003,N_1219);
nand U1697 (N_1697,N_1081,N_1447);
nand U1698 (N_1698,N_1474,N_1247);
and U1699 (N_1699,N_1302,N_1010);
nor U1700 (N_1700,N_1499,N_1266);
and U1701 (N_1701,N_1309,N_1242);
and U1702 (N_1702,N_1315,N_1059);
nand U1703 (N_1703,N_1042,N_1249);
nor U1704 (N_1704,N_1226,N_1026);
and U1705 (N_1705,N_1129,N_1337);
and U1706 (N_1706,N_1469,N_1076);
xnor U1707 (N_1707,N_1479,N_1227);
and U1708 (N_1708,N_1237,N_1358);
and U1709 (N_1709,N_1133,N_1394);
and U1710 (N_1710,N_1158,N_1055);
and U1711 (N_1711,N_1498,N_1320);
or U1712 (N_1712,N_1167,N_1030);
and U1713 (N_1713,N_1002,N_1332);
or U1714 (N_1714,N_1480,N_1452);
nand U1715 (N_1715,N_1464,N_1188);
and U1716 (N_1716,N_1166,N_1092);
xor U1717 (N_1717,N_1268,N_1183);
xor U1718 (N_1718,N_1044,N_1143);
and U1719 (N_1719,N_1034,N_1020);
nand U1720 (N_1720,N_1210,N_1287);
or U1721 (N_1721,N_1460,N_1111);
and U1722 (N_1722,N_1017,N_1011);
nor U1723 (N_1723,N_1199,N_1032);
nor U1724 (N_1724,N_1417,N_1161);
nor U1725 (N_1725,N_1015,N_1370);
nor U1726 (N_1726,N_1395,N_1316);
nor U1727 (N_1727,N_1330,N_1448);
nor U1728 (N_1728,N_1114,N_1236);
or U1729 (N_1729,N_1177,N_1387);
and U1730 (N_1730,N_1406,N_1179);
and U1731 (N_1731,N_1038,N_1137);
or U1732 (N_1732,N_1430,N_1321);
or U1733 (N_1733,N_1096,N_1175);
xor U1734 (N_1734,N_1380,N_1328);
xor U1735 (N_1735,N_1343,N_1298);
nor U1736 (N_1736,N_1182,N_1373);
nor U1737 (N_1737,N_1060,N_1482);
nand U1738 (N_1738,N_1035,N_1350);
nor U1739 (N_1739,N_1206,N_1368);
nand U1740 (N_1740,N_1493,N_1419);
nor U1741 (N_1741,N_1192,N_1097);
nand U1742 (N_1742,N_1165,N_1276);
xor U1743 (N_1743,N_1382,N_1389);
nor U1744 (N_1744,N_1187,N_1131);
xor U1745 (N_1745,N_1024,N_1434);
and U1746 (N_1746,N_1440,N_1127);
and U1747 (N_1747,N_1000,N_1473);
and U1748 (N_1748,N_1272,N_1391);
or U1749 (N_1749,N_1087,N_1025);
and U1750 (N_1750,N_1016,N_1159);
nand U1751 (N_1751,N_1479,N_1441);
or U1752 (N_1752,N_1090,N_1481);
nor U1753 (N_1753,N_1391,N_1042);
xor U1754 (N_1754,N_1411,N_1161);
or U1755 (N_1755,N_1387,N_1210);
and U1756 (N_1756,N_1355,N_1397);
nor U1757 (N_1757,N_1403,N_1332);
nand U1758 (N_1758,N_1269,N_1146);
and U1759 (N_1759,N_1237,N_1023);
nand U1760 (N_1760,N_1191,N_1123);
and U1761 (N_1761,N_1177,N_1278);
xnor U1762 (N_1762,N_1485,N_1007);
xor U1763 (N_1763,N_1488,N_1058);
or U1764 (N_1764,N_1251,N_1268);
or U1765 (N_1765,N_1028,N_1050);
nor U1766 (N_1766,N_1189,N_1165);
xor U1767 (N_1767,N_1364,N_1116);
xor U1768 (N_1768,N_1448,N_1152);
and U1769 (N_1769,N_1408,N_1410);
and U1770 (N_1770,N_1214,N_1451);
nand U1771 (N_1771,N_1166,N_1490);
nand U1772 (N_1772,N_1033,N_1221);
or U1773 (N_1773,N_1355,N_1179);
nor U1774 (N_1774,N_1381,N_1351);
nand U1775 (N_1775,N_1050,N_1072);
nor U1776 (N_1776,N_1222,N_1254);
or U1777 (N_1777,N_1135,N_1372);
or U1778 (N_1778,N_1295,N_1338);
or U1779 (N_1779,N_1433,N_1495);
nand U1780 (N_1780,N_1347,N_1274);
and U1781 (N_1781,N_1326,N_1060);
xnor U1782 (N_1782,N_1166,N_1468);
or U1783 (N_1783,N_1477,N_1221);
and U1784 (N_1784,N_1360,N_1059);
nand U1785 (N_1785,N_1325,N_1062);
nor U1786 (N_1786,N_1336,N_1046);
or U1787 (N_1787,N_1388,N_1277);
or U1788 (N_1788,N_1360,N_1270);
and U1789 (N_1789,N_1047,N_1285);
xnor U1790 (N_1790,N_1060,N_1335);
or U1791 (N_1791,N_1031,N_1334);
and U1792 (N_1792,N_1116,N_1290);
nand U1793 (N_1793,N_1022,N_1342);
nor U1794 (N_1794,N_1104,N_1368);
nor U1795 (N_1795,N_1394,N_1246);
nand U1796 (N_1796,N_1472,N_1192);
and U1797 (N_1797,N_1348,N_1415);
and U1798 (N_1798,N_1311,N_1449);
nand U1799 (N_1799,N_1136,N_1143);
nor U1800 (N_1800,N_1447,N_1064);
nand U1801 (N_1801,N_1202,N_1488);
xnor U1802 (N_1802,N_1028,N_1196);
or U1803 (N_1803,N_1045,N_1196);
or U1804 (N_1804,N_1030,N_1450);
xnor U1805 (N_1805,N_1025,N_1206);
and U1806 (N_1806,N_1129,N_1227);
nand U1807 (N_1807,N_1224,N_1201);
nor U1808 (N_1808,N_1471,N_1355);
and U1809 (N_1809,N_1182,N_1005);
nor U1810 (N_1810,N_1137,N_1451);
and U1811 (N_1811,N_1036,N_1401);
and U1812 (N_1812,N_1491,N_1262);
xor U1813 (N_1813,N_1321,N_1034);
nor U1814 (N_1814,N_1367,N_1089);
nor U1815 (N_1815,N_1479,N_1440);
and U1816 (N_1816,N_1003,N_1023);
or U1817 (N_1817,N_1399,N_1441);
nor U1818 (N_1818,N_1262,N_1103);
nand U1819 (N_1819,N_1340,N_1279);
nor U1820 (N_1820,N_1351,N_1094);
nor U1821 (N_1821,N_1184,N_1199);
nand U1822 (N_1822,N_1275,N_1102);
nand U1823 (N_1823,N_1452,N_1066);
or U1824 (N_1824,N_1453,N_1280);
or U1825 (N_1825,N_1319,N_1157);
xor U1826 (N_1826,N_1426,N_1185);
nor U1827 (N_1827,N_1378,N_1485);
nor U1828 (N_1828,N_1353,N_1086);
nor U1829 (N_1829,N_1339,N_1088);
and U1830 (N_1830,N_1174,N_1215);
or U1831 (N_1831,N_1129,N_1290);
xor U1832 (N_1832,N_1140,N_1109);
nand U1833 (N_1833,N_1389,N_1123);
nor U1834 (N_1834,N_1123,N_1462);
nand U1835 (N_1835,N_1252,N_1132);
and U1836 (N_1836,N_1475,N_1226);
or U1837 (N_1837,N_1298,N_1444);
or U1838 (N_1838,N_1039,N_1351);
nand U1839 (N_1839,N_1425,N_1073);
and U1840 (N_1840,N_1492,N_1024);
nor U1841 (N_1841,N_1129,N_1045);
nor U1842 (N_1842,N_1306,N_1401);
or U1843 (N_1843,N_1244,N_1353);
nand U1844 (N_1844,N_1416,N_1341);
nor U1845 (N_1845,N_1033,N_1015);
and U1846 (N_1846,N_1091,N_1286);
nor U1847 (N_1847,N_1261,N_1068);
nand U1848 (N_1848,N_1084,N_1275);
and U1849 (N_1849,N_1200,N_1161);
and U1850 (N_1850,N_1034,N_1134);
nand U1851 (N_1851,N_1410,N_1190);
or U1852 (N_1852,N_1078,N_1205);
or U1853 (N_1853,N_1377,N_1129);
or U1854 (N_1854,N_1433,N_1041);
nand U1855 (N_1855,N_1208,N_1160);
nand U1856 (N_1856,N_1078,N_1340);
nand U1857 (N_1857,N_1062,N_1272);
or U1858 (N_1858,N_1334,N_1147);
nor U1859 (N_1859,N_1124,N_1170);
or U1860 (N_1860,N_1495,N_1082);
nor U1861 (N_1861,N_1496,N_1423);
nor U1862 (N_1862,N_1341,N_1268);
nor U1863 (N_1863,N_1177,N_1204);
nand U1864 (N_1864,N_1077,N_1496);
and U1865 (N_1865,N_1374,N_1081);
or U1866 (N_1866,N_1484,N_1140);
nand U1867 (N_1867,N_1019,N_1452);
nand U1868 (N_1868,N_1102,N_1098);
or U1869 (N_1869,N_1015,N_1214);
or U1870 (N_1870,N_1142,N_1212);
and U1871 (N_1871,N_1274,N_1394);
xor U1872 (N_1872,N_1170,N_1122);
and U1873 (N_1873,N_1415,N_1256);
or U1874 (N_1874,N_1337,N_1294);
nand U1875 (N_1875,N_1265,N_1084);
or U1876 (N_1876,N_1064,N_1021);
nor U1877 (N_1877,N_1170,N_1393);
or U1878 (N_1878,N_1352,N_1117);
nand U1879 (N_1879,N_1359,N_1465);
nor U1880 (N_1880,N_1255,N_1379);
or U1881 (N_1881,N_1000,N_1188);
xor U1882 (N_1882,N_1379,N_1161);
and U1883 (N_1883,N_1043,N_1419);
nor U1884 (N_1884,N_1046,N_1018);
nor U1885 (N_1885,N_1011,N_1331);
nand U1886 (N_1886,N_1428,N_1340);
and U1887 (N_1887,N_1222,N_1250);
and U1888 (N_1888,N_1040,N_1216);
nand U1889 (N_1889,N_1184,N_1200);
nor U1890 (N_1890,N_1391,N_1053);
or U1891 (N_1891,N_1398,N_1112);
or U1892 (N_1892,N_1232,N_1381);
and U1893 (N_1893,N_1411,N_1239);
nand U1894 (N_1894,N_1316,N_1402);
nand U1895 (N_1895,N_1487,N_1481);
nand U1896 (N_1896,N_1013,N_1263);
and U1897 (N_1897,N_1423,N_1140);
or U1898 (N_1898,N_1281,N_1326);
nand U1899 (N_1899,N_1274,N_1471);
and U1900 (N_1900,N_1021,N_1132);
nand U1901 (N_1901,N_1063,N_1464);
nor U1902 (N_1902,N_1138,N_1371);
nand U1903 (N_1903,N_1477,N_1437);
xnor U1904 (N_1904,N_1074,N_1184);
nor U1905 (N_1905,N_1238,N_1471);
xnor U1906 (N_1906,N_1220,N_1355);
and U1907 (N_1907,N_1396,N_1365);
or U1908 (N_1908,N_1083,N_1412);
and U1909 (N_1909,N_1427,N_1105);
nor U1910 (N_1910,N_1176,N_1017);
nand U1911 (N_1911,N_1320,N_1094);
and U1912 (N_1912,N_1080,N_1103);
nor U1913 (N_1913,N_1127,N_1128);
or U1914 (N_1914,N_1258,N_1157);
xor U1915 (N_1915,N_1445,N_1077);
nor U1916 (N_1916,N_1242,N_1317);
xor U1917 (N_1917,N_1337,N_1453);
nor U1918 (N_1918,N_1412,N_1187);
nand U1919 (N_1919,N_1223,N_1311);
or U1920 (N_1920,N_1135,N_1023);
or U1921 (N_1921,N_1431,N_1165);
and U1922 (N_1922,N_1150,N_1166);
and U1923 (N_1923,N_1346,N_1254);
and U1924 (N_1924,N_1471,N_1117);
nor U1925 (N_1925,N_1112,N_1260);
and U1926 (N_1926,N_1230,N_1198);
and U1927 (N_1927,N_1227,N_1384);
nor U1928 (N_1928,N_1244,N_1174);
nand U1929 (N_1929,N_1448,N_1366);
nor U1930 (N_1930,N_1145,N_1212);
xor U1931 (N_1931,N_1431,N_1483);
or U1932 (N_1932,N_1452,N_1429);
nand U1933 (N_1933,N_1301,N_1395);
nand U1934 (N_1934,N_1205,N_1443);
or U1935 (N_1935,N_1122,N_1487);
and U1936 (N_1936,N_1478,N_1316);
or U1937 (N_1937,N_1274,N_1033);
xnor U1938 (N_1938,N_1034,N_1124);
and U1939 (N_1939,N_1365,N_1338);
or U1940 (N_1940,N_1339,N_1015);
nand U1941 (N_1941,N_1298,N_1050);
nand U1942 (N_1942,N_1152,N_1169);
and U1943 (N_1943,N_1125,N_1054);
and U1944 (N_1944,N_1439,N_1485);
or U1945 (N_1945,N_1059,N_1323);
nand U1946 (N_1946,N_1463,N_1489);
or U1947 (N_1947,N_1335,N_1475);
or U1948 (N_1948,N_1198,N_1118);
and U1949 (N_1949,N_1096,N_1321);
nor U1950 (N_1950,N_1446,N_1428);
nor U1951 (N_1951,N_1136,N_1096);
nand U1952 (N_1952,N_1210,N_1081);
or U1953 (N_1953,N_1322,N_1113);
or U1954 (N_1954,N_1274,N_1193);
nand U1955 (N_1955,N_1420,N_1346);
nand U1956 (N_1956,N_1203,N_1093);
nor U1957 (N_1957,N_1131,N_1211);
nor U1958 (N_1958,N_1408,N_1161);
nand U1959 (N_1959,N_1216,N_1399);
nor U1960 (N_1960,N_1159,N_1420);
or U1961 (N_1961,N_1141,N_1090);
or U1962 (N_1962,N_1173,N_1382);
or U1963 (N_1963,N_1132,N_1454);
and U1964 (N_1964,N_1257,N_1043);
nor U1965 (N_1965,N_1486,N_1114);
or U1966 (N_1966,N_1170,N_1279);
nor U1967 (N_1967,N_1397,N_1249);
nand U1968 (N_1968,N_1303,N_1048);
nor U1969 (N_1969,N_1123,N_1042);
nor U1970 (N_1970,N_1494,N_1257);
nand U1971 (N_1971,N_1356,N_1174);
and U1972 (N_1972,N_1093,N_1498);
or U1973 (N_1973,N_1035,N_1122);
and U1974 (N_1974,N_1261,N_1459);
or U1975 (N_1975,N_1069,N_1158);
xnor U1976 (N_1976,N_1095,N_1495);
nand U1977 (N_1977,N_1111,N_1134);
or U1978 (N_1978,N_1002,N_1089);
nor U1979 (N_1979,N_1362,N_1017);
or U1980 (N_1980,N_1409,N_1410);
xor U1981 (N_1981,N_1160,N_1090);
or U1982 (N_1982,N_1488,N_1095);
or U1983 (N_1983,N_1184,N_1233);
nand U1984 (N_1984,N_1380,N_1489);
nand U1985 (N_1985,N_1449,N_1091);
or U1986 (N_1986,N_1327,N_1259);
nand U1987 (N_1987,N_1053,N_1427);
xor U1988 (N_1988,N_1042,N_1407);
nand U1989 (N_1989,N_1113,N_1315);
and U1990 (N_1990,N_1233,N_1059);
and U1991 (N_1991,N_1113,N_1298);
and U1992 (N_1992,N_1463,N_1495);
nor U1993 (N_1993,N_1064,N_1095);
or U1994 (N_1994,N_1486,N_1379);
or U1995 (N_1995,N_1432,N_1419);
nand U1996 (N_1996,N_1059,N_1372);
or U1997 (N_1997,N_1096,N_1338);
or U1998 (N_1998,N_1157,N_1391);
and U1999 (N_1999,N_1462,N_1277);
nor U2000 (N_2000,N_1805,N_1524);
xor U2001 (N_2001,N_1967,N_1530);
nand U2002 (N_2002,N_1953,N_1681);
nor U2003 (N_2003,N_1818,N_1964);
nand U2004 (N_2004,N_1774,N_1770);
nand U2005 (N_2005,N_1769,N_1892);
or U2006 (N_2006,N_1725,N_1752);
or U2007 (N_2007,N_1811,N_1788);
nand U2008 (N_2008,N_1686,N_1763);
and U2009 (N_2009,N_1871,N_1834);
or U2010 (N_2010,N_1866,N_1697);
or U2011 (N_2011,N_1636,N_1747);
or U2012 (N_2012,N_1873,N_1927);
xor U2013 (N_2013,N_1813,N_1824);
nand U2014 (N_2014,N_1931,N_1629);
or U2015 (N_2015,N_1812,N_1921);
nand U2016 (N_2016,N_1977,N_1819);
or U2017 (N_2017,N_1573,N_1593);
nor U2018 (N_2018,N_1665,N_1878);
nor U2019 (N_2019,N_1862,N_1694);
xor U2020 (N_2020,N_1531,N_1858);
nor U2021 (N_2021,N_1876,N_1946);
nand U2022 (N_2022,N_1553,N_1614);
nor U2023 (N_2023,N_1500,N_1548);
xor U2024 (N_2024,N_1623,N_1900);
nand U2025 (N_2025,N_1962,N_1516);
nand U2026 (N_2026,N_1708,N_1838);
nor U2027 (N_2027,N_1569,N_1835);
nand U2028 (N_2028,N_1807,N_1670);
nor U2029 (N_2029,N_1658,N_1793);
nand U2030 (N_2030,N_1816,N_1800);
nand U2031 (N_2031,N_1933,N_1571);
and U2032 (N_2032,N_1863,N_1735);
or U2033 (N_2033,N_1579,N_1611);
and U2034 (N_2034,N_1621,N_1523);
nand U2035 (N_2035,N_1722,N_1625);
and U2036 (N_2036,N_1520,N_1856);
or U2037 (N_2037,N_1954,N_1973);
xor U2038 (N_2038,N_1705,N_1975);
or U2039 (N_2039,N_1837,N_1702);
and U2040 (N_2040,N_1624,N_1679);
and U2041 (N_2041,N_1791,N_1955);
or U2042 (N_2042,N_1581,N_1545);
or U2043 (N_2043,N_1675,N_1957);
and U2044 (N_2044,N_1560,N_1820);
and U2045 (N_2045,N_1910,N_1751);
nor U2046 (N_2046,N_1854,N_1959);
nor U2047 (N_2047,N_1999,N_1519);
or U2048 (N_2048,N_1794,N_1594);
xor U2049 (N_2049,N_1533,N_1896);
and U2050 (N_2050,N_1550,N_1653);
nand U2051 (N_2051,N_1993,N_1648);
and U2052 (N_2052,N_1626,N_1612);
or U2053 (N_2053,N_1916,N_1797);
nand U2054 (N_2054,N_1638,N_1828);
nand U2055 (N_2055,N_1897,N_1902);
nor U2056 (N_2056,N_1595,N_1898);
nor U2057 (N_2057,N_1689,N_1664);
nor U2058 (N_2058,N_1984,N_1552);
and U2059 (N_2059,N_1567,N_1982);
or U2060 (N_2060,N_1729,N_1660);
nand U2061 (N_2061,N_1591,N_1889);
and U2062 (N_2062,N_1724,N_1741);
nand U2063 (N_2063,N_1577,N_1869);
nor U2064 (N_2064,N_1960,N_1740);
nor U2065 (N_2065,N_1685,N_1888);
nand U2066 (N_2066,N_1965,N_1756);
nand U2067 (N_2067,N_1733,N_1590);
and U2068 (N_2068,N_1864,N_1908);
nor U2069 (N_2069,N_1559,N_1616);
nor U2070 (N_2070,N_1619,N_1654);
and U2071 (N_2071,N_1809,N_1842);
or U2072 (N_2072,N_1668,N_1720);
nor U2073 (N_2073,N_1731,N_1997);
nor U2074 (N_2074,N_1671,N_1572);
or U2075 (N_2075,N_1852,N_1502);
nand U2076 (N_2076,N_1586,N_1948);
or U2077 (N_2077,N_1757,N_1682);
or U2078 (N_2078,N_1749,N_1745);
nand U2079 (N_2079,N_1707,N_1996);
nand U2080 (N_2080,N_1564,N_1539);
and U2081 (N_2081,N_1817,N_1860);
nand U2082 (N_2082,N_1985,N_1883);
nand U2083 (N_2083,N_1678,N_1599);
nand U2084 (N_2084,N_1990,N_1775);
and U2085 (N_2085,N_1582,N_1557);
nor U2086 (N_2086,N_1727,N_1511);
nand U2087 (N_2087,N_1848,N_1949);
or U2088 (N_2088,N_1766,N_1806);
and U2089 (N_2089,N_1786,N_1692);
nand U2090 (N_2090,N_1872,N_1779);
nand U2091 (N_2091,N_1919,N_1696);
or U2092 (N_2092,N_1804,N_1723);
or U2093 (N_2093,N_1980,N_1526);
or U2094 (N_2094,N_1836,N_1887);
or U2095 (N_2095,N_1988,N_1978);
and U2096 (N_2096,N_1717,N_1968);
or U2097 (N_2097,N_1737,N_1995);
xor U2098 (N_2098,N_1913,N_1651);
nand U2099 (N_2099,N_1542,N_1998);
nor U2100 (N_2100,N_1632,N_1584);
or U2101 (N_2101,N_1983,N_1777);
and U2102 (N_2102,N_1547,N_1782);
nand U2103 (N_2103,N_1952,N_1754);
nor U2104 (N_2104,N_1849,N_1652);
xnor U2105 (N_2105,N_1903,N_1576);
or U2106 (N_2106,N_1534,N_1565);
nand U2107 (N_2107,N_1556,N_1918);
xnor U2108 (N_2108,N_1639,N_1691);
or U2109 (N_2109,N_1781,N_1503);
nor U2110 (N_2110,N_1840,N_1615);
nand U2111 (N_2111,N_1603,N_1914);
nand U2112 (N_2112,N_1522,N_1936);
or U2113 (N_2113,N_1833,N_1851);
or U2114 (N_2114,N_1891,N_1755);
xor U2115 (N_2115,N_1886,N_1767);
or U2116 (N_2116,N_1551,N_1801);
nand U2117 (N_2117,N_1610,N_1588);
nor U2118 (N_2118,N_1714,N_1938);
or U2119 (N_2119,N_1939,N_1620);
nand U2120 (N_2120,N_1792,N_1920);
nor U2121 (N_2121,N_1676,N_1969);
xor U2122 (N_2122,N_1554,N_1905);
or U2123 (N_2123,N_1855,N_1738);
xor U2124 (N_2124,N_1841,N_1950);
nand U2125 (N_2125,N_1808,N_1909);
nand U2126 (N_2126,N_1924,N_1859);
and U2127 (N_2127,N_1814,N_1570);
xor U2128 (N_2128,N_1881,N_1963);
nor U2129 (N_2129,N_1666,N_1945);
and U2130 (N_2130,N_1608,N_1901);
nor U2131 (N_2131,N_1944,N_1823);
and U2132 (N_2132,N_1613,N_1844);
and U2133 (N_2133,N_1875,N_1732);
nor U2134 (N_2134,N_1773,N_1958);
xnor U2135 (N_2135,N_1602,N_1701);
nand U2136 (N_2136,N_1663,N_1555);
and U2137 (N_2137,N_1687,N_1719);
or U2138 (N_2138,N_1537,N_1513);
and U2139 (N_2139,N_1600,N_1677);
nor U2140 (N_2140,N_1674,N_1865);
and U2141 (N_2141,N_1890,N_1821);
or U2142 (N_2142,N_1693,N_1704);
xor U2143 (N_2143,N_1605,N_1879);
and U2144 (N_2144,N_1847,N_1618);
nor U2145 (N_2145,N_1825,N_1987);
or U2146 (N_2146,N_1930,N_1885);
nand U2147 (N_2147,N_1877,N_1966);
and U2148 (N_2148,N_1748,N_1730);
or U2149 (N_2149,N_1937,N_1580);
and U2150 (N_2150,N_1597,N_1641);
nand U2151 (N_2151,N_1776,N_1672);
nand U2152 (N_2152,N_1830,N_1992);
nand U2153 (N_2153,N_1634,N_1647);
nand U2154 (N_2154,N_1839,N_1961);
and U2155 (N_2155,N_1540,N_1923);
and U2156 (N_2156,N_1867,N_1870);
and U2157 (N_2157,N_1649,N_1575);
xnor U2158 (N_2158,N_1832,N_1758);
nor U2159 (N_2159,N_1607,N_1562);
and U2160 (N_2160,N_1606,N_1785);
and U2161 (N_2161,N_1508,N_1906);
or U2162 (N_2162,N_1932,N_1661);
xnor U2163 (N_2163,N_1566,N_1911);
nor U2164 (N_2164,N_1994,N_1868);
nand U2165 (N_2165,N_1544,N_1831);
nand U2166 (N_2166,N_1667,N_1541);
or U2167 (N_2167,N_1784,N_1645);
and U2168 (N_2168,N_1922,N_1912);
xnor U2169 (N_2169,N_1631,N_1578);
or U2170 (N_2170,N_1587,N_1622);
and U2171 (N_2171,N_1635,N_1796);
or U2172 (N_2172,N_1604,N_1827);
and U2173 (N_2173,N_1907,N_1505);
or U2174 (N_2174,N_1771,N_1947);
or U2175 (N_2175,N_1713,N_1709);
xor U2176 (N_2176,N_1627,N_1650);
nand U2177 (N_2177,N_1787,N_1795);
or U2178 (N_2178,N_1934,N_1617);
xor U2179 (N_2179,N_1940,N_1515);
nor U2180 (N_2180,N_1643,N_1521);
nand U2181 (N_2181,N_1517,N_1514);
or U2182 (N_2182,N_1558,N_1899);
nor U2183 (N_2183,N_1504,N_1715);
and U2184 (N_2184,N_1549,N_1942);
nor U2185 (N_2185,N_1986,N_1706);
or U2186 (N_2186,N_1929,N_1759);
or U2187 (N_2187,N_1956,N_1857);
or U2188 (N_2188,N_1683,N_1972);
nand U2189 (N_2189,N_1935,N_1662);
nor U2190 (N_2190,N_1742,N_1532);
or U2191 (N_2191,N_1734,N_1861);
nand U2192 (N_2192,N_1989,N_1589);
nor U2193 (N_2193,N_1853,N_1790);
and U2194 (N_2194,N_1943,N_1760);
nor U2195 (N_2195,N_1761,N_1925);
or U2196 (N_2196,N_1543,N_1538);
nand U2197 (N_2197,N_1874,N_1970);
and U2198 (N_2198,N_1974,N_1768);
and U2199 (N_2199,N_1845,N_1574);
and U2200 (N_2200,N_1762,N_1506);
or U2201 (N_2201,N_1951,N_1765);
nand U2202 (N_2202,N_1716,N_1598);
or U2203 (N_2203,N_1633,N_1810);
and U2204 (N_2204,N_1640,N_1721);
and U2205 (N_2205,N_1846,N_1739);
nor U2206 (N_2206,N_1510,N_1815);
and U2207 (N_2207,N_1642,N_1711);
and U2208 (N_2208,N_1829,N_1525);
nor U2209 (N_2209,N_1802,N_1695);
or U2210 (N_2210,N_1981,N_1592);
or U2211 (N_2211,N_1798,N_1698);
xnor U2212 (N_2212,N_1882,N_1736);
nand U2213 (N_2213,N_1703,N_1991);
or U2214 (N_2214,N_1928,N_1710);
nor U2215 (N_2215,N_1780,N_1843);
nor U2216 (N_2216,N_1917,N_1583);
and U2217 (N_2217,N_1673,N_1601);
and U2218 (N_2218,N_1684,N_1563);
or U2219 (N_2219,N_1529,N_1743);
xor U2220 (N_2220,N_1528,N_1789);
or U2221 (N_2221,N_1728,N_1655);
xor U2222 (N_2222,N_1536,N_1753);
xor U2223 (N_2223,N_1726,N_1971);
or U2224 (N_2224,N_1746,N_1688);
nor U2225 (N_2225,N_1535,N_1630);
nand U2226 (N_2226,N_1657,N_1744);
and U2227 (N_2227,N_1764,N_1976);
nand U2228 (N_2228,N_1659,N_1656);
nor U2229 (N_2229,N_1637,N_1568);
or U2230 (N_2230,N_1527,N_1690);
xor U2231 (N_2231,N_1926,N_1904);
or U2232 (N_2232,N_1718,N_1915);
xnor U2233 (N_2233,N_1880,N_1822);
xor U2234 (N_2234,N_1507,N_1941);
and U2235 (N_2235,N_1509,N_1700);
or U2236 (N_2236,N_1596,N_1778);
and U2237 (N_2237,N_1585,N_1609);
nor U2238 (N_2238,N_1750,N_1850);
nor U2239 (N_2239,N_1680,N_1893);
and U2240 (N_2240,N_1501,N_1646);
nor U2241 (N_2241,N_1561,N_1699);
nand U2242 (N_2242,N_1518,N_1895);
or U2243 (N_2243,N_1712,N_1772);
xor U2244 (N_2244,N_1512,N_1669);
nand U2245 (N_2245,N_1803,N_1546);
xor U2246 (N_2246,N_1894,N_1783);
and U2247 (N_2247,N_1979,N_1799);
nand U2248 (N_2248,N_1628,N_1826);
nor U2249 (N_2249,N_1644,N_1884);
nor U2250 (N_2250,N_1804,N_1910);
or U2251 (N_2251,N_1716,N_1854);
or U2252 (N_2252,N_1849,N_1713);
or U2253 (N_2253,N_1878,N_1812);
nand U2254 (N_2254,N_1525,N_1564);
or U2255 (N_2255,N_1849,N_1955);
or U2256 (N_2256,N_1740,N_1642);
nand U2257 (N_2257,N_1738,N_1873);
nor U2258 (N_2258,N_1957,N_1996);
or U2259 (N_2259,N_1775,N_1859);
nand U2260 (N_2260,N_1733,N_1769);
nand U2261 (N_2261,N_1997,N_1671);
xnor U2262 (N_2262,N_1973,N_1608);
nand U2263 (N_2263,N_1742,N_1939);
or U2264 (N_2264,N_1846,N_1763);
or U2265 (N_2265,N_1834,N_1886);
nand U2266 (N_2266,N_1683,N_1728);
nor U2267 (N_2267,N_1724,N_1508);
nand U2268 (N_2268,N_1539,N_1891);
and U2269 (N_2269,N_1525,N_1681);
xnor U2270 (N_2270,N_1875,N_1670);
nand U2271 (N_2271,N_1650,N_1812);
or U2272 (N_2272,N_1749,N_1775);
and U2273 (N_2273,N_1979,N_1817);
nand U2274 (N_2274,N_1721,N_1538);
and U2275 (N_2275,N_1888,N_1518);
nand U2276 (N_2276,N_1690,N_1810);
or U2277 (N_2277,N_1541,N_1827);
nand U2278 (N_2278,N_1546,N_1705);
nor U2279 (N_2279,N_1575,N_1885);
and U2280 (N_2280,N_1579,N_1767);
nor U2281 (N_2281,N_1515,N_1523);
nand U2282 (N_2282,N_1815,N_1593);
nor U2283 (N_2283,N_1538,N_1638);
or U2284 (N_2284,N_1692,N_1777);
xnor U2285 (N_2285,N_1980,N_1951);
or U2286 (N_2286,N_1622,N_1703);
or U2287 (N_2287,N_1607,N_1516);
and U2288 (N_2288,N_1982,N_1557);
or U2289 (N_2289,N_1751,N_1879);
nor U2290 (N_2290,N_1935,N_1615);
nor U2291 (N_2291,N_1732,N_1551);
xor U2292 (N_2292,N_1954,N_1995);
or U2293 (N_2293,N_1753,N_1613);
and U2294 (N_2294,N_1958,N_1614);
or U2295 (N_2295,N_1521,N_1787);
nor U2296 (N_2296,N_1812,N_1877);
nor U2297 (N_2297,N_1806,N_1904);
or U2298 (N_2298,N_1612,N_1504);
or U2299 (N_2299,N_1783,N_1502);
or U2300 (N_2300,N_1794,N_1931);
or U2301 (N_2301,N_1620,N_1821);
or U2302 (N_2302,N_1696,N_1855);
and U2303 (N_2303,N_1545,N_1922);
and U2304 (N_2304,N_1979,N_1822);
nor U2305 (N_2305,N_1641,N_1738);
xnor U2306 (N_2306,N_1996,N_1788);
nor U2307 (N_2307,N_1828,N_1928);
xor U2308 (N_2308,N_1909,N_1899);
xnor U2309 (N_2309,N_1889,N_1648);
and U2310 (N_2310,N_1723,N_1666);
and U2311 (N_2311,N_1524,N_1793);
or U2312 (N_2312,N_1717,N_1952);
or U2313 (N_2313,N_1767,N_1681);
or U2314 (N_2314,N_1691,N_1919);
or U2315 (N_2315,N_1911,N_1551);
or U2316 (N_2316,N_1691,N_1596);
and U2317 (N_2317,N_1946,N_1817);
and U2318 (N_2318,N_1602,N_1725);
nand U2319 (N_2319,N_1904,N_1788);
or U2320 (N_2320,N_1994,N_1854);
nand U2321 (N_2321,N_1606,N_1882);
nor U2322 (N_2322,N_1971,N_1966);
or U2323 (N_2323,N_1845,N_1552);
nor U2324 (N_2324,N_1742,N_1935);
nand U2325 (N_2325,N_1666,N_1642);
nor U2326 (N_2326,N_1718,N_1857);
xnor U2327 (N_2327,N_1626,N_1778);
nor U2328 (N_2328,N_1726,N_1654);
xnor U2329 (N_2329,N_1746,N_1948);
and U2330 (N_2330,N_1963,N_1724);
or U2331 (N_2331,N_1600,N_1758);
or U2332 (N_2332,N_1506,N_1837);
or U2333 (N_2333,N_1733,N_1977);
xor U2334 (N_2334,N_1597,N_1708);
nor U2335 (N_2335,N_1943,N_1544);
nor U2336 (N_2336,N_1588,N_1612);
nand U2337 (N_2337,N_1621,N_1733);
nand U2338 (N_2338,N_1508,N_1813);
nand U2339 (N_2339,N_1543,N_1681);
nand U2340 (N_2340,N_1888,N_1791);
and U2341 (N_2341,N_1502,N_1907);
nand U2342 (N_2342,N_1986,N_1588);
or U2343 (N_2343,N_1589,N_1714);
nand U2344 (N_2344,N_1523,N_1576);
nand U2345 (N_2345,N_1821,N_1835);
or U2346 (N_2346,N_1744,N_1686);
or U2347 (N_2347,N_1835,N_1705);
nand U2348 (N_2348,N_1619,N_1918);
and U2349 (N_2349,N_1674,N_1930);
and U2350 (N_2350,N_1969,N_1514);
nor U2351 (N_2351,N_1653,N_1529);
or U2352 (N_2352,N_1743,N_1970);
and U2353 (N_2353,N_1901,N_1656);
or U2354 (N_2354,N_1610,N_1682);
nor U2355 (N_2355,N_1688,N_1676);
nor U2356 (N_2356,N_1503,N_1936);
or U2357 (N_2357,N_1703,N_1735);
xnor U2358 (N_2358,N_1657,N_1608);
or U2359 (N_2359,N_1929,N_1619);
and U2360 (N_2360,N_1946,N_1575);
nand U2361 (N_2361,N_1853,N_1910);
xor U2362 (N_2362,N_1969,N_1565);
nand U2363 (N_2363,N_1541,N_1747);
nor U2364 (N_2364,N_1526,N_1559);
nand U2365 (N_2365,N_1665,N_1545);
and U2366 (N_2366,N_1936,N_1794);
or U2367 (N_2367,N_1814,N_1864);
or U2368 (N_2368,N_1622,N_1629);
nor U2369 (N_2369,N_1558,N_1702);
nand U2370 (N_2370,N_1637,N_1837);
nor U2371 (N_2371,N_1587,N_1542);
nand U2372 (N_2372,N_1850,N_1790);
and U2373 (N_2373,N_1938,N_1993);
and U2374 (N_2374,N_1619,N_1580);
nor U2375 (N_2375,N_1826,N_1771);
nand U2376 (N_2376,N_1564,N_1946);
nand U2377 (N_2377,N_1864,N_1551);
and U2378 (N_2378,N_1702,N_1697);
nand U2379 (N_2379,N_1979,N_1633);
nand U2380 (N_2380,N_1871,N_1835);
and U2381 (N_2381,N_1856,N_1757);
nor U2382 (N_2382,N_1838,N_1861);
and U2383 (N_2383,N_1543,N_1670);
nand U2384 (N_2384,N_1656,N_1609);
or U2385 (N_2385,N_1610,N_1957);
and U2386 (N_2386,N_1648,N_1660);
and U2387 (N_2387,N_1897,N_1933);
nand U2388 (N_2388,N_1541,N_1670);
or U2389 (N_2389,N_1536,N_1576);
nand U2390 (N_2390,N_1640,N_1778);
nor U2391 (N_2391,N_1863,N_1574);
nor U2392 (N_2392,N_1808,N_1783);
and U2393 (N_2393,N_1989,N_1697);
nand U2394 (N_2394,N_1666,N_1937);
nor U2395 (N_2395,N_1651,N_1806);
nor U2396 (N_2396,N_1820,N_1953);
or U2397 (N_2397,N_1672,N_1869);
and U2398 (N_2398,N_1799,N_1922);
and U2399 (N_2399,N_1821,N_1613);
nand U2400 (N_2400,N_1779,N_1975);
nand U2401 (N_2401,N_1630,N_1678);
or U2402 (N_2402,N_1608,N_1967);
nor U2403 (N_2403,N_1887,N_1544);
or U2404 (N_2404,N_1907,N_1809);
nand U2405 (N_2405,N_1614,N_1823);
and U2406 (N_2406,N_1660,N_1670);
nor U2407 (N_2407,N_1857,N_1984);
nand U2408 (N_2408,N_1676,N_1637);
nor U2409 (N_2409,N_1645,N_1787);
and U2410 (N_2410,N_1531,N_1764);
nor U2411 (N_2411,N_1656,N_1965);
or U2412 (N_2412,N_1882,N_1775);
and U2413 (N_2413,N_1875,N_1545);
nand U2414 (N_2414,N_1573,N_1760);
nand U2415 (N_2415,N_1711,N_1597);
nand U2416 (N_2416,N_1938,N_1715);
or U2417 (N_2417,N_1736,N_1737);
or U2418 (N_2418,N_1722,N_1715);
xnor U2419 (N_2419,N_1618,N_1968);
xnor U2420 (N_2420,N_1547,N_1901);
and U2421 (N_2421,N_1947,N_1574);
or U2422 (N_2422,N_1822,N_1718);
or U2423 (N_2423,N_1811,N_1500);
nand U2424 (N_2424,N_1806,N_1625);
nor U2425 (N_2425,N_1868,N_1835);
or U2426 (N_2426,N_1505,N_1710);
nand U2427 (N_2427,N_1975,N_1531);
nand U2428 (N_2428,N_1860,N_1711);
xor U2429 (N_2429,N_1865,N_1806);
nor U2430 (N_2430,N_1973,N_1879);
and U2431 (N_2431,N_1807,N_1934);
nor U2432 (N_2432,N_1598,N_1712);
or U2433 (N_2433,N_1881,N_1975);
nand U2434 (N_2434,N_1648,N_1848);
or U2435 (N_2435,N_1732,N_1676);
nor U2436 (N_2436,N_1878,N_1594);
and U2437 (N_2437,N_1856,N_1582);
nor U2438 (N_2438,N_1618,N_1635);
and U2439 (N_2439,N_1810,N_1953);
nand U2440 (N_2440,N_1781,N_1521);
and U2441 (N_2441,N_1943,N_1880);
and U2442 (N_2442,N_1879,N_1913);
or U2443 (N_2443,N_1760,N_1534);
and U2444 (N_2444,N_1695,N_1932);
nand U2445 (N_2445,N_1612,N_1513);
nor U2446 (N_2446,N_1847,N_1877);
nand U2447 (N_2447,N_1610,N_1934);
nor U2448 (N_2448,N_1515,N_1652);
xnor U2449 (N_2449,N_1972,N_1588);
or U2450 (N_2450,N_1942,N_1761);
nand U2451 (N_2451,N_1940,N_1805);
or U2452 (N_2452,N_1532,N_1670);
and U2453 (N_2453,N_1509,N_1766);
or U2454 (N_2454,N_1724,N_1853);
nor U2455 (N_2455,N_1712,N_1720);
nor U2456 (N_2456,N_1929,N_1727);
or U2457 (N_2457,N_1728,N_1584);
nand U2458 (N_2458,N_1893,N_1984);
or U2459 (N_2459,N_1786,N_1854);
or U2460 (N_2460,N_1969,N_1555);
and U2461 (N_2461,N_1805,N_1907);
nor U2462 (N_2462,N_1621,N_1832);
and U2463 (N_2463,N_1924,N_1854);
and U2464 (N_2464,N_1744,N_1894);
and U2465 (N_2465,N_1743,N_1631);
and U2466 (N_2466,N_1736,N_1927);
and U2467 (N_2467,N_1645,N_1802);
nand U2468 (N_2468,N_1977,N_1582);
nor U2469 (N_2469,N_1915,N_1988);
nand U2470 (N_2470,N_1765,N_1822);
nand U2471 (N_2471,N_1560,N_1582);
nand U2472 (N_2472,N_1734,N_1922);
nor U2473 (N_2473,N_1879,N_1535);
and U2474 (N_2474,N_1973,N_1701);
xor U2475 (N_2475,N_1551,N_1754);
and U2476 (N_2476,N_1726,N_1713);
and U2477 (N_2477,N_1506,N_1913);
nor U2478 (N_2478,N_1561,N_1895);
and U2479 (N_2479,N_1772,N_1776);
nor U2480 (N_2480,N_1990,N_1654);
nand U2481 (N_2481,N_1875,N_1817);
nor U2482 (N_2482,N_1942,N_1585);
and U2483 (N_2483,N_1922,N_1913);
or U2484 (N_2484,N_1529,N_1506);
and U2485 (N_2485,N_1565,N_1829);
and U2486 (N_2486,N_1860,N_1762);
or U2487 (N_2487,N_1834,N_1738);
or U2488 (N_2488,N_1747,N_1785);
nand U2489 (N_2489,N_1698,N_1726);
nand U2490 (N_2490,N_1798,N_1935);
nand U2491 (N_2491,N_1865,N_1545);
and U2492 (N_2492,N_1713,N_1953);
xnor U2493 (N_2493,N_1616,N_1562);
nor U2494 (N_2494,N_1596,N_1573);
xnor U2495 (N_2495,N_1710,N_1943);
xor U2496 (N_2496,N_1576,N_1891);
or U2497 (N_2497,N_1534,N_1802);
nor U2498 (N_2498,N_1713,N_1826);
nor U2499 (N_2499,N_1841,N_1893);
or U2500 (N_2500,N_2059,N_2118);
or U2501 (N_2501,N_2254,N_2415);
nor U2502 (N_2502,N_2385,N_2367);
or U2503 (N_2503,N_2459,N_2463);
nor U2504 (N_2504,N_2216,N_2472);
nor U2505 (N_2505,N_2384,N_2190);
nor U2506 (N_2506,N_2184,N_2386);
nand U2507 (N_2507,N_2318,N_2012);
and U2508 (N_2508,N_2084,N_2471);
xor U2509 (N_2509,N_2414,N_2081);
xor U2510 (N_2510,N_2357,N_2293);
or U2511 (N_2511,N_2259,N_2372);
and U2512 (N_2512,N_2391,N_2202);
xnor U2513 (N_2513,N_2405,N_2133);
or U2514 (N_2514,N_2089,N_2140);
nor U2515 (N_2515,N_2148,N_2131);
nor U2516 (N_2516,N_2473,N_2319);
or U2517 (N_2517,N_2109,N_2295);
or U2518 (N_2518,N_2362,N_2365);
and U2519 (N_2519,N_2456,N_2086);
nor U2520 (N_2520,N_2182,N_2375);
nor U2521 (N_2521,N_2457,N_2045);
and U2522 (N_2522,N_2171,N_2040);
nand U2523 (N_2523,N_2031,N_2075);
or U2524 (N_2524,N_2345,N_2023);
nor U2525 (N_2525,N_2496,N_2007);
and U2526 (N_2526,N_2324,N_2066);
or U2527 (N_2527,N_2122,N_2379);
nor U2528 (N_2528,N_2433,N_2183);
nand U2529 (N_2529,N_2465,N_2177);
xor U2530 (N_2530,N_2240,N_2331);
nor U2531 (N_2531,N_2316,N_2296);
or U2532 (N_2532,N_2155,N_2169);
nor U2533 (N_2533,N_2033,N_2477);
or U2534 (N_2534,N_2020,N_2438);
and U2535 (N_2535,N_2279,N_2218);
or U2536 (N_2536,N_2154,N_2298);
nor U2537 (N_2537,N_2017,N_2111);
and U2538 (N_2538,N_2406,N_2399);
nand U2539 (N_2539,N_2490,N_2288);
nand U2540 (N_2540,N_2196,N_2371);
nand U2541 (N_2541,N_2241,N_2063);
nand U2542 (N_2542,N_2307,N_2359);
nor U2543 (N_2543,N_2201,N_2297);
and U2544 (N_2544,N_2360,N_2004);
or U2545 (N_2545,N_2139,N_2315);
or U2546 (N_2546,N_2046,N_2037);
or U2547 (N_2547,N_2132,N_2076);
nand U2548 (N_2548,N_2054,N_2071);
or U2549 (N_2549,N_2361,N_2260);
or U2550 (N_2550,N_2194,N_2016);
and U2551 (N_2551,N_2253,N_2166);
and U2552 (N_2552,N_2072,N_2058);
nor U2553 (N_2553,N_2096,N_2009);
or U2554 (N_2554,N_2080,N_2193);
nand U2555 (N_2555,N_2107,N_2393);
nand U2556 (N_2556,N_2369,N_2489);
nor U2557 (N_2557,N_2328,N_2083);
or U2558 (N_2558,N_2387,N_2018);
nand U2559 (N_2559,N_2085,N_2479);
nand U2560 (N_2560,N_2014,N_2492);
or U2561 (N_2561,N_2067,N_2181);
nand U2562 (N_2562,N_2113,N_2110);
and U2563 (N_2563,N_2255,N_2351);
and U2564 (N_2564,N_2310,N_2413);
and U2565 (N_2565,N_2127,N_2312);
nor U2566 (N_2566,N_2199,N_2238);
and U2567 (N_2567,N_2129,N_2205);
nand U2568 (N_2568,N_2325,N_2117);
nor U2569 (N_2569,N_2163,N_2236);
and U2570 (N_2570,N_2499,N_2250);
and U2571 (N_2571,N_2178,N_2374);
nor U2572 (N_2572,N_2243,N_2332);
nor U2573 (N_2573,N_2115,N_2093);
or U2574 (N_2574,N_2261,N_2130);
and U2575 (N_2575,N_2121,N_2273);
nand U2576 (N_2576,N_2207,N_2097);
and U2577 (N_2577,N_2388,N_2323);
and U2578 (N_2578,N_2334,N_2036);
nor U2579 (N_2579,N_2494,N_2431);
or U2580 (N_2580,N_2244,N_2120);
or U2581 (N_2581,N_2305,N_2398);
nand U2582 (N_2582,N_2150,N_2426);
nor U2583 (N_2583,N_2159,N_2057);
nand U2584 (N_2584,N_2348,N_2158);
and U2585 (N_2585,N_2397,N_2198);
or U2586 (N_2586,N_2137,N_2219);
xor U2587 (N_2587,N_2211,N_2002);
or U2588 (N_2588,N_2237,N_2454);
nor U2589 (N_2589,N_2247,N_2146);
nand U2590 (N_2590,N_2013,N_2252);
or U2591 (N_2591,N_2074,N_2460);
nand U2592 (N_2592,N_2000,N_2443);
nand U2593 (N_2593,N_2470,N_2149);
nand U2594 (N_2594,N_2088,N_2210);
and U2595 (N_2595,N_2336,N_2267);
nand U2596 (N_2596,N_2462,N_2466);
or U2597 (N_2597,N_2213,N_2491);
nor U2598 (N_2598,N_2095,N_2476);
nand U2599 (N_2599,N_2309,N_2100);
or U2600 (N_2600,N_2069,N_2151);
nand U2601 (N_2601,N_2223,N_2294);
and U2602 (N_2602,N_2061,N_2172);
nor U2603 (N_2603,N_2311,N_2314);
or U2604 (N_2604,N_2105,N_2440);
or U2605 (N_2605,N_2136,N_2073);
and U2606 (N_2606,N_2167,N_2390);
or U2607 (N_2607,N_2382,N_2419);
xor U2608 (N_2608,N_2200,N_2064);
or U2609 (N_2609,N_2246,N_2142);
or U2610 (N_2610,N_2153,N_2090);
xnor U2611 (N_2611,N_2432,N_2003);
and U2612 (N_2612,N_2354,N_2019);
nand U2613 (N_2613,N_2274,N_2157);
nand U2614 (N_2614,N_2444,N_2275);
nor U2615 (N_2615,N_2421,N_2481);
nor U2616 (N_2616,N_2428,N_2256);
nor U2617 (N_2617,N_2079,N_2068);
and U2618 (N_2618,N_2217,N_2168);
nor U2619 (N_2619,N_2344,N_2050);
nor U2620 (N_2620,N_2264,N_2226);
xor U2621 (N_2621,N_2497,N_2165);
and U2622 (N_2622,N_2049,N_2224);
and U2623 (N_2623,N_2436,N_2486);
nand U2624 (N_2624,N_2094,N_2484);
and U2625 (N_2625,N_2106,N_2227);
nand U2626 (N_2626,N_2333,N_2356);
nor U2627 (N_2627,N_2400,N_2292);
nor U2628 (N_2628,N_2349,N_2302);
nand U2629 (N_2629,N_2488,N_2102);
and U2630 (N_2630,N_2303,N_2478);
nor U2631 (N_2631,N_2078,N_2373);
and U2632 (N_2632,N_2425,N_2407);
nor U2633 (N_2633,N_2366,N_2383);
nor U2634 (N_2634,N_2416,N_2378);
or U2635 (N_2635,N_2412,N_2034);
nor U2636 (N_2636,N_2185,N_2268);
nand U2637 (N_2637,N_2022,N_2041);
nand U2638 (N_2638,N_2437,N_2424);
or U2639 (N_2639,N_2343,N_2204);
and U2640 (N_2640,N_2179,N_2364);
or U2641 (N_2641,N_2006,N_2266);
nor U2642 (N_2642,N_2317,N_2104);
nand U2643 (N_2643,N_2103,N_2212);
or U2644 (N_2644,N_2304,N_2475);
xnor U2645 (N_2645,N_2082,N_2152);
nor U2646 (N_2646,N_2162,N_2186);
nand U2647 (N_2647,N_2192,N_2353);
or U2648 (N_2648,N_2270,N_2376);
and U2649 (N_2649,N_2269,N_2143);
and U2650 (N_2650,N_2394,N_2234);
xnor U2651 (N_2651,N_2147,N_2164);
and U2652 (N_2652,N_2287,N_2430);
nand U2653 (N_2653,N_2188,N_2209);
xor U2654 (N_2654,N_2232,N_2215);
or U2655 (N_2655,N_2119,N_2285);
nand U2656 (N_2656,N_2469,N_2039);
nand U2657 (N_2657,N_2156,N_2480);
and U2658 (N_2658,N_2487,N_2035);
and U2659 (N_2659,N_2320,N_2145);
nand U2660 (N_2660,N_2441,N_2409);
nand U2661 (N_2661,N_2467,N_2427);
nand U2662 (N_2662,N_2498,N_2144);
xor U2663 (N_2663,N_2283,N_2429);
nor U2664 (N_2664,N_2235,N_2474);
nor U2665 (N_2665,N_2187,N_2442);
nand U2666 (N_2666,N_2423,N_2026);
nor U2667 (N_2667,N_2380,N_2308);
and U2668 (N_2668,N_2126,N_2134);
nand U2669 (N_2669,N_2338,N_2485);
nand U2670 (N_2670,N_2180,N_2214);
or U2671 (N_2671,N_2245,N_2203);
nand U2672 (N_2672,N_2249,N_2220);
xnor U2673 (N_2673,N_2321,N_2493);
xor U2674 (N_2674,N_2191,N_2322);
and U2675 (N_2675,N_2025,N_2077);
nand U2676 (N_2676,N_2233,N_2087);
and U2677 (N_2677,N_2197,N_2055);
xor U2678 (N_2678,N_2053,N_2042);
and U2679 (N_2679,N_2251,N_2173);
nor U2680 (N_2680,N_2434,N_2483);
and U2681 (N_2681,N_2482,N_2160);
and U2682 (N_2682,N_2008,N_2263);
xnor U2683 (N_2683,N_2029,N_2141);
nand U2684 (N_2684,N_2138,N_2028);
or U2685 (N_2685,N_2449,N_2352);
nand U2686 (N_2686,N_2346,N_2300);
nor U2687 (N_2687,N_2229,N_2370);
nand U2688 (N_2688,N_2340,N_2060);
nand U2689 (N_2689,N_2411,N_2044);
and U2690 (N_2690,N_2389,N_2450);
nor U2691 (N_2691,N_2281,N_2221);
nor U2692 (N_2692,N_2170,N_2306);
and U2693 (N_2693,N_2001,N_2329);
nand U2694 (N_2694,N_2402,N_2065);
nor U2695 (N_2695,N_2410,N_2447);
nor U2696 (N_2696,N_2278,N_2418);
xnor U2697 (N_2697,N_2092,N_2291);
nand U2698 (N_2698,N_2358,N_2404);
and U2699 (N_2699,N_2101,N_2038);
nand U2700 (N_2700,N_2257,N_2368);
and U2701 (N_2701,N_2056,N_2455);
or U2702 (N_2702,N_2091,N_2231);
or U2703 (N_2703,N_2286,N_2271);
or U2704 (N_2704,N_2228,N_2128);
and U2705 (N_2705,N_2052,N_2070);
and U2706 (N_2706,N_2341,N_2377);
nor U2707 (N_2707,N_2242,N_2272);
nor U2708 (N_2708,N_2299,N_2439);
or U2709 (N_2709,N_2258,N_2381);
nor U2710 (N_2710,N_2123,N_2363);
nor U2711 (N_2711,N_2024,N_2337);
nand U2712 (N_2712,N_2051,N_2448);
and U2713 (N_2713,N_2032,N_2048);
and U2714 (N_2714,N_2420,N_2021);
and U2715 (N_2715,N_2208,N_2125);
nor U2716 (N_2716,N_2284,N_2265);
nand U2717 (N_2717,N_2230,N_2047);
nor U2718 (N_2718,N_2495,N_2248);
nor U2719 (N_2719,N_2445,N_2195);
nand U2720 (N_2720,N_2010,N_2453);
or U2721 (N_2721,N_2451,N_2301);
nor U2722 (N_2722,N_2290,N_2464);
and U2723 (N_2723,N_2114,N_2262);
or U2724 (N_2724,N_2395,N_2161);
or U2725 (N_2725,N_2175,N_2350);
or U2726 (N_2726,N_2176,N_2401);
and U2727 (N_2727,N_2174,N_2396);
or U2728 (N_2728,N_2435,N_2392);
and U2729 (N_2729,N_2116,N_2043);
or U2730 (N_2730,N_2112,N_2189);
and U2731 (N_2731,N_2011,N_2124);
or U2732 (N_2732,N_2339,N_2417);
xor U2733 (N_2733,N_2452,N_2099);
and U2734 (N_2734,N_2446,N_2030);
nor U2735 (N_2735,N_2206,N_2015);
or U2736 (N_2736,N_2108,N_2225);
or U2737 (N_2737,N_2347,N_2277);
and U2738 (N_2738,N_2342,N_2355);
nand U2739 (N_2739,N_2327,N_2098);
nand U2740 (N_2740,N_2062,N_2280);
nand U2741 (N_2741,N_2422,N_2403);
or U2742 (N_2742,N_2326,N_2135);
or U2743 (N_2743,N_2282,N_2330);
or U2744 (N_2744,N_2458,N_2289);
xor U2745 (N_2745,N_2239,N_2335);
nand U2746 (N_2746,N_2222,N_2313);
and U2747 (N_2747,N_2027,N_2468);
nand U2748 (N_2748,N_2461,N_2276);
nand U2749 (N_2749,N_2408,N_2005);
nor U2750 (N_2750,N_2171,N_2213);
nand U2751 (N_2751,N_2275,N_2271);
and U2752 (N_2752,N_2109,N_2389);
nor U2753 (N_2753,N_2198,N_2394);
or U2754 (N_2754,N_2103,N_2327);
and U2755 (N_2755,N_2398,N_2419);
nand U2756 (N_2756,N_2083,N_2177);
or U2757 (N_2757,N_2078,N_2220);
nor U2758 (N_2758,N_2404,N_2309);
nor U2759 (N_2759,N_2008,N_2161);
nor U2760 (N_2760,N_2421,N_2430);
and U2761 (N_2761,N_2257,N_2349);
nor U2762 (N_2762,N_2370,N_2487);
and U2763 (N_2763,N_2310,N_2226);
nand U2764 (N_2764,N_2020,N_2299);
nand U2765 (N_2765,N_2087,N_2335);
nor U2766 (N_2766,N_2444,N_2161);
xnor U2767 (N_2767,N_2416,N_2215);
or U2768 (N_2768,N_2067,N_2198);
nor U2769 (N_2769,N_2234,N_2299);
xnor U2770 (N_2770,N_2297,N_2319);
nor U2771 (N_2771,N_2496,N_2087);
nand U2772 (N_2772,N_2478,N_2231);
nor U2773 (N_2773,N_2432,N_2100);
nand U2774 (N_2774,N_2331,N_2242);
nor U2775 (N_2775,N_2344,N_2428);
nand U2776 (N_2776,N_2231,N_2193);
or U2777 (N_2777,N_2002,N_2338);
nor U2778 (N_2778,N_2281,N_2393);
and U2779 (N_2779,N_2270,N_2101);
nand U2780 (N_2780,N_2477,N_2291);
nor U2781 (N_2781,N_2246,N_2062);
or U2782 (N_2782,N_2010,N_2059);
or U2783 (N_2783,N_2338,N_2379);
or U2784 (N_2784,N_2044,N_2186);
and U2785 (N_2785,N_2334,N_2344);
nor U2786 (N_2786,N_2113,N_2328);
or U2787 (N_2787,N_2147,N_2391);
nand U2788 (N_2788,N_2405,N_2058);
and U2789 (N_2789,N_2221,N_2282);
xor U2790 (N_2790,N_2281,N_2159);
nor U2791 (N_2791,N_2149,N_2465);
nor U2792 (N_2792,N_2045,N_2218);
nor U2793 (N_2793,N_2142,N_2034);
nand U2794 (N_2794,N_2084,N_2049);
or U2795 (N_2795,N_2148,N_2374);
or U2796 (N_2796,N_2313,N_2239);
nand U2797 (N_2797,N_2355,N_2104);
or U2798 (N_2798,N_2492,N_2221);
or U2799 (N_2799,N_2482,N_2360);
and U2800 (N_2800,N_2204,N_2234);
nand U2801 (N_2801,N_2243,N_2284);
nand U2802 (N_2802,N_2290,N_2190);
nand U2803 (N_2803,N_2180,N_2480);
and U2804 (N_2804,N_2371,N_2273);
and U2805 (N_2805,N_2089,N_2293);
nand U2806 (N_2806,N_2248,N_2168);
or U2807 (N_2807,N_2378,N_2450);
or U2808 (N_2808,N_2497,N_2441);
nor U2809 (N_2809,N_2376,N_2260);
xnor U2810 (N_2810,N_2138,N_2274);
nand U2811 (N_2811,N_2245,N_2157);
or U2812 (N_2812,N_2369,N_2071);
or U2813 (N_2813,N_2258,N_2323);
nor U2814 (N_2814,N_2283,N_2098);
nor U2815 (N_2815,N_2055,N_2284);
and U2816 (N_2816,N_2461,N_2410);
nand U2817 (N_2817,N_2287,N_2296);
and U2818 (N_2818,N_2075,N_2270);
xor U2819 (N_2819,N_2470,N_2476);
xor U2820 (N_2820,N_2212,N_2017);
and U2821 (N_2821,N_2357,N_2255);
nor U2822 (N_2822,N_2350,N_2147);
or U2823 (N_2823,N_2014,N_2052);
nand U2824 (N_2824,N_2154,N_2384);
nor U2825 (N_2825,N_2442,N_2087);
nand U2826 (N_2826,N_2474,N_2047);
nand U2827 (N_2827,N_2327,N_2030);
nand U2828 (N_2828,N_2046,N_2124);
nand U2829 (N_2829,N_2228,N_2250);
nor U2830 (N_2830,N_2404,N_2053);
xnor U2831 (N_2831,N_2053,N_2185);
nand U2832 (N_2832,N_2081,N_2385);
xor U2833 (N_2833,N_2026,N_2170);
and U2834 (N_2834,N_2250,N_2092);
or U2835 (N_2835,N_2270,N_2429);
nor U2836 (N_2836,N_2145,N_2253);
nand U2837 (N_2837,N_2172,N_2404);
or U2838 (N_2838,N_2133,N_2089);
or U2839 (N_2839,N_2212,N_2048);
nor U2840 (N_2840,N_2365,N_2125);
nor U2841 (N_2841,N_2273,N_2000);
or U2842 (N_2842,N_2337,N_2049);
and U2843 (N_2843,N_2486,N_2422);
nand U2844 (N_2844,N_2499,N_2178);
and U2845 (N_2845,N_2275,N_2374);
nand U2846 (N_2846,N_2480,N_2444);
and U2847 (N_2847,N_2336,N_2348);
and U2848 (N_2848,N_2044,N_2180);
and U2849 (N_2849,N_2364,N_2395);
or U2850 (N_2850,N_2089,N_2379);
nand U2851 (N_2851,N_2085,N_2193);
or U2852 (N_2852,N_2373,N_2210);
nor U2853 (N_2853,N_2160,N_2255);
nand U2854 (N_2854,N_2041,N_2184);
and U2855 (N_2855,N_2439,N_2312);
nand U2856 (N_2856,N_2334,N_2156);
or U2857 (N_2857,N_2245,N_2068);
nor U2858 (N_2858,N_2235,N_2117);
nor U2859 (N_2859,N_2379,N_2195);
xnor U2860 (N_2860,N_2147,N_2169);
nand U2861 (N_2861,N_2216,N_2448);
and U2862 (N_2862,N_2417,N_2138);
nor U2863 (N_2863,N_2335,N_2495);
or U2864 (N_2864,N_2032,N_2175);
or U2865 (N_2865,N_2134,N_2497);
or U2866 (N_2866,N_2400,N_2090);
nand U2867 (N_2867,N_2271,N_2357);
or U2868 (N_2868,N_2161,N_2466);
xnor U2869 (N_2869,N_2064,N_2273);
nand U2870 (N_2870,N_2361,N_2280);
and U2871 (N_2871,N_2044,N_2477);
nor U2872 (N_2872,N_2347,N_2214);
nand U2873 (N_2873,N_2160,N_2213);
and U2874 (N_2874,N_2090,N_2253);
nand U2875 (N_2875,N_2388,N_2357);
and U2876 (N_2876,N_2320,N_2210);
nor U2877 (N_2877,N_2079,N_2050);
nor U2878 (N_2878,N_2396,N_2426);
xor U2879 (N_2879,N_2391,N_2342);
or U2880 (N_2880,N_2123,N_2452);
and U2881 (N_2881,N_2115,N_2344);
and U2882 (N_2882,N_2034,N_2443);
nor U2883 (N_2883,N_2103,N_2427);
xor U2884 (N_2884,N_2208,N_2441);
nor U2885 (N_2885,N_2433,N_2313);
nand U2886 (N_2886,N_2389,N_2471);
nor U2887 (N_2887,N_2094,N_2493);
nand U2888 (N_2888,N_2266,N_2428);
and U2889 (N_2889,N_2025,N_2071);
and U2890 (N_2890,N_2321,N_2473);
nor U2891 (N_2891,N_2413,N_2260);
and U2892 (N_2892,N_2005,N_2023);
nand U2893 (N_2893,N_2132,N_2244);
or U2894 (N_2894,N_2222,N_2296);
or U2895 (N_2895,N_2050,N_2211);
and U2896 (N_2896,N_2007,N_2366);
nand U2897 (N_2897,N_2202,N_2418);
nand U2898 (N_2898,N_2028,N_2406);
xnor U2899 (N_2899,N_2275,N_2198);
and U2900 (N_2900,N_2447,N_2464);
nor U2901 (N_2901,N_2475,N_2233);
xnor U2902 (N_2902,N_2080,N_2140);
nand U2903 (N_2903,N_2441,N_2010);
nand U2904 (N_2904,N_2039,N_2329);
or U2905 (N_2905,N_2058,N_2426);
or U2906 (N_2906,N_2014,N_2005);
and U2907 (N_2907,N_2267,N_2428);
nor U2908 (N_2908,N_2323,N_2315);
nand U2909 (N_2909,N_2092,N_2277);
nor U2910 (N_2910,N_2416,N_2249);
nand U2911 (N_2911,N_2042,N_2093);
nor U2912 (N_2912,N_2120,N_2479);
nand U2913 (N_2913,N_2112,N_2485);
and U2914 (N_2914,N_2091,N_2262);
nor U2915 (N_2915,N_2417,N_2428);
nand U2916 (N_2916,N_2347,N_2400);
and U2917 (N_2917,N_2424,N_2403);
or U2918 (N_2918,N_2302,N_2173);
nor U2919 (N_2919,N_2074,N_2161);
nor U2920 (N_2920,N_2111,N_2238);
or U2921 (N_2921,N_2406,N_2313);
nand U2922 (N_2922,N_2104,N_2012);
or U2923 (N_2923,N_2075,N_2152);
nand U2924 (N_2924,N_2357,N_2102);
xnor U2925 (N_2925,N_2241,N_2490);
xnor U2926 (N_2926,N_2363,N_2173);
xor U2927 (N_2927,N_2476,N_2030);
and U2928 (N_2928,N_2005,N_2463);
nor U2929 (N_2929,N_2010,N_2362);
xnor U2930 (N_2930,N_2195,N_2248);
and U2931 (N_2931,N_2026,N_2314);
nand U2932 (N_2932,N_2275,N_2197);
nor U2933 (N_2933,N_2415,N_2433);
or U2934 (N_2934,N_2263,N_2260);
and U2935 (N_2935,N_2340,N_2199);
nor U2936 (N_2936,N_2278,N_2372);
or U2937 (N_2937,N_2050,N_2451);
nand U2938 (N_2938,N_2128,N_2348);
nand U2939 (N_2939,N_2136,N_2043);
or U2940 (N_2940,N_2462,N_2319);
xnor U2941 (N_2941,N_2484,N_2195);
nand U2942 (N_2942,N_2427,N_2346);
or U2943 (N_2943,N_2119,N_2040);
nor U2944 (N_2944,N_2318,N_2088);
or U2945 (N_2945,N_2256,N_2478);
or U2946 (N_2946,N_2094,N_2239);
nand U2947 (N_2947,N_2455,N_2383);
or U2948 (N_2948,N_2305,N_2375);
and U2949 (N_2949,N_2021,N_2276);
and U2950 (N_2950,N_2497,N_2443);
nor U2951 (N_2951,N_2078,N_2485);
and U2952 (N_2952,N_2014,N_2270);
nand U2953 (N_2953,N_2313,N_2424);
and U2954 (N_2954,N_2293,N_2487);
xnor U2955 (N_2955,N_2237,N_2122);
nand U2956 (N_2956,N_2068,N_2123);
nand U2957 (N_2957,N_2071,N_2490);
and U2958 (N_2958,N_2317,N_2122);
nand U2959 (N_2959,N_2069,N_2177);
and U2960 (N_2960,N_2077,N_2055);
nand U2961 (N_2961,N_2195,N_2221);
nor U2962 (N_2962,N_2270,N_2042);
nor U2963 (N_2963,N_2138,N_2144);
nand U2964 (N_2964,N_2183,N_2422);
nand U2965 (N_2965,N_2350,N_2209);
nor U2966 (N_2966,N_2438,N_2369);
xor U2967 (N_2967,N_2446,N_2109);
xor U2968 (N_2968,N_2029,N_2061);
or U2969 (N_2969,N_2479,N_2438);
or U2970 (N_2970,N_2477,N_2386);
xnor U2971 (N_2971,N_2436,N_2324);
nand U2972 (N_2972,N_2177,N_2188);
nor U2973 (N_2973,N_2309,N_2080);
and U2974 (N_2974,N_2051,N_2326);
or U2975 (N_2975,N_2079,N_2289);
or U2976 (N_2976,N_2335,N_2447);
nor U2977 (N_2977,N_2385,N_2426);
nand U2978 (N_2978,N_2379,N_2336);
nor U2979 (N_2979,N_2056,N_2285);
nor U2980 (N_2980,N_2327,N_2471);
and U2981 (N_2981,N_2369,N_2127);
nand U2982 (N_2982,N_2357,N_2116);
nor U2983 (N_2983,N_2337,N_2327);
or U2984 (N_2984,N_2230,N_2334);
or U2985 (N_2985,N_2205,N_2201);
nand U2986 (N_2986,N_2450,N_2146);
or U2987 (N_2987,N_2016,N_2109);
nand U2988 (N_2988,N_2433,N_2076);
nor U2989 (N_2989,N_2236,N_2231);
nand U2990 (N_2990,N_2137,N_2106);
or U2991 (N_2991,N_2153,N_2279);
nor U2992 (N_2992,N_2343,N_2300);
nor U2993 (N_2993,N_2324,N_2405);
nor U2994 (N_2994,N_2284,N_2166);
nor U2995 (N_2995,N_2125,N_2354);
nor U2996 (N_2996,N_2383,N_2454);
nor U2997 (N_2997,N_2394,N_2417);
xor U2998 (N_2998,N_2215,N_2451);
nand U2999 (N_2999,N_2256,N_2413);
nor U3000 (N_3000,N_2578,N_2745);
or U3001 (N_3001,N_2866,N_2896);
nand U3002 (N_3002,N_2945,N_2953);
or U3003 (N_3003,N_2799,N_2765);
or U3004 (N_3004,N_2822,N_2545);
nor U3005 (N_3005,N_2861,N_2814);
and U3006 (N_3006,N_2942,N_2825);
nand U3007 (N_3007,N_2719,N_2725);
or U3008 (N_3008,N_2510,N_2950);
or U3009 (N_3009,N_2877,N_2702);
and U3010 (N_3010,N_2947,N_2742);
or U3011 (N_3011,N_2559,N_2837);
nand U3012 (N_3012,N_2900,N_2606);
nand U3013 (N_3013,N_2812,N_2603);
or U3014 (N_3014,N_2983,N_2671);
or U3015 (N_3015,N_2675,N_2576);
xor U3016 (N_3016,N_2818,N_2723);
nand U3017 (N_3017,N_2922,N_2705);
nand U3018 (N_3018,N_2733,N_2797);
nand U3019 (N_3019,N_2806,N_2616);
xor U3020 (N_3020,N_2557,N_2573);
nor U3021 (N_3021,N_2787,N_2928);
nand U3022 (N_3022,N_2568,N_2650);
or U3023 (N_3023,N_2832,N_2630);
nor U3024 (N_3024,N_2701,N_2612);
nor U3025 (N_3025,N_2501,N_2644);
and U3026 (N_3026,N_2770,N_2854);
or U3027 (N_3027,N_2524,N_2810);
and U3028 (N_3028,N_2535,N_2869);
nand U3029 (N_3029,N_2871,N_2727);
xnor U3030 (N_3030,N_2722,N_2566);
xnor U3031 (N_3031,N_2564,N_2767);
xor U3032 (N_3032,N_2631,N_2561);
and U3033 (N_3033,N_2614,N_2919);
and U3034 (N_3034,N_2632,N_2562);
xor U3035 (N_3035,N_2639,N_2528);
and U3036 (N_3036,N_2542,N_2514);
nor U3037 (N_3037,N_2527,N_2899);
nand U3038 (N_3038,N_2581,N_2623);
nand U3039 (N_3039,N_2776,N_2629);
nor U3040 (N_3040,N_2683,N_2613);
or U3041 (N_3041,N_2696,N_2763);
xor U3042 (N_3042,N_2918,N_2716);
or U3043 (N_3043,N_2887,N_2815);
and U3044 (N_3044,N_2661,N_2688);
and U3045 (N_3045,N_2657,N_2924);
nor U3046 (N_3046,N_2969,N_2570);
and U3047 (N_3047,N_2802,N_2707);
nor U3048 (N_3048,N_2646,N_2740);
nand U3049 (N_3049,N_2758,N_2941);
xnor U3050 (N_3050,N_2826,N_2820);
nor U3051 (N_3051,N_2749,N_2540);
or U3052 (N_3052,N_2883,N_2714);
and U3053 (N_3053,N_2638,N_2793);
nor U3054 (N_3054,N_2778,N_2584);
or U3055 (N_3055,N_2615,N_2952);
nor U3056 (N_3056,N_2626,N_2914);
and U3057 (N_3057,N_2656,N_2951);
nor U3058 (N_3058,N_2607,N_2841);
and U3059 (N_3059,N_2890,N_2731);
and U3060 (N_3060,N_2968,N_2715);
and U3061 (N_3061,N_2577,N_2721);
and U3062 (N_3062,N_2990,N_2582);
nand U3063 (N_3063,N_2682,N_2588);
xor U3064 (N_3064,N_2999,N_2687);
nor U3065 (N_3065,N_2912,N_2549);
or U3066 (N_3066,N_2594,N_2788);
xnor U3067 (N_3067,N_2816,N_2930);
nand U3068 (N_3068,N_2591,N_2959);
or U3069 (N_3069,N_2773,N_2590);
or U3070 (N_3070,N_2936,N_2636);
and U3071 (N_3071,N_2972,N_2686);
xnor U3072 (N_3072,N_2658,N_2921);
nor U3073 (N_3073,N_2592,N_2800);
nor U3074 (N_3074,N_2691,N_2779);
or U3075 (N_3075,N_2766,N_2505);
or U3076 (N_3076,N_2823,N_2830);
nor U3077 (N_3077,N_2597,N_2729);
and U3078 (N_3078,N_2831,N_2531);
and U3079 (N_3079,N_2599,N_2637);
or U3080 (N_3080,N_2543,N_2500);
nor U3081 (N_3081,N_2579,N_2610);
nand U3082 (N_3082,N_2813,N_2619);
or U3083 (N_3083,N_2509,N_2625);
and U3084 (N_3084,N_2840,N_2943);
nand U3085 (N_3085,N_2709,N_2875);
nand U3086 (N_3086,N_2670,N_2911);
and U3087 (N_3087,N_2991,N_2835);
or U3088 (N_3088,N_2586,N_2673);
nor U3089 (N_3089,N_2621,N_2885);
or U3090 (N_3090,N_2624,N_2906);
and U3091 (N_3091,N_2640,N_2532);
or U3092 (N_3092,N_2734,N_2583);
or U3093 (N_3093,N_2774,N_2751);
nand U3094 (N_3094,N_2703,N_2664);
nor U3095 (N_3095,N_2992,N_2595);
and U3096 (N_3096,N_2667,N_2781);
xor U3097 (N_3097,N_2771,N_2975);
nand U3098 (N_3098,N_2746,N_2934);
nor U3099 (N_3099,N_2865,N_2948);
and U3100 (N_3100,N_2873,N_2757);
nor U3101 (N_3101,N_2717,N_2651);
and U3102 (N_3102,N_2989,N_2548);
xor U3103 (N_3103,N_2805,N_2986);
nand U3104 (N_3104,N_2889,N_2756);
nand U3105 (N_3105,N_2768,N_2710);
nand U3106 (N_3106,N_2694,N_2801);
nor U3107 (N_3107,N_2539,N_2518);
nand U3108 (N_3108,N_2507,N_2849);
and U3109 (N_3109,N_2519,N_2598);
nor U3110 (N_3110,N_2609,N_2931);
nand U3111 (N_3111,N_2777,N_2977);
nand U3112 (N_3112,N_2556,N_2970);
nor U3113 (N_3113,N_2876,N_2792);
and U3114 (N_3114,N_2760,N_2649);
nor U3115 (N_3115,N_2834,N_2958);
nor U3116 (N_3116,N_2563,N_2713);
and U3117 (N_3117,N_2523,N_2521);
or U3118 (N_3118,N_2574,N_2516);
nor U3119 (N_3119,N_2726,N_2888);
nand U3120 (N_3120,N_2659,N_2971);
nor U3121 (N_3121,N_2672,N_2753);
nor U3122 (N_3122,N_2907,N_2735);
nor U3123 (N_3123,N_2522,N_2634);
xnor U3124 (N_3124,N_2937,N_2819);
and U3125 (N_3125,N_2844,N_2796);
and U3126 (N_3126,N_2700,N_2593);
or U3127 (N_3127,N_2909,N_2994);
or U3128 (N_3128,N_2738,N_2600);
or U3129 (N_3129,N_2571,N_2517);
nor U3130 (N_3130,N_2782,N_2643);
and U3131 (N_3131,N_2962,N_2580);
or U3132 (N_3132,N_2917,N_2935);
and U3133 (N_3133,N_2957,N_2515);
and U3134 (N_3134,N_2836,N_2784);
nor U3135 (N_3135,N_2905,N_2620);
nor U3136 (N_3136,N_2652,N_2504);
xor U3137 (N_3137,N_2602,N_2698);
and U3138 (N_3138,N_2979,N_2882);
nor U3139 (N_3139,N_2622,N_2827);
nor U3140 (N_3140,N_2647,N_2526);
nand U3141 (N_3141,N_2982,N_2685);
and U3142 (N_3142,N_2926,N_2569);
nor U3143 (N_3143,N_2891,N_2892);
or U3144 (N_3144,N_2728,N_2886);
nor U3145 (N_3145,N_2920,N_2572);
and U3146 (N_3146,N_2944,N_2544);
and U3147 (N_3147,N_2674,N_2856);
and U3148 (N_3148,N_2839,N_2974);
nor U3149 (N_3149,N_2684,N_2536);
nor U3150 (N_3150,N_2976,N_2993);
or U3151 (N_3151,N_2681,N_2967);
xor U3152 (N_3152,N_2870,N_2963);
nor U3153 (N_3153,N_2955,N_2772);
xor U3154 (N_3154,N_2965,N_2828);
or U3155 (N_3155,N_2803,N_2748);
or U3156 (N_3156,N_2791,N_2699);
nor U3157 (N_3157,N_2884,N_2858);
and U3158 (N_3158,N_2711,N_2833);
xnor U3159 (N_3159,N_2995,N_2933);
nand U3160 (N_3160,N_2966,N_2680);
and U3161 (N_3161,N_2712,N_2601);
nor U3162 (N_3162,N_2956,N_2985);
or U3163 (N_3163,N_2927,N_2857);
nor U3164 (N_3164,N_2940,N_2642);
xor U3165 (N_3165,N_2506,N_2736);
or U3166 (N_3166,N_2704,N_2904);
nor U3167 (N_3167,N_2775,N_2786);
and U3168 (N_3168,N_2783,N_2874);
and U3169 (N_3169,N_2520,N_2817);
nor U3170 (N_3170,N_2750,N_2916);
and U3171 (N_3171,N_2508,N_2860);
nor U3172 (N_3172,N_2648,N_2554);
nand U3173 (N_3173,N_2973,N_2780);
or U3174 (N_3174,N_2737,N_2880);
or U3175 (N_3175,N_2910,N_2850);
nand U3176 (N_3176,N_2903,N_2628);
nor U3177 (N_3177,N_2747,N_2752);
nor U3178 (N_3178,N_2997,N_2879);
and U3179 (N_3179,N_2895,N_2808);
xor U3180 (N_3180,N_2795,N_2961);
xnor U3181 (N_3181,N_2980,N_2503);
xnor U3182 (N_3182,N_2732,N_2862);
nor U3183 (N_3183,N_2692,N_2764);
or U3184 (N_3184,N_2938,N_2996);
nand U3185 (N_3185,N_2718,N_2635);
or U3186 (N_3186,N_2617,N_2641);
nand U3187 (N_3187,N_2987,N_2811);
or U3188 (N_3188,N_2847,N_2533);
or U3189 (N_3189,N_2878,N_2541);
nor U3190 (N_3190,N_2852,N_2960);
nor U3191 (N_3191,N_2894,N_2845);
and U3192 (N_3192,N_2925,N_2846);
nor U3193 (N_3193,N_2645,N_2998);
nand U3194 (N_3194,N_2575,N_2537);
and U3195 (N_3195,N_2678,N_2853);
nor U3196 (N_3196,N_2690,N_2502);
or U3197 (N_3197,N_2720,N_2739);
nand U3198 (N_3198,N_2868,N_2789);
nor U3199 (N_3199,N_2618,N_2913);
or U3200 (N_3200,N_2743,N_2538);
nor U3201 (N_3201,N_2534,N_2693);
nor U3202 (N_3202,N_2908,N_2949);
nand U3203 (N_3203,N_2550,N_2964);
xor U3204 (N_3204,N_2859,N_2724);
nand U3205 (N_3205,N_2754,N_2755);
and U3206 (N_3206,N_2513,N_2633);
nor U3207 (N_3207,N_2843,N_2668);
nor U3208 (N_3208,N_2842,N_2558);
and U3209 (N_3209,N_2662,N_2984);
and U3210 (N_3210,N_2863,N_2798);
nand U3211 (N_3211,N_2653,N_2676);
nand U3212 (N_3212,N_2848,N_2530);
and U3213 (N_3213,N_2585,N_2730);
xor U3214 (N_3214,N_2851,N_2829);
nand U3215 (N_3215,N_2589,N_2855);
nor U3216 (N_3216,N_2669,N_2665);
or U3217 (N_3217,N_2769,N_2872);
nand U3218 (N_3218,N_2547,N_2596);
or U3219 (N_3219,N_2915,N_2978);
nand U3220 (N_3220,N_2654,N_2804);
nand U3221 (N_3221,N_2565,N_2807);
and U3222 (N_3222,N_2525,N_2660);
or U3223 (N_3223,N_2809,N_2655);
nand U3224 (N_3224,N_2611,N_2902);
and U3225 (N_3225,N_2864,N_2666);
and U3226 (N_3226,N_2511,N_2794);
xor U3227 (N_3227,N_2923,N_2546);
xor U3228 (N_3228,N_2679,N_2677);
nor U3229 (N_3229,N_2587,N_2838);
nand U3230 (N_3230,N_2608,N_2954);
nand U3231 (N_3231,N_2560,N_2785);
nor U3232 (N_3232,N_2689,N_2708);
nor U3233 (N_3233,N_2939,N_2605);
and U3234 (N_3234,N_2762,N_2761);
nand U3235 (N_3235,N_2932,N_2604);
nor U3236 (N_3236,N_2555,N_2790);
nor U3237 (N_3237,N_2821,N_2929);
or U3238 (N_3238,N_2897,N_2627);
and U3239 (N_3239,N_2988,N_2551);
nand U3240 (N_3240,N_2981,N_2553);
and U3241 (N_3241,N_2567,N_2706);
nor U3242 (N_3242,N_2898,N_2881);
nand U3243 (N_3243,N_2697,N_2901);
or U3244 (N_3244,N_2744,N_2893);
nand U3245 (N_3245,N_2663,N_2695);
or U3246 (N_3246,N_2759,N_2946);
xnor U3247 (N_3247,N_2552,N_2867);
nand U3248 (N_3248,N_2824,N_2512);
or U3249 (N_3249,N_2741,N_2529);
or U3250 (N_3250,N_2816,N_2735);
or U3251 (N_3251,N_2512,N_2887);
nand U3252 (N_3252,N_2977,N_2655);
or U3253 (N_3253,N_2947,N_2968);
or U3254 (N_3254,N_2793,N_2852);
and U3255 (N_3255,N_2716,N_2783);
xor U3256 (N_3256,N_2797,N_2928);
nor U3257 (N_3257,N_2546,N_2538);
and U3258 (N_3258,N_2993,N_2956);
nand U3259 (N_3259,N_2898,N_2562);
or U3260 (N_3260,N_2836,N_2886);
nand U3261 (N_3261,N_2753,N_2961);
nand U3262 (N_3262,N_2810,N_2536);
and U3263 (N_3263,N_2858,N_2916);
nor U3264 (N_3264,N_2884,N_2941);
nor U3265 (N_3265,N_2756,N_2553);
and U3266 (N_3266,N_2940,N_2710);
or U3267 (N_3267,N_2960,N_2821);
nand U3268 (N_3268,N_2740,N_2916);
xnor U3269 (N_3269,N_2631,N_2957);
nor U3270 (N_3270,N_2638,N_2864);
and U3271 (N_3271,N_2772,N_2754);
or U3272 (N_3272,N_2886,N_2985);
or U3273 (N_3273,N_2929,N_2646);
nand U3274 (N_3274,N_2828,N_2704);
nor U3275 (N_3275,N_2524,N_2803);
xnor U3276 (N_3276,N_2579,N_2947);
nor U3277 (N_3277,N_2932,N_2720);
or U3278 (N_3278,N_2592,N_2900);
nand U3279 (N_3279,N_2929,N_2942);
nor U3280 (N_3280,N_2524,N_2916);
nor U3281 (N_3281,N_2730,N_2866);
nor U3282 (N_3282,N_2831,N_2722);
or U3283 (N_3283,N_2882,N_2895);
nand U3284 (N_3284,N_2965,N_2619);
nor U3285 (N_3285,N_2680,N_2513);
and U3286 (N_3286,N_2647,N_2700);
nand U3287 (N_3287,N_2937,N_2915);
nand U3288 (N_3288,N_2634,N_2858);
and U3289 (N_3289,N_2666,N_2619);
and U3290 (N_3290,N_2924,N_2745);
nand U3291 (N_3291,N_2792,N_2591);
xnor U3292 (N_3292,N_2762,N_2978);
nor U3293 (N_3293,N_2517,N_2988);
and U3294 (N_3294,N_2977,N_2983);
or U3295 (N_3295,N_2619,N_2685);
xor U3296 (N_3296,N_2680,N_2934);
or U3297 (N_3297,N_2544,N_2613);
or U3298 (N_3298,N_2703,N_2940);
or U3299 (N_3299,N_2874,N_2599);
nand U3300 (N_3300,N_2541,N_2617);
xnor U3301 (N_3301,N_2753,N_2821);
nor U3302 (N_3302,N_2560,N_2966);
nand U3303 (N_3303,N_2956,N_2518);
and U3304 (N_3304,N_2550,N_2619);
and U3305 (N_3305,N_2823,N_2820);
nand U3306 (N_3306,N_2620,N_2635);
nor U3307 (N_3307,N_2651,N_2997);
nor U3308 (N_3308,N_2693,N_2815);
or U3309 (N_3309,N_2872,N_2901);
or U3310 (N_3310,N_2700,N_2722);
nand U3311 (N_3311,N_2933,N_2699);
nor U3312 (N_3312,N_2899,N_2801);
nor U3313 (N_3313,N_2547,N_2965);
nor U3314 (N_3314,N_2827,N_2514);
or U3315 (N_3315,N_2906,N_2768);
nand U3316 (N_3316,N_2917,N_2730);
xor U3317 (N_3317,N_2796,N_2657);
nor U3318 (N_3318,N_2689,N_2717);
nor U3319 (N_3319,N_2566,N_2530);
nor U3320 (N_3320,N_2873,N_2966);
or U3321 (N_3321,N_2906,N_2597);
or U3322 (N_3322,N_2747,N_2577);
and U3323 (N_3323,N_2572,N_2859);
nor U3324 (N_3324,N_2982,N_2547);
nor U3325 (N_3325,N_2629,N_2895);
and U3326 (N_3326,N_2959,N_2528);
and U3327 (N_3327,N_2655,N_2933);
nand U3328 (N_3328,N_2747,N_2688);
or U3329 (N_3329,N_2925,N_2917);
or U3330 (N_3330,N_2720,N_2911);
or U3331 (N_3331,N_2513,N_2975);
and U3332 (N_3332,N_2761,N_2735);
and U3333 (N_3333,N_2743,N_2920);
xor U3334 (N_3334,N_2608,N_2713);
or U3335 (N_3335,N_2765,N_2875);
or U3336 (N_3336,N_2766,N_2647);
and U3337 (N_3337,N_2832,N_2559);
or U3338 (N_3338,N_2793,N_2856);
and U3339 (N_3339,N_2632,N_2884);
nor U3340 (N_3340,N_2658,N_2952);
and U3341 (N_3341,N_2612,N_2693);
nand U3342 (N_3342,N_2800,N_2602);
or U3343 (N_3343,N_2957,N_2757);
or U3344 (N_3344,N_2559,N_2568);
nor U3345 (N_3345,N_2541,N_2584);
nor U3346 (N_3346,N_2906,N_2518);
or U3347 (N_3347,N_2878,N_2647);
nand U3348 (N_3348,N_2964,N_2937);
or U3349 (N_3349,N_2747,N_2842);
nand U3350 (N_3350,N_2886,N_2617);
xnor U3351 (N_3351,N_2632,N_2576);
nor U3352 (N_3352,N_2766,N_2623);
and U3353 (N_3353,N_2748,N_2972);
nand U3354 (N_3354,N_2997,N_2936);
nand U3355 (N_3355,N_2735,N_2770);
nand U3356 (N_3356,N_2642,N_2971);
nor U3357 (N_3357,N_2778,N_2797);
and U3358 (N_3358,N_2551,N_2876);
nor U3359 (N_3359,N_2710,N_2688);
nand U3360 (N_3360,N_2622,N_2822);
nand U3361 (N_3361,N_2642,N_2915);
or U3362 (N_3362,N_2927,N_2745);
nand U3363 (N_3363,N_2514,N_2844);
and U3364 (N_3364,N_2580,N_2657);
nand U3365 (N_3365,N_2784,N_2746);
nand U3366 (N_3366,N_2745,N_2664);
nor U3367 (N_3367,N_2896,N_2829);
or U3368 (N_3368,N_2940,N_2707);
nand U3369 (N_3369,N_2518,N_2691);
xnor U3370 (N_3370,N_2967,N_2608);
nand U3371 (N_3371,N_2720,N_2986);
or U3372 (N_3372,N_2706,N_2792);
or U3373 (N_3373,N_2978,N_2557);
nor U3374 (N_3374,N_2531,N_2706);
or U3375 (N_3375,N_2903,N_2683);
xnor U3376 (N_3376,N_2566,N_2510);
xnor U3377 (N_3377,N_2579,N_2802);
nor U3378 (N_3378,N_2888,N_2667);
nand U3379 (N_3379,N_2955,N_2565);
nand U3380 (N_3380,N_2574,N_2846);
nor U3381 (N_3381,N_2738,N_2596);
or U3382 (N_3382,N_2638,N_2568);
and U3383 (N_3383,N_2639,N_2566);
or U3384 (N_3384,N_2919,N_2580);
xnor U3385 (N_3385,N_2569,N_2705);
or U3386 (N_3386,N_2666,N_2541);
and U3387 (N_3387,N_2796,N_2705);
or U3388 (N_3388,N_2500,N_2787);
and U3389 (N_3389,N_2771,N_2942);
nand U3390 (N_3390,N_2992,N_2800);
nor U3391 (N_3391,N_2799,N_2846);
nor U3392 (N_3392,N_2928,N_2513);
nand U3393 (N_3393,N_2809,N_2737);
xor U3394 (N_3394,N_2729,N_2504);
or U3395 (N_3395,N_2861,N_2518);
nor U3396 (N_3396,N_2793,N_2572);
nand U3397 (N_3397,N_2706,N_2901);
nor U3398 (N_3398,N_2938,N_2797);
nand U3399 (N_3399,N_2692,N_2924);
and U3400 (N_3400,N_2921,N_2734);
nor U3401 (N_3401,N_2588,N_2629);
nand U3402 (N_3402,N_2574,N_2787);
nand U3403 (N_3403,N_2653,N_2710);
xnor U3404 (N_3404,N_2818,N_2901);
and U3405 (N_3405,N_2517,N_2771);
nand U3406 (N_3406,N_2981,N_2681);
and U3407 (N_3407,N_2956,N_2570);
nand U3408 (N_3408,N_2675,N_2597);
or U3409 (N_3409,N_2513,N_2752);
nor U3410 (N_3410,N_2833,N_2795);
xnor U3411 (N_3411,N_2756,N_2926);
and U3412 (N_3412,N_2823,N_2685);
nor U3413 (N_3413,N_2780,N_2878);
nor U3414 (N_3414,N_2693,N_2724);
nand U3415 (N_3415,N_2563,N_2613);
nand U3416 (N_3416,N_2865,N_2690);
nor U3417 (N_3417,N_2642,N_2751);
and U3418 (N_3418,N_2595,N_2986);
or U3419 (N_3419,N_2854,N_2925);
nand U3420 (N_3420,N_2931,N_2788);
nor U3421 (N_3421,N_2914,N_2820);
and U3422 (N_3422,N_2862,N_2924);
or U3423 (N_3423,N_2665,N_2744);
and U3424 (N_3424,N_2706,N_2615);
or U3425 (N_3425,N_2685,N_2911);
or U3426 (N_3426,N_2615,N_2943);
and U3427 (N_3427,N_2501,N_2536);
and U3428 (N_3428,N_2852,N_2754);
nand U3429 (N_3429,N_2669,N_2551);
or U3430 (N_3430,N_2940,N_2755);
nand U3431 (N_3431,N_2696,N_2838);
nor U3432 (N_3432,N_2840,N_2945);
or U3433 (N_3433,N_2940,N_2721);
nor U3434 (N_3434,N_2586,N_2820);
and U3435 (N_3435,N_2894,N_2708);
or U3436 (N_3436,N_2516,N_2770);
nor U3437 (N_3437,N_2575,N_2805);
xor U3438 (N_3438,N_2808,N_2503);
nor U3439 (N_3439,N_2753,N_2863);
nand U3440 (N_3440,N_2523,N_2752);
nand U3441 (N_3441,N_2885,N_2588);
nand U3442 (N_3442,N_2879,N_2706);
and U3443 (N_3443,N_2846,N_2743);
xor U3444 (N_3444,N_2557,N_2897);
nand U3445 (N_3445,N_2535,N_2782);
nor U3446 (N_3446,N_2888,N_2642);
nor U3447 (N_3447,N_2866,N_2868);
nor U3448 (N_3448,N_2568,N_2760);
or U3449 (N_3449,N_2720,N_2859);
nand U3450 (N_3450,N_2826,N_2692);
or U3451 (N_3451,N_2576,N_2860);
and U3452 (N_3452,N_2805,N_2682);
nor U3453 (N_3453,N_2806,N_2729);
nor U3454 (N_3454,N_2718,N_2734);
xor U3455 (N_3455,N_2621,N_2517);
nand U3456 (N_3456,N_2928,N_2589);
nor U3457 (N_3457,N_2749,N_2677);
nor U3458 (N_3458,N_2628,N_2977);
and U3459 (N_3459,N_2707,N_2530);
nand U3460 (N_3460,N_2939,N_2745);
nand U3461 (N_3461,N_2662,N_2856);
nand U3462 (N_3462,N_2707,N_2935);
nand U3463 (N_3463,N_2840,N_2779);
or U3464 (N_3464,N_2885,N_2716);
or U3465 (N_3465,N_2994,N_2579);
nand U3466 (N_3466,N_2511,N_2562);
nand U3467 (N_3467,N_2741,N_2696);
nor U3468 (N_3468,N_2587,N_2775);
and U3469 (N_3469,N_2647,N_2549);
nor U3470 (N_3470,N_2570,N_2770);
and U3471 (N_3471,N_2732,N_2573);
nor U3472 (N_3472,N_2527,N_2635);
nand U3473 (N_3473,N_2844,N_2551);
xor U3474 (N_3474,N_2848,N_2581);
nor U3475 (N_3475,N_2697,N_2770);
nor U3476 (N_3476,N_2850,N_2804);
and U3477 (N_3477,N_2510,N_2868);
nand U3478 (N_3478,N_2712,N_2653);
and U3479 (N_3479,N_2968,N_2560);
xor U3480 (N_3480,N_2644,N_2755);
nand U3481 (N_3481,N_2626,N_2564);
nor U3482 (N_3482,N_2680,N_2582);
or U3483 (N_3483,N_2965,N_2689);
nor U3484 (N_3484,N_2870,N_2508);
or U3485 (N_3485,N_2656,N_2510);
or U3486 (N_3486,N_2633,N_2876);
nor U3487 (N_3487,N_2624,N_2739);
and U3488 (N_3488,N_2956,N_2774);
or U3489 (N_3489,N_2668,N_2540);
and U3490 (N_3490,N_2878,N_2734);
or U3491 (N_3491,N_2621,N_2920);
nor U3492 (N_3492,N_2726,N_2825);
or U3493 (N_3493,N_2515,N_2893);
or U3494 (N_3494,N_2558,N_2976);
and U3495 (N_3495,N_2971,N_2873);
and U3496 (N_3496,N_2953,N_2776);
and U3497 (N_3497,N_2513,N_2603);
nor U3498 (N_3498,N_2896,N_2990);
nor U3499 (N_3499,N_2726,N_2588);
nor U3500 (N_3500,N_3013,N_3138);
nand U3501 (N_3501,N_3272,N_3172);
and U3502 (N_3502,N_3025,N_3405);
or U3503 (N_3503,N_3200,N_3166);
or U3504 (N_3504,N_3391,N_3477);
or U3505 (N_3505,N_3457,N_3120);
nand U3506 (N_3506,N_3462,N_3180);
or U3507 (N_3507,N_3413,N_3182);
nand U3508 (N_3508,N_3194,N_3400);
nor U3509 (N_3509,N_3156,N_3312);
or U3510 (N_3510,N_3011,N_3398);
or U3511 (N_3511,N_3291,N_3484);
xor U3512 (N_3512,N_3237,N_3455);
nand U3513 (N_3513,N_3043,N_3419);
nand U3514 (N_3514,N_3203,N_3224);
and U3515 (N_3515,N_3229,N_3289);
or U3516 (N_3516,N_3357,N_3451);
nor U3517 (N_3517,N_3481,N_3275);
or U3518 (N_3518,N_3044,N_3360);
nand U3519 (N_3519,N_3217,N_3000);
nand U3520 (N_3520,N_3458,N_3049);
nor U3521 (N_3521,N_3308,N_3428);
xor U3522 (N_3522,N_3082,N_3062);
and U3523 (N_3523,N_3454,N_3397);
nor U3524 (N_3524,N_3252,N_3209);
nand U3525 (N_3525,N_3205,N_3113);
or U3526 (N_3526,N_3157,N_3035);
nor U3527 (N_3527,N_3117,N_3039);
nand U3528 (N_3528,N_3336,N_3263);
nor U3529 (N_3529,N_3257,N_3358);
and U3530 (N_3530,N_3173,N_3068);
and U3531 (N_3531,N_3111,N_3202);
nand U3532 (N_3532,N_3109,N_3052);
nor U3533 (N_3533,N_3161,N_3486);
or U3534 (N_3534,N_3430,N_3235);
nor U3535 (N_3535,N_3073,N_3404);
nor U3536 (N_3536,N_3315,N_3163);
and U3537 (N_3537,N_3331,N_3136);
or U3538 (N_3538,N_3438,N_3219);
nor U3539 (N_3539,N_3348,N_3036);
xor U3540 (N_3540,N_3145,N_3086);
nor U3541 (N_3541,N_3305,N_3223);
or U3542 (N_3542,N_3241,N_3239);
nand U3543 (N_3543,N_3393,N_3242);
nand U3544 (N_3544,N_3273,N_3016);
and U3545 (N_3545,N_3048,N_3444);
nand U3546 (N_3546,N_3147,N_3142);
or U3547 (N_3547,N_3485,N_3148);
and U3548 (N_3548,N_3187,N_3078);
xor U3549 (N_3549,N_3302,N_3411);
or U3550 (N_3550,N_3018,N_3283);
or U3551 (N_3551,N_3421,N_3255);
and U3552 (N_3552,N_3055,N_3488);
and U3553 (N_3553,N_3338,N_3352);
nand U3554 (N_3554,N_3318,N_3408);
or U3555 (N_3555,N_3435,N_3406);
nor U3556 (N_3556,N_3079,N_3096);
nor U3557 (N_3557,N_3080,N_3297);
or U3558 (N_3558,N_3323,N_3403);
and U3559 (N_3559,N_3159,N_3285);
nor U3560 (N_3560,N_3464,N_3350);
nand U3561 (N_3561,N_3063,N_3115);
or U3562 (N_3562,N_3045,N_3014);
or U3563 (N_3563,N_3456,N_3066);
and U3564 (N_3564,N_3005,N_3046);
and U3565 (N_3565,N_3491,N_3232);
nand U3566 (N_3566,N_3024,N_3377);
xnor U3567 (N_3567,N_3296,N_3245);
nand U3568 (N_3568,N_3123,N_3058);
nand U3569 (N_3569,N_3056,N_3480);
or U3570 (N_3570,N_3425,N_3370);
or U3571 (N_3571,N_3069,N_3322);
or U3572 (N_3572,N_3216,N_3470);
nand U3573 (N_3573,N_3121,N_3333);
or U3574 (N_3574,N_3437,N_3294);
xnor U3575 (N_3575,N_3231,N_3251);
nor U3576 (N_3576,N_3290,N_3204);
or U3577 (N_3577,N_3375,N_3385);
nand U3578 (N_3578,N_3309,N_3335);
or U3579 (N_3579,N_3211,N_3093);
and U3580 (N_3580,N_3353,N_3116);
nand U3581 (N_3581,N_3114,N_3284);
nor U3582 (N_3582,N_3206,N_3372);
nand U3583 (N_3583,N_3198,N_3442);
or U3584 (N_3584,N_3483,N_3139);
nor U3585 (N_3585,N_3171,N_3426);
nor U3586 (N_3586,N_3065,N_3339);
xnor U3587 (N_3587,N_3461,N_3356);
and U3588 (N_3588,N_3416,N_3320);
and U3589 (N_3589,N_3299,N_3394);
nand U3590 (N_3590,N_3432,N_3351);
nand U3591 (N_3591,N_3327,N_3012);
or U3592 (N_3592,N_3176,N_3498);
nor U3593 (N_3593,N_3310,N_3247);
and U3594 (N_3594,N_3193,N_3174);
xnor U3595 (N_3595,N_3183,N_3029);
and U3596 (N_3596,N_3420,N_3050);
nor U3597 (N_3597,N_3033,N_3101);
and U3598 (N_3598,N_3190,N_3369);
nand U3599 (N_3599,N_3077,N_3249);
and U3600 (N_3600,N_3246,N_3152);
and U3601 (N_3601,N_3020,N_3164);
nand U3602 (N_3602,N_3165,N_3402);
nand U3603 (N_3603,N_3053,N_3155);
xor U3604 (N_3604,N_3207,N_3493);
nand U3605 (N_3605,N_3060,N_3149);
xnor U3606 (N_3606,N_3466,N_3003);
nor U3607 (N_3607,N_3441,N_3074);
xnor U3608 (N_3608,N_3355,N_3220);
xor U3609 (N_3609,N_3316,N_3445);
nor U3610 (N_3610,N_3340,N_3017);
or U3611 (N_3611,N_3097,N_3192);
nand U3612 (N_3612,N_3407,N_3343);
nor U3613 (N_3613,N_3324,N_3387);
and U3614 (N_3614,N_3112,N_3081);
nor U3615 (N_3615,N_3179,N_3042);
or U3616 (N_3616,N_3492,N_3459);
or U3617 (N_3617,N_3474,N_3233);
xnor U3618 (N_3618,N_3363,N_3143);
or U3619 (N_3619,N_3361,N_3104);
and U3620 (N_3620,N_3095,N_3282);
and U3621 (N_3621,N_3376,N_3390);
nor U3622 (N_3622,N_3278,N_3325);
or U3623 (N_3623,N_3041,N_3276);
and U3624 (N_3624,N_3258,N_3424);
or U3625 (N_3625,N_3307,N_3448);
and U3626 (N_3626,N_3076,N_3141);
nor U3627 (N_3627,N_3134,N_3218);
or U3628 (N_3628,N_3250,N_3383);
nand U3629 (N_3629,N_3450,N_3146);
and U3630 (N_3630,N_3191,N_3021);
xor U3631 (N_3631,N_3059,N_3479);
nor U3632 (N_3632,N_3128,N_3215);
nor U3633 (N_3633,N_3061,N_3449);
nor U3634 (N_3634,N_3034,N_3422);
nor U3635 (N_3635,N_3471,N_3364);
nor U3636 (N_3636,N_3099,N_3040);
nand U3637 (N_3637,N_3015,N_3254);
and U3638 (N_3638,N_3195,N_3395);
or U3639 (N_3639,N_3277,N_3085);
and U3640 (N_3640,N_3381,N_3184);
or U3641 (N_3641,N_3022,N_3108);
or U3642 (N_3642,N_3349,N_3100);
nand U3643 (N_3643,N_3177,N_3047);
and U3644 (N_3644,N_3067,N_3468);
nor U3645 (N_3645,N_3368,N_3197);
nand U3646 (N_3646,N_3135,N_3140);
nor U3647 (N_3647,N_3433,N_3286);
nor U3648 (N_3648,N_3124,N_3279);
nand U3649 (N_3649,N_3359,N_3399);
nand U3650 (N_3650,N_3160,N_3170);
nand U3651 (N_3651,N_3472,N_3482);
or U3652 (N_3652,N_3303,N_3269);
nor U3653 (N_3653,N_3465,N_3027);
xor U3654 (N_3654,N_3181,N_3270);
or U3655 (N_3655,N_3409,N_3329);
nor U3656 (N_3656,N_3092,N_3064);
and U3657 (N_3657,N_3083,N_3446);
or U3658 (N_3658,N_3230,N_3330);
nor U3659 (N_3659,N_3280,N_3344);
nand U3660 (N_3660,N_3119,N_3028);
nand U3661 (N_3661,N_3214,N_3354);
or U3662 (N_3662,N_3168,N_3261);
nand U3663 (N_3663,N_3264,N_3019);
xor U3664 (N_3664,N_3337,N_3362);
or U3665 (N_3665,N_3389,N_3071);
and U3666 (N_3666,N_3396,N_3098);
nand U3667 (N_3667,N_3007,N_3130);
nor U3668 (N_3668,N_3127,N_3102);
or U3669 (N_3669,N_3497,N_3133);
or U3670 (N_3670,N_3495,N_3415);
and U3671 (N_3671,N_3281,N_3201);
nand U3672 (N_3672,N_3371,N_3439);
and U3673 (N_3673,N_3225,N_3301);
nor U3674 (N_3674,N_3401,N_3030);
and U3675 (N_3675,N_3378,N_3158);
xor U3676 (N_3676,N_3431,N_3228);
and U3677 (N_3677,N_3188,N_3494);
nor U3678 (N_3678,N_3208,N_3392);
and U3679 (N_3679,N_3010,N_3256);
xor U3680 (N_3680,N_3434,N_3189);
and U3681 (N_3681,N_3463,N_3326);
and U3682 (N_3682,N_3153,N_3057);
nand U3683 (N_3683,N_3167,N_3221);
and U3684 (N_3684,N_3185,N_3380);
or U3685 (N_3685,N_3346,N_3103);
nor U3686 (N_3686,N_3473,N_3126);
and U3687 (N_3687,N_3196,N_3089);
nand U3688 (N_3688,N_3210,N_3265);
nor U3689 (N_3689,N_3162,N_3332);
xnor U3690 (N_3690,N_3287,N_3447);
and U3691 (N_3691,N_3427,N_3125);
nand U3692 (N_3692,N_3418,N_3137);
nor U3693 (N_3693,N_3429,N_3212);
nand U3694 (N_3694,N_3150,N_3260);
and U3695 (N_3695,N_3293,N_3496);
nand U3696 (N_3696,N_3091,N_3118);
and U3697 (N_3697,N_3213,N_3094);
xor U3698 (N_3698,N_3366,N_3051);
xor U3699 (N_3699,N_3499,N_3259);
or U3700 (N_3700,N_3106,N_3075);
or U3701 (N_3701,N_3410,N_3379);
xnor U3702 (N_3702,N_3026,N_3298);
nand U3703 (N_3703,N_3002,N_3388);
nor U3704 (N_3704,N_3006,N_3154);
nor U3705 (N_3705,N_3382,N_3417);
nor U3706 (N_3706,N_3341,N_3151);
xor U3707 (N_3707,N_3088,N_3453);
xnor U3708 (N_3708,N_3412,N_3414);
and U3709 (N_3709,N_3084,N_3373);
or U3710 (N_3710,N_3244,N_3266);
or U3711 (N_3711,N_3031,N_3271);
nor U3712 (N_3712,N_3090,N_3132);
nand U3713 (N_3713,N_3070,N_3365);
or U3714 (N_3714,N_3268,N_3313);
nor U3715 (N_3715,N_3009,N_3469);
and U3716 (N_3716,N_3238,N_3436);
nand U3717 (N_3717,N_3476,N_3008);
or U3718 (N_3718,N_3234,N_3248);
nor U3719 (N_3719,N_3334,N_3131);
nor U3720 (N_3720,N_3374,N_3317);
nor U3721 (N_3721,N_3240,N_3328);
or U3722 (N_3722,N_3226,N_3110);
nor U3723 (N_3723,N_3490,N_3032);
nor U3724 (N_3724,N_3443,N_3023);
nor U3725 (N_3725,N_3087,N_3262);
nor U3726 (N_3726,N_3440,N_3243);
or U3727 (N_3727,N_3295,N_3253);
or U3728 (N_3728,N_3300,N_3452);
and U3729 (N_3729,N_3169,N_3054);
xnor U3730 (N_3730,N_3222,N_3178);
nor U3731 (N_3731,N_3175,N_3107);
nor U3732 (N_3732,N_3227,N_3342);
xnor U3733 (N_3733,N_3478,N_3037);
and U3734 (N_3734,N_3314,N_3467);
and U3735 (N_3735,N_3304,N_3274);
and U3736 (N_3736,N_3475,N_3292);
nor U3737 (N_3737,N_3423,N_3186);
nand U3738 (N_3738,N_3321,N_3384);
nand U3739 (N_3739,N_3345,N_3001);
and U3740 (N_3740,N_3004,N_3122);
nand U3741 (N_3741,N_3386,N_3460);
xor U3742 (N_3742,N_3347,N_3319);
nor U3743 (N_3743,N_3288,N_3306);
or U3744 (N_3744,N_3144,N_3199);
nand U3745 (N_3745,N_3072,N_3487);
nor U3746 (N_3746,N_3038,N_3489);
nor U3747 (N_3747,N_3267,N_3367);
xnor U3748 (N_3748,N_3105,N_3311);
nor U3749 (N_3749,N_3236,N_3129);
nand U3750 (N_3750,N_3224,N_3250);
nor U3751 (N_3751,N_3277,N_3274);
nor U3752 (N_3752,N_3142,N_3011);
xor U3753 (N_3753,N_3168,N_3363);
or U3754 (N_3754,N_3054,N_3157);
or U3755 (N_3755,N_3372,N_3247);
nor U3756 (N_3756,N_3223,N_3251);
nor U3757 (N_3757,N_3263,N_3126);
xnor U3758 (N_3758,N_3460,N_3145);
nor U3759 (N_3759,N_3275,N_3331);
and U3760 (N_3760,N_3129,N_3052);
and U3761 (N_3761,N_3360,N_3126);
xnor U3762 (N_3762,N_3059,N_3226);
nor U3763 (N_3763,N_3061,N_3008);
nor U3764 (N_3764,N_3269,N_3097);
or U3765 (N_3765,N_3392,N_3496);
xnor U3766 (N_3766,N_3399,N_3156);
nand U3767 (N_3767,N_3345,N_3479);
or U3768 (N_3768,N_3106,N_3453);
and U3769 (N_3769,N_3466,N_3099);
xnor U3770 (N_3770,N_3115,N_3489);
and U3771 (N_3771,N_3385,N_3020);
and U3772 (N_3772,N_3223,N_3429);
nor U3773 (N_3773,N_3014,N_3188);
and U3774 (N_3774,N_3035,N_3070);
and U3775 (N_3775,N_3297,N_3427);
nor U3776 (N_3776,N_3036,N_3035);
xnor U3777 (N_3777,N_3413,N_3395);
nand U3778 (N_3778,N_3333,N_3046);
nor U3779 (N_3779,N_3085,N_3313);
xor U3780 (N_3780,N_3432,N_3073);
nand U3781 (N_3781,N_3476,N_3455);
or U3782 (N_3782,N_3235,N_3252);
and U3783 (N_3783,N_3133,N_3196);
nor U3784 (N_3784,N_3492,N_3441);
nand U3785 (N_3785,N_3290,N_3330);
and U3786 (N_3786,N_3243,N_3435);
or U3787 (N_3787,N_3267,N_3005);
and U3788 (N_3788,N_3433,N_3424);
xor U3789 (N_3789,N_3152,N_3183);
and U3790 (N_3790,N_3033,N_3475);
or U3791 (N_3791,N_3207,N_3100);
or U3792 (N_3792,N_3115,N_3260);
or U3793 (N_3793,N_3375,N_3244);
or U3794 (N_3794,N_3312,N_3089);
and U3795 (N_3795,N_3304,N_3346);
nand U3796 (N_3796,N_3160,N_3440);
or U3797 (N_3797,N_3362,N_3136);
nor U3798 (N_3798,N_3490,N_3190);
nor U3799 (N_3799,N_3334,N_3053);
nor U3800 (N_3800,N_3371,N_3249);
xor U3801 (N_3801,N_3319,N_3320);
or U3802 (N_3802,N_3043,N_3013);
xor U3803 (N_3803,N_3154,N_3379);
or U3804 (N_3804,N_3018,N_3250);
nand U3805 (N_3805,N_3033,N_3395);
and U3806 (N_3806,N_3395,N_3346);
or U3807 (N_3807,N_3243,N_3475);
nor U3808 (N_3808,N_3097,N_3056);
or U3809 (N_3809,N_3426,N_3490);
nor U3810 (N_3810,N_3191,N_3076);
nand U3811 (N_3811,N_3398,N_3016);
xor U3812 (N_3812,N_3409,N_3352);
nor U3813 (N_3813,N_3414,N_3142);
and U3814 (N_3814,N_3302,N_3198);
or U3815 (N_3815,N_3404,N_3054);
nor U3816 (N_3816,N_3204,N_3009);
or U3817 (N_3817,N_3350,N_3338);
or U3818 (N_3818,N_3328,N_3048);
or U3819 (N_3819,N_3309,N_3111);
nor U3820 (N_3820,N_3352,N_3035);
and U3821 (N_3821,N_3353,N_3395);
xnor U3822 (N_3822,N_3266,N_3443);
nor U3823 (N_3823,N_3091,N_3042);
and U3824 (N_3824,N_3477,N_3416);
or U3825 (N_3825,N_3344,N_3112);
nor U3826 (N_3826,N_3008,N_3077);
or U3827 (N_3827,N_3338,N_3169);
xor U3828 (N_3828,N_3335,N_3080);
nand U3829 (N_3829,N_3180,N_3327);
or U3830 (N_3830,N_3246,N_3302);
xnor U3831 (N_3831,N_3153,N_3371);
or U3832 (N_3832,N_3195,N_3307);
or U3833 (N_3833,N_3201,N_3198);
or U3834 (N_3834,N_3487,N_3133);
nand U3835 (N_3835,N_3168,N_3054);
or U3836 (N_3836,N_3004,N_3324);
xnor U3837 (N_3837,N_3403,N_3380);
and U3838 (N_3838,N_3435,N_3381);
xnor U3839 (N_3839,N_3389,N_3140);
nor U3840 (N_3840,N_3334,N_3492);
and U3841 (N_3841,N_3364,N_3059);
and U3842 (N_3842,N_3349,N_3218);
xnor U3843 (N_3843,N_3225,N_3486);
nand U3844 (N_3844,N_3111,N_3356);
xnor U3845 (N_3845,N_3371,N_3072);
nor U3846 (N_3846,N_3306,N_3187);
and U3847 (N_3847,N_3438,N_3400);
nor U3848 (N_3848,N_3361,N_3306);
or U3849 (N_3849,N_3131,N_3280);
nand U3850 (N_3850,N_3339,N_3188);
and U3851 (N_3851,N_3367,N_3431);
nand U3852 (N_3852,N_3370,N_3127);
nand U3853 (N_3853,N_3149,N_3051);
xnor U3854 (N_3854,N_3136,N_3025);
and U3855 (N_3855,N_3109,N_3386);
xnor U3856 (N_3856,N_3449,N_3241);
nand U3857 (N_3857,N_3140,N_3390);
xnor U3858 (N_3858,N_3018,N_3191);
nor U3859 (N_3859,N_3238,N_3282);
nand U3860 (N_3860,N_3165,N_3196);
nor U3861 (N_3861,N_3487,N_3114);
or U3862 (N_3862,N_3249,N_3480);
or U3863 (N_3863,N_3078,N_3150);
or U3864 (N_3864,N_3033,N_3267);
or U3865 (N_3865,N_3319,N_3384);
or U3866 (N_3866,N_3170,N_3250);
nand U3867 (N_3867,N_3048,N_3185);
and U3868 (N_3868,N_3074,N_3080);
nand U3869 (N_3869,N_3436,N_3499);
nand U3870 (N_3870,N_3068,N_3367);
nand U3871 (N_3871,N_3260,N_3459);
xnor U3872 (N_3872,N_3368,N_3233);
nand U3873 (N_3873,N_3287,N_3215);
and U3874 (N_3874,N_3271,N_3383);
nor U3875 (N_3875,N_3328,N_3273);
and U3876 (N_3876,N_3205,N_3019);
nor U3877 (N_3877,N_3403,N_3363);
nor U3878 (N_3878,N_3112,N_3432);
nor U3879 (N_3879,N_3296,N_3161);
nor U3880 (N_3880,N_3010,N_3002);
or U3881 (N_3881,N_3288,N_3113);
or U3882 (N_3882,N_3107,N_3200);
nand U3883 (N_3883,N_3174,N_3195);
nor U3884 (N_3884,N_3377,N_3112);
nor U3885 (N_3885,N_3044,N_3435);
nor U3886 (N_3886,N_3300,N_3188);
nand U3887 (N_3887,N_3189,N_3474);
or U3888 (N_3888,N_3081,N_3080);
and U3889 (N_3889,N_3365,N_3469);
xnor U3890 (N_3890,N_3041,N_3289);
xor U3891 (N_3891,N_3427,N_3114);
and U3892 (N_3892,N_3097,N_3197);
or U3893 (N_3893,N_3047,N_3018);
nand U3894 (N_3894,N_3499,N_3458);
and U3895 (N_3895,N_3152,N_3393);
xor U3896 (N_3896,N_3138,N_3380);
or U3897 (N_3897,N_3113,N_3471);
and U3898 (N_3898,N_3326,N_3055);
or U3899 (N_3899,N_3048,N_3409);
or U3900 (N_3900,N_3098,N_3376);
nand U3901 (N_3901,N_3270,N_3335);
or U3902 (N_3902,N_3332,N_3192);
and U3903 (N_3903,N_3291,N_3015);
nor U3904 (N_3904,N_3137,N_3201);
nand U3905 (N_3905,N_3426,N_3306);
or U3906 (N_3906,N_3315,N_3235);
or U3907 (N_3907,N_3001,N_3399);
nor U3908 (N_3908,N_3241,N_3076);
or U3909 (N_3909,N_3265,N_3380);
xor U3910 (N_3910,N_3246,N_3286);
or U3911 (N_3911,N_3433,N_3185);
nor U3912 (N_3912,N_3182,N_3189);
nor U3913 (N_3913,N_3207,N_3162);
nor U3914 (N_3914,N_3477,N_3024);
nor U3915 (N_3915,N_3457,N_3181);
nor U3916 (N_3916,N_3266,N_3497);
xor U3917 (N_3917,N_3308,N_3213);
or U3918 (N_3918,N_3032,N_3104);
nand U3919 (N_3919,N_3495,N_3305);
nand U3920 (N_3920,N_3278,N_3478);
nand U3921 (N_3921,N_3425,N_3222);
nor U3922 (N_3922,N_3269,N_3201);
nand U3923 (N_3923,N_3276,N_3288);
nand U3924 (N_3924,N_3384,N_3478);
nor U3925 (N_3925,N_3330,N_3320);
and U3926 (N_3926,N_3085,N_3331);
nor U3927 (N_3927,N_3176,N_3401);
xor U3928 (N_3928,N_3206,N_3293);
or U3929 (N_3929,N_3481,N_3185);
or U3930 (N_3930,N_3477,N_3226);
nand U3931 (N_3931,N_3189,N_3370);
or U3932 (N_3932,N_3049,N_3142);
or U3933 (N_3933,N_3184,N_3168);
nand U3934 (N_3934,N_3496,N_3412);
nand U3935 (N_3935,N_3349,N_3115);
nor U3936 (N_3936,N_3347,N_3131);
nor U3937 (N_3937,N_3089,N_3378);
nor U3938 (N_3938,N_3069,N_3139);
or U3939 (N_3939,N_3128,N_3089);
nand U3940 (N_3940,N_3215,N_3019);
and U3941 (N_3941,N_3347,N_3016);
nand U3942 (N_3942,N_3050,N_3315);
nand U3943 (N_3943,N_3189,N_3043);
or U3944 (N_3944,N_3452,N_3189);
nor U3945 (N_3945,N_3249,N_3334);
nand U3946 (N_3946,N_3490,N_3059);
nand U3947 (N_3947,N_3000,N_3201);
xor U3948 (N_3948,N_3334,N_3096);
or U3949 (N_3949,N_3195,N_3460);
and U3950 (N_3950,N_3117,N_3273);
or U3951 (N_3951,N_3442,N_3280);
xor U3952 (N_3952,N_3242,N_3191);
nand U3953 (N_3953,N_3155,N_3431);
nand U3954 (N_3954,N_3213,N_3369);
nand U3955 (N_3955,N_3309,N_3162);
xor U3956 (N_3956,N_3070,N_3451);
and U3957 (N_3957,N_3344,N_3100);
nand U3958 (N_3958,N_3149,N_3413);
and U3959 (N_3959,N_3404,N_3082);
nor U3960 (N_3960,N_3492,N_3130);
nand U3961 (N_3961,N_3477,N_3435);
nor U3962 (N_3962,N_3184,N_3202);
and U3963 (N_3963,N_3424,N_3205);
or U3964 (N_3964,N_3438,N_3295);
xnor U3965 (N_3965,N_3453,N_3178);
nand U3966 (N_3966,N_3489,N_3270);
nand U3967 (N_3967,N_3038,N_3369);
or U3968 (N_3968,N_3145,N_3441);
and U3969 (N_3969,N_3207,N_3006);
nor U3970 (N_3970,N_3415,N_3210);
nor U3971 (N_3971,N_3245,N_3197);
nor U3972 (N_3972,N_3068,N_3258);
and U3973 (N_3973,N_3410,N_3015);
nor U3974 (N_3974,N_3404,N_3213);
nand U3975 (N_3975,N_3329,N_3078);
nor U3976 (N_3976,N_3401,N_3451);
and U3977 (N_3977,N_3407,N_3023);
nor U3978 (N_3978,N_3056,N_3115);
and U3979 (N_3979,N_3160,N_3434);
and U3980 (N_3980,N_3330,N_3011);
nor U3981 (N_3981,N_3341,N_3174);
and U3982 (N_3982,N_3193,N_3296);
nor U3983 (N_3983,N_3466,N_3461);
or U3984 (N_3984,N_3192,N_3308);
nand U3985 (N_3985,N_3256,N_3228);
nor U3986 (N_3986,N_3132,N_3342);
or U3987 (N_3987,N_3408,N_3136);
and U3988 (N_3988,N_3009,N_3489);
and U3989 (N_3989,N_3078,N_3265);
nand U3990 (N_3990,N_3100,N_3306);
nand U3991 (N_3991,N_3336,N_3476);
or U3992 (N_3992,N_3160,N_3419);
nor U3993 (N_3993,N_3268,N_3324);
nand U3994 (N_3994,N_3248,N_3433);
xnor U3995 (N_3995,N_3063,N_3244);
xor U3996 (N_3996,N_3098,N_3246);
or U3997 (N_3997,N_3287,N_3016);
xnor U3998 (N_3998,N_3127,N_3232);
or U3999 (N_3999,N_3016,N_3231);
and U4000 (N_4000,N_3792,N_3715);
or U4001 (N_4001,N_3742,N_3837);
and U4002 (N_4002,N_3842,N_3761);
nor U4003 (N_4003,N_3689,N_3936);
or U4004 (N_4004,N_3789,N_3935);
and U4005 (N_4005,N_3802,N_3850);
nor U4006 (N_4006,N_3696,N_3815);
nand U4007 (N_4007,N_3757,N_3708);
nor U4008 (N_4008,N_3739,N_3680);
nor U4009 (N_4009,N_3740,N_3533);
nor U4010 (N_4010,N_3748,N_3526);
and U4011 (N_4011,N_3623,N_3738);
and U4012 (N_4012,N_3671,N_3774);
and U4013 (N_4013,N_3885,N_3890);
or U4014 (N_4014,N_3556,N_3867);
and U4015 (N_4015,N_3956,N_3636);
nand U4016 (N_4016,N_3955,N_3871);
nand U4017 (N_4017,N_3522,N_3627);
or U4018 (N_4018,N_3690,N_3781);
nor U4019 (N_4019,N_3506,N_3662);
or U4020 (N_4020,N_3787,N_3704);
or U4021 (N_4021,N_3967,N_3628);
nor U4022 (N_4022,N_3863,N_3713);
nand U4023 (N_4023,N_3812,N_3679);
nor U4024 (N_4024,N_3992,N_3917);
nor U4025 (N_4025,N_3879,N_3737);
nand U4026 (N_4026,N_3640,N_3675);
nand U4027 (N_4027,N_3509,N_3869);
nor U4028 (N_4028,N_3559,N_3818);
nand U4029 (N_4029,N_3809,N_3805);
xor U4030 (N_4030,N_3940,N_3898);
nor U4031 (N_4031,N_3540,N_3843);
and U4032 (N_4032,N_3702,N_3845);
nor U4033 (N_4033,N_3865,N_3545);
or U4034 (N_4034,N_3548,N_3839);
nor U4035 (N_4035,N_3648,N_3614);
nand U4036 (N_4036,N_3693,N_3705);
or U4037 (N_4037,N_3606,N_3771);
nand U4038 (N_4038,N_3797,N_3870);
nand U4039 (N_4039,N_3767,N_3510);
nand U4040 (N_4040,N_3605,N_3560);
and U4041 (N_4041,N_3552,N_3999);
and U4042 (N_4042,N_3504,N_3663);
xor U4043 (N_4043,N_3562,N_3779);
and U4044 (N_4044,N_3905,N_3523);
and U4045 (N_4045,N_3672,N_3727);
xor U4046 (N_4046,N_3983,N_3601);
and U4047 (N_4047,N_3951,N_3794);
nand U4048 (N_4048,N_3859,N_3777);
and U4049 (N_4049,N_3883,N_3884);
or U4050 (N_4050,N_3546,N_3827);
nand U4051 (N_4051,N_3780,N_3950);
and U4052 (N_4052,N_3847,N_3961);
xnor U4053 (N_4053,N_3946,N_3891);
nor U4054 (N_4054,N_3996,N_3778);
or U4055 (N_4055,N_3635,N_3751);
nand U4056 (N_4056,N_3590,N_3563);
nand U4057 (N_4057,N_3800,N_3776);
or U4058 (N_4058,N_3927,N_3531);
and U4059 (N_4059,N_3592,N_3821);
xor U4060 (N_4060,N_3529,N_3993);
and U4061 (N_4061,N_3834,N_3527);
nand U4062 (N_4062,N_3670,N_3652);
xor U4063 (N_4063,N_3989,N_3581);
and U4064 (N_4064,N_3641,N_3997);
nand U4065 (N_4065,N_3906,N_3622);
nand U4066 (N_4066,N_3939,N_3578);
nor U4067 (N_4067,N_3889,N_3991);
nor U4068 (N_4068,N_3784,N_3686);
nand U4069 (N_4069,N_3613,N_3788);
or U4070 (N_4070,N_3785,N_3550);
nand U4071 (N_4071,N_3579,N_3571);
or U4072 (N_4072,N_3979,N_3683);
nor U4073 (N_4073,N_3593,N_3897);
nor U4074 (N_4074,N_3574,N_3920);
nor U4075 (N_4075,N_3799,N_3942);
or U4076 (N_4076,N_3624,N_3908);
and U4077 (N_4077,N_3512,N_3654);
nand U4078 (N_4078,N_3911,N_3912);
nor U4079 (N_4079,N_3749,N_3852);
and U4080 (N_4080,N_3882,N_3822);
or U4081 (N_4081,N_3710,N_3820);
nand U4082 (N_4082,N_3895,N_3591);
and U4083 (N_4083,N_3669,N_3975);
or U4084 (N_4084,N_3611,N_3846);
or U4085 (N_4085,N_3528,N_3625);
nand U4086 (N_4086,N_3661,N_3549);
or U4087 (N_4087,N_3734,N_3832);
xnor U4088 (N_4088,N_3860,N_3568);
nand U4089 (N_4089,N_3658,N_3602);
xor U4090 (N_4090,N_3886,N_3730);
nor U4091 (N_4091,N_3765,N_3947);
nor U4092 (N_4092,N_3914,N_3646);
and U4093 (N_4093,N_3970,N_3726);
and U4094 (N_4094,N_3915,N_3577);
and U4095 (N_4095,N_3554,N_3985);
nor U4096 (N_4096,N_3618,N_3828);
nor U4097 (N_4097,N_3925,N_3616);
nor U4098 (N_4098,N_3836,N_3513);
nor U4099 (N_4099,N_3877,N_3644);
or U4100 (N_4100,N_3878,N_3651);
nand U4101 (N_4101,N_3858,N_3630);
and U4102 (N_4102,N_3535,N_3746);
or U4103 (N_4103,N_3678,N_3698);
nand U4104 (N_4104,N_3561,N_3755);
xor U4105 (N_4105,N_3586,N_3995);
nor U4106 (N_4106,N_3949,N_3733);
nor U4107 (N_4107,N_3638,N_3724);
and U4108 (N_4108,N_3501,N_3966);
nor U4109 (N_4109,N_3524,N_3544);
nand U4110 (N_4110,N_3539,N_3933);
nand U4111 (N_4111,N_3918,N_3609);
xor U4112 (N_4112,N_3823,N_3572);
and U4113 (N_4113,N_3584,N_3945);
or U4114 (N_4114,N_3982,N_3600);
or U4115 (N_4115,N_3718,N_3875);
or U4116 (N_4116,N_3538,N_3758);
nand U4117 (N_4117,N_3585,N_3928);
and U4118 (N_4118,N_3866,N_3987);
or U4119 (N_4119,N_3965,N_3876);
or U4120 (N_4120,N_3707,N_3807);
nor U4121 (N_4121,N_3768,N_3924);
and U4122 (N_4122,N_3634,N_3954);
and U4123 (N_4123,N_3732,N_3854);
nand U4124 (N_4124,N_3717,N_3621);
nor U4125 (N_4125,N_3864,N_3551);
and U4126 (N_4126,N_3682,N_3676);
nand U4127 (N_4127,N_3811,N_3608);
or U4128 (N_4128,N_3804,N_3857);
xnor U4129 (N_4129,N_3547,N_3824);
nor U4130 (N_4130,N_3971,N_3555);
and U4131 (N_4131,N_3931,N_3597);
nand U4132 (N_4132,N_3753,N_3817);
or U4133 (N_4133,N_3957,N_3507);
xor U4134 (N_4134,N_3830,N_3849);
and U4135 (N_4135,N_3673,N_3813);
or U4136 (N_4136,N_3716,N_3786);
nor U4137 (N_4137,N_3534,N_3791);
nand U4138 (N_4138,N_3978,N_3626);
nor U4139 (N_4139,N_3948,N_3720);
nor U4140 (N_4140,N_3894,N_3903);
xor U4141 (N_4141,N_3964,N_3573);
nor U4142 (N_4142,N_3750,N_3969);
nor U4143 (N_4143,N_3731,N_3598);
or U4144 (N_4144,N_3582,N_3632);
and U4145 (N_4145,N_3566,N_3976);
nor U4146 (N_4146,N_3580,N_3760);
or U4147 (N_4147,N_3610,N_3517);
nand U4148 (N_4148,N_3902,N_3612);
nand U4149 (N_4149,N_3576,N_3930);
or U4150 (N_4150,N_3503,N_3831);
xor U4151 (N_4151,N_3943,N_3844);
nor U4152 (N_4152,N_3558,N_3639);
nor U4153 (N_4153,N_3694,N_3688);
and U4154 (N_4154,N_3910,N_3629);
nor U4155 (N_4155,N_3922,N_3505);
and U4156 (N_4156,N_3773,N_3667);
and U4157 (N_4157,N_3692,N_3594);
or U4158 (N_4158,N_3806,N_3620);
nor U4159 (N_4159,N_3656,N_3814);
and U4160 (N_4160,N_3972,N_3793);
or U4161 (N_4161,N_3981,N_3744);
nor U4162 (N_4162,N_3599,N_3783);
or U4163 (N_4163,N_3596,N_3557);
or U4164 (N_4164,N_3685,N_3570);
nand U4165 (N_4165,N_3643,N_3988);
xnor U4166 (N_4166,N_3838,N_3714);
nor U4167 (N_4167,N_3994,N_3699);
nand U4168 (N_4168,N_3703,N_3500);
or U4169 (N_4169,N_3722,N_3587);
and U4170 (N_4170,N_3650,N_3901);
or U4171 (N_4171,N_3665,N_3808);
and U4172 (N_4172,N_3926,N_3937);
and U4173 (N_4173,N_3615,N_3759);
and U4174 (N_4174,N_3681,N_3769);
xnor U4175 (N_4175,N_3916,N_3896);
or U4176 (N_4176,N_3525,N_3923);
nand U4177 (N_4177,N_3810,N_3941);
or U4178 (N_4178,N_3677,N_3874);
xnor U4179 (N_4179,N_3893,N_3660);
or U4180 (N_4180,N_3984,N_3511);
nor U4181 (N_4181,N_3856,N_3973);
or U4182 (N_4182,N_3762,N_3655);
nor U4183 (N_4183,N_3887,N_3537);
or U4184 (N_4184,N_3633,N_3960);
or U4185 (N_4185,N_3674,N_3637);
and U4186 (N_4186,N_3723,N_3645);
and U4187 (N_4187,N_3521,N_3795);
nor U4188 (N_4188,N_3881,N_3880);
nand U4189 (N_4189,N_3900,N_3701);
and U4190 (N_4190,N_3861,N_3706);
nand U4191 (N_4191,N_3642,N_3790);
xnor U4192 (N_4192,N_3841,N_3873);
nor U4193 (N_4193,N_3741,N_3607);
xor U4194 (N_4194,N_3711,N_3721);
nor U4195 (N_4195,N_3938,N_3868);
nand U4196 (N_4196,N_3929,N_3958);
or U4197 (N_4197,N_3803,N_3668);
or U4198 (N_4198,N_3840,N_3653);
nor U4199 (N_4199,N_3588,N_3567);
nand U4200 (N_4200,N_3855,N_3801);
nand U4201 (N_4201,N_3743,N_3872);
and U4202 (N_4202,N_3959,N_3819);
nor U4203 (N_4203,N_3968,N_3709);
xnor U4204 (N_4204,N_3649,N_3853);
and U4205 (N_4205,N_3775,N_3851);
nand U4206 (N_4206,N_3745,N_3664);
or U4207 (N_4207,N_3536,N_3725);
nor U4208 (N_4208,N_3617,N_3862);
nor U4209 (N_4209,N_3729,N_3833);
nor U4210 (N_4210,N_3691,N_3892);
nor U4211 (N_4211,N_3754,N_3520);
and U4212 (N_4212,N_3974,N_3657);
nor U4213 (N_4213,N_3532,N_3909);
nand U4214 (N_4214,N_3565,N_3595);
nor U4215 (N_4215,N_3583,N_3932);
and U4216 (N_4216,N_3604,N_3747);
nor U4217 (N_4217,N_3719,N_3603);
or U4218 (N_4218,N_3904,N_3763);
xnor U4219 (N_4219,N_3921,N_3736);
nand U4220 (N_4220,N_3835,N_3515);
nor U4221 (N_4221,N_3728,N_3756);
and U4222 (N_4222,N_3953,N_3919);
or U4223 (N_4223,N_3772,N_3508);
or U4224 (N_4224,N_3543,N_3986);
and U4225 (N_4225,N_3735,N_3564);
and U4226 (N_4226,N_3825,N_3990);
nand U4227 (N_4227,N_3829,N_3687);
and U4228 (N_4228,N_3944,N_3766);
or U4229 (N_4229,N_3977,N_3848);
or U4230 (N_4230,N_3619,N_3659);
xnor U4231 (N_4231,N_3575,N_3569);
nand U4232 (N_4232,N_3518,N_3684);
nor U4233 (N_4233,N_3782,N_3695);
nor U4234 (N_4234,N_3963,N_3952);
and U4235 (N_4235,N_3516,N_3796);
and U4236 (N_4236,N_3980,N_3700);
or U4237 (N_4237,N_3764,N_3553);
or U4238 (N_4238,N_3752,N_3712);
nand U4239 (N_4239,N_3998,N_3647);
nor U4240 (N_4240,N_3888,N_3530);
nand U4241 (N_4241,N_3913,N_3798);
nand U4242 (N_4242,N_3934,N_3666);
or U4243 (N_4243,N_3697,N_3899);
nor U4244 (N_4244,N_3542,N_3907);
nand U4245 (N_4245,N_3589,N_3816);
nor U4246 (N_4246,N_3826,N_3962);
nor U4247 (N_4247,N_3770,N_3631);
and U4248 (N_4248,N_3514,N_3502);
or U4249 (N_4249,N_3541,N_3519);
or U4250 (N_4250,N_3963,N_3572);
nor U4251 (N_4251,N_3849,N_3804);
nor U4252 (N_4252,N_3852,N_3874);
and U4253 (N_4253,N_3693,N_3930);
and U4254 (N_4254,N_3915,N_3728);
or U4255 (N_4255,N_3829,N_3895);
or U4256 (N_4256,N_3614,N_3852);
nor U4257 (N_4257,N_3953,N_3718);
and U4258 (N_4258,N_3642,N_3529);
nor U4259 (N_4259,N_3995,N_3675);
or U4260 (N_4260,N_3936,N_3865);
and U4261 (N_4261,N_3761,N_3718);
or U4262 (N_4262,N_3759,N_3519);
and U4263 (N_4263,N_3617,N_3681);
xnor U4264 (N_4264,N_3879,N_3565);
nor U4265 (N_4265,N_3778,N_3695);
and U4266 (N_4266,N_3751,N_3514);
or U4267 (N_4267,N_3523,N_3619);
nand U4268 (N_4268,N_3668,N_3880);
nor U4269 (N_4269,N_3527,N_3565);
and U4270 (N_4270,N_3507,N_3704);
xnor U4271 (N_4271,N_3633,N_3675);
and U4272 (N_4272,N_3573,N_3750);
nand U4273 (N_4273,N_3552,N_3637);
and U4274 (N_4274,N_3698,N_3918);
or U4275 (N_4275,N_3989,N_3709);
and U4276 (N_4276,N_3914,N_3718);
nand U4277 (N_4277,N_3624,N_3786);
xor U4278 (N_4278,N_3944,N_3856);
nor U4279 (N_4279,N_3756,N_3892);
nor U4280 (N_4280,N_3671,N_3616);
and U4281 (N_4281,N_3924,N_3998);
nor U4282 (N_4282,N_3681,N_3646);
nand U4283 (N_4283,N_3553,N_3651);
or U4284 (N_4284,N_3763,N_3996);
nor U4285 (N_4285,N_3594,N_3655);
nand U4286 (N_4286,N_3971,N_3631);
nor U4287 (N_4287,N_3873,N_3705);
nor U4288 (N_4288,N_3576,N_3917);
nor U4289 (N_4289,N_3961,N_3951);
and U4290 (N_4290,N_3636,N_3600);
nand U4291 (N_4291,N_3846,N_3527);
and U4292 (N_4292,N_3577,N_3971);
nand U4293 (N_4293,N_3965,N_3668);
or U4294 (N_4294,N_3958,N_3985);
or U4295 (N_4295,N_3648,N_3533);
nand U4296 (N_4296,N_3592,N_3600);
nor U4297 (N_4297,N_3524,N_3782);
or U4298 (N_4298,N_3598,N_3748);
and U4299 (N_4299,N_3961,N_3647);
and U4300 (N_4300,N_3824,N_3871);
nand U4301 (N_4301,N_3712,N_3605);
xnor U4302 (N_4302,N_3989,N_3995);
nand U4303 (N_4303,N_3680,N_3658);
and U4304 (N_4304,N_3939,N_3692);
xnor U4305 (N_4305,N_3624,N_3651);
nand U4306 (N_4306,N_3626,N_3727);
nor U4307 (N_4307,N_3658,N_3598);
and U4308 (N_4308,N_3648,N_3967);
nand U4309 (N_4309,N_3900,N_3555);
and U4310 (N_4310,N_3713,N_3583);
or U4311 (N_4311,N_3965,N_3977);
nor U4312 (N_4312,N_3858,N_3879);
nand U4313 (N_4313,N_3536,N_3841);
and U4314 (N_4314,N_3997,N_3559);
xnor U4315 (N_4315,N_3652,N_3565);
nand U4316 (N_4316,N_3893,N_3553);
nor U4317 (N_4317,N_3603,N_3787);
nand U4318 (N_4318,N_3661,N_3648);
xor U4319 (N_4319,N_3525,N_3538);
nor U4320 (N_4320,N_3885,N_3948);
or U4321 (N_4321,N_3721,N_3914);
xnor U4322 (N_4322,N_3576,N_3718);
nor U4323 (N_4323,N_3539,N_3964);
and U4324 (N_4324,N_3924,N_3999);
nand U4325 (N_4325,N_3912,N_3724);
nor U4326 (N_4326,N_3862,N_3930);
nand U4327 (N_4327,N_3770,N_3526);
or U4328 (N_4328,N_3990,N_3965);
nor U4329 (N_4329,N_3979,N_3922);
nor U4330 (N_4330,N_3585,N_3838);
or U4331 (N_4331,N_3675,N_3521);
nor U4332 (N_4332,N_3510,N_3615);
xnor U4333 (N_4333,N_3900,N_3657);
nor U4334 (N_4334,N_3977,N_3916);
or U4335 (N_4335,N_3939,N_3638);
nand U4336 (N_4336,N_3799,N_3780);
nand U4337 (N_4337,N_3606,N_3531);
and U4338 (N_4338,N_3753,N_3799);
xnor U4339 (N_4339,N_3596,N_3641);
nor U4340 (N_4340,N_3631,N_3757);
nor U4341 (N_4341,N_3965,N_3738);
nand U4342 (N_4342,N_3682,N_3816);
or U4343 (N_4343,N_3816,N_3982);
nor U4344 (N_4344,N_3997,N_3678);
and U4345 (N_4345,N_3529,N_3882);
or U4346 (N_4346,N_3703,N_3646);
or U4347 (N_4347,N_3937,N_3503);
xnor U4348 (N_4348,N_3579,N_3975);
nor U4349 (N_4349,N_3586,N_3993);
and U4350 (N_4350,N_3586,N_3566);
xor U4351 (N_4351,N_3598,N_3673);
nor U4352 (N_4352,N_3550,N_3906);
xnor U4353 (N_4353,N_3697,N_3647);
and U4354 (N_4354,N_3945,N_3844);
or U4355 (N_4355,N_3552,N_3731);
or U4356 (N_4356,N_3581,N_3585);
and U4357 (N_4357,N_3955,N_3896);
nor U4358 (N_4358,N_3784,N_3993);
nand U4359 (N_4359,N_3509,N_3741);
nor U4360 (N_4360,N_3625,N_3898);
and U4361 (N_4361,N_3631,N_3613);
or U4362 (N_4362,N_3842,N_3845);
xnor U4363 (N_4363,N_3767,N_3806);
xor U4364 (N_4364,N_3804,N_3924);
or U4365 (N_4365,N_3979,N_3853);
and U4366 (N_4366,N_3730,N_3622);
nor U4367 (N_4367,N_3833,N_3755);
and U4368 (N_4368,N_3537,N_3703);
nand U4369 (N_4369,N_3710,N_3974);
or U4370 (N_4370,N_3820,N_3907);
nor U4371 (N_4371,N_3920,N_3747);
and U4372 (N_4372,N_3572,N_3777);
nand U4373 (N_4373,N_3630,N_3685);
and U4374 (N_4374,N_3822,N_3826);
xor U4375 (N_4375,N_3963,N_3696);
nor U4376 (N_4376,N_3731,N_3829);
or U4377 (N_4377,N_3815,N_3699);
nor U4378 (N_4378,N_3704,N_3655);
nor U4379 (N_4379,N_3756,N_3747);
and U4380 (N_4380,N_3655,N_3854);
nand U4381 (N_4381,N_3845,N_3569);
nor U4382 (N_4382,N_3915,N_3774);
nand U4383 (N_4383,N_3849,N_3988);
xor U4384 (N_4384,N_3807,N_3927);
nor U4385 (N_4385,N_3862,N_3840);
and U4386 (N_4386,N_3709,N_3531);
or U4387 (N_4387,N_3785,N_3852);
or U4388 (N_4388,N_3660,N_3706);
nand U4389 (N_4389,N_3812,N_3897);
or U4390 (N_4390,N_3585,N_3543);
or U4391 (N_4391,N_3581,N_3923);
or U4392 (N_4392,N_3736,N_3955);
and U4393 (N_4393,N_3898,N_3548);
nor U4394 (N_4394,N_3838,N_3776);
nor U4395 (N_4395,N_3682,N_3907);
or U4396 (N_4396,N_3933,N_3782);
nand U4397 (N_4397,N_3872,N_3693);
and U4398 (N_4398,N_3960,N_3690);
nor U4399 (N_4399,N_3675,N_3843);
xnor U4400 (N_4400,N_3931,N_3917);
and U4401 (N_4401,N_3538,N_3969);
and U4402 (N_4402,N_3506,N_3557);
and U4403 (N_4403,N_3802,N_3522);
nand U4404 (N_4404,N_3940,N_3836);
nor U4405 (N_4405,N_3647,N_3790);
and U4406 (N_4406,N_3785,N_3716);
or U4407 (N_4407,N_3740,N_3546);
or U4408 (N_4408,N_3982,N_3568);
xnor U4409 (N_4409,N_3512,N_3710);
and U4410 (N_4410,N_3867,N_3665);
nor U4411 (N_4411,N_3766,N_3784);
nand U4412 (N_4412,N_3714,N_3901);
nand U4413 (N_4413,N_3945,N_3674);
nor U4414 (N_4414,N_3540,N_3663);
and U4415 (N_4415,N_3602,N_3918);
or U4416 (N_4416,N_3763,N_3865);
and U4417 (N_4417,N_3870,N_3722);
nor U4418 (N_4418,N_3543,N_3538);
nand U4419 (N_4419,N_3592,N_3578);
and U4420 (N_4420,N_3960,N_3934);
nand U4421 (N_4421,N_3868,N_3503);
and U4422 (N_4422,N_3732,N_3519);
xor U4423 (N_4423,N_3517,N_3655);
and U4424 (N_4424,N_3810,N_3791);
nor U4425 (N_4425,N_3963,N_3922);
and U4426 (N_4426,N_3909,N_3791);
xor U4427 (N_4427,N_3890,N_3947);
and U4428 (N_4428,N_3528,N_3907);
or U4429 (N_4429,N_3579,N_3651);
xnor U4430 (N_4430,N_3588,N_3793);
nor U4431 (N_4431,N_3833,N_3530);
or U4432 (N_4432,N_3578,N_3786);
and U4433 (N_4433,N_3787,N_3600);
and U4434 (N_4434,N_3516,N_3792);
and U4435 (N_4435,N_3716,N_3934);
nor U4436 (N_4436,N_3568,N_3729);
xor U4437 (N_4437,N_3867,N_3537);
xnor U4438 (N_4438,N_3675,N_3913);
or U4439 (N_4439,N_3995,N_3964);
or U4440 (N_4440,N_3678,N_3660);
nand U4441 (N_4441,N_3960,N_3794);
or U4442 (N_4442,N_3813,N_3626);
nor U4443 (N_4443,N_3858,N_3654);
xnor U4444 (N_4444,N_3541,N_3910);
or U4445 (N_4445,N_3892,N_3616);
nor U4446 (N_4446,N_3893,N_3984);
and U4447 (N_4447,N_3756,N_3727);
nor U4448 (N_4448,N_3924,N_3597);
and U4449 (N_4449,N_3958,N_3746);
xor U4450 (N_4450,N_3936,N_3506);
and U4451 (N_4451,N_3832,N_3923);
and U4452 (N_4452,N_3520,N_3929);
nand U4453 (N_4453,N_3922,N_3640);
and U4454 (N_4454,N_3580,N_3531);
nor U4455 (N_4455,N_3809,N_3709);
xnor U4456 (N_4456,N_3935,N_3805);
nand U4457 (N_4457,N_3965,N_3550);
or U4458 (N_4458,N_3721,N_3876);
or U4459 (N_4459,N_3546,N_3588);
or U4460 (N_4460,N_3838,N_3923);
nor U4461 (N_4461,N_3574,N_3938);
nand U4462 (N_4462,N_3788,N_3717);
nand U4463 (N_4463,N_3854,N_3819);
or U4464 (N_4464,N_3673,N_3543);
nor U4465 (N_4465,N_3738,N_3749);
and U4466 (N_4466,N_3893,N_3512);
nor U4467 (N_4467,N_3669,N_3759);
or U4468 (N_4468,N_3916,N_3772);
xnor U4469 (N_4469,N_3540,N_3613);
or U4470 (N_4470,N_3689,N_3849);
nand U4471 (N_4471,N_3565,N_3959);
and U4472 (N_4472,N_3905,N_3725);
and U4473 (N_4473,N_3545,N_3656);
or U4474 (N_4474,N_3651,N_3996);
and U4475 (N_4475,N_3913,N_3648);
nand U4476 (N_4476,N_3792,N_3934);
nand U4477 (N_4477,N_3925,N_3835);
nor U4478 (N_4478,N_3709,N_3958);
nor U4479 (N_4479,N_3744,N_3507);
nand U4480 (N_4480,N_3591,N_3734);
or U4481 (N_4481,N_3892,N_3696);
or U4482 (N_4482,N_3893,N_3867);
nand U4483 (N_4483,N_3988,N_3776);
and U4484 (N_4484,N_3878,N_3590);
nor U4485 (N_4485,N_3639,N_3672);
and U4486 (N_4486,N_3553,N_3778);
and U4487 (N_4487,N_3957,N_3881);
xnor U4488 (N_4488,N_3876,N_3880);
nor U4489 (N_4489,N_3568,N_3567);
nor U4490 (N_4490,N_3614,N_3703);
xor U4491 (N_4491,N_3623,N_3753);
nor U4492 (N_4492,N_3805,N_3996);
and U4493 (N_4493,N_3995,N_3706);
nor U4494 (N_4494,N_3848,N_3766);
nand U4495 (N_4495,N_3912,N_3881);
and U4496 (N_4496,N_3966,N_3575);
and U4497 (N_4497,N_3778,N_3878);
nand U4498 (N_4498,N_3856,N_3967);
or U4499 (N_4499,N_3695,N_3571);
xor U4500 (N_4500,N_4135,N_4349);
and U4501 (N_4501,N_4194,N_4422);
nor U4502 (N_4502,N_4230,N_4131);
or U4503 (N_4503,N_4165,N_4168);
and U4504 (N_4504,N_4035,N_4495);
and U4505 (N_4505,N_4247,N_4221);
and U4506 (N_4506,N_4460,N_4033);
or U4507 (N_4507,N_4401,N_4493);
and U4508 (N_4508,N_4072,N_4242);
xnor U4509 (N_4509,N_4152,N_4477);
or U4510 (N_4510,N_4442,N_4408);
nand U4511 (N_4511,N_4410,N_4086);
and U4512 (N_4512,N_4406,N_4133);
or U4513 (N_4513,N_4284,N_4001);
nor U4514 (N_4514,N_4107,N_4464);
and U4515 (N_4515,N_4210,N_4379);
nor U4516 (N_4516,N_4146,N_4262);
nand U4517 (N_4517,N_4090,N_4458);
nor U4518 (N_4518,N_4261,N_4164);
or U4519 (N_4519,N_4371,N_4491);
or U4520 (N_4520,N_4307,N_4201);
nand U4521 (N_4521,N_4157,N_4448);
nor U4522 (N_4522,N_4283,N_4323);
nor U4523 (N_4523,N_4004,N_4122);
and U4524 (N_4524,N_4063,N_4309);
or U4525 (N_4525,N_4368,N_4471);
or U4526 (N_4526,N_4002,N_4332);
nor U4527 (N_4527,N_4171,N_4330);
nor U4528 (N_4528,N_4156,N_4255);
xor U4529 (N_4529,N_4338,N_4182);
nor U4530 (N_4530,N_4314,N_4263);
nand U4531 (N_4531,N_4075,N_4336);
nand U4532 (N_4532,N_4062,N_4183);
nor U4533 (N_4533,N_4029,N_4364);
and U4534 (N_4534,N_4178,N_4275);
nor U4535 (N_4535,N_4048,N_4313);
nand U4536 (N_4536,N_4279,N_4097);
nand U4537 (N_4537,N_4318,N_4130);
and U4538 (N_4538,N_4119,N_4016);
nor U4539 (N_4539,N_4227,N_4038);
nor U4540 (N_4540,N_4294,N_4073);
or U4541 (N_4541,N_4274,N_4042);
nor U4542 (N_4542,N_4025,N_4374);
nor U4543 (N_4543,N_4414,N_4228);
nor U4544 (N_4544,N_4434,N_4200);
nand U4545 (N_4545,N_4158,N_4101);
nor U4546 (N_4546,N_4193,N_4118);
or U4547 (N_4547,N_4149,N_4478);
nand U4548 (N_4548,N_4304,N_4249);
nor U4549 (N_4549,N_4267,N_4077);
nor U4550 (N_4550,N_4487,N_4356);
or U4551 (N_4551,N_4189,N_4259);
and U4552 (N_4552,N_4093,N_4206);
or U4553 (N_4553,N_4079,N_4049);
or U4554 (N_4554,N_4302,N_4325);
and U4555 (N_4555,N_4316,N_4211);
and U4556 (N_4556,N_4469,N_4184);
nor U4557 (N_4557,N_4236,N_4468);
nand U4558 (N_4558,N_4011,N_4369);
nand U4559 (N_4559,N_4053,N_4328);
and U4560 (N_4560,N_4081,N_4012);
or U4561 (N_4561,N_4240,N_4306);
and U4562 (N_4562,N_4060,N_4253);
or U4563 (N_4563,N_4244,N_4040);
nand U4564 (N_4564,N_4078,N_4454);
nand U4565 (N_4565,N_4465,N_4346);
or U4566 (N_4566,N_4186,N_4098);
nor U4567 (N_4567,N_4102,N_4017);
or U4568 (N_4568,N_4494,N_4199);
and U4569 (N_4569,N_4473,N_4250);
nor U4570 (N_4570,N_4428,N_4147);
or U4571 (N_4571,N_4087,N_4455);
xor U4572 (N_4572,N_4136,N_4172);
or U4573 (N_4573,N_4169,N_4481);
xor U4574 (N_4574,N_4407,N_4257);
nor U4575 (N_4575,N_4112,N_4051);
xor U4576 (N_4576,N_4376,N_4363);
nor U4577 (N_4577,N_4266,N_4334);
nor U4578 (N_4578,N_4030,N_4387);
xor U4579 (N_4579,N_4345,N_4065);
and U4580 (N_4580,N_4396,N_4344);
nand U4581 (N_4581,N_4142,N_4339);
and U4582 (N_4582,N_4181,N_4020);
nand U4583 (N_4583,N_4427,N_4394);
or U4584 (N_4584,N_4044,N_4365);
or U4585 (N_4585,N_4238,N_4397);
and U4586 (N_4586,N_4289,N_4089);
nand U4587 (N_4587,N_4483,N_4202);
nand U4588 (N_4588,N_4014,N_4319);
nand U4589 (N_4589,N_4237,N_4174);
or U4590 (N_4590,N_4282,N_4034);
nand U4591 (N_4591,N_4067,N_4446);
nand U4592 (N_4592,N_4404,N_4050);
and U4593 (N_4593,N_4281,N_4411);
nand U4594 (N_4594,N_4461,N_4343);
nand U4595 (N_4595,N_4231,N_4132);
or U4596 (N_4596,N_4085,N_4399);
and U4597 (N_4597,N_4393,N_4324);
nand U4598 (N_4598,N_4254,N_4204);
or U4599 (N_4599,N_4443,N_4362);
nor U4600 (N_4600,N_4166,N_4175);
nor U4601 (N_4601,N_4456,N_4269);
nand U4602 (N_4602,N_4459,N_4492);
nand U4603 (N_4603,N_4214,N_4441);
nand U4604 (N_4604,N_4398,N_4288);
and U4605 (N_4605,N_4179,N_4335);
nor U4606 (N_4606,N_4191,N_4153);
nand U4607 (N_4607,N_4245,N_4366);
nor U4608 (N_4608,N_4046,N_4452);
and U4609 (N_4609,N_4177,N_4110);
nand U4610 (N_4610,N_4084,N_4351);
nand U4611 (N_4611,N_4497,N_4280);
and U4612 (N_4612,N_4232,N_4248);
or U4613 (N_4613,N_4392,N_4064);
nand U4614 (N_4614,N_4217,N_4117);
nand U4615 (N_4615,N_4121,N_4485);
and U4616 (N_4616,N_4056,N_4092);
xor U4617 (N_4617,N_4161,N_4276);
or U4618 (N_4618,N_4273,N_4252);
nor U4619 (N_4619,N_4239,N_4488);
nor U4620 (N_4620,N_4074,N_4145);
or U4621 (N_4621,N_4403,N_4195);
or U4622 (N_4622,N_4192,N_4241);
and U4623 (N_4623,N_4449,N_4315);
nor U4624 (N_4624,N_4061,N_4439);
xnor U4625 (N_4625,N_4450,N_4099);
and U4626 (N_4626,N_4287,N_4312);
or U4627 (N_4627,N_4111,N_4482);
nand U4628 (N_4628,N_4278,N_4140);
or U4629 (N_4629,N_4367,N_4032);
or U4630 (N_4630,N_4384,N_4126);
and U4631 (N_4631,N_4355,N_4385);
or U4632 (N_4632,N_4331,N_4021);
and U4633 (N_4633,N_4484,N_4337);
nor U4634 (N_4634,N_4160,N_4197);
nor U4635 (N_4635,N_4486,N_4120);
or U4636 (N_4636,N_4297,N_4419);
or U4637 (N_4637,N_4383,N_4027);
and U4638 (N_4638,N_4036,N_4045);
and U4639 (N_4639,N_4474,N_4018);
and U4640 (N_4640,N_4358,N_4436);
xnor U4641 (N_4641,N_4321,N_4251);
nor U4642 (N_4642,N_4463,N_4006);
nor U4643 (N_4643,N_4170,N_4402);
or U4644 (N_4644,N_4317,N_4003);
nand U4645 (N_4645,N_4423,N_4303);
nor U4646 (N_4646,N_4322,N_4354);
and U4647 (N_4647,N_4472,N_4475);
nand U4648 (N_4648,N_4347,N_4489);
or U4649 (N_4649,N_4047,N_4148);
and U4650 (N_4650,N_4270,N_4068);
nand U4651 (N_4651,N_4310,N_4219);
xor U4652 (N_4652,N_4352,N_4496);
nand U4653 (N_4653,N_4139,N_4415);
nand U4654 (N_4654,N_4215,N_4080);
or U4655 (N_4655,N_4476,N_4076);
or U4656 (N_4656,N_4176,N_4286);
nand U4657 (N_4657,N_4440,N_4188);
nor U4658 (N_4658,N_4190,N_4069);
or U4659 (N_4659,N_4059,N_4100);
or U4660 (N_4660,N_4432,N_4370);
and U4661 (N_4661,N_4348,N_4445);
and U4662 (N_4662,N_4447,N_4083);
and U4663 (N_4663,N_4405,N_4425);
and U4664 (N_4664,N_4070,N_4435);
nand U4665 (N_4665,N_4203,N_4420);
nor U4666 (N_4666,N_4479,N_4341);
nor U4667 (N_4667,N_4498,N_4375);
nand U4668 (N_4668,N_4426,N_4417);
nand U4669 (N_4669,N_4155,N_4388);
and U4670 (N_4670,N_4416,N_4088);
nand U4671 (N_4671,N_4071,N_4413);
xnor U4672 (N_4672,N_4225,N_4127);
nand U4673 (N_4673,N_4433,N_4389);
and U4674 (N_4674,N_4391,N_4150);
nand U4675 (N_4675,N_4360,N_4058);
nand U4676 (N_4676,N_4031,N_4378);
nor U4677 (N_4677,N_4421,N_4381);
nor U4678 (N_4678,N_4305,N_4395);
and U4679 (N_4679,N_4128,N_4094);
nand U4680 (N_4680,N_4342,N_4327);
nor U4681 (N_4681,N_4019,N_4115);
nor U4682 (N_4682,N_4359,N_4180);
nand U4683 (N_4683,N_4429,N_4052);
nor U4684 (N_4684,N_4167,N_4213);
or U4685 (N_4685,N_4187,N_4185);
or U4686 (N_4686,N_4466,N_4470);
nor U4687 (N_4687,N_4124,N_4437);
and U4688 (N_4688,N_4041,N_4308);
nor U4689 (N_4689,N_4260,N_4296);
nor U4690 (N_4690,N_4005,N_4224);
nor U4691 (N_4691,N_4380,N_4022);
and U4692 (N_4692,N_4235,N_4114);
or U4693 (N_4693,N_4285,N_4300);
nand U4694 (N_4694,N_4196,N_4007);
and U4695 (N_4695,N_4226,N_4438);
nor U4696 (N_4696,N_4096,N_4104);
nor U4697 (N_4697,N_4462,N_4277);
or U4698 (N_4698,N_4125,N_4229);
and U4699 (N_4699,N_4424,N_4023);
nand U4700 (N_4700,N_4151,N_4386);
nor U4701 (N_4701,N_4295,N_4026);
nor U4702 (N_4702,N_4216,N_4028);
nor U4703 (N_4703,N_4008,N_4141);
nand U4704 (N_4704,N_4418,N_4123);
or U4705 (N_4705,N_4015,N_4066);
or U4706 (N_4706,N_4212,N_4037);
and U4707 (N_4707,N_4361,N_4000);
nor U4708 (N_4708,N_4326,N_4431);
nand U4709 (N_4709,N_4246,N_4159);
or U4710 (N_4710,N_4451,N_4292);
nor U4711 (N_4711,N_4243,N_4143);
and U4712 (N_4712,N_4412,N_4264);
xor U4713 (N_4713,N_4091,N_4301);
and U4714 (N_4714,N_4299,N_4009);
nor U4715 (N_4715,N_4173,N_4134);
or U4716 (N_4716,N_4162,N_4108);
nor U4717 (N_4717,N_4223,N_4154);
and U4718 (N_4718,N_4329,N_4082);
and U4719 (N_4719,N_4208,N_4467);
or U4720 (N_4720,N_4207,N_4010);
nor U4721 (N_4721,N_4137,N_4054);
and U4722 (N_4722,N_4373,N_4057);
or U4723 (N_4723,N_4209,N_4055);
xor U4724 (N_4724,N_4095,N_4013);
nor U4725 (N_4725,N_4444,N_4105);
nand U4726 (N_4726,N_4390,N_4039);
and U4727 (N_4727,N_4372,N_4233);
nand U4728 (N_4728,N_4268,N_4400);
or U4729 (N_4729,N_4353,N_4453);
nand U4730 (N_4730,N_4382,N_4198);
nand U4731 (N_4731,N_4499,N_4024);
nand U4732 (N_4732,N_4377,N_4220);
or U4733 (N_4733,N_4144,N_4234);
and U4734 (N_4734,N_4271,N_4258);
or U4735 (N_4735,N_4291,N_4256);
and U4736 (N_4736,N_4043,N_4457);
xor U4737 (N_4737,N_4205,N_4340);
nand U4738 (N_4738,N_4357,N_4298);
nand U4739 (N_4739,N_4222,N_4293);
or U4740 (N_4740,N_4113,N_4106);
and U4741 (N_4741,N_4129,N_4350);
or U4742 (N_4742,N_4265,N_4103);
nand U4743 (N_4743,N_4311,N_4109);
nand U4744 (N_4744,N_4480,N_4138);
nor U4745 (N_4745,N_4409,N_4320);
nand U4746 (N_4746,N_4430,N_4272);
and U4747 (N_4747,N_4333,N_4163);
nor U4748 (N_4748,N_4490,N_4218);
nand U4749 (N_4749,N_4116,N_4290);
and U4750 (N_4750,N_4342,N_4063);
nor U4751 (N_4751,N_4230,N_4065);
and U4752 (N_4752,N_4196,N_4162);
and U4753 (N_4753,N_4327,N_4031);
and U4754 (N_4754,N_4312,N_4051);
or U4755 (N_4755,N_4170,N_4471);
or U4756 (N_4756,N_4488,N_4104);
or U4757 (N_4757,N_4466,N_4015);
and U4758 (N_4758,N_4013,N_4106);
or U4759 (N_4759,N_4245,N_4389);
and U4760 (N_4760,N_4307,N_4261);
nand U4761 (N_4761,N_4316,N_4091);
nand U4762 (N_4762,N_4375,N_4140);
or U4763 (N_4763,N_4220,N_4348);
or U4764 (N_4764,N_4497,N_4135);
xor U4765 (N_4765,N_4092,N_4264);
xnor U4766 (N_4766,N_4374,N_4433);
xor U4767 (N_4767,N_4428,N_4305);
nand U4768 (N_4768,N_4453,N_4491);
or U4769 (N_4769,N_4252,N_4081);
and U4770 (N_4770,N_4011,N_4371);
nor U4771 (N_4771,N_4083,N_4467);
nand U4772 (N_4772,N_4203,N_4302);
nor U4773 (N_4773,N_4092,N_4484);
and U4774 (N_4774,N_4385,N_4266);
nand U4775 (N_4775,N_4114,N_4393);
and U4776 (N_4776,N_4353,N_4237);
nand U4777 (N_4777,N_4465,N_4065);
nor U4778 (N_4778,N_4031,N_4022);
and U4779 (N_4779,N_4415,N_4427);
xnor U4780 (N_4780,N_4263,N_4055);
nand U4781 (N_4781,N_4310,N_4168);
nor U4782 (N_4782,N_4316,N_4373);
nand U4783 (N_4783,N_4449,N_4314);
nand U4784 (N_4784,N_4318,N_4221);
or U4785 (N_4785,N_4010,N_4222);
or U4786 (N_4786,N_4439,N_4025);
and U4787 (N_4787,N_4476,N_4482);
nor U4788 (N_4788,N_4444,N_4346);
and U4789 (N_4789,N_4168,N_4326);
nand U4790 (N_4790,N_4468,N_4128);
nor U4791 (N_4791,N_4275,N_4357);
xor U4792 (N_4792,N_4138,N_4291);
and U4793 (N_4793,N_4052,N_4479);
and U4794 (N_4794,N_4015,N_4163);
nor U4795 (N_4795,N_4370,N_4241);
or U4796 (N_4796,N_4254,N_4371);
xnor U4797 (N_4797,N_4156,N_4428);
or U4798 (N_4798,N_4494,N_4122);
and U4799 (N_4799,N_4334,N_4022);
nand U4800 (N_4800,N_4229,N_4223);
or U4801 (N_4801,N_4363,N_4253);
nand U4802 (N_4802,N_4014,N_4067);
or U4803 (N_4803,N_4221,N_4289);
nand U4804 (N_4804,N_4493,N_4184);
and U4805 (N_4805,N_4363,N_4472);
nand U4806 (N_4806,N_4012,N_4140);
and U4807 (N_4807,N_4323,N_4473);
nor U4808 (N_4808,N_4453,N_4013);
xor U4809 (N_4809,N_4013,N_4400);
or U4810 (N_4810,N_4231,N_4347);
or U4811 (N_4811,N_4032,N_4144);
or U4812 (N_4812,N_4126,N_4127);
or U4813 (N_4813,N_4038,N_4151);
nand U4814 (N_4814,N_4097,N_4133);
nor U4815 (N_4815,N_4023,N_4239);
and U4816 (N_4816,N_4242,N_4192);
or U4817 (N_4817,N_4426,N_4291);
nor U4818 (N_4818,N_4202,N_4414);
xnor U4819 (N_4819,N_4007,N_4106);
nand U4820 (N_4820,N_4074,N_4429);
nand U4821 (N_4821,N_4206,N_4119);
nand U4822 (N_4822,N_4111,N_4266);
nor U4823 (N_4823,N_4184,N_4295);
xor U4824 (N_4824,N_4185,N_4260);
nor U4825 (N_4825,N_4040,N_4192);
and U4826 (N_4826,N_4108,N_4102);
or U4827 (N_4827,N_4214,N_4192);
or U4828 (N_4828,N_4283,N_4112);
and U4829 (N_4829,N_4026,N_4344);
and U4830 (N_4830,N_4366,N_4202);
nor U4831 (N_4831,N_4085,N_4251);
nand U4832 (N_4832,N_4434,N_4002);
and U4833 (N_4833,N_4395,N_4398);
or U4834 (N_4834,N_4229,N_4121);
and U4835 (N_4835,N_4195,N_4398);
xor U4836 (N_4836,N_4158,N_4134);
or U4837 (N_4837,N_4415,N_4222);
and U4838 (N_4838,N_4074,N_4379);
or U4839 (N_4839,N_4069,N_4312);
nand U4840 (N_4840,N_4462,N_4372);
and U4841 (N_4841,N_4094,N_4032);
xor U4842 (N_4842,N_4348,N_4192);
and U4843 (N_4843,N_4265,N_4446);
nor U4844 (N_4844,N_4409,N_4338);
nor U4845 (N_4845,N_4243,N_4367);
or U4846 (N_4846,N_4435,N_4299);
nand U4847 (N_4847,N_4264,N_4241);
or U4848 (N_4848,N_4277,N_4005);
nor U4849 (N_4849,N_4421,N_4369);
and U4850 (N_4850,N_4251,N_4035);
or U4851 (N_4851,N_4091,N_4287);
xnor U4852 (N_4852,N_4388,N_4395);
nand U4853 (N_4853,N_4211,N_4370);
or U4854 (N_4854,N_4052,N_4037);
nand U4855 (N_4855,N_4152,N_4363);
xnor U4856 (N_4856,N_4141,N_4320);
and U4857 (N_4857,N_4343,N_4094);
and U4858 (N_4858,N_4201,N_4485);
or U4859 (N_4859,N_4162,N_4003);
or U4860 (N_4860,N_4483,N_4194);
xor U4861 (N_4861,N_4071,N_4141);
xnor U4862 (N_4862,N_4447,N_4337);
and U4863 (N_4863,N_4490,N_4007);
or U4864 (N_4864,N_4037,N_4233);
nand U4865 (N_4865,N_4406,N_4279);
and U4866 (N_4866,N_4157,N_4431);
and U4867 (N_4867,N_4211,N_4034);
and U4868 (N_4868,N_4168,N_4490);
nand U4869 (N_4869,N_4192,N_4224);
nor U4870 (N_4870,N_4281,N_4014);
nor U4871 (N_4871,N_4254,N_4472);
nor U4872 (N_4872,N_4150,N_4397);
nand U4873 (N_4873,N_4037,N_4041);
and U4874 (N_4874,N_4378,N_4476);
nand U4875 (N_4875,N_4053,N_4243);
or U4876 (N_4876,N_4164,N_4480);
xnor U4877 (N_4877,N_4224,N_4167);
nand U4878 (N_4878,N_4451,N_4297);
or U4879 (N_4879,N_4324,N_4190);
and U4880 (N_4880,N_4209,N_4433);
or U4881 (N_4881,N_4171,N_4150);
nand U4882 (N_4882,N_4234,N_4217);
nor U4883 (N_4883,N_4046,N_4463);
or U4884 (N_4884,N_4339,N_4385);
nand U4885 (N_4885,N_4370,N_4264);
and U4886 (N_4886,N_4326,N_4090);
nor U4887 (N_4887,N_4273,N_4158);
and U4888 (N_4888,N_4156,N_4157);
nor U4889 (N_4889,N_4152,N_4487);
nor U4890 (N_4890,N_4392,N_4203);
nor U4891 (N_4891,N_4144,N_4232);
xnor U4892 (N_4892,N_4187,N_4423);
nand U4893 (N_4893,N_4190,N_4320);
nor U4894 (N_4894,N_4339,N_4340);
or U4895 (N_4895,N_4248,N_4494);
nor U4896 (N_4896,N_4445,N_4335);
xnor U4897 (N_4897,N_4454,N_4309);
or U4898 (N_4898,N_4104,N_4152);
or U4899 (N_4899,N_4081,N_4150);
or U4900 (N_4900,N_4032,N_4192);
and U4901 (N_4901,N_4205,N_4351);
nor U4902 (N_4902,N_4495,N_4113);
nor U4903 (N_4903,N_4129,N_4090);
and U4904 (N_4904,N_4256,N_4233);
or U4905 (N_4905,N_4224,N_4318);
xor U4906 (N_4906,N_4235,N_4478);
xnor U4907 (N_4907,N_4314,N_4207);
and U4908 (N_4908,N_4112,N_4209);
and U4909 (N_4909,N_4059,N_4287);
nand U4910 (N_4910,N_4347,N_4499);
or U4911 (N_4911,N_4177,N_4017);
nor U4912 (N_4912,N_4094,N_4331);
nor U4913 (N_4913,N_4290,N_4289);
or U4914 (N_4914,N_4131,N_4052);
nand U4915 (N_4915,N_4392,N_4273);
and U4916 (N_4916,N_4328,N_4150);
nand U4917 (N_4917,N_4301,N_4161);
nor U4918 (N_4918,N_4359,N_4334);
and U4919 (N_4919,N_4419,N_4107);
or U4920 (N_4920,N_4259,N_4451);
nor U4921 (N_4921,N_4115,N_4159);
nand U4922 (N_4922,N_4412,N_4186);
and U4923 (N_4923,N_4273,N_4218);
or U4924 (N_4924,N_4147,N_4405);
nand U4925 (N_4925,N_4490,N_4354);
or U4926 (N_4926,N_4091,N_4436);
and U4927 (N_4927,N_4396,N_4439);
or U4928 (N_4928,N_4188,N_4359);
or U4929 (N_4929,N_4382,N_4413);
and U4930 (N_4930,N_4165,N_4445);
xnor U4931 (N_4931,N_4230,N_4209);
nand U4932 (N_4932,N_4359,N_4495);
or U4933 (N_4933,N_4176,N_4263);
or U4934 (N_4934,N_4384,N_4467);
nand U4935 (N_4935,N_4175,N_4130);
nand U4936 (N_4936,N_4133,N_4011);
or U4937 (N_4937,N_4054,N_4298);
and U4938 (N_4938,N_4462,N_4007);
nand U4939 (N_4939,N_4406,N_4403);
and U4940 (N_4940,N_4125,N_4260);
or U4941 (N_4941,N_4080,N_4348);
and U4942 (N_4942,N_4187,N_4077);
or U4943 (N_4943,N_4191,N_4412);
nor U4944 (N_4944,N_4424,N_4031);
or U4945 (N_4945,N_4089,N_4457);
or U4946 (N_4946,N_4398,N_4120);
and U4947 (N_4947,N_4219,N_4393);
nor U4948 (N_4948,N_4466,N_4394);
nor U4949 (N_4949,N_4255,N_4376);
nor U4950 (N_4950,N_4203,N_4349);
nor U4951 (N_4951,N_4069,N_4451);
or U4952 (N_4952,N_4435,N_4102);
nand U4953 (N_4953,N_4405,N_4469);
and U4954 (N_4954,N_4233,N_4002);
nand U4955 (N_4955,N_4237,N_4239);
xor U4956 (N_4956,N_4137,N_4382);
nor U4957 (N_4957,N_4423,N_4487);
nand U4958 (N_4958,N_4338,N_4098);
and U4959 (N_4959,N_4122,N_4037);
xor U4960 (N_4960,N_4217,N_4418);
nand U4961 (N_4961,N_4459,N_4030);
nor U4962 (N_4962,N_4459,N_4363);
and U4963 (N_4963,N_4340,N_4306);
xor U4964 (N_4964,N_4258,N_4025);
and U4965 (N_4965,N_4192,N_4031);
nand U4966 (N_4966,N_4484,N_4327);
and U4967 (N_4967,N_4237,N_4010);
or U4968 (N_4968,N_4082,N_4247);
xnor U4969 (N_4969,N_4239,N_4220);
xnor U4970 (N_4970,N_4255,N_4382);
or U4971 (N_4971,N_4139,N_4130);
and U4972 (N_4972,N_4341,N_4369);
nor U4973 (N_4973,N_4064,N_4468);
and U4974 (N_4974,N_4249,N_4276);
nand U4975 (N_4975,N_4261,N_4291);
nand U4976 (N_4976,N_4064,N_4285);
nor U4977 (N_4977,N_4233,N_4395);
nand U4978 (N_4978,N_4055,N_4081);
and U4979 (N_4979,N_4029,N_4028);
nand U4980 (N_4980,N_4040,N_4480);
and U4981 (N_4981,N_4489,N_4353);
nor U4982 (N_4982,N_4468,N_4428);
and U4983 (N_4983,N_4114,N_4291);
nor U4984 (N_4984,N_4469,N_4219);
or U4985 (N_4985,N_4275,N_4369);
or U4986 (N_4986,N_4087,N_4282);
nor U4987 (N_4987,N_4136,N_4016);
or U4988 (N_4988,N_4242,N_4255);
nor U4989 (N_4989,N_4098,N_4238);
nor U4990 (N_4990,N_4266,N_4309);
and U4991 (N_4991,N_4149,N_4072);
nand U4992 (N_4992,N_4163,N_4346);
or U4993 (N_4993,N_4074,N_4481);
or U4994 (N_4994,N_4264,N_4304);
nand U4995 (N_4995,N_4146,N_4125);
xnor U4996 (N_4996,N_4021,N_4036);
nor U4997 (N_4997,N_4200,N_4467);
and U4998 (N_4998,N_4477,N_4180);
nand U4999 (N_4999,N_4494,N_4048);
or U5000 (N_5000,N_4766,N_4771);
or U5001 (N_5001,N_4551,N_4696);
nor U5002 (N_5002,N_4978,N_4684);
nand U5003 (N_5003,N_4977,N_4794);
and U5004 (N_5004,N_4951,N_4922);
nand U5005 (N_5005,N_4719,N_4909);
and U5006 (N_5006,N_4941,N_4688);
xor U5007 (N_5007,N_4830,N_4575);
nand U5008 (N_5008,N_4752,N_4526);
xor U5009 (N_5009,N_4962,N_4541);
xnor U5010 (N_5010,N_4736,N_4809);
nor U5011 (N_5011,N_4864,N_4923);
nand U5012 (N_5012,N_4993,N_4981);
xor U5013 (N_5013,N_4553,N_4964);
and U5014 (N_5014,N_4595,N_4834);
nand U5015 (N_5015,N_4742,N_4516);
or U5016 (N_5016,N_4972,N_4792);
or U5017 (N_5017,N_4732,N_4798);
or U5018 (N_5018,N_4645,N_4643);
nor U5019 (N_5019,N_4974,N_4799);
nand U5020 (N_5020,N_4698,N_4695);
nand U5021 (N_5021,N_4904,N_4940);
and U5022 (N_5022,N_4802,N_4765);
and U5023 (N_5023,N_4928,N_4926);
nor U5024 (N_5024,N_4673,N_4915);
nor U5025 (N_5025,N_4775,N_4814);
or U5026 (N_5026,N_4670,N_4801);
and U5027 (N_5027,N_4681,N_4669);
or U5028 (N_5028,N_4674,N_4729);
nor U5029 (N_5029,N_4519,N_4697);
and U5030 (N_5030,N_4524,N_4743);
nand U5031 (N_5031,N_4581,N_4818);
or U5032 (N_5032,N_4758,N_4877);
xor U5033 (N_5033,N_4957,N_4892);
nand U5034 (N_5034,N_4852,N_4590);
nor U5035 (N_5035,N_4689,N_4651);
nand U5036 (N_5036,N_4896,N_4550);
or U5037 (N_5037,N_4829,N_4745);
nand U5038 (N_5038,N_4756,N_4931);
or U5039 (N_5039,N_4703,N_4539);
or U5040 (N_5040,N_4726,N_4582);
nand U5041 (N_5041,N_4841,N_4855);
nor U5042 (N_5042,N_4984,N_4800);
or U5043 (N_5043,N_4911,N_4889);
nor U5044 (N_5044,N_4881,N_4639);
nand U5045 (N_5045,N_4867,N_4947);
nand U5046 (N_5046,N_4712,N_4883);
nor U5047 (N_5047,N_4784,N_4568);
and U5048 (N_5048,N_4733,N_4515);
or U5049 (N_5049,N_4634,N_4598);
nor U5050 (N_5050,N_4603,N_4523);
or U5051 (N_5051,N_4822,N_4907);
xor U5052 (N_5052,N_4737,N_4930);
nand U5053 (N_5053,N_4584,N_4608);
and U5054 (N_5054,N_4837,N_4810);
and U5055 (N_5055,N_4586,N_4805);
and U5056 (N_5056,N_4648,N_4715);
or U5057 (N_5057,N_4969,N_4546);
nor U5058 (N_5058,N_4630,N_4606);
nand U5059 (N_5059,N_4537,N_4549);
nand U5060 (N_5060,N_4916,N_4876);
and U5061 (N_5061,N_4796,N_4649);
or U5062 (N_5062,N_4990,N_4835);
or U5063 (N_5063,N_4569,N_4567);
nor U5064 (N_5064,N_4936,N_4777);
or U5065 (N_5065,N_4768,N_4533);
or U5066 (N_5066,N_4716,N_4543);
and U5067 (N_5067,N_4913,N_4518);
nor U5068 (N_5068,N_4991,N_4657);
nor U5069 (N_5069,N_4629,N_4843);
nor U5070 (N_5070,N_4788,N_4601);
nand U5071 (N_5071,N_4885,N_4908);
and U5072 (N_5072,N_4833,N_4793);
xor U5073 (N_5073,N_4987,N_4979);
nor U5074 (N_5074,N_4740,N_4520);
nor U5075 (N_5075,N_4986,N_4556);
or U5076 (N_5076,N_4783,N_4866);
nor U5077 (N_5077,N_4536,N_4682);
or U5078 (N_5078,N_4613,N_4845);
or U5079 (N_5079,N_4791,N_4786);
or U5080 (N_5080,N_4659,N_4751);
or U5081 (N_5081,N_4735,N_4741);
or U5082 (N_5082,N_4849,N_4778);
and U5083 (N_5083,N_4500,N_4680);
nand U5084 (N_5084,N_4637,N_4787);
nor U5085 (N_5085,N_4760,N_4868);
and U5086 (N_5086,N_4874,N_4683);
nor U5087 (N_5087,N_4548,N_4609);
nand U5088 (N_5088,N_4624,N_4699);
xnor U5089 (N_5089,N_4824,N_4522);
nand U5090 (N_5090,N_4966,N_4985);
nand U5091 (N_5091,N_4627,N_4970);
nand U5092 (N_5092,N_4812,N_4815);
or U5093 (N_5093,N_4617,N_4547);
nand U5094 (N_5094,N_4717,N_4646);
or U5095 (N_5095,N_4508,N_4517);
nand U5096 (N_5096,N_4917,N_4538);
nand U5097 (N_5097,N_4789,N_4755);
and U5098 (N_5098,N_4621,N_4655);
nor U5099 (N_5099,N_4934,N_4501);
nor U5100 (N_5100,N_4555,N_4754);
nor U5101 (N_5101,N_4708,N_4811);
and U5102 (N_5102,N_4975,N_4713);
nand U5103 (N_5103,N_4865,N_4946);
or U5104 (N_5104,N_4857,N_4502);
xor U5105 (N_5105,N_4847,N_4906);
nor U5106 (N_5106,N_4544,N_4579);
xor U5107 (N_5107,N_4999,N_4825);
nor U5108 (N_5108,N_4509,N_4589);
nand U5109 (N_5109,N_4563,N_4914);
and U5110 (N_5110,N_4514,N_4738);
nor U5111 (N_5111,N_4540,N_4562);
or U5112 (N_5112,N_4678,N_4846);
or U5113 (N_5113,N_4968,N_4641);
or U5114 (N_5114,N_4510,N_4869);
nand U5115 (N_5115,N_4512,N_4620);
or U5116 (N_5116,N_4631,N_4618);
and U5117 (N_5117,N_4943,N_4694);
and U5118 (N_5118,N_4894,N_4827);
and U5119 (N_5119,N_4529,N_4723);
nor U5120 (N_5120,N_4761,N_4570);
nand U5121 (N_5121,N_4616,N_4956);
xnor U5122 (N_5122,N_4728,N_4583);
or U5123 (N_5123,N_4658,N_4939);
and U5124 (N_5124,N_4554,N_4714);
and U5125 (N_5125,N_4654,N_4823);
and U5126 (N_5126,N_4503,N_4961);
nand U5127 (N_5127,N_4779,N_4856);
or U5128 (N_5128,N_4781,N_4672);
nor U5129 (N_5129,N_4893,N_4587);
nor U5130 (N_5130,N_4691,N_4594);
nor U5131 (N_5131,N_4666,N_4880);
and U5132 (N_5132,N_4886,N_4901);
or U5133 (N_5133,N_4782,N_4954);
and U5134 (N_5134,N_4638,N_4776);
nand U5135 (N_5135,N_4711,N_4636);
and U5136 (N_5136,N_4535,N_4832);
nor U5137 (N_5137,N_4900,N_4965);
and U5138 (N_5138,N_4642,N_4588);
nor U5139 (N_5139,N_4710,N_4602);
xnor U5140 (N_5140,N_4804,N_4844);
nor U5141 (N_5141,N_4808,N_4619);
and U5142 (N_5142,N_4953,N_4903);
nand U5143 (N_5143,N_4942,N_4722);
or U5144 (N_5144,N_4872,N_4566);
or U5145 (N_5145,N_4692,N_4534);
and U5146 (N_5146,N_4918,N_4924);
and U5147 (N_5147,N_4851,N_4706);
and U5148 (N_5148,N_4593,N_4763);
and U5149 (N_5149,N_4836,N_4933);
nor U5150 (N_5150,N_4967,N_4675);
nand U5151 (N_5151,N_4727,N_4817);
nor U5152 (N_5152,N_4705,N_4938);
nor U5153 (N_5153,N_4898,N_4560);
or U5154 (N_5154,N_4744,N_4826);
nor U5155 (N_5155,N_4653,N_4944);
or U5156 (N_5156,N_4925,N_4772);
and U5157 (N_5157,N_4973,N_4821);
nand U5158 (N_5158,N_4660,N_4599);
or U5159 (N_5159,N_4596,N_4718);
nand U5160 (N_5160,N_4559,N_4511);
nor U5161 (N_5161,N_4757,N_4773);
nor U5162 (N_5162,N_4607,N_4960);
nand U5163 (N_5163,N_4959,N_4640);
and U5164 (N_5164,N_4693,N_4937);
and U5165 (N_5165,N_4828,N_4950);
and U5166 (N_5166,N_4532,N_4963);
nand U5167 (N_5167,N_4668,N_4875);
nor U5168 (N_5168,N_4803,N_4665);
and U5169 (N_5169,N_4888,N_4912);
and U5170 (N_5170,N_4870,N_4677);
and U5171 (N_5171,N_4679,N_4667);
xor U5172 (N_5172,N_4955,N_4685);
or U5173 (N_5173,N_4605,N_4610);
nor U5174 (N_5174,N_4612,N_4615);
nor U5175 (N_5175,N_4611,N_4806);
nand U5176 (N_5176,N_4861,N_4785);
or U5177 (N_5177,N_4650,N_4592);
and U5178 (N_5178,N_4921,N_4790);
and U5179 (N_5179,N_4949,N_4573);
or U5180 (N_5180,N_4873,N_4988);
xnor U5181 (N_5181,N_4840,N_4687);
nand U5182 (N_5182,N_4513,N_4895);
nor U5183 (N_5183,N_4850,N_4995);
and U5184 (N_5184,N_4734,N_4730);
or U5185 (N_5185,N_4557,N_4644);
nand U5186 (N_5186,N_4720,N_4848);
nand U5187 (N_5187,N_4625,N_4797);
xnor U5188 (N_5188,N_4702,N_4527);
or U5189 (N_5189,N_4564,N_4597);
and U5190 (N_5190,N_4748,N_4614);
or U5191 (N_5191,N_4528,N_4819);
and U5192 (N_5192,N_4747,N_4769);
or U5193 (N_5193,N_4558,N_4971);
nand U5194 (N_5194,N_4635,N_4853);
or U5195 (N_5195,N_4525,N_4725);
nand U5196 (N_5196,N_4552,N_4762);
nor U5197 (N_5197,N_4591,N_4565);
or U5198 (N_5198,N_4746,N_4676);
or U5199 (N_5199,N_4577,N_4749);
or U5200 (N_5200,N_4879,N_4753);
nor U5201 (N_5201,N_4632,N_4671);
and U5202 (N_5202,N_4952,N_4996);
nand U5203 (N_5203,N_4838,N_4686);
nor U5204 (N_5204,N_4504,N_4750);
nand U5205 (N_5205,N_4759,N_4932);
or U5206 (N_5206,N_4983,N_4647);
xor U5207 (N_5207,N_4731,N_4600);
and U5208 (N_5208,N_4576,N_4507);
xor U5209 (N_5209,N_4531,N_4989);
or U5210 (N_5210,N_4795,N_4704);
nand U5211 (N_5211,N_4628,N_4767);
xnor U5212 (N_5212,N_4920,N_4664);
and U5213 (N_5213,N_4816,N_4905);
and U5214 (N_5214,N_4807,N_4842);
or U5215 (N_5215,N_4623,N_4839);
nor U5216 (N_5216,N_4780,N_4831);
or U5217 (N_5217,N_4871,N_4902);
and U5218 (N_5218,N_4663,N_4948);
or U5219 (N_5219,N_4813,N_4604);
and U5220 (N_5220,N_4884,N_4709);
nand U5221 (N_5221,N_4882,N_4958);
nand U5222 (N_5222,N_4998,N_4572);
nor U5223 (N_5223,N_4633,N_4820);
nand U5224 (N_5224,N_4994,N_4945);
xor U5225 (N_5225,N_4980,N_4530);
nand U5226 (N_5226,N_4887,N_4910);
or U5227 (N_5227,N_4585,N_4542);
nand U5228 (N_5228,N_4770,N_4545);
or U5229 (N_5229,N_4859,N_4721);
nor U5230 (N_5230,N_4899,N_4724);
nand U5231 (N_5231,N_4574,N_4707);
nor U5232 (N_5232,N_4858,N_4580);
nand U5233 (N_5233,N_4561,N_4982);
nand U5234 (N_5234,N_4863,N_4701);
and U5235 (N_5235,N_4927,N_4878);
or U5236 (N_5236,N_4578,N_4661);
nand U5237 (N_5237,N_4626,N_4860);
or U5238 (N_5238,N_4976,N_4764);
or U5239 (N_5239,N_4919,N_4652);
nor U5240 (N_5240,N_4521,N_4656);
and U5241 (N_5241,N_4890,N_4935);
nor U5242 (N_5242,N_4739,N_4505);
and U5243 (N_5243,N_4571,N_4929);
nand U5244 (N_5244,N_4891,N_4862);
or U5245 (N_5245,N_4662,N_4622);
or U5246 (N_5246,N_4897,N_4997);
nand U5247 (N_5247,N_4992,N_4506);
and U5248 (N_5248,N_4774,N_4690);
nor U5249 (N_5249,N_4700,N_4854);
nand U5250 (N_5250,N_4750,N_4757);
or U5251 (N_5251,N_4531,N_4976);
nand U5252 (N_5252,N_4609,N_4552);
xnor U5253 (N_5253,N_4906,N_4607);
nand U5254 (N_5254,N_4507,N_4619);
nand U5255 (N_5255,N_4916,N_4713);
or U5256 (N_5256,N_4929,N_4836);
and U5257 (N_5257,N_4657,N_4553);
and U5258 (N_5258,N_4775,N_4807);
nand U5259 (N_5259,N_4776,N_4524);
nor U5260 (N_5260,N_4994,N_4944);
and U5261 (N_5261,N_4786,N_4631);
and U5262 (N_5262,N_4970,N_4794);
or U5263 (N_5263,N_4904,N_4740);
or U5264 (N_5264,N_4625,N_4823);
nand U5265 (N_5265,N_4584,N_4966);
and U5266 (N_5266,N_4735,N_4882);
or U5267 (N_5267,N_4898,N_4706);
xor U5268 (N_5268,N_4585,N_4810);
nand U5269 (N_5269,N_4577,N_4551);
or U5270 (N_5270,N_4883,N_4980);
or U5271 (N_5271,N_4534,N_4868);
or U5272 (N_5272,N_4794,N_4716);
nor U5273 (N_5273,N_4634,N_4524);
and U5274 (N_5274,N_4777,N_4841);
and U5275 (N_5275,N_4629,N_4512);
or U5276 (N_5276,N_4683,N_4854);
and U5277 (N_5277,N_4862,N_4898);
nor U5278 (N_5278,N_4837,N_4582);
or U5279 (N_5279,N_4669,N_4710);
and U5280 (N_5280,N_4748,N_4581);
nor U5281 (N_5281,N_4567,N_4988);
or U5282 (N_5282,N_4783,N_4990);
and U5283 (N_5283,N_4686,N_4771);
nor U5284 (N_5284,N_4654,N_4975);
nand U5285 (N_5285,N_4859,N_4510);
and U5286 (N_5286,N_4663,N_4730);
or U5287 (N_5287,N_4942,N_4969);
nor U5288 (N_5288,N_4967,N_4817);
or U5289 (N_5289,N_4908,N_4751);
nand U5290 (N_5290,N_4943,N_4584);
nor U5291 (N_5291,N_4662,N_4698);
and U5292 (N_5292,N_4892,N_4634);
nor U5293 (N_5293,N_4744,N_4971);
or U5294 (N_5294,N_4506,N_4859);
or U5295 (N_5295,N_4674,N_4673);
nand U5296 (N_5296,N_4764,N_4523);
nor U5297 (N_5297,N_4703,N_4533);
nand U5298 (N_5298,N_4507,N_4501);
or U5299 (N_5299,N_4931,N_4792);
and U5300 (N_5300,N_4533,N_4583);
nand U5301 (N_5301,N_4701,N_4539);
nand U5302 (N_5302,N_4623,N_4944);
or U5303 (N_5303,N_4800,N_4845);
and U5304 (N_5304,N_4978,N_4977);
and U5305 (N_5305,N_4549,N_4574);
or U5306 (N_5306,N_4818,N_4573);
or U5307 (N_5307,N_4564,N_4942);
and U5308 (N_5308,N_4671,N_4914);
nand U5309 (N_5309,N_4997,N_4848);
nand U5310 (N_5310,N_4629,N_4743);
nor U5311 (N_5311,N_4960,N_4510);
xor U5312 (N_5312,N_4988,N_4999);
and U5313 (N_5313,N_4514,N_4971);
or U5314 (N_5314,N_4989,N_4877);
nand U5315 (N_5315,N_4559,N_4745);
nand U5316 (N_5316,N_4857,N_4987);
or U5317 (N_5317,N_4673,N_4953);
or U5318 (N_5318,N_4804,N_4580);
xnor U5319 (N_5319,N_4932,N_4733);
nand U5320 (N_5320,N_4649,N_4946);
or U5321 (N_5321,N_4530,N_4796);
nand U5322 (N_5322,N_4625,N_4719);
or U5323 (N_5323,N_4840,N_4591);
nor U5324 (N_5324,N_4988,N_4586);
and U5325 (N_5325,N_4823,N_4650);
nand U5326 (N_5326,N_4698,N_4753);
nor U5327 (N_5327,N_4636,N_4788);
nor U5328 (N_5328,N_4790,N_4998);
nor U5329 (N_5329,N_4784,N_4534);
or U5330 (N_5330,N_4513,N_4788);
nand U5331 (N_5331,N_4919,N_4673);
or U5332 (N_5332,N_4824,N_4889);
nor U5333 (N_5333,N_4992,N_4584);
nand U5334 (N_5334,N_4912,N_4629);
nand U5335 (N_5335,N_4804,N_4992);
xnor U5336 (N_5336,N_4514,N_4942);
or U5337 (N_5337,N_4739,N_4968);
and U5338 (N_5338,N_4776,N_4582);
and U5339 (N_5339,N_4979,N_4883);
xor U5340 (N_5340,N_4524,N_4746);
nor U5341 (N_5341,N_4998,N_4626);
nand U5342 (N_5342,N_4692,N_4742);
xnor U5343 (N_5343,N_4824,N_4871);
nor U5344 (N_5344,N_4775,N_4797);
nand U5345 (N_5345,N_4947,N_4543);
and U5346 (N_5346,N_4574,N_4836);
nand U5347 (N_5347,N_4901,N_4696);
nor U5348 (N_5348,N_4845,N_4808);
nand U5349 (N_5349,N_4788,N_4913);
or U5350 (N_5350,N_4781,N_4964);
nand U5351 (N_5351,N_4652,N_4921);
and U5352 (N_5352,N_4815,N_4668);
nand U5353 (N_5353,N_4825,N_4821);
and U5354 (N_5354,N_4905,N_4885);
nand U5355 (N_5355,N_4903,N_4513);
and U5356 (N_5356,N_4796,N_4767);
nor U5357 (N_5357,N_4838,N_4644);
and U5358 (N_5358,N_4762,N_4691);
and U5359 (N_5359,N_4592,N_4776);
and U5360 (N_5360,N_4523,N_4594);
nand U5361 (N_5361,N_4884,N_4772);
nor U5362 (N_5362,N_4513,N_4610);
or U5363 (N_5363,N_4988,N_4724);
nand U5364 (N_5364,N_4697,N_4993);
or U5365 (N_5365,N_4622,N_4648);
nand U5366 (N_5366,N_4945,N_4831);
nand U5367 (N_5367,N_4787,N_4862);
or U5368 (N_5368,N_4996,N_4943);
nand U5369 (N_5369,N_4561,N_4823);
nand U5370 (N_5370,N_4893,N_4923);
or U5371 (N_5371,N_4564,N_4838);
xnor U5372 (N_5372,N_4591,N_4991);
xnor U5373 (N_5373,N_4902,N_4737);
nor U5374 (N_5374,N_4604,N_4906);
nor U5375 (N_5375,N_4874,N_4604);
nor U5376 (N_5376,N_4753,N_4626);
nor U5377 (N_5377,N_4628,N_4596);
nand U5378 (N_5378,N_4959,N_4830);
nand U5379 (N_5379,N_4550,N_4923);
xor U5380 (N_5380,N_4988,N_4588);
nand U5381 (N_5381,N_4765,N_4994);
nor U5382 (N_5382,N_4611,N_4967);
nand U5383 (N_5383,N_4782,N_4820);
nand U5384 (N_5384,N_4684,N_4589);
xnor U5385 (N_5385,N_4560,N_4658);
and U5386 (N_5386,N_4502,N_4607);
nor U5387 (N_5387,N_4942,N_4622);
or U5388 (N_5388,N_4597,N_4796);
nand U5389 (N_5389,N_4780,N_4775);
nor U5390 (N_5390,N_4838,N_4701);
and U5391 (N_5391,N_4965,N_4679);
nand U5392 (N_5392,N_4936,N_4960);
and U5393 (N_5393,N_4692,N_4626);
nand U5394 (N_5394,N_4706,N_4809);
and U5395 (N_5395,N_4763,N_4953);
nor U5396 (N_5396,N_4848,N_4519);
nand U5397 (N_5397,N_4832,N_4674);
or U5398 (N_5398,N_4969,N_4808);
nor U5399 (N_5399,N_4966,N_4802);
nor U5400 (N_5400,N_4582,N_4946);
or U5401 (N_5401,N_4846,N_4761);
nor U5402 (N_5402,N_4613,N_4658);
and U5403 (N_5403,N_4689,N_4728);
or U5404 (N_5404,N_4890,N_4796);
nor U5405 (N_5405,N_4571,N_4705);
nor U5406 (N_5406,N_4571,N_4594);
xnor U5407 (N_5407,N_4942,N_4846);
or U5408 (N_5408,N_4655,N_4920);
xor U5409 (N_5409,N_4793,N_4588);
or U5410 (N_5410,N_4868,N_4939);
or U5411 (N_5411,N_4629,N_4752);
and U5412 (N_5412,N_4832,N_4515);
nor U5413 (N_5413,N_4777,N_4599);
and U5414 (N_5414,N_4959,N_4636);
or U5415 (N_5415,N_4741,N_4806);
and U5416 (N_5416,N_4735,N_4688);
nand U5417 (N_5417,N_4741,N_4662);
xor U5418 (N_5418,N_4825,N_4693);
and U5419 (N_5419,N_4984,N_4790);
and U5420 (N_5420,N_4800,N_4597);
and U5421 (N_5421,N_4599,N_4809);
and U5422 (N_5422,N_4764,N_4848);
nand U5423 (N_5423,N_4681,N_4985);
or U5424 (N_5424,N_4523,N_4914);
or U5425 (N_5425,N_4507,N_4691);
nand U5426 (N_5426,N_4974,N_4703);
xor U5427 (N_5427,N_4760,N_4959);
nor U5428 (N_5428,N_4902,N_4742);
and U5429 (N_5429,N_4848,N_4864);
and U5430 (N_5430,N_4675,N_4969);
nor U5431 (N_5431,N_4595,N_4730);
nand U5432 (N_5432,N_4876,N_4863);
nor U5433 (N_5433,N_4962,N_4949);
nor U5434 (N_5434,N_4729,N_4526);
and U5435 (N_5435,N_4826,N_4902);
or U5436 (N_5436,N_4817,N_4590);
or U5437 (N_5437,N_4506,N_4914);
nand U5438 (N_5438,N_4828,N_4855);
or U5439 (N_5439,N_4951,N_4607);
or U5440 (N_5440,N_4747,N_4735);
or U5441 (N_5441,N_4760,N_4916);
and U5442 (N_5442,N_4676,N_4807);
or U5443 (N_5443,N_4728,N_4924);
nor U5444 (N_5444,N_4620,N_4573);
nor U5445 (N_5445,N_4540,N_4945);
nor U5446 (N_5446,N_4571,N_4628);
nor U5447 (N_5447,N_4724,N_4560);
nand U5448 (N_5448,N_4882,N_4974);
or U5449 (N_5449,N_4729,N_4903);
xnor U5450 (N_5450,N_4835,N_4834);
and U5451 (N_5451,N_4768,N_4724);
or U5452 (N_5452,N_4629,N_4815);
or U5453 (N_5453,N_4799,N_4856);
and U5454 (N_5454,N_4753,N_4887);
nand U5455 (N_5455,N_4662,N_4908);
nand U5456 (N_5456,N_4622,N_4715);
and U5457 (N_5457,N_4732,N_4552);
xor U5458 (N_5458,N_4700,N_4955);
nor U5459 (N_5459,N_4773,N_4797);
and U5460 (N_5460,N_4607,N_4725);
nand U5461 (N_5461,N_4918,N_4966);
nand U5462 (N_5462,N_4615,N_4695);
nor U5463 (N_5463,N_4688,N_4573);
and U5464 (N_5464,N_4979,N_4743);
nor U5465 (N_5465,N_4966,N_4818);
or U5466 (N_5466,N_4891,N_4999);
or U5467 (N_5467,N_4562,N_4736);
and U5468 (N_5468,N_4555,N_4936);
nor U5469 (N_5469,N_4652,N_4845);
and U5470 (N_5470,N_4927,N_4993);
and U5471 (N_5471,N_4584,N_4728);
xnor U5472 (N_5472,N_4503,N_4867);
nor U5473 (N_5473,N_4581,N_4691);
nand U5474 (N_5474,N_4975,N_4755);
and U5475 (N_5475,N_4506,N_4714);
nor U5476 (N_5476,N_4710,N_4859);
and U5477 (N_5477,N_4663,N_4693);
nand U5478 (N_5478,N_4684,N_4577);
nor U5479 (N_5479,N_4897,N_4854);
and U5480 (N_5480,N_4942,N_4693);
nor U5481 (N_5481,N_4561,N_4639);
nor U5482 (N_5482,N_4506,N_4656);
nand U5483 (N_5483,N_4684,N_4691);
or U5484 (N_5484,N_4837,N_4960);
or U5485 (N_5485,N_4961,N_4573);
nor U5486 (N_5486,N_4823,N_4716);
nor U5487 (N_5487,N_4654,N_4658);
or U5488 (N_5488,N_4649,N_4690);
nand U5489 (N_5489,N_4729,N_4800);
or U5490 (N_5490,N_4831,N_4603);
and U5491 (N_5491,N_4567,N_4738);
xor U5492 (N_5492,N_4684,N_4605);
nor U5493 (N_5493,N_4892,N_4573);
nand U5494 (N_5494,N_4718,N_4786);
xor U5495 (N_5495,N_4913,N_4958);
xnor U5496 (N_5496,N_4587,N_4830);
nand U5497 (N_5497,N_4618,N_4952);
nand U5498 (N_5498,N_4950,N_4800);
nand U5499 (N_5499,N_4764,N_4996);
xor U5500 (N_5500,N_5437,N_5059);
nand U5501 (N_5501,N_5291,N_5126);
nand U5502 (N_5502,N_5380,N_5283);
nand U5503 (N_5503,N_5333,N_5486);
or U5504 (N_5504,N_5496,N_5371);
xnor U5505 (N_5505,N_5260,N_5325);
nor U5506 (N_5506,N_5293,N_5206);
nor U5507 (N_5507,N_5472,N_5422);
and U5508 (N_5508,N_5363,N_5247);
nor U5509 (N_5509,N_5439,N_5300);
nand U5510 (N_5510,N_5008,N_5473);
or U5511 (N_5511,N_5424,N_5379);
nor U5512 (N_5512,N_5197,N_5401);
nand U5513 (N_5513,N_5382,N_5184);
and U5514 (N_5514,N_5235,N_5296);
nand U5515 (N_5515,N_5031,N_5007);
or U5516 (N_5516,N_5030,N_5451);
nor U5517 (N_5517,N_5043,N_5114);
nand U5518 (N_5518,N_5049,N_5110);
nor U5519 (N_5519,N_5324,N_5236);
xnor U5520 (N_5520,N_5376,N_5109);
and U5521 (N_5521,N_5116,N_5183);
and U5522 (N_5522,N_5447,N_5285);
or U5523 (N_5523,N_5090,N_5394);
and U5524 (N_5524,N_5240,N_5017);
nand U5525 (N_5525,N_5212,N_5431);
xnor U5526 (N_5526,N_5028,N_5051);
and U5527 (N_5527,N_5281,N_5050);
nor U5528 (N_5528,N_5024,N_5493);
nand U5529 (N_5529,N_5163,N_5067);
and U5530 (N_5530,N_5080,N_5270);
or U5531 (N_5531,N_5432,N_5266);
or U5532 (N_5532,N_5057,N_5341);
and U5533 (N_5533,N_5357,N_5471);
nor U5534 (N_5534,N_5046,N_5182);
and U5535 (N_5535,N_5275,N_5087);
and U5536 (N_5536,N_5315,N_5048);
or U5537 (N_5537,N_5054,N_5117);
nor U5538 (N_5538,N_5263,N_5053);
and U5539 (N_5539,N_5309,N_5223);
and U5540 (N_5540,N_5244,N_5360);
nor U5541 (N_5541,N_5129,N_5414);
or U5542 (N_5542,N_5016,N_5278);
nor U5543 (N_5543,N_5100,N_5156);
nand U5544 (N_5544,N_5257,N_5326);
or U5545 (N_5545,N_5108,N_5130);
nor U5546 (N_5546,N_5288,N_5128);
nand U5547 (N_5547,N_5176,N_5137);
nand U5548 (N_5548,N_5061,N_5345);
and U5549 (N_5549,N_5218,N_5179);
xor U5550 (N_5550,N_5340,N_5430);
nand U5551 (N_5551,N_5454,N_5011);
and U5552 (N_5552,N_5194,N_5417);
or U5553 (N_5553,N_5416,N_5354);
or U5554 (N_5554,N_5413,N_5083);
xor U5555 (N_5555,N_5045,N_5072);
nor U5556 (N_5556,N_5005,N_5224);
xor U5557 (N_5557,N_5252,N_5427);
nand U5558 (N_5558,N_5042,N_5077);
and U5559 (N_5559,N_5167,N_5032);
or U5560 (N_5560,N_5151,N_5464);
and U5561 (N_5561,N_5243,N_5407);
and U5562 (N_5562,N_5242,N_5264);
nor U5563 (N_5563,N_5286,N_5081);
nor U5564 (N_5564,N_5457,N_5289);
xor U5565 (N_5565,N_5238,N_5180);
and U5566 (N_5566,N_5148,N_5466);
and U5567 (N_5567,N_5138,N_5041);
nor U5568 (N_5568,N_5111,N_5409);
nand U5569 (N_5569,N_5455,N_5175);
or U5570 (N_5570,N_5265,N_5085);
and U5571 (N_5571,N_5115,N_5095);
xnor U5572 (N_5572,N_5356,N_5458);
and U5573 (N_5573,N_5461,N_5034);
and U5574 (N_5574,N_5322,N_5298);
and U5575 (N_5575,N_5143,N_5284);
nor U5576 (N_5576,N_5144,N_5406);
nor U5577 (N_5577,N_5075,N_5029);
or U5578 (N_5578,N_5255,N_5127);
or U5579 (N_5579,N_5348,N_5249);
xnor U5580 (N_5580,N_5062,N_5153);
and U5581 (N_5581,N_5217,N_5490);
and U5582 (N_5582,N_5230,N_5359);
or U5583 (N_5583,N_5372,N_5010);
nor U5584 (N_5584,N_5392,N_5489);
or U5585 (N_5585,N_5344,N_5463);
nand U5586 (N_5586,N_5303,N_5171);
nor U5587 (N_5587,N_5155,N_5462);
nand U5588 (N_5588,N_5316,N_5311);
nand U5589 (N_5589,N_5159,N_5410);
nand U5590 (N_5590,N_5203,N_5301);
and U5591 (N_5591,N_5297,N_5202);
xor U5592 (N_5592,N_5004,N_5273);
or U5593 (N_5593,N_5377,N_5052);
nor U5594 (N_5594,N_5477,N_5207);
nor U5595 (N_5595,N_5211,N_5334);
and U5596 (N_5596,N_5400,N_5122);
nand U5597 (N_5597,N_5146,N_5027);
nand U5598 (N_5598,N_5200,N_5039);
nand U5599 (N_5599,N_5078,N_5441);
or U5600 (N_5600,N_5036,N_5113);
or U5601 (N_5601,N_5358,N_5459);
or U5602 (N_5602,N_5272,N_5346);
and U5603 (N_5603,N_5438,N_5139);
or U5604 (N_5604,N_5436,N_5295);
or U5605 (N_5605,N_5119,N_5373);
nor U5606 (N_5606,N_5302,N_5329);
and U5607 (N_5607,N_5313,N_5019);
and U5608 (N_5608,N_5418,N_5412);
or U5609 (N_5609,N_5259,N_5369);
nor U5610 (N_5610,N_5003,N_5251);
or U5611 (N_5611,N_5395,N_5399);
or U5612 (N_5612,N_5187,N_5076);
nor U5613 (N_5613,N_5483,N_5403);
and U5614 (N_5614,N_5349,N_5221);
and U5615 (N_5615,N_5445,N_5443);
and U5616 (N_5616,N_5158,N_5415);
nand U5617 (N_5617,N_5215,N_5446);
and U5618 (N_5618,N_5071,N_5089);
nor U5619 (N_5619,N_5262,N_5419);
nor U5620 (N_5620,N_5166,N_5185);
nor U5621 (N_5621,N_5140,N_5368);
or U5622 (N_5622,N_5352,N_5168);
or U5623 (N_5623,N_5258,N_5219);
and U5624 (N_5624,N_5105,N_5231);
nand U5625 (N_5625,N_5481,N_5460);
nand U5626 (N_5626,N_5411,N_5320);
nor U5627 (N_5627,N_5101,N_5210);
or U5628 (N_5628,N_5063,N_5404);
nor U5629 (N_5629,N_5339,N_5145);
and U5630 (N_5630,N_5009,N_5064);
nand U5631 (N_5631,N_5305,N_5191);
nand U5632 (N_5632,N_5389,N_5118);
and U5633 (N_5633,N_5213,N_5169);
nor U5634 (N_5634,N_5226,N_5121);
and U5635 (N_5635,N_5012,N_5013);
or U5636 (N_5636,N_5038,N_5170);
nand U5637 (N_5637,N_5035,N_5290);
nand U5638 (N_5638,N_5103,N_5181);
and U5639 (N_5639,N_5025,N_5323);
or U5640 (N_5640,N_5201,N_5269);
nand U5641 (N_5641,N_5331,N_5245);
nand U5642 (N_5642,N_5435,N_5044);
and U5643 (N_5643,N_5040,N_5307);
nor U5644 (N_5644,N_5361,N_5174);
nand U5645 (N_5645,N_5469,N_5364);
nand U5646 (N_5646,N_5375,N_5492);
nor U5647 (N_5647,N_5189,N_5299);
and U5648 (N_5648,N_5006,N_5020);
or U5649 (N_5649,N_5274,N_5001);
nor U5650 (N_5650,N_5332,N_5246);
xnor U5651 (N_5651,N_5342,N_5271);
or U5652 (N_5652,N_5237,N_5021);
or U5653 (N_5653,N_5442,N_5147);
or U5654 (N_5654,N_5190,N_5397);
or U5655 (N_5655,N_5487,N_5425);
or U5656 (N_5656,N_5058,N_5152);
or U5657 (N_5657,N_5088,N_5094);
nor U5658 (N_5658,N_5287,N_5378);
nor U5659 (N_5659,N_5141,N_5456);
xnor U5660 (N_5660,N_5385,N_5222);
nor U5661 (N_5661,N_5216,N_5276);
nor U5662 (N_5662,N_5306,N_5099);
nor U5663 (N_5663,N_5070,N_5254);
xnor U5664 (N_5664,N_5069,N_5093);
nor U5665 (N_5665,N_5253,N_5267);
or U5666 (N_5666,N_5068,N_5350);
or U5667 (N_5667,N_5106,N_5037);
and U5668 (N_5668,N_5026,N_5304);
and U5669 (N_5669,N_5355,N_5336);
and U5670 (N_5670,N_5188,N_5172);
nor U5671 (N_5671,N_5157,N_5091);
xnor U5672 (N_5672,N_5092,N_5277);
nand U5673 (N_5673,N_5383,N_5123);
nand U5674 (N_5674,N_5002,N_5241);
or U5675 (N_5675,N_5381,N_5136);
nand U5676 (N_5676,N_5018,N_5014);
or U5677 (N_5677,N_5480,N_5429);
and U5678 (N_5678,N_5314,N_5374);
xor U5679 (N_5679,N_5388,N_5239);
and U5680 (N_5680,N_5097,N_5112);
and U5681 (N_5681,N_5452,N_5065);
xnor U5682 (N_5682,N_5468,N_5227);
or U5683 (N_5683,N_5494,N_5449);
nor U5684 (N_5684,N_5467,N_5261);
nand U5685 (N_5685,N_5150,N_5124);
nor U5686 (N_5686,N_5402,N_5022);
and U5687 (N_5687,N_5351,N_5328);
and U5688 (N_5688,N_5327,N_5135);
and U5689 (N_5689,N_5335,N_5084);
and U5690 (N_5690,N_5292,N_5131);
xnor U5691 (N_5691,N_5465,N_5149);
xnor U5692 (N_5692,N_5476,N_5102);
nand U5693 (N_5693,N_5015,N_5484);
or U5694 (N_5694,N_5066,N_5338);
and U5695 (N_5695,N_5470,N_5023);
or U5696 (N_5696,N_5164,N_5120);
and U5697 (N_5697,N_5162,N_5370);
and U5698 (N_5698,N_5198,N_5423);
and U5699 (N_5699,N_5033,N_5308);
or U5700 (N_5700,N_5228,N_5485);
nor U5701 (N_5701,N_5256,N_5362);
or U5702 (N_5702,N_5433,N_5421);
nand U5703 (N_5703,N_5347,N_5428);
or U5704 (N_5704,N_5000,N_5186);
nor U5705 (N_5705,N_5312,N_5160);
xnor U5706 (N_5706,N_5199,N_5475);
and U5707 (N_5707,N_5125,N_5498);
or U5708 (N_5708,N_5384,N_5074);
or U5709 (N_5709,N_5386,N_5229);
xor U5710 (N_5710,N_5250,N_5233);
nor U5711 (N_5711,N_5209,N_5330);
xnor U5712 (N_5712,N_5499,N_5390);
and U5713 (N_5713,N_5391,N_5234);
nor U5714 (N_5714,N_5474,N_5134);
or U5715 (N_5715,N_5319,N_5178);
or U5716 (N_5716,N_5491,N_5205);
nand U5717 (N_5717,N_5426,N_5387);
or U5718 (N_5718,N_5107,N_5232);
nand U5719 (N_5719,N_5060,N_5154);
xnor U5720 (N_5720,N_5321,N_5353);
xor U5721 (N_5721,N_5367,N_5279);
and U5722 (N_5722,N_5405,N_5133);
nor U5723 (N_5723,N_5343,N_5444);
and U5724 (N_5724,N_5195,N_5408);
nand U5725 (N_5725,N_5056,N_5310);
xnor U5726 (N_5726,N_5365,N_5220);
or U5727 (N_5727,N_5453,N_5104);
nand U5728 (N_5728,N_5497,N_5073);
or U5729 (N_5729,N_5440,N_5317);
and U5730 (N_5730,N_5337,N_5208);
and U5731 (N_5731,N_5047,N_5393);
and U5732 (N_5732,N_5225,N_5161);
nor U5733 (N_5733,N_5204,N_5142);
or U5734 (N_5734,N_5398,N_5248);
and U5735 (N_5735,N_5282,N_5098);
xnor U5736 (N_5736,N_5495,N_5132);
and U5737 (N_5737,N_5420,N_5280);
nand U5738 (N_5738,N_5450,N_5079);
and U5739 (N_5739,N_5479,N_5318);
nand U5740 (N_5740,N_5366,N_5173);
and U5741 (N_5741,N_5434,N_5082);
nor U5742 (N_5742,N_5096,N_5192);
or U5743 (N_5743,N_5193,N_5294);
nand U5744 (N_5744,N_5488,N_5478);
or U5745 (N_5745,N_5177,N_5055);
nor U5746 (N_5746,N_5396,N_5268);
nor U5747 (N_5747,N_5196,N_5482);
nand U5748 (N_5748,N_5086,N_5448);
nor U5749 (N_5749,N_5214,N_5165);
nor U5750 (N_5750,N_5290,N_5127);
or U5751 (N_5751,N_5010,N_5067);
nand U5752 (N_5752,N_5347,N_5224);
xnor U5753 (N_5753,N_5384,N_5371);
or U5754 (N_5754,N_5452,N_5262);
xor U5755 (N_5755,N_5124,N_5246);
nor U5756 (N_5756,N_5118,N_5045);
and U5757 (N_5757,N_5220,N_5466);
xor U5758 (N_5758,N_5496,N_5476);
nor U5759 (N_5759,N_5323,N_5113);
nor U5760 (N_5760,N_5453,N_5477);
nand U5761 (N_5761,N_5413,N_5027);
and U5762 (N_5762,N_5266,N_5368);
or U5763 (N_5763,N_5367,N_5127);
xnor U5764 (N_5764,N_5319,N_5067);
nand U5765 (N_5765,N_5418,N_5119);
and U5766 (N_5766,N_5391,N_5308);
nand U5767 (N_5767,N_5161,N_5092);
nor U5768 (N_5768,N_5045,N_5179);
and U5769 (N_5769,N_5137,N_5117);
or U5770 (N_5770,N_5467,N_5019);
and U5771 (N_5771,N_5441,N_5233);
or U5772 (N_5772,N_5042,N_5370);
and U5773 (N_5773,N_5312,N_5214);
or U5774 (N_5774,N_5416,N_5342);
nor U5775 (N_5775,N_5189,N_5081);
xnor U5776 (N_5776,N_5180,N_5208);
nor U5777 (N_5777,N_5071,N_5375);
or U5778 (N_5778,N_5336,N_5220);
nand U5779 (N_5779,N_5015,N_5176);
and U5780 (N_5780,N_5244,N_5341);
or U5781 (N_5781,N_5384,N_5385);
and U5782 (N_5782,N_5417,N_5321);
xnor U5783 (N_5783,N_5390,N_5088);
nand U5784 (N_5784,N_5048,N_5489);
and U5785 (N_5785,N_5078,N_5029);
or U5786 (N_5786,N_5219,N_5004);
and U5787 (N_5787,N_5244,N_5186);
or U5788 (N_5788,N_5404,N_5192);
nand U5789 (N_5789,N_5300,N_5160);
or U5790 (N_5790,N_5161,N_5369);
xnor U5791 (N_5791,N_5150,N_5194);
or U5792 (N_5792,N_5399,N_5444);
nand U5793 (N_5793,N_5337,N_5142);
and U5794 (N_5794,N_5474,N_5418);
nor U5795 (N_5795,N_5496,N_5058);
nor U5796 (N_5796,N_5109,N_5076);
nor U5797 (N_5797,N_5454,N_5372);
xnor U5798 (N_5798,N_5445,N_5354);
nand U5799 (N_5799,N_5069,N_5058);
or U5800 (N_5800,N_5121,N_5481);
or U5801 (N_5801,N_5218,N_5267);
nor U5802 (N_5802,N_5141,N_5190);
xnor U5803 (N_5803,N_5185,N_5083);
or U5804 (N_5804,N_5327,N_5268);
nand U5805 (N_5805,N_5110,N_5317);
nand U5806 (N_5806,N_5426,N_5254);
nor U5807 (N_5807,N_5380,N_5196);
and U5808 (N_5808,N_5156,N_5086);
nand U5809 (N_5809,N_5186,N_5223);
and U5810 (N_5810,N_5470,N_5145);
nor U5811 (N_5811,N_5487,N_5321);
or U5812 (N_5812,N_5469,N_5408);
nor U5813 (N_5813,N_5187,N_5154);
or U5814 (N_5814,N_5121,N_5183);
and U5815 (N_5815,N_5373,N_5384);
nand U5816 (N_5816,N_5131,N_5006);
or U5817 (N_5817,N_5228,N_5054);
or U5818 (N_5818,N_5219,N_5388);
nand U5819 (N_5819,N_5223,N_5133);
or U5820 (N_5820,N_5419,N_5488);
xor U5821 (N_5821,N_5299,N_5381);
nand U5822 (N_5822,N_5265,N_5092);
xnor U5823 (N_5823,N_5463,N_5008);
or U5824 (N_5824,N_5279,N_5439);
nor U5825 (N_5825,N_5199,N_5205);
nor U5826 (N_5826,N_5223,N_5122);
nand U5827 (N_5827,N_5350,N_5214);
nand U5828 (N_5828,N_5115,N_5276);
nand U5829 (N_5829,N_5307,N_5354);
or U5830 (N_5830,N_5370,N_5449);
nor U5831 (N_5831,N_5365,N_5180);
nand U5832 (N_5832,N_5357,N_5440);
and U5833 (N_5833,N_5361,N_5283);
or U5834 (N_5834,N_5061,N_5084);
and U5835 (N_5835,N_5111,N_5407);
nand U5836 (N_5836,N_5497,N_5243);
and U5837 (N_5837,N_5063,N_5024);
nand U5838 (N_5838,N_5056,N_5015);
and U5839 (N_5839,N_5125,N_5050);
nor U5840 (N_5840,N_5100,N_5430);
or U5841 (N_5841,N_5079,N_5048);
nor U5842 (N_5842,N_5093,N_5486);
xnor U5843 (N_5843,N_5178,N_5276);
xor U5844 (N_5844,N_5226,N_5127);
nand U5845 (N_5845,N_5272,N_5050);
nor U5846 (N_5846,N_5457,N_5201);
or U5847 (N_5847,N_5495,N_5051);
nand U5848 (N_5848,N_5303,N_5218);
and U5849 (N_5849,N_5002,N_5434);
or U5850 (N_5850,N_5028,N_5487);
nand U5851 (N_5851,N_5385,N_5014);
nor U5852 (N_5852,N_5099,N_5480);
nand U5853 (N_5853,N_5408,N_5431);
or U5854 (N_5854,N_5139,N_5165);
and U5855 (N_5855,N_5262,N_5260);
nand U5856 (N_5856,N_5440,N_5336);
and U5857 (N_5857,N_5294,N_5082);
nor U5858 (N_5858,N_5355,N_5066);
nand U5859 (N_5859,N_5051,N_5397);
nand U5860 (N_5860,N_5139,N_5454);
or U5861 (N_5861,N_5488,N_5150);
or U5862 (N_5862,N_5256,N_5453);
or U5863 (N_5863,N_5057,N_5246);
nor U5864 (N_5864,N_5461,N_5448);
nor U5865 (N_5865,N_5258,N_5263);
nand U5866 (N_5866,N_5327,N_5425);
or U5867 (N_5867,N_5118,N_5221);
nand U5868 (N_5868,N_5057,N_5228);
nand U5869 (N_5869,N_5043,N_5375);
and U5870 (N_5870,N_5178,N_5457);
and U5871 (N_5871,N_5239,N_5016);
or U5872 (N_5872,N_5279,N_5300);
xor U5873 (N_5873,N_5444,N_5156);
nor U5874 (N_5874,N_5406,N_5314);
and U5875 (N_5875,N_5189,N_5253);
and U5876 (N_5876,N_5189,N_5481);
and U5877 (N_5877,N_5298,N_5241);
and U5878 (N_5878,N_5273,N_5076);
nor U5879 (N_5879,N_5071,N_5470);
nand U5880 (N_5880,N_5297,N_5486);
or U5881 (N_5881,N_5327,N_5454);
nor U5882 (N_5882,N_5400,N_5228);
or U5883 (N_5883,N_5351,N_5382);
nor U5884 (N_5884,N_5289,N_5417);
and U5885 (N_5885,N_5183,N_5357);
nand U5886 (N_5886,N_5445,N_5236);
and U5887 (N_5887,N_5246,N_5122);
and U5888 (N_5888,N_5427,N_5196);
and U5889 (N_5889,N_5272,N_5195);
and U5890 (N_5890,N_5090,N_5495);
xnor U5891 (N_5891,N_5033,N_5441);
or U5892 (N_5892,N_5263,N_5208);
and U5893 (N_5893,N_5367,N_5291);
and U5894 (N_5894,N_5449,N_5366);
xnor U5895 (N_5895,N_5077,N_5398);
and U5896 (N_5896,N_5159,N_5328);
nor U5897 (N_5897,N_5277,N_5362);
nand U5898 (N_5898,N_5063,N_5204);
nor U5899 (N_5899,N_5415,N_5046);
nor U5900 (N_5900,N_5390,N_5315);
nor U5901 (N_5901,N_5061,N_5470);
or U5902 (N_5902,N_5464,N_5256);
nor U5903 (N_5903,N_5082,N_5103);
nand U5904 (N_5904,N_5350,N_5042);
and U5905 (N_5905,N_5189,N_5022);
nand U5906 (N_5906,N_5241,N_5191);
nor U5907 (N_5907,N_5404,N_5049);
or U5908 (N_5908,N_5398,N_5145);
xnor U5909 (N_5909,N_5058,N_5414);
nor U5910 (N_5910,N_5204,N_5246);
xnor U5911 (N_5911,N_5332,N_5108);
and U5912 (N_5912,N_5174,N_5118);
or U5913 (N_5913,N_5016,N_5049);
or U5914 (N_5914,N_5280,N_5275);
nor U5915 (N_5915,N_5253,N_5037);
or U5916 (N_5916,N_5304,N_5250);
nand U5917 (N_5917,N_5132,N_5215);
and U5918 (N_5918,N_5336,N_5466);
nor U5919 (N_5919,N_5159,N_5058);
and U5920 (N_5920,N_5480,N_5094);
nor U5921 (N_5921,N_5444,N_5281);
and U5922 (N_5922,N_5188,N_5116);
nand U5923 (N_5923,N_5017,N_5455);
or U5924 (N_5924,N_5430,N_5390);
and U5925 (N_5925,N_5252,N_5471);
nor U5926 (N_5926,N_5088,N_5413);
nand U5927 (N_5927,N_5110,N_5104);
or U5928 (N_5928,N_5453,N_5176);
nand U5929 (N_5929,N_5426,N_5340);
nor U5930 (N_5930,N_5175,N_5248);
nand U5931 (N_5931,N_5112,N_5080);
nand U5932 (N_5932,N_5229,N_5222);
nand U5933 (N_5933,N_5213,N_5102);
nor U5934 (N_5934,N_5139,N_5411);
and U5935 (N_5935,N_5486,N_5226);
and U5936 (N_5936,N_5000,N_5169);
and U5937 (N_5937,N_5300,N_5028);
xor U5938 (N_5938,N_5490,N_5375);
and U5939 (N_5939,N_5117,N_5078);
or U5940 (N_5940,N_5060,N_5137);
nor U5941 (N_5941,N_5046,N_5388);
xnor U5942 (N_5942,N_5295,N_5437);
nor U5943 (N_5943,N_5111,N_5266);
or U5944 (N_5944,N_5436,N_5240);
nor U5945 (N_5945,N_5392,N_5266);
or U5946 (N_5946,N_5165,N_5014);
or U5947 (N_5947,N_5195,N_5301);
or U5948 (N_5948,N_5384,N_5029);
and U5949 (N_5949,N_5175,N_5029);
or U5950 (N_5950,N_5286,N_5346);
and U5951 (N_5951,N_5032,N_5489);
nor U5952 (N_5952,N_5493,N_5219);
or U5953 (N_5953,N_5104,N_5125);
and U5954 (N_5954,N_5218,N_5301);
or U5955 (N_5955,N_5330,N_5191);
nand U5956 (N_5956,N_5362,N_5282);
nand U5957 (N_5957,N_5227,N_5263);
xnor U5958 (N_5958,N_5351,N_5060);
nor U5959 (N_5959,N_5279,N_5184);
or U5960 (N_5960,N_5435,N_5316);
or U5961 (N_5961,N_5280,N_5477);
or U5962 (N_5962,N_5101,N_5050);
or U5963 (N_5963,N_5151,N_5137);
nor U5964 (N_5964,N_5415,N_5318);
or U5965 (N_5965,N_5045,N_5456);
nor U5966 (N_5966,N_5118,N_5099);
or U5967 (N_5967,N_5087,N_5230);
and U5968 (N_5968,N_5177,N_5013);
and U5969 (N_5969,N_5030,N_5416);
xor U5970 (N_5970,N_5137,N_5309);
and U5971 (N_5971,N_5484,N_5117);
xnor U5972 (N_5972,N_5364,N_5324);
nor U5973 (N_5973,N_5407,N_5499);
and U5974 (N_5974,N_5113,N_5218);
and U5975 (N_5975,N_5381,N_5352);
or U5976 (N_5976,N_5399,N_5218);
nor U5977 (N_5977,N_5134,N_5251);
xor U5978 (N_5978,N_5249,N_5366);
xnor U5979 (N_5979,N_5266,N_5472);
nand U5980 (N_5980,N_5396,N_5140);
nand U5981 (N_5981,N_5197,N_5404);
and U5982 (N_5982,N_5186,N_5384);
nand U5983 (N_5983,N_5174,N_5473);
nand U5984 (N_5984,N_5281,N_5172);
or U5985 (N_5985,N_5218,N_5077);
nor U5986 (N_5986,N_5113,N_5481);
xor U5987 (N_5987,N_5350,N_5163);
or U5988 (N_5988,N_5463,N_5301);
nor U5989 (N_5989,N_5171,N_5036);
nand U5990 (N_5990,N_5023,N_5076);
nor U5991 (N_5991,N_5415,N_5240);
and U5992 (N_5992,N_5208,N_5128);
or U5993 (N_5993,N_5482,N_5152);
or U5994 (N_5994,N_5141,N_5094);
and U5995 (N_5995,N_5120,N_5404);
xor U5996 (N_5996,N_5284,N_5315);
nand U5997 (N_5997,N_5063,N_5098);
or U5998 (N_5998,N_5183,N_5345);
nor U5999 (N_5999,N_5114,N_5049);
nand U6000 (N_6000,N_5922,N_5635);
nor U6001 (N_6001,N_5529,N_5742);
nor U6002 (N_6002,N_5897,N_5915);
or U6003 (N_6003,N_5599,N_5739);
nor U6004 (N_6004,N_5910,N_5592);
nand U6005 (N_6005,N_5824,N_5993);
nor U6006 (N_6006,N_5530,N_5821);
and U6007 (N_6007,N_5947,N_5532);
nor U6008 (N_6008,N_5655,N_5623);
and U6009 (N_6009,N_5698,N_5841);
and U6010 (N_6010,N_5856,N_5893);
or U6011 (N_6011,N_5810,N_5773);
nand U6012 (N_6012,N_5694,N_5997);
nor U6013 (N_6013,N_5878,N_5836);
or U6014 (N_6014,N_5746,N_5781);
or U6015 (N_6015,N_5526,N_5958);
nand U6016 (N_6016,N_5525,N_5660);
nand U6017 (N_6017,N_5743,N_5653);
and U6018 (N_6018,N_5617,N_5735);
and U6019 (N_6019,N_5516,N_5760);
nand U6020 (N_6020,N_5846,N_5828);
xor U6021 (N_6021,N_5757,N_5896);
and U6022 (N_6022,N_5848,N_5785);
or U6023 (N_6023,N_5511,N_5581);
nand U6024 (N_6024,N_5590,N_5789);
nor U6025 (N_6025,N_5942,N_5974);
and U6026 (N_6026,N_5800,N_5969);
xnor U6027 (N_6027,N_5827,N_5538);
nand U6028 (N_6028,N_5798,N_5913);
or U6029 (N_6029,N_5718,N_5555);
and U6030 (N_6030,N_5920,N_5933);
and U6031 (N_6031,N_5730,N_5895);
or U6032 (N_6032,N_5639,N_5971);
or U6033 (N_6033,N_5570,N_5979);
xnor U6034 (N_6034,N_5713,N_5531);
nor U6035 (N_6035,N_5797,N_5952);
nand U6036 (N_6036,N_5954,N_5812);
nor U6037 (N_6037,N_5731,N_5962);
nand U6038 (N_6038,N_5948,N_5792);
nand U6039 (N_6039,N_5700,N_5990);
nand U6040 (N_6040,N_5680,N_5949);
and U6041 (N_6041,N_5862,N_5884);
nand U6042 (N_6042,N_5683,N_5647);
or U6043 (N_6043,N_5692,N_5833);
xor U6044 (N_6044,N_5853,N_5507);
nand U6045 (N_6045,N_5543,N_5609);
or U6046 (N_6046,N_5972,N_5927);
or U6047 (N_6047,N_5634,N_5811);
nor U6048 (N_6048,N_5867,N_5665);
or U6049 (N_6049,N_5989,N_5726);
and U6050 (N_6050,N_5957,N_5676);
or U6051 (N_6051,N_5766,N_5500);
or U6052 (N_6052,N_5548,N_5638);
nor U6053 (N_6053,N_5956,N_5847);
nor U6054 (N_6054,N_5747,N_5835);
nor U6055 (N_6055,N_5780,N_5807);
nor U6056 (N_6056,N_5549,N_5678);
nand U6057 (N_6057,N_5541,N_5759);
nand U6058 (N_6058,N_5652,N_5911);
and U6059 (N_6059,N_5783,N_5980);
and U6060 (N_6060,N_5691,N_5641);
and U6061 (N_6061,N_5814,N_5578);
nor U6062 (N_6062,N_5805,N_5734);
or U6063 (N_6063,N_5615,N_5685);
or U6064 (N_6064,N_5951,N_5554);
or U6065 (N_6065,N_5955,N_5898);
nand U6066 (N_6066,N_5575,N_5918);
and U6067 (N_6067,N_5518,N_5619);
nand U6068 (N_6068,N_5630,N_5673);
and U6069 (N_6069,N_5816,N_5857);
nand U6070 (N_6070,N_5544,N_5854);
and U6071 (N_6071,N_5813,N_5715);
nand U6072 (N_6072,N_5991,N_5968);
nor U6073 (N_6073,N_5697,N_5642);
and U6074 (N_6074,N_5565,N_5643);
or U6075 (N_6075,N_5782,N_5964);
nor U6076 (N_6076,N_5690,N_5926);
or U6077 (N_6077,N_5901,N_5605);
nor U6078 (N_6078,N_5576,N_5675);
nor U6079 (N_6079,N_5902,N_5657);
and U6080 (N_6080,N_5719,N_5745);
or U6081 (N_6081,N_5618,N_5784);
nor U6082 (N_6082,N_5880,N_5793);
nand U6083 (N_6083,N_5999,N_5596);
xor U6084 (N_6084,N_5661,N_5706);
or U6085 (N_6085,N_5716,N_5855);
nor U6086 (N_6086,N_5899,N_5961);
nor U6087 (N_6087,N_5817,N_5629);
nor U6088 (N_6088,N_5737,N_5662);
xor U6089 (N_6089,N_5561,N_5975);
nand U6090 (N_6090,N_5939,N_5936);
or U6091 (N_6091,N_5876,N_5869);
nor U6092 (N_6092,N_5912,N_5754);
nand U6093 (N_6093,N_5938,N_5625);
nor U6094 (N_6094,N_5967,N_5577);
nand U6095 (N_6095,N_5602,N_5668);
nand U6096 (N_6096,N_5900,N_5996);
and U6097 (N_6097,N_5689,N_5574);
or U6098 (N_6098,N_5527,N_5707);
and U6099 (N_6099,N_5891,N_5935);
and U6100 (N_6100,N_5520,N_5654);
or U6101 (N_6101,N_5904,N_5571);
and U6102 (N_6102,N_5658,N_5567);
nor U6103 (N_6103,N_5569,N_5748);
and U6104 (N_6104,N_5677,N_5708);
or U6105 (N_6105,N_5514,N_5723);
and U6106 (N_6106,N_5950,N_5981);
and U6107 (N_6107,N_5681,N_5553);
nor U6108 (N_6108,N_5725,N_5883);
nor U6109 (N_6109,N_5998,N_5732);
xnor U6110 (N_6110,N_5589,N_5930);
nand U6111 (N_6111,N_5579,N_5542);
and U6112 (N_6112,N_5551,N_5533);
or U6113 (N_6113,N_5843,N_5712);
nand U6114 (N_6114,N_5545,N_5872);
xor U6115 (N_6115,N_5562,N_5776);
xor U6116 (N_6116,N_5838,N_5837);
or U6117 (N_6117,N_5767,N_5803);
and U6118 (N_6118,N_5907,N_5744);
and U6119 (N_6119,N_5620,N_5585);
and U6120 (N_6120,N_5830,N_5870);
and U6121 (N_6121,N_5818,N_5995);
nand U6122 (N_6122,N_5953,N_5674);
nor U6123 (N_6123,N_5563,N_5916);
and U6124 (N_6124,N_5945,N_5826);
nor U6125 (N_6125,N_5963,N_5510);
nand U6126 (N_6126,N_5842,N_5977);
nand U6127 (N_6127,N_5850,N_5779);
and U6128 (N_6128,N_5517,N_5566);
nor U6129 (N_6129,N_5670,N_5769);
or U6130 (N_6130,N_5909,N_5886);
xnor U6131 (N_6131,N_5502,N_5787);
nand U6132 (N_6132,N_5522,N_5573);
nand U6133 (N_6133,N_5931,N_5663);
and U6134 (N_6134,N_5687,N_5626);
and U6135 (N_6135,N_5671,N_5628);
nand U6136 (N_6136,N_5815,N_5705);
xnor U6137 (N_6137,N_5774,N_5925);
nor U6138 (N_6138,N_5515,N_5825);
and U6139 (N_6139,N_5940,N_5840);
or U6140 (N_6140,N_5829,N_5651);
nor U6141 (N_6141,N_5863,N_5908);
or U6142 (N_6142,N_5921,N_5738);
nor U6143 (N_6143,N_5688,N_5831);
and U6144 (N_6144,N_5944,N_5582);
nand U6145 (N_6145,N_5640,N_5546);
nand U6146 (N_6146,N_5804,N_5636);
and U6147 (N_6147,N_5859,N_5959);
and U6148 (N_6148,N_5988,N_5729);
nor U6149 (N_6149,N_5695,N_5875);
nand U6150 (N_6150,N_5888,N_5524);
nor U6151 (N_6151,N_5976,N_5994);
and U6152 (N_6152,N_5978,N_5604);
and U6153 (N_6153,N_5984,N_5645);
and U6154 (N_6154,N_5598,N_5871);
or U6155 (N_6155,N_5568,N_5986);
nand U6156 (N_6156,N_5672,N_5889);
or U6157 (N_6157,N_5597,N_5905);
and U6158 (N_6158,N_5556,N_5664);
and U6159 (N_6159,N_5914,N_5591);
nand U6160 (N_6160,N_5801,N_5616);
xnor U6161 (N_6161,N_5970,N_5627);
nand U6162 (N_6162,N_5540,N_5513);
and U6163 (N_6163,N_5584,N_5587);
nor U6164 (N_6164,N_5868,N_5644);
and U6165 (N_6165,N_5865,N_5667);
or U6166 (N_6166,N_5777,N_5666);
nand U6167 (N_6167,N_5560,N_5758);
or U6168 (N_6168,N_5761,N_5637);
and U6169 (N_6169,N_5534,N_5874);
or U6170 (N_6170,N_5822,N_5771);
nand U6171 (N_6171,N_5682,N_5608);
and U6172 (N_6172,N_5588,N_5937);
nand U6173 (N_6173,N_5832,N_5790);
nor U6174 (N_6174,N_5523,N_5621);
nor U6175 (N_6175,N_5794,N_5704);
nand U6176 (N_6176,N_5946,N_5844);
or U6177 (N_6177,N_5547,N_5923);
nor U6178 (N_6178,N_5624,N_5508);
or U6179 (N_6179,N_5504,N_5686);
nor U6180 (N_6180,N_5772,N_5966);
nor U6181 (N_6181,N_5752,N_5903);
or U6182 (N_6182,N_5756,N_5802);
nand U6183 (N_6183,N_5724,N_5786);
or U6184 (N_6184,N_5834,N_5808);
nor U6185 (N_6185,N_5890,N_5934);
nor U6186 (N_6186,N_5528,N_5762);
or U6187 (N_6187,N_5750,N_5509);
nor U6188 (N_6188,N_5741,N_5659);
and U6189 (N_6189,N_5572,N_5506);
and U6190 (N_6190,N_5535,N_5632);
xor U6191 (N_6191,N_5932,N_5985);
and U6192 (N_6192,N_5894,N_5613);
and U6193 (N_6193,N_5823,N_5622);
nand U6194 (N_6194,N_5631,N_5799);
nor U6195 (N_6195,N_5722,N_5558);
nand U6196 (N_6196,N_5603,N_5879);
and U6197 (N_6197,N_5749,N_5648);
nor U6198 (N_6198,N_5633,N_5877);
and U6199 (N_6199,N_5965,N_5650);
and U6200 (N_6200,N_5649,N_5564);
and U6201 (N_6201,N_5537,N_5882);
nand U6202 (N_6202,N_5796,N_5519);
nor U6203 (N_6203,N_5924,N_5768);
and U6204 (N_6204,N_5881,N_5646);
nor U6205 (N_6205,N_5552,N_5987);
or U6206 (N_6206,N_5791,N_5607);
or U6207 (N_6207,N_5941,N_5806);
or U6208 (N_6208,N_5919,N_5559);
nand U6209 (N_6209,N_5736,N_5550);
or U6210 (N_6210,N_5778,N_5819);
nand U6211 (N_6211,N_5892,N_5885);
nand U6212 (N_6212,N_5610,N_5536);
and U6213 (N_6213,N_5714,N_5809);
or U6214 (N_6214,N_5765,N_5611);
or U6215 (N_6215,N_5727,N_5866);
or U6216 (N_6216,N_5612,N_5860);
nor U6217 (N_6217,N_5770,N_5928);
nand U6218 (N_6218,N_5852,N_5594);
nor U6219 (N_6219,N_5503,N_5788);
xnor U6220 (N_6220,N_5693,N_5539);
nand U6221 (N_6221,N_5557,N_5764);
nor U6222 (N_6222,N_5600,N_5728);
nor U6223 (N_6223,N_5669,N_5703);
xor U6224 (N_6224,N_5709,N_5861);
xnor U6225 (N_6225,N_5753,N_5795);
and U6226 (N_6226,N_5501,N_5614);
and U6227 (N_6227,N_5858,N_5906);
nand U6228 (N_6228,N_5721,N_5755);
or U6229 (N_6229,N_5586,N_5717);
or U6230 (N_6230,N_5943,N_5580);
xor U6231 (N_6231,N_5505,N_5701);
nor U6232 (N_6232,N_5820,N_5851);
nand U6233 (N_6233,N_5702,N_5595);
and U6234 (N_6234,N_5696,N_5711);
nand U6235 (N_6235,N_5720,N_5751);
and U6236 (N_6236,N_5992,N_5929);
nand U6237 (N_6237,N_5775,N_5960);
nand U6238 (N_6238,N_5873,N_5512);
nand U6239 (N_6239,N_5740,N_5763);
nor U6240 (N_6240,N_5887,N_5521);
nor U6241 (N_6241,N_5684,N_5845);
xor U6242 (N_6242,N_5699,N_5849);
xor U6243 (N_6243,N_5733,N_5656);
nand U6244 (N_6244,N_5679,N_5983);
nor U6245 (N_6245,N_5864,N_5973);
nor U6246 (N_6246,N_5710,N_5606);
nand U6247 (N_6247,N_5982,N_5839);
nor U6248 (N_6248,N_5583,N_5917);
nor U6249 (N_6249,N_5593,N_5601);
and U6250 (N_6250,N_5674,N_5858);
nor U6251 (N_6251,N_5767,N_5859);
nor U6252 (N_6252,N_5642,N_5803);
or U6253 (N_6253,N_5611,N_5820);
nand U6254 (N_6254,N_5991,N_5762);
nand U6255 (N_6255,N_5561,N_5820);
and U6256 (N_6256,N_5551,N_5526);
or U6257 (N_6257,N_5717,N_5707);
nor U6258 (N_6258,N_5861,N_5722);
nand U6259 (N_6259,N_5845,N_5824);
xor U6260 (N_6260,N_5923,N_5573);
nor U6261 (N_6261,N_5502,N_5536);
and U6262 (N_6262,N_5805,N_5898);
or U6263 (N_6263,N_5809,N_5633);
and U6264 (N_6264,N_5976,N_5879);
and U6265 (N_6265,N_5967,N_5817);
or U6266 (N_6266,N_5817,N_5822);
nor U6267 (N_6267,N_5959,N_5829);
or U6268 (N_6268,N_5805,N_5753);
or U6269 (N_6269,N_5932,N_5753);
nand U6270 (N_6270,N_5575,N_5513);
and U6271 (N_6271,N_5710,N_5922);
nor U6272 (N_6272,N_5738,N_5963);
and U6273 (N_6273,N_5941,N_5705);
xnor U6274 (N_6274,N_5870,N_5854);
xor U6275 (N_6275,N_5589,N_5944);
nor U6276 (N_6276,N_5955,N_5892);
nor U6277 (N_6277,N_5627,N_5654);
or U6278 (N_6278,N_5561,N_5526);
nor U6279 (N_6279,N_5840,N_5806);
nor U6280 (N_6280,N_5528,N_5586);
and U6281 (N_6281,N_5642,N_5886);
nor U6282 (N_6282,N_5636,N_5795);
xnor U6283 (N_6283,N_5691,N_5723);
xor U6284 (N_6284,N_5833,N_5613);
xnor U6285 (N_6285,N_5542,N_5891);
nand U6286 (N_6286,N_5917,N_5960);
nor U6287 (N_6287,N_5758,N_5539);
nand U6288 (N_6288,N_5673,N_5961);
nor U6289 (N_6289,N_5767,N_5515);
and U6290 (N_6290,N_5646,N_5764);
nor U6291 (N_6291,N_5714,N_5524);
xnor U6292 (N_6292,N_5649,N_5972);
or U6293 (N_6293,N_5889,N_5750);
or U6294 (N_6294,N_5501,N_5588);
nand U6295 (N_6295,N_5559,N_5870);
or U6296 (N_6296,N_5751,N_5923);
nor U6297 (N_6297,N_5885,N_5729);
and U6298 (N_6298,N_5978,N_5677);
nand U6299 (N_6299,N_5580,N_5876);
and U6300 (N_6300,N_5551,N_5725);
xnor U6301 (N_6301,N_5658,N_5653);
nor U6302 (N_6302,N_5767,N_5762);
and U6303 (N_6303,N_5789,N_5512);
nand U6304 (N_6304,N_5562,N_5655);
nor U6305 (N_6305,N_5892,N_5995);
nand U6306 (N_6306,N_5813,N_5878);
nor U6307 (N_6307,N_5632,N_5798);
and U6308 (N_6308,N_5790,N_5559);
nand U6309 (N_6309,N_5619,N_5902);
and U6310 (N_6310,N_5956,N_5881);
and U6311 (N_6311,N_5698,N_5826);
and U6312 (N_6312,N_5641,N_5518);
or U6313 (N_6313,N_5662,N_5632);
nor U6314 (N_6314,N_5802,N_5744);
nor U6315 (N_6315,N_5959,N_5878);
or U6316 (N_6316,N_5634,N_5802);
nand U6317 (N_6317,N_5929,N_5546);
or U6318 (N_6318,N_5771,N_5690);
nand U6319 (N_6319,N_5847,N_5733);
nand U6320 (N_6320,N_5647,N_5977);
or U6321 (N_6321,N_5878,N_5891);
or U6322 (N_6322,N_5868,N_5699);
nand U6323 (N_6323,N_5902,N_5926);
nor U6324 (N_6324,N_5916,N_5796);
nand U6325 (N_6325,N_5794,N_5910);
and U6326 (N_6326,N_5785,N_5907);
nor U6327 (N_6327,N_5609,N_5722);
or U6328 (N_6328,N_5611,N_5614);
and U6329 (N_6329,N_5800,N_5920);
nand U6330 (N_6330,N_5736,N_5571);
nand U6331 (N_6331,N_5835,N_5976);
and U6332 (N_6332,N_5762,N_5830);
or U6333 (N_6333,N_5659,N_5813);
nor U6334 (N_6334,N_5568,N_5801);
xor U6335 (N_6335,N_5861,N_5833);
xor U6336 (N_6336,N_5877,N_5926);
and U6337 (N_6337,N_5811,N_5739);
xor U6338 (N_6338,N_5834,N_5984);
and U6339 (N_6339,N_5848,N_5892);
or U6340 (N_6340,N_5930,N_5522);
nor U6341 (N_6341,N_5658,N_5642);
nand U6342 (N_6342,N_5980,N_5745);
nand U6343 (N_6343,N_5733,N_5514);
and U6344 (N_6344,N_5703,N_5667);
or U6345 (N_6345,N_5836,N_5630);
nand U6346 (N_6346,N_5735,N_5925);
and U6347 (N_6347,N_5885,N_5970);
nor U6348 (N_6348,N_5905,N_5654);
nor U6349 (N_6349,N_5970,N_5869);
nor U6350 (N_6350,N_5954,N_5675);
nand U6351 (N_6351,N_5567,N_5783);
nand U6352 (N_6352,N_5984,N_5822);
and U6353 (N_6353,N_5972,N_5568);
nor U6354 (N_6354,N_5628,N_5632);
nor U6355 (N_6355,N_5703,N_5602);
nand U6356 (N_6356,N_5759,N_5686);
nor U6357 (N_6357,N_5733,N_5630);
and U6358 (N_6358,N_5886,N_5790);
or U6359 (N_6359,N_5812,N_5789);
nand U6360 (N_6360,N_5929,N_5597);
nor U6361 (N_6361,N_5548,N_5806);
nand U6362 (N_6362,N_5838,N_5699);
nor U6363 (N_6363,N_5888,N_5520);
or U6364 (N_6364,N_5710,N_5759);
and U6365 (N_6365,N_5702,N_5510);
nand U6366 (N_6366,N_5751,N_5730);
and U6367 (N_6367,N_5633,N_5862);
nand U6368 (N_6368,N_5806,N_5656);
xor U6369 (N_6369,N_5746,N_5665);
nand U6370 (N_6370,N_5770,N_5649);
or U6371 (N_6371,N_5978,N_5903);
and U6372 (N_6372,N_5857,N_5528);
nand U6373 (N_6373,N_5629,N_5501);
nand U6374 (N_6374,N_5657,N_5845);
and U6375 (N_6375,N_5874,N_5709);
or U6376 (N_6376,N_5839,N_5561);
nor U6377 (N_6377,N_5855,N_5624);
nand U6378 (N_6378,N_5860,N_5963);
nor U6379 (N_6379,N_5739,N_5675);
nand U6380 (N_6380,N_5787,N_5542);
nor U6381 (N_6381,N_5606,N_5503);
nor U6382 (N_6382,N_5670,N_5530);
nand U6383 (N_6383,N_5680,N_5990);
nor U6384 (N_6384,N_5941,N_5640);
and U6385 (N_6385,N_5586,N_5864);
and U6386 (N_6386,N_5667,N_5898);
nor U6387 (N_6387,N_5760,N_5755);
and U6388 (N_6388,N_5761,N_5670);
nand U6389 (N_6389,N_5569,N_5795);
or U6390 (N_6390,N_5651,N_5962);
and U6391 (N_6391,N_5676,N_5751);
and U6392 (N_6392,N_5647,N_5881);
and U6393 (N_6393,N_5738,N_5619);
nor U6394 (N_6394,N_5664,N_5861);
or U6395 (N_6395,N_5892,N_5521);
nand U6396 (N_6396,N_5666,N_5967);
nor U6397 (N_6397,N_5647,N_5791);
and U6398 (N_6398,N_5664,N_5518);
nand U6399 (N_6399,N_5680,N_5873);
nor U6400 (N_6400,N_5985,N_5918);
nand U6401 (N_6401,N_5711,N_5875);
or U6402 (N_6402,N_5792,N_5895);
nor U6403 (N_6403,N_5889,N_5712);
and U6404 (N_6404,N_5886,N_5645);
and U6405 (N_6405,N_5998,N_5725);
and U6406 (N_6406,N_5812,N_5736);
or U6407 (N_6407,N_5936,N_5814);
nand U6408 (N_6408,N_5549,N_5635);
and U6409 (N_6409,N_5510,N_5761);
and U6410 (N_6410,N_5504,N_5545);
or U6411 (N_6411,N_5540,N_5968);
nand U6412 (N_6412,N_5972,N_5936);
and U6413 (N_6413,N_5687,N_5746);
or U6414 (N_6414,N_5848,N_5910);
xor U6415 (N_6415,N_5899,N_5533);
or U6416 (N_6416,N_5875,N_5934);
nand U6417 (N_6417,N_5537,N_5621);
xor U6418 (N_6418,N_5918,N_5688);
xor U6419 (N_6419,N_5801,N_5885);
nor U6420 (N_6420,N_5800,N_5905);
xnor U6421 (N_6421,N_5940,N_5816);
or U6422 (N_6422,N_5966,N_5716);
and U6423 (N_6423,N_5924,N_5566);
and U6424 (N_6424,N_5553,N_5618);
xnor U6425 (N_6425,N_5721,N_5799);
or U6426 (N_6426,N_5566,N_5597);
or U6427 (N_6427,N_5930,N_5513);
nor U6428 (N_6428,N_5636,N_5544);
or U6429 (N_6429,N_5542,N_5669);
and U6430 (N_6430,N_5715,N_5758);
nand U6431 (N_6431,N_5661,N_5819);
and U6432 (N_6432,N_5842,N_5677);
and U6433 (N_6433,N_5695,N_5828);
and U6434 (N_6434,N_5613,N_5862);
nand U6435 (N_6435,N_5774,N_5539);
nand U6436 (N_6436,N_5559,N_5603);
nand U6437 (N_6437,N_5905,N_5906);
nand U6438 (N_6438,N_5521,N_5503);
nand U6439 (N_6439,N_5910,N_5741);
or U6440 (N_6440,N_5500,N_5546);
nand U6441 (N_6441,N_5736,N_5872);
nand U6442 (N_6442,N_5584,N_5980);
or U6443 (N_6443,N_5733,N_5688);
nand U6444 (N_6444,N_5722,N_5928);
or U6445 (N_6445,N_5752,N_5839);
nand U6446 (N_6446,N_5651,N_5804);
and U6447 (N_6447,N_5854,N_5729);
and U6448 (N_6448,N_5790,N_5517);
xor U6449 (N_6449,N_5713,N_5914);
nor U6450 (N_6450,N_5783,N_5762);
and U6451 (N_6451,N_5593,N_5855);
or U6452 (N_6452,N_5556,N_5500);
xor U6453 (N_6453,N_5819,N_5582);
nor U6454 (N_6454,N_5660,N_5889);
nor U6455 (N_6455,N_5982,N_5762);
or U6456 (N_6456,N_5762,N_5611);
nand U6457 (N_6457,N_5519,N_5548);
nor U6458 (N_6458,N_5625,N_5607);
and U6459 (N_6459,N_5637,N_5643);
nor U6460 (N_6460,N_5604,N_5960);
and U6461 (N_6461,N_5937,N_5513);
and U6462 (N_6462,N_5813,N_5611);
xnor U6463 (N_6463,N_5712,N_5657);
nand U6464 (N_6464,N_5766,N_5981);
and U6465 (N_6465,N_5950,N_5832);
and U6466 (N_6466,N_5576,N_5940);
nand U6467 (N_6467,N_5647,N_5835);
or U6468 (N_6468,N_5571,N_5751);
nand U6469 (N_6469,N_5834,N_5966);
xor U6470 (N_6470,N_5785,N_5711);
nor U6471 (N_6471,N_5522,N_5628);
and U6472 (N_6472,N_5698,N_5504);
nand U6473 (N_6473,N_5963,N_5909);
nand U6474 (N_6474,N_5925,N_5710);
nor U6475 (N_6475,N_5935,N_5861);
nand U6476 (N_6476,N_5519,N_5615);
and U6477 (N_6477,N_5620,N_5613);
nor U6478 (N_6478,N_5566,N_5742);
and U6479 (N_6479,N_5596,N_5818);
nand U6480 (N_6480,N_5660,N_5555);
nor U6481 (N_6481,N_5626,N_5806);
nand U6482 (N_6482,N_5603,N_5866);
and U6483 (N_6483,N_5507,N_5598);
nand U6484 (N_6484,N_5947,N_5803);
or U6485 (N_6485,N_5690,N_5915);
nor U6486 (N_6486,N_5732,N_5521);
and U6487 (N_6487,N_5913,N_5721);
nand U6488 (N_6488,N_5598,N_5554);
nand U6489 (N_6489,N_5716,N_5856);
or U6490 (N_6490,N_5915,N_5903);
or U6491 (N_6491,N_5827,N_5841);
or U6492 (N_6492,N_5872,N_5925);
or U6493 (N_6493,N_5738,N_5909);
nor U6494 (N_6494,N_5784,N_5500);
xor U6495 (N_6495,N_5763,N_5664);
or U6496 (N_6496,N_5882,N_5900);
or U6497 (N_6497,N_5823,N_5922);
and U6498 (N_6498,N_5590,N_5642);
xor U6499 (N_6499,N_5775,N_5569);
xnor U6500 (N_6500,N_6361,N_6133);
xnor U6501 (N_6501,N_6107,N_6355);
nand U6502 (N_6502,N_6138,N_6165);
and U6503 (N_6503,N_6073,N_6384);
nand U6504 (N_6504,N_6452,N_6425);
nand U6505 (N_6505,N_6345,N_6113);
nand U6506 (N_6506,N_6144,N_6053);
nor U6507 (N_6507,N_6310,N_6221);
nand U6508 (N_6508,N_6022,N_6397);
or U6509 (N_6509,N_6434,N_6206);
nand U6510 (N_6510,N_6489,N_6088);
nor U6511 (N_6511,N_6120,N_6481);
nand U6512 (N_6512,N_6150,N_6155);
or U6513 (N_6513,N_6328,N_6395);
or U6514 (N_6514,N_6400,N_6075);
or U6515 (N_6515,N_6391,N_6202);
nand U6516 (N_6516,N_6068,N_6339);
nor U6517 (N_6517,N_6371,N_6314);
or U6518 (N_6518,N_6366,N_6326);
xor U6519 (N_6519,N_6055,N_6082);
nand U6520 (N_6520,N_6454,N_6418);
or U6521 (N_6521,N_6365,N_6143);
nand U6522 (N_6522,N_6278,N_6207);
nor U6523 (N_6523,N_6252,N_6342);
or U6524 (N_6524,N_6478,N_6367);
nor U6525 (N_6525,N_6200,N_6448);
nor U6526 (N_6526,N_6049,N_6389);
nand U6527 (N_6527,N_6069,N_6432);
and U6528 (N_6528,N_6370,N_6187);
or U6529 (N_6529,N_6343,N_6374);
or U6530 (N_6530,N_6334,N_6110);
nor U6531 (N_6531,N_6281,N_6080);
or U6532 (N_6532,N_6161,N_6424);
or U6533 (N_6533,N_6182,N_6014);
nor U6534 (N_6534,N_6316,N_6309);
and U6535 (N_6535,N_6140,N_6402);
or U6536 (N_6536,N_6231,N_6405);
nand U6537 (N_6537,N_6219,N_6387);
and U6538 (N_6538,N_6232,N_6142);
nor U6539 (N_6539,N_6280,N_6139);
nand U6540 (N_6540,N_6225,N_6214);
or U6541 (N_6541,N_6275,N_6290);
or U6542 (N_6542,N_6344,N_6050);
xnor U6543 (N_6543,N_6479,N_6490);
and U6544 (N_6544,N_6171,N_6153);
nor U6545 (N_6545,N_6018,N_6117);
nor U6546 (N_6546,N_6047,N_6054);
nor U6547 (N_6547,N_6414,N_6222);
and U6548 (N_6548,N_6484,N_6408);
nor U6549 (N_6549,N_6455,N_6060);
nor U6550 (N_6550,N_6382,N_6357);
nor U6551 (N_6551,N_6185,N_6091);
and U6552 (N_6552,N_6305,N_6295);
and U6553 (N_6553,N_6306,N_6460);
nand U6554 (N_6554,N_6026,N_6498);
nor U6555 (N_6555,N_6360,N_6246);
xor U6556 (N_6556,N_6058,N_6476);
nor U6557 (N_6557,N_6486,N_6495);
nor U6558 (N_6558,N_6488,N_6215);
and U6559 (N_6559,N_6103,N_6259);
or U6560 (N_6560,N_6403,N_6218);
or U6561 (N_6561,N_6304,N_6381);
nand U6562 (N_6562,N_6449,N_6040);
and U6563 (N_6563,N_6464,N_6429);
or U6564 (N_6564,N_6067,N_6065);
nor U6565 (N_6565,N_6390,N_6186);
or U6566 (N_6566,N_6427,N_6444);
nor U6567 (N_6567,N_6172,N_6205);
nand U6568 (N_6568,N_6269,N_6146);
nand U6569 (N_6569,N_6363,N_6124);
or U6570 (N_6570,N_6465,N_6019);
or U6571 (N_6571,N_6235,N_6213);
nor U6572 (N_6572,N_6072,N_6409);
nor U6573 (N_6573,N_6227,N_6028);
or U6574 (N_6574,N_6070,N_6102);
nor U6575 (N_6575,N_6445,N_6007);
xor U6576 (N_6576,N_6148,N_6496);
nand U6577 (N_6577,N_6000,N_6052);
or U6578 (N_6578,N_6211,N_6043);
nand U6579 (N_6579,N_6372,N_6085);
or U6580 (N_6580,N_6433,N_6106);
and U6581 (N_6581,N_6011,N_6201);
or U6582 (N_6582,N_6137,N_6272);
and U6583 (N_6583,N_6020,N_6157);
xor U6584 (N_6584,N_6356,N_6292);
and U6585 (N_6585,N_6216,N_6122);
nand U6586 (N_6586,N_6285,N_6482);
nand U6587 (N_6587,N_6288,N_6192);
or U6588 (N_6588,N_6457,N_6164);
and U6589 (N_6589,N_6025,N_6188);
or U6590 (N_6590,N_6181,N_6362);
and U6591 (N_6591,N_6447,N_6412);
nor U6592 (N_6592,N_6443,N_6034);
nand U6593 (N_6593,N_6430,N_6220);
nor U6594 (N_6594,N_6179,N_6250);
nor U6595 (N_6595,N_6112,N_6035);
nor U6596 (N_6596,N_6271,N_6475);
xnor U6597 (N_6597,N_6061,N_6247);
or U6598 (N_6598,N_6237,N_6251);
and U6599 (N_6599,N_6458,N_6262);
nor U6600 (N_6600,N_6287,N_6089);
and U6601 (N_6601,N_6123,N_6173);
nand U6602 (N_6602,N_6353,N_6062);
and U6603 (N_6603,N_6254,N_6177);
or U6604 (N_6604,N_6210,N_6036);
and U6605 (N_6605,N_6386,N_6266);
or U6606 (N_6606,N_6041,N_6168);
or U6607 (N_6607,N_6325,N_6086);
nor U6608 (N_6608,N_6166,N_6184);
and U6609 (N_6609,N_6337,N_6174);
or U6610 (N_6610,N_6241,N_6003);
nand U6611 (N_6611,N_6136,N_6079);
xnor U6612 (N_6612,N_6236,N_6493);
nand U6613 (N_6613,N_6456,N_6477);
and U6614 (N_6614,N_6491,N_6346);
nand U6615 (N_6615,N_6471,N_6422);
nand U6616 (N_6616,N_6240,N_6037);
xor U6617 (N_6617,N_6098,N_6135);
nand U6618 (N_6618,N_6063,N_6239);
or U6619 (N_6619,N_6300,N_6261);
nand U6620 (N_6620,N_6015,N_6027);
or U6621 (N_6621,N_6059,N_6109);
xor U6622 (N_6622,N_6335,N_6273);
nand U6623 (N_6623,N_6128,N_6466);
and U6624 (N_6624,N_6436,N_6338);
nor U6625 (N_6625,N_6132,N_6283);
xnor U6626 (N_6626,N_6212,N_6230);
or U6627 (N_6627,N_6039,N_6416);
or U6628 (N_6628,N_6031,N_6078);
and U6629 (N_6629,N_6233,N_6330);
and U6630 (N_6630,N_6291,N_6111);
nand U6631 (N_6631,N_6004,N_6130);
nand U6632 (N_6632,N_6198,N_6255);
or U6633 (N_6633,N_6263,N_6013);
or U6634 (N_6634,N_6473,N_6264);
nor U6635 (N_6635,N_6094,N_6302);
or U6636 (N_6636,N_6242,N_6324);
or U6637 (N_6637,N_6118,N_6322);
or U6638 (N_6638,N_6159,N_6497);
or U6639 (N_6639,N_6415,N_6125);
and U6640 (N_6640,N_6435,N_6327);
nor U6641 (N_6641,N_6190,N_6450);
or U6642 (N_6642,N_6394,N_6453);
nand U6643 (N_6643,N_6048,N_6413);
nor U6644 (N_6644,N_6289,N_6244);
and U6645 (N_6645,N_6101,N_6010);
nor U6646 (N_6646,N_6191,N_6196);
nand U6647 (N_6647,N_6317,N_6045);
nor U6648 (N_6648,N_6487,N_6340);
or U6649 (N_6649,N_6277,N_6284);
nor U6650 (N_6650,N_6468,N_6131);
and U6651 (N_6651,N_6392,N_6193);
or U6652 (N_6652,N_6379,N_6176);
or U6653 (N_6653,N_6152,N_6199);
or U6654 (N_6654,N_6350,N_6293);
or U6655 (N_6655,N_6162,N_6462);
and U6656 (N_6656,N_6396,N_6358);
nand U6657 (N_6657,N_6002,N_6141);
nand U6658 (N_6658,N_6352,N_6156);
nand U6659 (N_6659,N_6194,N_6294);
xor U6660 (N_6660,N_6319,N_6407);
and U6661 (N_6661,N_6223,N_6224);
or U6662 (N_6662,N_6204,N_6459);
nand U6663 (N_6663,N_6084,N_6467);
nor U6664 (N_6664,N_6099,N_6209);
and U6665 (N_6665,N_6437,N_6299);
nor U6666 (N_6666,N_6296,N_6175);
or U6667 (N_6667,N_6313,N_6017);
or U6668 (N_6668,N_6238,N_6134);
nor U6669 (N_6669,N_6105,N_6461);
nor U6670 (N_6670,N_6032,N_6170);
nor U6671 (N_6671,N_6243,N_6178);
nand U6672 (N_6672,N_6151,N_6354);
xnor U6673 (N_6673,N_6114,N_6393);
or U6674 (N_6674,N_6348,N_6248);
xor U6675 (N_6675,N_6228,N_6349);
nand U6676 (N_6676,N_6006,N_6419);
nand U6677 (N_6677,N_6286,N_6127);
and U6678 (N_6678,N_6021,N_6116);
or U6679 (N_6679,N_6428,N_6038);
and U6680 (N_6680,N_6009,N_6108);
and U6681 (N_6681,N_6485,N_6426);
or U6682 (N_6682,N_6197,N_6404);
or U6683 (N_6683,N_6149,N_6158);
or U6684 (N_6684,N_6267,N_6042);
or U6685 (N_6685,N_6208,N_6442);
or U6686 (N_6686,N_6311,N_6249);
nor U6687 (N_6687,N_6217,N_6057);
or U6688 (N_6688,N_6129,N_6411);
nor U6689 (N_6689,N_6347,N_6451);
or U6690 (N_6690,N_6029,N_6033);
or U6691 (N_6691,N_6093,N_6377);
nand U6692 (N_6692,N_6410,N_6332);
or U6693 (N_6693,N_6030,N_6115);
and U6694 (N_6694,N_6323,N_6090);
xor U6695 (N_6695,N_6016,N_6195);
nor U6696 (N_6696,N_6480,N_6147);
nand U6697 (N_6697,N_6100,N_6472);
nor U6698 (N_6698,N_6051,N_6044);
and U6699 (N_6699,N_6297,N_6083);
and U6700 (N_6700,N_6469,N_6097);
and U6701 (N_6701,N_6315,N_6376);
nor U6702 (N_6702,N_6440,N_6245);
and U6703 (N_6703,N_6441,N_6321);
nor U6704 (N_6704,N_6092,N_6388);
nand U6705 (N_6705,N_6257,N_6298);
or U6706 (N_6706,N_6470,N_6368);
and U6707 (N_6707,N_6256,N_6163);
nand U6708 (N_6708,N_6183,N_6483);
nand U6709 (N_6709,N_6253,N_6001);
nor U6710 (N_6710,N_6104,N_6378);
nand U6711 (N_6711,N_6066,N_6234);
nor U6712 (N_6712,N_6375,N_6406);
and U6713 (N_6713,N_6203,N_6154);
xor U6714 (N_6714,N_6081,N_6270);
and U6715 (N_6715,N_6126,N_6274);
xor U6716 (N_6716,N_6420,N_6303);
and U6717 (N_6717,N_6494,N_6383);
and U6718 (N_6718,N_6380,N_6359);
or U6719 (N_6719,N_6096,N_6421);
nand U6720 (N_6720,N_6145,N_6071);
nor U6721 (N_6721,N_6301,N_6074);
nor U6722 (N_6722,N_6331,N_6446);
nor U6723 (N_6723,N_6474,N_6336);
nand U6724 (N_6724,N_6024,N_6265);
or U6725 (N_6725,N_6229,N_6369);
xnor U6726 (N_6726,N_6318,N_6398);
or U6727 (N_6727,N_6056,N_6260);
and U6728 (N_6728,N_6046,N_6012);
and U6729 (N_6729,N_6385,N_6023);
xnor U6730 (N_6730,N_6167,N_6008);
xor U6731 (N_6731,N_6282,N_6431);
and U6732 (N_6732,N_6341,N_6077);
nand U6733 (N_6733,N_6439,N_6121);
or U6734 (N_6734,N_6258,N_6307);
xor U6735 (N_6735,N_6492,N_6312);
and U6736 (N_6736,N_6119,N_6005);
and U6737 (N_6737,N_6417,N_6279);
nor U6738 (N_6738,N_6160,N_6276);
nor U6739 (N_6739,N_6364,N_6308);
or U6740 (N_6740,N_6189,N_6333);
and U6741 (N_6741,N_6351,N_6268);
nor U6742 (N_6742,N_6438,N_6401);
and U6743 (N_6743,N_6329,N_6087);
nor U6744 (N_6744,N_6373,N_6076);
nor U6745 (N_6745,N_6226,N_6499);
or U6746 (N_6746,N_6463,N_6399);
nor U6747 (N_6747,N_6064,N_6169);
and U6748 (N_6748,N_6095,N_6423);
nor U6749 (N_6749,N_6180,N_6320);
xor U6750 (N_6750,N_6019,N_6180);
nor U6751 (N_6751,N_6351,N_6360);
nand U6752 (N_6752,N_6456,N_6229);
nor U6753 (N_6753,N_6082,N_6329);
nand U6754 (N_6754,N_6174,N_6431);
and U6755 (N_6755,N_6145,N_6478);
or U6756 (N_6756,N_6010,N_6347);
xnor U6757 (N_6757,N_6348,N_6256);
or U6758 (N_6758,N_6100,N_6477);
xor U6759 (N_6759,N_6164,N_6154);
xor U6760 (N_6760,N_6385,N_6216);
xnor U6761 (N_6761,N_6460,N_6001);
and U6762 (N_6762,N_6355,N_6072);
and U6763 (N_6763,N_6300,N_6443);
nand U6764 (N_6764,N_6370,N_6467);
and U6765 (N_6765,N_6234,N_6405);
nand U6766 (N_6766,N_6130,N_6426);
xnor U6767 (N_6767,N_6282,N_6140);
nor U6768 (N_6768,N_6298,N_6397);
nor U6769 (N_6769,N_6469,N_6062);
nand U6770 (N_6770,N_6078,N_6451);
or U6771 (N_6771,N_6452,N_6128);
or U6772 (N_6772,N_6456,N_6079);
nor U6773 (N_6773,N_6045,N_6207);
and U6774 (N_6774,N_6324,N_6215);
and U6775 (N_6775,N_6160,N_6426);
and U6776 (N_6776,N_6110,N_6384);
nand U6777 (N_6777,N_6218,N_6242);
nor U6778 (N_6778,N_6426,N_6184);
nor U6779 (N_6779,N_6075,N_6376);
or U6780 (N_6780,N_6173,N_6460);
nor U6781 (N_6781,N_6410,N_6153);
xnor U6782 (N_6782,N_6298,N_6140);
or U6783 (N_6783,N_6449,N_6465);
or U6784 (N_6784,N_6081,N_6210);
and U6785 (N_6785,N_6399,N_6042);
nand U6786 (N_6786,N_6283,N_6091);
nor U6787 (N_6787,N_6449,N_6251);
nor U6788 (N_6788,N_6472,N_6154);
and U6789 (N_6789,N_6211,N_6273);
nand U6790 (N_6790,N_6013,N_6213);
and U6791 (N_6791,N_6166,N_6200);
nand U6792 (N_6792,N_6379,N_6484);
or U6793 (N_6793,N_6170,N_6082);
and U6794 (N_6794,N_6401,N_6095);
nand U6795 (N_6795,N_6226,N_6209);
nor U6796 (N_6796,N_6424,N_6341);
or U6797 (N_6797,N_6066,N_6284);
or U6798 (N_6798,N_6468,N_6455);
nor U6799 (N_6799,N_6146,N_6249);
nor U6800 (N_6800,N_6422,N_6263);
xor U6801 (N_6801,N_6427,N_6149);
nand U6802 (N_6802,N_6181,N_6482);
nand U6803 (N_6803,N_6019,N_6321);
nand U6804 (N_6804,N_6494,N_6209);
and U6805 (N_6805,N_6324,N_6361);
and U6806 (N_6806,N_6038,N_6085);
nor U6807 (N_6807,N_6000,N_6437);
and U6808 (N_6808,N_6347,N_6376);
or U6809 (N_6809,N_6264,N_6186);
or U6810 (N_6810,N_6298,N_6252);
or U6811 (N_6811,N_6458,N_6017);
or U6812 (N_6812,N_6340,N_6078);
nand U6813 (N_6813,N_6132,N_6340);
nand U6814 (N_6814,N_6163,N_6338);
nand U6815 (N_6815,N_6409,N_6097);
or U6816 (N_6816,N_6215,N_6355);
nor U6817 (N_6817,N_6088,N_6429);
or U6818 (N_6818,N_6409,N_6367);
nand U6819 (N_6819,N_6273,N_6140);
nand U6820 (N_6820,N_6086,N_6481);
nor U6821 (N_6821,N_6280,N_6216);
nor U6822 (N_6822,N_6276,N_6090);
nand U6823 (N_6823,N_6084,N_6334);
nand U6824 (N_6824,N_6446,N_6353);
xnor U6825 (N_6825,N_6164,N_6462);
nor U6826 (N_6826,N_6493,N_6070);
and U6827 (N_6827,N_6467,N_6156);
or U6828 (N_6828,N_6330,N_6132);
and U6829 (N_6829,N_6255,N_6023);
nor U6830 (N_6830,N_6234,N_6431);
nand U6831 (N_6831,N_6131,N_6285);
nand U6832 (N_6832,N_6129,N_6207);
and U6833 (N_6833,N_6181,N_6364);
nand U6834 (N_6834,N_6132,N_6022);
and U6835 (N_6835,N_6109,N_6132);
or U6836 (N_6836,N_6301,N_6231);
nor U6837 (N_6837,N_6199,N_6080);
nand U6838 (N_6838,N_6264,N_6203);
and U6839 (N_6839,N_6366,N_6447);
and U6840 (N_6840,N_6029,N_6048);
or U6841 (N_6841,N_6459,N_6151);
nor U6842 (N_6842,N_6264,N_6204);
and U6843 (N_6843,N_6308,N_6292);
or U6844 (N_6844,N_6065,N_6122);
nor U6845 (N_6845,N_6071,N_6076);
nand U6846 (N_6846,N_6031,N_6244);
xor U6847 (N_6847,N_6146,N_6438);
nor U6848 (N_6848,N_6053,N_6360);
or U6849 (N_6849,N_6455,N_6205);
and U6850 (N_6850,N_6319,N_6443);
and U6851 (N_6851,N_6069,N_6488);
nand U6852 (N_6852,N_6262,N_6080);
and U6853 (N_6853,N_6206,N_6390);
nor U6854 (N_6854,N_6310,N_6424);
nor U6855 (N_6855,N_6247,N_6241);
or U6856 (N_6856,N_6388,N_6059);
nor U6857 (N_6857,N_6215,N_6307);
nor U6858 (N_6858,N_6344,N_6033);
and U6859 (N_6859,N_6246,N_6188);
nor U6860 (N_6860,N_6167,N_6225);
xnor U6861 (N_6861,N_6477,N_6025);
nor U6862 (N_6862,N_6468,N_6405);
and U6863 (N_6863,N_6416,N_6414);
nor U6864 (N_6864,N_6212,N_6296);
nor U6865 (N_6865,N_6027,N_6047);
xnor U6866 (N_6866,N_6339,N_6326);
nor U6867 (N_6867,N_6228,N_6082);
and U6868 (N_6868,N_6416,N_6031);
and U6869 (N_6869,N_6335,N_6492);
or U6870 (N_6870,N_6090,N_6065);
or U6871 (N_6871,N_6102,N_6055);
xnor U6872 (N_6872,N_6456,N_6358);
nand U6873 (N_6873,N_6140,N_6135);
and U6874 (N_6874,N_6060,N_6052);
and U6875 (N_6875,N_6266,N_6236);
and U6876 (N_6876,N_6497,N_6225);
nand U6877 (N_6877,N_6370,N_6360);
or U6878 (N_6878,N_6100,N_6488);
and U6879 (N_6879,N_6497,N_6112);
nand U6880 (N_6880,N_6318,N_6155);
nor U6881 (N_6881,N_6176,N_6305);
and U6882 (N_6882,N_6325,N_6067);
nor U6883 (N_6883,N_6487,N_6125);
and U6884 (N_6884,N_6439,N_6208);
nand U6885 (N_6885,N_6439,N_6219);
nor U6886 (N_6886,N_6219,N_6440);
or U6887 (N_6887,N_6423,N_6280);
nor U6888 (N_6888,N_6277,N_6342);
nand U6889 (N_6889,N_6169,N_6065);
or U6890 (N_6890,N_6136,N_6259);
nor U6891 (N_6891,N_6306,N_6416);
or U6892 (N_6892,N_6213,N_6112);
or U6893 (N_6893,N_6245,N_6468);
or U6894 (N_6894,N_6261,N_6251);
nand U6895 (N_6895,N_6184,N_6135);
nor U6896 (N_6896,N_6113,N_6350);
or U6897 (N_6897,N_6272,N_6277);
nor U6898 (N_6898,N_6166,N_6312);
nand U6899 (N_6899,N_6303,N_6000);
nor U6900 (N_6900,N_6008,N_6116);
nand U6901 (N_6901,N_6436,N_6357);
nor U6902 (N_6902,N_6036,N_6449);
xnor U6903 (N_6903,N_6100,N_6416);
and U6904 (N_6904,N_6440,N_6446);
and U6905 (N_6905,N_6010,N_6451);
nand U6906 (N_6906,N_6111,N_6397);
and U6907 (N_6907,N_6402,N_6103);
nor U6908 (N_6908,N_6166,N_6017);
nor U6909 (N_6909,N_6464,N_6119);
nand U6910 (N_6910,N_6061,N_6209);
xor U6911 (N_6911,N_6083,N_6038);
nand U6912 (N_6912,N_6487,N_6438);
nor U6913 (N_6913,N_6149,N_6245);
xor U6914 (N_6914,N_6006,N_6381);
or U6915 (N_6915,N_6260,N_6127);
nor U6916 (N_6916,N_6354,N_6437);
and U6917 (N_6917,N_6081,N_6310);
nand U6918 (N_6918,N_6283,N_6439);
nor U6919 (N_6919,N_6314,N_6454);
nand U6920 (N_6920,N_6071,N_6420);
and U6921 (N_6921,N_6222,N_6437);
nor U6922 (N_6922,N_6084,N_6135);
nand U6923 (N_6923,N_6440,N_6002);
nand U6924 (N_6924,N_6392,N_6290);
nor U6925 (N_6925,N_6414,N_6437);
nand U6926 (N_6926,N_6399,N_6100);
nand U6927 (N_6927,N_6069,N_6352);
nand U6928 (N_6928,N_6214,N_6357);
nor U6929 (N_6929,N_6246,N_6020);
nand U6930 (N_6930,N_6329,N_6042);
nand U6931 (N_6931,N_6125,N_6489);
nand U6932 (N_6932,N_6196,N_6175);
nor U6933 (N_6933,N_6092,N_6006);
nand U6934 (N_6934,N_6187,N_6017);
nand U6935 (N_6935,N_6161,N_6052);
and U6936 (N_6936,N_6390,N_6130);
nor U6937 (N_6937,N_6226,N_6219);
and U6938 (N_6938,N_6262,N_6448);
and U6939 (N_6939,N_6492,N_6251);
and U6940 (N_6940,N_6291,N_6236);
and U6941 (N_6941,N_6402,N_6399);
nand U6942 (N_6942,N_6372,N_6126);
or U6943 (N_6943,N_6417,N_6232);
and U6944 (N_6944,N_6335,N_6088);
or U6945 (N_6945,N_6347,N_6168);
nand U6946 (N_6946,N_6075,N_6348);
and U6947 (N_6947,N_6386,N_6081);
or U6948 (N_6948,N_6138,N_6437);
nor U6949 (N_6949,N_6049,N_6183);
nor U6950 (N_6950,N_6035,N_6463);
and U6951 (N_6951,N_6434,N_6344);
or U6952 (N_6952,N_6095,N_6218);
xnor U6953 (N_6953,N_6007,N_6408);
or U6954 (N_6954,N_6021,N_6428);
nor U6955 (N_6955,N_6400,N_6093);
and U6956 (N_6956,N_6159,N_6164);
and U6957 (N_6957,N_6345,N_6394);
xnor U6958 (N_6958,N_6421,N_6285);
or U6959 (N_6959,N_6066,N_6020);
nand U6960 (N_6960,N_6258,N_6208);
or U6961 (N_6961,N_6248,N_6015);
and U6962 (N_6962,N_6109,N_6317);
or U6963 (N_6963,N_6098,N_6036);
or U6964 (N_6964,N_6435,N_6476);
nor U6965 (N_6965,N_6351,N_6341);
nand U6966 (N_6966,N_6000,N_6147);
nor U6967 (N_6967,N_6460,N_6312);
and U6968 (N_6968,N_6236,N_6099);
and U6969 (N_6969,N_6085,N_6490);
nand U6970 (N_6970,N_6009,N_6164);
or U6971 (N_6971,N_6259,N_6377);
xor U6972 (N_6972,N_6012,N_6076);
nor U6973 (N_6973,N_6488,N_6016);
nor U6974 (N_6974,N_6035,N_6038);
nor U6975 (N_6975,N_6333,N_6291);
or U6976 (N_6976,N_6125,N_6256);
nand U6977 (N_6977,N_6201,N_6060);
or U6978 (N_6978,N_6279,N_6369);
and U6979 (N_6979,N_6148,N_6190);
nor U6980 (N_6980,N_6146,N_6303);
nand U6981 (N_6981,N_6094,N_6194);
and U6982 (N_6982,N_6181,N_6007);
or U6983 (N_6983,N_6387,N_6023);
xor U6984 (N_6984,N_6069,N_6208);
and U6985 (N_6985,N_6215,N_6182);
and U6986 (N_6986,N_6308,N_6178);
nand U6987 (N_6987,N_6285,N_6494);
and U6988 (N_6988,N_6342,N_6408);
and U6989 (N_6989,N_6371,N_6169);
or U6990 (N_6990,N_6421,N_6023);
nand U6991 (N_6991,N_6319,N_6159);
nor U6992 (N_6992,N_6197,N_6318);
or U6993 (N_6993,N_6162,N_6078);
xnor U6994 (N_6994,N_6129,N_6313);
xor U6995 (N_6995,N_6282,N_6260);
or U6996 (N_6996,N_6268,N_6423);
or U6997 (N_6997,N_6145,N_6448);
or U6998 (N_6998,N_6107,N_6294);
xnor U6999 (N_6999,N_6226,N_6307);
or U7000 (N_7000,N_6786,N_6684);
and U7001 (N_7001,N_6896,N_6781);
nand U7002 (N_7002,N_6898,N_6914);
nor U7003 (N_7003,N_6511,N_6952);
and U7004 (N_7004,N_6856,N_6912);
and U7005 (N_7005,N_6860,N_6531);
or U7006 (N_7006,N_6879,N_6549);
and U7007 (N_7007,N_6576,N_6908);
or U7008 (N_7008,N_6548,N_6866);
nand U7009 (N_7009,N_6774,N_6739);
or U7010 (N_7010,N_6832,N_6975);
and U7011 (N_7011,N_6698,N_6997);
nor U7012 (N_7012,N_6841,N_6513);
nor U7013 (N_7013,N_6568,N_6803);
or U7014 (N_7014,N_6569,N_6710);
or U7015 (N_7015,N_6543,N_6905);
nand U7016 (N_7016,N_6565,N_6536);
xnor U7017 (N_7017,N_6618,N_6572);
nor U7018 (N_7018,N_6923,N_6933);
nand U7019 (N_7019,N_6883,N_6737);
nand U7020 (N_7020,N_6628,N_6944);
nand U7021 (N_7021,N_6849,N_6502);
xor U7022 (N_7022,N_6943,N_6974);
or U7023 (N_7023,N_6953,N_6514);
or U7024 (N_7024,N_6509,N_6740);
or U7025 (N_7025,N_6695,N_6816);
and U7026 (N_7026,N_6960,N_6985);
or U7027 (N_7027,N_6718,N_6983);
nand U7028 (N_7028,N_6515,N_6779);
and U7029 (N_7029,N_6920,N_6998);
nor U7030 (N_7030,N_6916,N_6609);
xnor U7031 (N_7031,N_6909,N_6873);
xor U7032 (N_7032,N_6720,N_6717);
nand U7033 (N_7033,N_6969,N_6527);
or U7034 (N_7034,N_6968,N_6725);
nand U7035 (N_7035,N_6627,N_6506);
nor U7036 (N_7036,N_6801,N_6980);
and U7037 (N_7037,N_6693,N_6654);
nor U7038 (N_7038,N_6673,N_6743);
nor U7039 (N_7039,N_6523,N_6554);
nand U7040 (N_7040,N_6624,N_6656);
nand U7041 (N_7041,N_6604,N_6962);
nand U7042 (N_7042,N_6669,N_6823);
and U7043 (N_7043,N_6868,N_6761);
xor U7044 (N_7044,N_6675,N_6963);
nor U7045 (N_7045,N_6540,N_6731);
or U7046 (N_7046,N_6723,N_6903);
or U7047 (N_7047,N_6704,N_6804);
or U7048 (N_7048,N_6735,N_6713);
nor U7049 (N_7049,N_6680,N_6508);
and U7050 (N_7050,N_6929,N_6537);
nand U7051 (N_7051,N_6907,N_6639);
or U7052 (N_7052,N_6794,N_6505);
nand U7053 (N_7053,N_6844,N_6575);
nand U7054 (N_7054,N_6864,N_6876);
nor U7055 (N_7055,N_6857,N_6555);
or U7056 (N_7056,N_6754,N_6707);
or U7057 (N_7057,N_6696,N_6521);
xnor U7058 (N_7058,N_6899,N_6994);
or U7059 (N_7059,N_6776,N_6783);
xnor U7060 (N_7060,N_6660,N_6677);
or U7061 (N_7061,N_6981,N_6749);
and U7062 (N_7062,N_6799,N_6995);
or U7063 (N_7063,N_6818,N_6588);
or U7064 (N_7064,N_6959,N_6692);
nor U7065 (N_7065,N_6825,N_6989);
and U7066 (N_7066,N_6579,N_6854);
and U7067 (N_7067,N_6798,N_6805);
or U7068 (N_7068,N_6941,N_6577);
nor U7069 (N_7069,N_6758,N_6770);
or U7070 (N_7070,N_6500,N_6766);
xor U7071 (N_7071,N_6910,N_6733);
and U7072 (N_7072,N_6711,N_6587);
xor U7073 (N_7073,N_6842,N_6926);
and U7074 (N_7074,N_6780,N_6788);
nand U7075 (N_7075,N_6890,N_6778);
nor U7076 (N_7076,N_6745,N_6746);
nor U7077 (N_7077,N_6951,N_6824);
and U7078 (N_7078,N_6672,N_6752);
or U7079 (N_7079,N_6571,N_6751);
and U7080 (N_7080,N_6978,N_6626);
xor U7081 (N_7081,N_6875,N_6886);
nor U7082 (N_7082,N_6853,N_6900);
or U7083 (N_7083,N_6881,N_6831);
nor U7084 (N_7084,N_6796,N_6719);
or U7085 (N_7085,N_6690,N_6694);
nor U7086 (N_7086,N_6593,N_6855);
nand U7087 (N_7087,N_6691,N_6889);
or U7088 (N_7088,N_6651,N_6615);
or U7089 (N_7089,N_6556,N_6946);
nand U7090 (N_7090,N_6620,N_6906);
and U7091 (N_7091,N_6802,N_6646);
xnor U7092 (N_7092,N_6728,N_6644);
nor U7093 (N_7093,N_6867,N_6918);
nor U7094 (N_7094,N_6819,N_6773);
or U7095 (N_7095,N_6659,N_6534);
or U7096 (N_7096,N_6822,N_6701);
or U7097 (N_7097,N_6870,N_6837);
xnor U7098 (N_7098,N_6964,N_6605);
or U7099 (N_7099,N_6580,N_6880);
nor U7100 (N_7100,N_6670,N_6629);
or U7101 (N_7101,N_6817,N_6631);
and U7102 (N_7102,N_6750,N_6949);
nor U7103 (N_7103,N_6595,N_6851);
nor U7104 (N_7104,N_6747,N_6991);
and U7105 (N_7105,N_6520,N_6785);
xnor U7106 (N_7106,N_6524,N_6501);
or U7107 (N_7107,N_6538,N_6871);
nand U7108 (N_7108,N_6662,N_6947);
and U7109 (N_7109,N_6700,N_6667);
nand U7110 (N_7110,N_6843,N_6999);
nor U7111 (N_7111,N_6679,N_6760);
xor U7112 (N_7112,N_6955,N_6744);
or U7113 (N_7113,N_6621,N_6793);
nand U7114 (N_7114,N_6563,N_6800);
nand U7115 (N_7115,N_6767,N_6703);
xor U7116 (N_7116,N_6573,N_6858);
nor U7117 (N_7117,N_6863,N_6996);
and U7118 (N_7118,N_6901,N_6708);
and U7119 (N_7119,N_6567,N_6652);
nor U7120 (N_7120,N_6932,N_6558);
or U7121 (N_7121,N_6777,N_6546);
nor U7122 (N_7122,N_6782,N_6967);
or U7123 (N_7123,N_6674,N_6810);
or U7124 (N_7124,N_6834,N_6594);
nand U7125 (N_7125,N_6560,N_6535);
nand U7126 (N_7126,N_6602,N_6736);
nor U7127 (N_7127,N_6795,N_6619);
and U7128 (N_7128,N_6924,N_6552);
nor U7129 (N_7129,N_6665,N_6519);
nand U7130 (N_7130,N_6882,N_6574);
nand U7131 (N_7131,N_6977,N_6623);
nor U7132 (N_7132,N_6525,N_6765);
nand U7133 (N_7133,N_6862,N_6729);
nor U7134 (N_7134,N_6990,N_6657);
nor U7135 (N_7135,N_6714,N_6811);
and U7136 (N_7136,N_6922,N_6820);
xor U7137 (N_7137,N_6861,N_6902);
nor U7138 (N_7138,N_6836,N_6592);
and U7139 (N_7139,N_6727,N_6894);
nand U7140 (N_7140,N_6597,N_6547);
nor U7141 (N_7141,N_6763,N_6610);
and U7142 (N_7142,N_6895,N_6650);
nand U7143 (N_7143,N_6833,N_6529);
or U7144 (N_7144,N_6771,N_6636);
and U7145 (N_7145,N_6869,N_6581);
or U7146 (N_7146,N_6504,N_6539);
nand U7147 (N_7147,N_6884,N_6913);
or U7148 (N_7148,N_6954,N_6755);
or U7149 (N_7149,N_6828,N_6682);
nand U7150 (N_7150,N_6601,N_6958);
and U7151 (N_7151,N_6607,N_6756);
and U7152 (N_7152,N_6848,N_6550);
nor U7153 (N_7153,N_6835,N_6641);
or U7154 (N_7154,N_6784,N_6653);
nand U7155 (N_7155,N_6516,N_6789);
nand U7156 (N_7156,N_6925,N_6937);
nor U7157 (N_7157,N_6561,N_6965);
and U7158 (N_7158,N_6570,N_6812);
or U7159 (N_7159,N_6721,N_6753);
xnor U7160 (N_7160,N_6772,N_6988);
and U7161 (N_7161,N_6510,N_6915);
nor U7162 (N_7162,N_6809,N_6970);
or U7163 (N_7163,N_6808,N_6877);
nor U7164 (N_7164,N_6512,N_6892);
and U7165 (N_7165,N_6613,N_6878);
and U7166 (N_7166,N_6839,N_6530);
or U7167 (N_7167,N_6961,N_6663);
and U7168 (N_7168,N_6813,N_6671);
nand U7169 (N_7169,N_6689,N_6971);
xnor U7170 (N_7170,N_6865,N_6716);
nor U7171 (N_7171,N_6685,N_6688);
nor U7172 (N_7172,N_6526,N_6838);
nor U7173 (N_7173,N_6935,N_6642);
nor U7174 (N_7174,N_6919,N_6706);
nand U7175 (N_7175,N_6874,N_6608);
nand U7176 (N_7176,N_6564,N_6562);
and U7177 (N_7177,N_6829,N_6541);
xor U7178 (N_7178,N_6936,N_6726);
nand U7179 (N_7179,N_6606,N_6806);
nand U7180 (N_7180,N_6775,N_6634);
nand U7181 (N_7181,N_6791,N_6625);
nor U7182 (N_7182,N_6972,N_6840);
xor U7183 (N_7183,N_6846,N_6681);
or U7184 (N_7184,N_6940,N_6887);
or U7185 (N_7185,N_6640,N_6827);
nor U7186 (N_7186,N_6732,N_6709);
or U7187 (N_7187,N_6611,N_6528);
nand U7188 (N_7188,N_6522,N_6950);
and U7189 (N_7189,N_6635,N_6614);
and U7190 (N_7190,N_6589,N_6850);
nor U7191 (N_7191,N_6585,N_6697);
or U7192 (N_7192,N_6648,N_6518);
nand U7193 (N_7193,N_6742,N_6712);
nand U7194 (N_7194,N_6715,N_6655);
nor U7195 (N_7195,N_6661,N_6930);
nand U7196 (N_7196,N_6676,N_6938);
nand U7197 (N_7197,N_6598,N_6591);
or U7198 (N_7198,N_6993,N_6957);
nand U7199 (N_7199,N_6845,N_6814);
and U7200 (N_7200,N_6738,N_6927);
nor U7201 (N_7201,N_6664,N_6699);
nor U7202 (N_7202,N_6643,N_6815);
nor U7203 (N_7203,N_6931,N_6921);
and U7204 (N_7204,N_6559,N_6533);
or U7205 (N_7205,N_6544,N_6645);
nand U7206 (N_7206,N_6852,N_6764);
or U7207 (N_7207,N_6658,N_6934);
and U7208 (N_7208,N_6583,N_6928);
nor U7209 (N_7209,N_6787,N_6622);
xnor U7210 (N_7210,N_6762,N_6939);
and U7211 (N_7211,N_6638,N_6724);
nand U7212 (N_7212,N_6633,N_6807);
nand U7213 (N_7213,N_6722,N_6945);
or U7214 (N_7214,N_6911,N_6668);
and U7215 (N_7215,N_6847,N_6830);
nand U7216 (N_7216,N_6599,N_6956);
and U7217 (N_7217,N_6649,N_6893);
and U7218 (N_7218,N_6942,N_6600);
nor U7219 (N_7219,N_6966,N_6578);
xnor U7220 (N_7220,N_6630,N_6917);
and U7221 (N_7221,N_6557,N_6979);
xnor U7222 (N_7222,N_6617,N_6821);
or U7223 (N_7223,N_6702,N_6590);
and U7224 (N_7224,N_6730,N_6553);
nor U7225 (N_7225,N_6986,N_6705);
nand U7226 (N_7226,N_6686,N_6992);
or U7227 (N_7227,N_6637,N_6741);
or U7228 (N_7228,N_6734,N_6632);
nand U7229 (N_7229,N_6566,N_6987);
nor U7230 (N_7230,N_6872,N_6897);
nand U7231 (N_7231,N_6984,N_6507);
or U7232 (N_7232,N_6666,N_6687);
or U7233 (N_7233,N_6532,N_6888);
xor U7234 (N_7234,N_6582,N_6948);
nand U7235 (N_7235,N_6826,N_6683);
nand U7236 (N_7236,N_6982,N_6757);
nor U7237 (N_7237,N_6973,N_6551);
nor U7238 (N_7238,N_6769,N_6678);
and U7239 (N_7239,N_6647,N_6748);
and U7240 (N_7240,N_6542,N_6596);
or U7241 (N_7241,N_6503,N_6603);
or U7242 (N_7242,N_6790,N_6759);
and U7243 (N_7243,N_6768,N_6586);
nand U7244 (N_7244,N_6976,N_6517);
and U7245 (N_7245,N_6797,N_6885);
nor U7246 (N_7246,N_6792,N_6612);
nor U7247 (N_7247,N_6904,N_6859);
xor U7248 (N_7248,N_6545,N_6616);
nand U7249 (N_7249,N_6584,N_6891);
or U7250 (N_7250,N_6879,N_6900);
nand U7251 (N_7251,N_6953,N_6609);
or U7252 (N_7252,N_6671,N_6577);
and U7253 (N_7253,N_6617,N_6689);
nor U7254 (N_7254,N_6779,N_6911);
and U7255 (N_7255,N_6942,N_6657);
nand U7256 (N_7256,N_6631,N_6971);
nor U7257 (N_7257,N_6699,N_6790);
nand U7258 (N_7258,N_6896,N_6643);
or U7259 (N_7259,N_6585,N_6958);
or U7260 (N_7260,N_6942,N_6646);
or U7261 (N_7261,N_6621,N_6611);
nor U7262 (N_7262,N_6635,N_6548);
xor U7263 (N_7263,N_6571,N_6991);
and U7264 (N_7264,N_6649,N_6673);
nor U7265 (N_7265,N_6549,N_6988);
or U7266 (N_7266,N_6821,N_6941);
xor U7267 (N_7267,N_6927,N_6967);
nor U7268 (N_7268,N_6736,N_6925);
nor U7269 (N_7269,N_6694,N_6983);
xnor U7270 (N_7270,N_6826,N_6737);
xnor U7271 (N_7271,N_6582,N_6805);
nor U7272 (N_7272,N_6529,N_6859);
and U7273 (N_7273,N_6564,N_6965);
nand U7274 (N_7274,N_6729,N_6736);
or U7275 (N_7275,N_6664,N_6971);
and U7276 (N_7276,N_6945,N_6710);
or U7277 (N_7277,N_6741,N_6851);
or U7278 (N_7278,N_6581,N_6854);
or U7279 (N_7279,N_6509,N_6590);
or U7280 (N_7280,N_6675,N_6548);
and U7281 (N_7281,N_6611,N_6531);
xor U7282 (N_7282,N_6603,N_6541);
and U7283 (N_7283,N_6722,N_6666);
and U7284 (N_7284,N_6503,N_6900);
or U7285 (N_7285,N_6653,N_6894);
nor U7286 (N_7286,N_6920,N_6926);
xnor U7287 (N_7287,N_6950,N_6542);
or U7288 (N_7288,N_6540,N_6754);
and U7289 (N_7289,N_6716,N_6717);
or U7290 (N_7290,N_6792,N_6646);
nand U7291 (N_7291,N_6765,N_6670);
nand U7292 (N_7292,N_6800,N_6618);
nor U7293 (N_7293,N_6508,N_6688);
nand U7294 (N_7294,N_6636,N_6850);
or U7295 (N_7295,N_6966,N_6910);
nor U7296 (N_7296,N_6793,N_6875);
nand U7297 (N_7297,N_6919,N_6504);
nand U7298 (N_7298,N_6871,N_6915);
and U7299 (N_7299,N_6870,N_6787);
nand U7300 (N_7300,N_6790,N_6896);
nand U7301 (N_7301,N_6892,N_6668);
nand U7302 (N_7302,N_6922,N_6873);
nand U7303 (N_7303,N_6740,N_6883);
nand U7304 (N_7304,N_6745,N_6693);
xnor U7305 (N_7305,N_6782,N_6800);
or U7306 (N_7306,N_6832,N_6906);
nand U7307 (N_7307,N_6682,N_6788);
nor U7308 (N_7308,N_6538,N_6862);
and U7309 (N_7309,N_6751,N_6794);
nand U7310 (N_7310,N_6710,N_6507);
or U7311 (N_7311,N_6627,N_6976);
or U7312 (N_7312,N_6543,N_6515);
xor U7313 (N_7313,N_6948,N_6697);
nand U7314 (N_7314,N_6944,N_6811);
nor U7315 (N_7315,N_6558,N_6951);
and U7316 (N_7316,N_6502,N_6821);
nor U7317 (N_7317,N_6919,N_6850);
nand U7318 (N_7318,N_6766,N_6822);
nand U7319 (N_7319,N_6735,N_6600);
or U7320 (N_7320,N_6518,N_6692);
or U7321 (N_7321,N_6970,N_6998);
xnor U7322 (N_7322,N_6646,N_6841);
or U7323 (N_7323,N_6986,N_6883);
or U7324 (N_7324,N_6773,N_6947);
or U7325 (N_7325,N_6837,N_6763);
and U7326 (N_7326,N_6519,N_6959);
or U7327 (N_7327,N_6919,N_6869);
and U7328 (N_7328,N_6980,N_6615);
xnor U7329 (N_7329,N_6560,N_6537);
or U7330 (N_7330,N_6732,N_6989);
nand U7331 (N_7331,N_6504,N_6979);
or U7332 (N_7332,N_6734,N_6624);
nor U7333 (N_7333,N_6873,N_6562);
nand U7334 (N_7334,N_6921,N_6674);
xnor U7335 (N_7335,N_6822,N_6618);
and U7336 (N_7336,N_6879,N_6625);
and U7337 (N_7337,N_6995,N_6562);
xnor U7338 (N_7338,N_6650,N_6600);
and U7339 (N_7339,N_6890,N_6867);
nor U7340 (N_7340,N_6608,N_6803);
and U7341 (N_7341,N_6962,N_6923);
nand U7342 (N_7342,N_6845,N_6558);
nand U7343 (N_7343,N_6616,N_6762);
nor U7344 (N_7344,N_6983,N_6993);
or U7345 (N_7345,N_6717,N_6762);
and U7346 (N_7346,N_6740,N_6914);
and U7347 (N_7347,N_6513,N_6921);
nand U7348 (N_7348,N_6872,N_6773);
xor U7349 (N_7349,N_6865,N_6584);
xnor U7350 (N_7350,N_6829,N_6932);
nand U7351 (N_7351,N_6729,N_6896);
xor U7352 (N_7352,N_6893,N_6758);
nor U7353 (N_7353,N_6727,N_6790);
xnor U7354 (N_7354,N_6745,N_6737);
nor U7355 (N_7355,N_6636,N_6960);
or U7356 (N_7356,N_6758,N_6751);
nand U7357 (N_7357,N_6596,N_6840);
xor U7358 (N_7358,N_6810,N_6951);
or U7359 (N_7359,N_6982,N_6748);
and U7360 (N_7360,N_6804,N_6676);
nand U7361 (N_7361,N_6646,N_6662);
nand U7362 (N_7362,N_6832,N_6976);
xor U7363 (N_7363,N_6771,N_6919);
or U7364 (N_7364,N_6939,N_6719);
and U7365 (N_7365,N_6971,N_6947);
xor U7366 (N_7366,N_6534,N_6932);
xnor U7367 (N_7367,N_6805,N_6912);
or U7368 (N_7368,N_6573,N_6707);
nand U7369 (N_7369,N_6681,N_6716);
or U7370 (N_7370,N_6714,N_6536);
nand U7371 (N_7371,N_6835,N_6943);
nand U7372 (N_7372,N_6679,N_6815);
and U7373 (N_7373,N_6520,N_6897);
xnor U7374 (N_7374,N_6778,N_6599);
xnor U7375 (N_7375,N_6637,N_6946);
and U7376 (N_7376,N_6994,N_6787);
nand U7377 (N_7377,N_6828,N_6560);
nor U7378 (N_7378,N_6794,N_6922);
or U7379 (N_7379,N_6723,N_6868);
nor U7380 (N_7380,N_6925,N_6773);
and U7381 (N_7381,N_6992,N_6601);
xor U7382 (N_7382,N_6771,N_6606);
xor U7383 (N_7383,N_6505,N_6924);
and U7384 (N_7384,N_6613,N_6681);
nand U7385 (N_7385,N_6992,N_6699);
nor U7386 (N_7386,N_6917,N_6659);
nand U7387 (N_7387,N_6936,N_6760);
and U7388 (N_7388,N_6767,N_6771);
and U7389 (N_7389,N_6617,N_6563);
and U7390 (N_7390,N_6576,N_6560);
and U7391 (N_7391,N_6710,N_6834);
or U7392 (N_7392,N_6576,N_6886);
or U7393 (N_7393,N_6510,N_6523);
xnor U7394 (N_7394,N_6600,N_6536);
or U7395 (N_7395,N_6616,N_6700);
or U7396 (N_7396,N_6709,N_6555);
and U7397 (N_7397,N_6775,N_6531);
nor U7398 (N_7398,N_6535,N_6779);
or U7399 (N_7399,N_6726,N_6583);
nand U7400 (N_7400,N_6750,N_6612);
and U7401 (N_7401,N_6574,N_6825);
nor U7402 (N_7402,N_6999,N_6816);
nand U7403 (N_7403,N_6951,N_6814);
or U7404 (N_7404,N_6551,N_6629);
xnor U7405 (N_7405,N_6867,N_6572);
and U7406 (N_7406,N_6976,N_6746);
nor U7407 (N_7407,N_6644,N_6539);
xnor U7408 (N_7408,N_6994,N_6608);
and U7409 (N_7409,N_6902,N_6609);
xor U7410 (N_7410,N_6950,N_6786);
nor U7411 (N_7411,N_6936,N_6589);
nor U7412 (N_7412,N_6559,N_6963);
and U7413 (N_7413,N_6627,N_6805);
or U7414 (N_7414,N_6639,N_6851);
nand U7415 (N_7415,N_6867,N_6718);
and U7416 (N_7416,N_6560,N_6778);
or U7417 (N_7417,N_6543,N_6983);
nand U7418 (N_7418,N_6660,N_6647);
nand U7419 (N_7419,N_6835,N_6968);
nand U7420 (N_7420,N_6966,N_6517);
nand U7421 (N_7421,N_6770,N_6546);
nand U7422 (N_7422,N_6897,N_6870);
nor U7423 (N_7423,N_6507,N_6773);
nor U7424 (N_7424,N_6980,N_6905);
nor U7425 (N_7425,N_6867,N_6632);
nor U7426 (N_7426,N_6597,N_6958);
xor U7427 (N_7427,N_6500,N_6626);
or U7428 (N_7428,N_6600,N_6520);
or U7429 (N_7429,N_6725,N_6973);
nor U7430 (N_7430,N_6684,N_6733);
or U7431 (N_7431,N_6794,N_6799);
xnor U7432 (N_7432,N_6953,N_6636);
nand U7433 (N_7433,N_6642,N_6848);
nor U7434 (N_7434,N_6643,N_6917);
or U7435 (N_7435,N_6596,N_6746);
or U7436 (N_7436,N_6982,N_6834);
or U7437 (N_7437,N_6714,N_6668);
nand U7438 (N_7438,N_6772,N_6887);
and U7439 (N_7439,N_6941,N_6894);
nand U7440 (N_7440,N_6995,N_6956);
nor U7441 (N_7441,N_6525,N_6740);
xnor U7442 (N_7442,N_6695,N_6500);
and U7443 (N_7443,N_6831,N_6670);
or U7444 (N_7444,N_6880,N_6885);
or U7445 (N_7445,N_6563,N_6770);
nand U7446 (N_7446,N_6680,N_6685);
nor U7447 (N_7447,N_6750,N_6516);
nand U7448 (N_7448,N_6774,N_6834);
or U7449 (N_7449,N_6537,N_6888);
nand U7450 (N_7450,N_6976,N_6507);
xnor U7451 (N_7451,N_6903,N_6522);
and U7452 (N_7452,N_6754,N_6614);
nor U7453 (N_7453,N_6833,N_6568);
or U7454 (N_7454,N_6890,N_6632);
and U7455 (N_7455,N_6709,N_6567);
nand U7456 (N_7456,N_6905,N_6799);
nand U7457 (N_7457,N_6700,N_6998);
nand U7458 (N_7458,N_6826,N_6745);
or U7459 (N_7459,N_6524,N_6588);
nand U7460 (N_7460,N_6514,N_6976);
nor U7461 (N_7461,N_6967,N_6848);
and U7462 (N_7462,N_6902,N_6907);
nand U7463 (N_7463,N_6935,N_6552);
xor U7464 (N_7464,N_6617,N_6567);
or U7465 (N_7465,N_6533,N_6554);
and U7466 (N_7466,N_6730,N_6505);
or U7467 (N_7467,N_6606,N_6820);
nor U7468 (N_7468,N_6848,N_6769);
or U7469 (N_7469,N_6947,N_6711);
nand U7470 (N_7470,N_6583,N_6546);
and U7471 (N_7471,N_6968,N_6786);
nand U7472 (N_7472,N_6760,N_6651);
xor U7473 (N_7473,N_6647,N_6537);
and U7474 (N_7474,N_6681,N_6855);
and U7475 (N_7475,N_6852,N_6883);
nand U7476 (N_7476,N_6592,N_6556);
or U7477 (N_7477,N_6863,N_6604);
nor U7478 (N_7478,N_6660,N_6612);
nand U7479 (N_7479,N_6826,N_6700);
or U7480 (N_7480,N_6761,N_6692);
or U7481 (N_7481,N_6866,N_6847);
nand U7482 (N_7482,N_6637,N_6688);
nand U7483 (N_7483,N_6668,N_6588);
nor U7484 (N_7484,N_6994,N_6594);
nor U7485 (N_7485,N_6621,N_6852);
nor U7486 (N_7486,N_6909,N_6915);
or U7487 (N_7487,N_6830,N_6675);
nor U7488 (N_7488,N_6874,N_6970);
xnor U7489 (N_7489,N_6849,N_6529);
and U7490 (N_7490,N_6861,N_6864);
nor U7491 (N_7491,N_6771,N_6790);
nand U7492 (N_7492,N_6952,N_6710);
or U7493 (N_7493,N_6853,N_6759);
nand U7494 (N_7494,N_6549,N_6857);
xor U7495 (N_7495,N_6514,N_6989);
nand U7496 (N_7496,N_6765,N_6551);
nor U7497 (N_7497,N_6673,N_6637);
or U7498 (N_7498,N_6601,N_6971);
xnor U7499 (N_7499,N_6763,N_6645);
and U7500 (N_7500,N_7374,N_7403);
nor U7501 (N_7501,N_7058,N_7410);
or U7502 (N_7502,N_7172,N_7224);
nor U7503 (N_7503,N_7479,N_7472);
nand U7504 (N_7504,N_7034,N_7400);
nor U7505 (N_7505,N_7320,N_7312);
or U7506 (N_7506,N_7071,N_7061);
and U7507 (N_7507,N_7168,N_7185);
nor U7508 (N_7508,N_7226,N_7268);
nand U7509 (N_7509,N_7392,N_7029);
nor U7510 (N_7510,N_7093,N_7489);
nand U7511 (N_7511,N_7076,N_7349);
or U7512 (N_7512,N_7255,N_7084);
nand U7513 (N_7513,N_7330,N_7345);
nand U7514 (N_7514,N_7462,N_7324);
and U7515 (N_7515,N_7144,N_7298);
or U7516 (N_7516,N_7015,N_7316);
and U7517 (N_7517,N_7340,N_7087);
nor U7518 (N_7518,N_7492,N_7277);
nand U7519 (N_7519,N_7220,N_7456);
nand U7520 (N_7520,N_7395,N_7066);
and U7521 (N_7521,N_7122,N_7287);
nand U7522 (N_7522,N_7259,N_7473);
or U7523 (N_7523,N_7482,N_7008);
nor U7524 (N_7524,N_7191,N_7091);
or U7525 (N_7525,N_7496,N_7202);
nand U7526 (N_7526,N_7193,N_7411);
nor U7527 (N_7527,N_7329,N_7267);
xnor U7528 (N_7528,N_7003,N_7274);
nand U7529 (N_7529,N_7326,N_7189);
nor U7530 (N_7530,N_7219,N_7363);
and U7531 (N_7531,N_7052,N_7152);
or U7532 (N_7532,N_7205,N_7444);
or U7533 (N_7533,N_7151,N_7460);
or U7534 (N_7534,N_7421,N_7368);
nor U7535 (N_7535,N_7306,N_7317);
nand U7536 (N_7536,N_7105,N_7040);
and U7537 (N_7537,N_7389,N_7470);
nor U7538 (N_7538,N_7433,N_7141);
xor U7539 (N_7539,N_7090,N_7399);
nor U7540 (N_7540,N_7404,N_7490);
xor U7541 (N_7541,N_7384,N_7390);
nor U7542 (N_7542,N_7092,N_7406);
nor U7543 (N_7543,N_7007,N_7212);
nor U7544 (N_7544,N_7222,N_7116);
or U7545 (N_7545,N_7258,N_7109);
and U7546 (N_7546,N_7165,N_7254);
and U7547 (N_7547,N_7211,N_7332);
and U7548 (N_7548,N_7104,N_7325);
and U7549 (N_7549,N_7438,N_7037);
and U7550 (N_7550,N_7278,N_7292);
or U7551 (N_7551,N_7108,N_7497);
or U7552 (N_7552,N_7049,N_7327);
xnor U7553 (N_7553,N_7286,N_7159);
nor U7554 (N_7554,N_7471,N_7130);
nand U7555 (N_7555,N_7143,N_7239);
or U7556 (N_7556,N_7214,N_7230);
nand U7557 (N_7557,N_7055,N_7194);
nor U7558 (N_7558,N_7081,N_7088);
or U7559 (N_7559,N_7469,N_7441);
nor U7560 (N_7560,N_7132,N_7361);
or U7561 (N_7561,N_7458,N_7256);
or U7562 (N_7562,N_7266,N_7017);
and U7563 (N_7563,N_7373,N_7032);
or U7564 (N_7564,N_7459,N_7260);
xnor U7565 (N_7565,N_7275,N_7199);
nand U7566 (N_7566,N_7112,N_7311);
or U7567 (N_7567,N_7270,N_7367);
xnor U7568 (N_7568,N_7225,N_7026);
or U7569 (N_7569,N_7234,N_7059);
nor U7570 (N_7570,N_7269,N_7209);
nand U7571 (N_7571,N_7377,N_7171);
nor U7572 (N_7572,N_7419,N_7414);
and U7573 (N_7573,N_7195,N_7436);
and U7574 (N_7574,N_7494,N_7321);
nor U7575 (N_7575,N_7023,N_7429);
nand U7576 (N_7576,N_7481,N_7253);
nand U7577 (N_7577,N_7094,N_7356);
and U7578 (N_7578,N_7177,N_7315);
nand U7579 (N_7579,N_7158,N_7028);
and U7580 (N_7580,N_7449,N_7282);
or U7581 (N_7581,N_7001,N_7378);
nor U7582 (N_7582,N_7068,N_7393);
nand U7583 (N_7583,N_7382,N_7450);
or U7584 (N_7584,N_7498,N_7475);
nand U7585 (N_7585,N_7207,N_7319);
nor U7586 (N_7586,N_7430,N_7206);
and U7587 (N_7587,N_7110,N_7290);
nand U7588 (N_7588,N_7417,N_7022);
or U7589 (N_7589,N_7050,N_7103);
or U7590 (N_7590,N_7153,N_7499);
or U7591 (N_7591,N_7121,N_7183);
and U7592 (N_7592,N_7204,N_7346);
or U7593 (N_7593,N_7101,N_7294);
nor U7594 (N_7594,N_7082,N_7301);
nor U7595 (N_7595,N_7333,N_7237);
or U7596 (N_7596,N_7263,N_7228);
or U7597 (N_7597,N_7054,N_7048);
or U7598 (N_7598,N_7432,N_7412);
and U7599 (N_7599,N_7283,N_7273);
nand U7600 (N_7600,N_7435,N_7407);
and U7601 (N_7601,N_7145,N_7201);
nor U7602 (N_7602,N_7147,N_7218);
and U7603 (N_7603,N_7437,N_7047);
and U7604 (N_7604,N_7451,N_7369);
nor U7605 (N_7605,N_7344,N_7073);
nor U7606 (N_7606,N_7339,N_7215);
nand U7607 (N_7607,N_7394,N_7370);
and U7608 (N_7608,N_7100,N_7495);
nor U7609 (N_7609,N_7457,N_7196);
or U7610 (N_7610,N_7466,N_7004);
nor U7611 (N_7611,N_7396,N_7120);
nand U7612 (N_7612,N_7376,N_7186);
nor U7613 (N_7613,N_7129,N_7099);
nand U7614 (N_7614,N_7272,N_7416);
or U7615 (N_7615,N_7408,N_7210);
xor U7616 (N_7616,N_7453,N_7123);
xnor U7617 (N_7617,N_7271,N_7423);
xnor U7618 (N_7618,N_7284,N_7425);
xor U7619 (N_7619,N_7231,N_7448);
and U7620 (N_7620,N_7262,N_7309);
and U7621 (N_7621,N_7197,N_7227);
xor U7622 (N_7622,N_7030,N_7488);
nand U7623 (N_7623,N_7013,N_7166);
or U7624 (N_7624,N_7486,N_7308);
nor U7625 (N_7625,N_7304,N_7035);
and U7626 (N_7626,N_7223,N_7245);
or U7627 (N_7627,N_7086,N_7235);
and U7628 (N_7628,N_7178,N_7322);
nor U7629 (N_7629,N_7420,N_7305);
and U7630 (N_7630,N_7426,N_7401);
xor U7631 (N_7631,N_7276,N_7351);
nand U7632 (N_7632,N_7163,N_7043);
or U7633 (N_7633,N_7440,N_7280);
nor U7634 (N_7634,N_7203,N_7478);
nor U7635 (N_7635,N_7251,N_7247);
or U7636 (N_7636,N_7250,N_7075);
and U7637 (N_7637,N_7042,N_7175);
nand U7638 (N_7638,N_7372,N_7447);
xor U7639 (N_7639,N_7160,N_7338);
and U7640 (N_7640,N_7487,N_7257);
or U7641 (N_7641,N_7057,N_7386);
xor U7642 (N_7642,N_7138,N_7474);
or U7643 (N_7643,N_7480,N_7118);
xnor U7644 (N_7644,N_7036,N_7375);
and U7645 (N_7645,N_7167,N_7485);
or U7646 (N_7646,N_7463,N_7115);
nand U7647 (N_7647,N_7455,N_7261);
and U7648 (N_7648,N_7221,N_7302);
nand U7649 (N_7649,N_7025,N_7174);
nand U7650 (N_7650,N_7347,N_7011);
nand U7651 (N_7651,N_7300,N_7134);
nor U7652 (N_7652,N_7442,N_7019);
nor U7653 (N_7653,N_7187,N_7006);
nand U7654 (N_7654,N_7359,N_7288);
nand U7655 (N_7655,N_7446,N_7249);
and U7656 (N_7656,N_7111,N_7184);
xnor U7657 (N_7657,N_7461,N_7065);
and U7658 (N_7658,N_7358,N_7079);
and U7659 (N_7659,N_7080,N_7014);
xnor U7660 (N_7660,N_7364,N_7281);
nor U7661 (N_7661,N_7360,N_7044);
nor U7662 (N_7662,N_7181,N_7062);
xor U7663 (N_7663,N_7162,N_7337);
and U7664 (N_7664,N_7096,N_7126);
and U7665 (N_7665,N_7016,N_7136);
or U7666 (N_7666,N_7354,N_7310);
nor U7667 (N_7667,N_7379,N_7169);
or U7668 (N_7668,N_7000,N_7216);
nand U7669 (N_7669,N_7350,N_7341);
or U7670 (N_7670,N_7434,N_7119);
xor U7671 (N_7671,N_7009,N_7156);
or U7672 (N_7672,N_7279,N_7095);
nor U7673 (N_7673,N_7038,N_7385);
and U7674 (N_7674,N_7137,N_7074);
nor U7675 (N_7675,N_7297,N_7021);
xnor U7676 (N_7676,N_7039,N_7056);
or U7677 (N_7677,N_7125,N_7484);
or U7678 (N_7678,N_7452,N_7493);
or U7679 (N_7679,N_7102,N_7217);
nor U7680 (N_7680,N_7142,N_7293);
or U7681 (N_7681,N_7117,N_7180);
nand U7682 (N_7682,N_7176,N_7366);
and U7683 (N_7683,N_7238,N_7069);
nand U7684 (N_7684,N_7198,N_7097);
and U7685 (N_7685,N_7033,N_7133);
and U7686 (N_7686,N_7307,N_7241);
and U7687 (N_7687,N_7467,N_7380);
and U7688 (N_7688,N_7208,N_7296);
or U7689 (N_7689,N_7422,N_7173);
nor U7690 (N_7690,N_7246,N_7018);
nand U7691 (N_7691,N_7465,N_7140);
nor U7692 (N_7692,N_7342,N_7365);
and U7693 (N_7693,N_7010,N_7331);
and U7694 (N_7694,N_7264,N_7343);
nor U7695 (N_7695,N_7314,N_7031);
nor U7696 (N_7696,N_7170,N_7157);
and U7697 (N_7697,N_7439,N_7213);
nand U7698 (N_7698,N_7418,N_7128);
nand U7699 (N_7699,N_7295,N_7371);
or U7700 (N_7700,N_7402,N_7085);
and U7701 (N_7701,N_7318,N_7002);
nor U7702 (N_7702,N_7483,N_7313);
nor U7703 (N_7703,N_7353,N_7024);
and U7704 (N_7704,N_7053,N_7188);
and U7705 (N_7705,N_7233,N_7182);
nand U7706 (N_7706,N_7005,N_7362);
or U7707 (N_7707,N_7192,N_7107);
nor U7708 (N_7708,N_7424,N_7323);
xor U7709 (N_7709,N_7291,N_7243);
nor U7710 (N_7710,N_7491,N_7355);
nor U7711 (N_7711,N_7063,N_7135);
nand U7712 (N_7712,N_7381,N_7303);
and U7713 (N_7713,N_7078,N_7200);
and U7714 (N_7714,N_7072,N_7299);
nand U7715 (N_7715,N_7445,N_7012);
and U7716 (N_7716,N_7265,N_7443);
nor U7717 (N_7717,N_7248,N_7106);
or U7718 (N_7718,N_7336,N_7348);
and U7719 (N_7719,N_7020,N_7244);
and U7720 (N_7720,N_7391,N_7113);
or U7721 (N_7721,N_7164,N_7179);
nand U7722 (N_7722,N_7229,N_7027);
xor U7723 (N_7723,N_7328,N_7150);
nor U7724 (N_7724,N_7252,N_7352);
xnor U7725 (N_7725,N_7335,N_7131);
nor U7726 (N_7726,N_7387,N_7454);
and U7727 (N_7727,N_7190,N_7236);
nor U7728 (N_7728,N_7041,N_7139);
xnor U7729 (N_7729,N_7146,N_7415);
nor U7730 (N_7730,N_7114,N_7161);
nand U7731 (N_7731,N_7240,N_7070);
and U7732 (N_7732,N_7334,N_7127);
and U7733 (N_7733,N_7383,N_7155);
xor U7734 (N_7734,N_7398,N_7148);
nor U7735 (N_7735,N_7285,N_7427);
and U7736 (N_7736,N_7397,N_7083);
nor U7737 (N_7737,N_7405,N_7289);
or U7738 (N_7738,N_7067,N_7089);
and U7739 (N_7739,N_7154,N_7232);
nor U7740 (N_7740,N_7413,N_7124);
nor U7741 (N_7741,N_7046,N_7468);
nor U7742 (N_7742,N_7064,N_7357);
nor U7743 (N_7743,N_7476,N_7477);
and U7744 (N_7744,N_7428,N_7388);
and U7745 (N_7745,N_7051,N_7045);
nor U7746 (N_7746,N_7242,N_7060);
nand U7747 (N_7747,N_7431,N_7464);
or U7748 (N_7748,N_7409,N_7149);
nor U7749 (N_7749,N_7077,N_7098);
nand U7750 (N_7750,N_7103,N_7106);
xor U7751 (N_7751,N_7251,N_7420);
or U7752 (N_7752,N_7134,N_7164);
and U7753 (N_7753,N_7129,N_7056);
or U7754 (N_7754,N_7374,N_7318);
or U7755 (N_7755,N_7240,N_7106);
nor U7756 (N_7756,N_7130,N_7346);
nor U7757 (N_7757,N_7011,N_7466);
and U7758 (N_7758,N_7062,N_7213);
nand U7759 (N_7759,N_7300,N_7218);
and U7760 (N_7760,N_7328,N_7368);
or U7761 (N_7761,N_7107,N_7098);
and U7762 (N_7762,N_7024,N_7167);
nor U7763 (N_7763,N_7487,N_7433);
and U7764 (N_7764,N_7120,N_7150);
nand U7765 (N_7765,N_7292,N_7395);
and U7766 (N_7766,N_7021,N_7060);
or U7767 (N_7767,N_7270,N_7165);
nand U7768 (N_7768,N_7045,N_7353);
or U7769 (N_7769,N_7233,N_7154);
and U7770 (N_7770,N_7159,N_7368);
and U7771 (N_7771,N_7469,N_7433);
and U7772 (N_7772,N_7274,N_7448);
nand U7773 (N_7773,N_7020,N_7120);
nand U7774 (N_7774,N_7199,N_7136);
xnor U7775 (N_7775,N_7059,N_7020);
or U7776 (N_7776,N_7176,N_7222);
and U7777 (N_7777,N_7365,N_7277);
or U7778 (N_7778,N_7272,N_7372);
nand U7779 (N_7779,N_7108,N_7237);
and U7780 (N_7780,N_7470,N_7319);
nand U7781 (N_7781,N_7047,N_7424);
nand U7782 (N_7782,N_7087,N_7372);
xor U7783 (N_7783,N_7313,N_7324);
or U7784 (N_7784,N_7404,N_7385);
nand U7785 (N_7785,N_7029,N_7326);
or U7786 (N_7786,N_7260,N_7041);
nand U7787 (N_7787,N_7409,N_7118);
or U7788 (N_7788,N_7253,N_7413);
and U7789 (N_7789,N_7412,N_7068);
nand U7790 (N_7790,N_7262,N_7107);
nor U7791 (N_7791,N_7189,N_7376);
and U7792 (N_7792,N_7448,N_7222);
or U7793 (N_7793,N_7097,N_7076);
or U7794 (N_7794,N_7496,N_7043);
nor U7795 (N_7795,N_7334,N_7363);
nand U7796 (N_7796,N_7485,N_7131);
xnor U7797 (N_7797,N_7451,N_7109);
nand U7798 (N_7798,N_7000,N_7201);
or U7799 (N_7799,N_7137,N_7376);
and U7800 (N_7800,N_7245,N_7438);
and U7801 (N_7801,N_7039,N_7199);
nor U7802 (N_7802,N_7420,N_7073);
nor U7803 (N_7803,N_7217,N_7203);
and U7804 (N_7804,N_7010,N_7202);
nor U7805 (N_7805,N_7446,N_7200);
and U7806 (N_7806,N_7419,N_7373);
or U7807 (N_7807,N_7187,N_7331);
nand U7808 (N_7808,N_7327,N_7129);
and U7809 (N_7809,N_7183,N_7453);
or U7810 (N_7810,N_7429,N_7370);
or U7811 (N_7811,N_7499,N_7049);
nand U7812 (N_7812,N_7310,N_7409);
xnor U7813 (N_7813,N_7139,N_7276);
nor U7814 (N_7814,N_7356,N_7498);
xnor U7815 (N_7815,N_7325,N_7445);
or U7816 (N_7816,N_7282,N_7004);
and U7817 (N_7817,N_7411,N_7423);
or U7818 (N_7818,N_7242,N_7433);
and U7819 (N_7819,N_7462,N_7059);
nor U7820 (N_7820,N_7315,N_7033);
nand U7821 (N_7821,N_7355,N_7297);
nor U7822 (N_7822,N_7428,N_7384);
nor U7823 (N_7823,N_7105,N_7167);
xor U7824 (N_7824,N_7203,N_7364);
nor U7825 (N_7825,N_7006,N_7149);
or U7826 (N_7826,N_7373,N_7043);
and U7827 (N_7827,N_7094,N_7048);
nand U7828 (N_7828,N_7393,N_7016);
or U7829 (N_7829,N_7225,N_7128);
or U7830 (N_7830,N_7488,N_7199);
nand U7831 (N_7831,N_7343,N_7359);
nand U7832 (N_7832,N_7147,N_7099);
nand U7833 (N_7833,N_7122,N_7488);
nor U7834 (N_7834,N_7295,N_7474);
nand U7835 (N_7835,N_7257,N_7049);
xor U7836 (N_7836,N_7386,N_7479);
and U7837 (N_7837,N_7223,N_7450);
nand U7838 (N_7838,N_7190,N_7201);
nand U7839 (N_7839,N_7341,N_7119);
or U7840 (N_7840,N_7309,N_7412);
nand U7841 (N_7841,N_7329,N_7010);
nor U7842 (N_7842,N_7391,N_7154);
and U7843 (N_7843,N_7065,N_7085);
nand U7844 (N_7844,N_7200,N_7240);
nor U7845 (N_7845,N_7333,N_7293);
or U7846 (N_7846,N_7131,N_7319);
or U7847 (N_7847,N_7005,N_7231);
or U7848 (N_7848,N_7023,N_7240);
nand U7849 (N_7849,N_7273,N_7480);
or U7850 (N_7850,N_7324,N_7416);
nor U7851 (N_7851,N_7497,N_7338);
nand U7852 (N_7852,N_7253,N_7073);
nor U7853 (N_7853,N_7285,N_7268);
nand U7854 (N_7854,N_7132,N_7021);
or U7855 (N_7855,N_7135,N_7341);
nand U7856 (N_7856,N_7440,N_7433);
or U7857 (N_7857,N_7126,N_7055);
xnor U7858 (N_7858,N_7219,N_7357);
and U7859 (N_7859,N_7151,N_7173);
nor U7860 (N_7860,N_7047,N_7321);
nor U7861 (N_7861,N_7223,N_7168);
nand U7862 (N_7862,N_7138,N_7036);
or U7863 (N_7863,N_7398,N_7063);
xor U7864 (N_7864,N_7147,N_7375);
nand U7865 (N_7865,N_7209,N_7338);
xnor U7866 (N_7866,N_7095,N_7427);
nor U7867 (N_7867,N_7463,N_7338);
nand U7868 (N_7868,N_7497,N_7491);
nand U7869 (N_7869,N_7020,N_7384);
nor U7870 (N_7870,N_7051,N_7010);
and U7871 (N_7871,N_7421,N_7135);
xnor U7872 (N_7872,N_7453,N_7320);
nand U7873 (N_7873,N_7186,N_7432);
nand U7874 (N_7874,N_7463,N_7034);
or U7875 (N_7875,N_7054,N_7128);
nor U7876 (N_7876,N_7074,N_7395);
nand U7877 (N_7877,N_7348,N_7176);
and U7878 (N_7878,N_7154,N_7177);
xor U7879 (N_7879,N_7024,N_7359);
nand U7880 (N_7880,N_7051,N_7232);
nor U7881 (N_7881,N_7322,N_7130);
nor U7882 (N_7882,N_7475,N_7441);
nand U7883 (N_7883,N_7281,N_7292);
nand U7884 (N_7884,N_7313,N_7163);
and U7885 (N_7885,N_7093,N_7438);
xor U7886 (N_7886,N_7223,N_7070);
or U7887 (N_7887,N_7302,N_7014);
or U7888 (N_7888,N_7190,N_7276);
nand U7889 (N_7889,N_7123,N_7214);
and U7890 (N_7890,N_7284,N_7450);
or U7891 (N_7891,N_7143,N_7096);
nand U7892 (N_7892,N_7289,N_7211);
nor U7893 (N_7893,N_7372,N_7340);
nor U7894 (N_7894,N_7436,N_7096);
or U7895 (N_7895,N_7005,N_7207);
nand U7896 (N_7896,N_7484,N_7384);
and U7897 (N_7897,N_7472,N_7169);
nand U7898 (N_7898,N_7160,N_7269);
nor U7899 (N_7899,N_7333,N_7048);
or U7900 (N_7900,N_7366,N_7409);
or U7901 (N_7901,N_7157,N_7021);
nand U7902 (N_7902,N_7014,N_7083);
nand U7903 (N_7903,N_7333,N_7112);
nor U7904 (N_7904,N_7311,N_7192);
or U7905 (N_7905,N_7221,N_7315);
and U7906 (N_7906,N_7465,N_7435);
or U7907 (N_7907,N_7276,N_7164);
nor U7908 (N_7908,N_7331,N_7247);
and U7909 (N_7909,N_7060,N_7286);
xnor U7910 (N_7910,N_7052,N_7407);
nor U7911 (N_7911,N_7035,N_7479);
and U7912 (N_7912,N_7078,N_7383);
and U7913 (N_7913,N_7463,N_7152);
and U7914 (N_7914,N_7211,N_7392);
or U7915 (N_7915,N_7485,N_7302);
and U7916 (N_7916,N_7386,N_7155);
xor U7917 (N_7917,N_7477,N_7277);
and U7918 (N_7918,N_7102,N_7353);
and U7919 (N_7919,N_7474,N_7013);
or U7920 (N_7920,N_7101,N_7271);
nand U7921 (N_7921,N_7459,N_7208);
nor U7922 (N_7922,N_7020,N_7052);
nand U7923 (N_7923,N_7337,N_7422);
nand U7924 (N_7924,N_7021,N_7472);
or U7925 (N_7925,N_7397,N_7106);
nor U7926 (N_7926,N_7165,N_7256);
nand U7927 (N_7927,N_7492,N_7464);
nand U7928 (N_7928,N_7379,N_7142);
and U7929 (N_7929,N_7386,N_7248);
nor U7930 (N_7930,N_7463,N_7465);
xnor U7931 (N_7931,N_7155,N_7019);
and U7932 (N_7932,N_7052,N_7468);
and U7933 (N_7933,N_7178,N_7245);
or U7934 (N_7934,N_7079,N_7454);
nand U7935 (N_7935,N_7305,N_7243);
nor U7936 (N_7936,N_7342,N_7489);
nand U7937 (N_7937,N_7099,N_7181);
or U7938 (N_7938,N_7073,N_7410);
or U7939 (N_7939,N_7294,N_7398);
nor U7940 (N_7940,N_7431,N_7191);
nand U7941 (N_7941,N_7265,N_7382);
nand U7942 (N_7942,N_7024,N_7110);
nor U7943 (N_7943,N_7168,N_7267);
nor U7944 (N_7944,N_7097,N_7430);
or U7945 (N_7945,N_7100,N_7050);
or U7946 (N_7946,N_7360,N_7350);
nand U7947 (N_7947,N_7094,N_7438);
nor U7948 (N_7948,N_7211,N_7069);
nor U7949 (N_7949,N_7314,N_7398);
and U7950 (N_7950,N_7095,N_7391);
nand U7951 (N_7951,N_7238,N_7191);
xnor U7952 (N_7952,N_7394,N_7307);
or U7953 (N_7953,N_7485,N_7276);
xor U7954 (N_7954,N_7435,N_7401);
nor U7955 (N_7955,N_7439,N_7207);
or U7956 (N_7956,N_7122,N_7162);
or U7957 (N_7957,N_7282,N_7337);
and U7958 (N_7958,N_7377,N_7336);
nor U7959 (N_7959,N_7107,N_7498);
or U7960 (N_7960,N_7173,N_7161);
or U7961 (N_7961,N_7327,N_7387);
nor U7962 (N_7962,N_7104,N_7298);
xnor U7963 (N_7963,N_7082,N_7486);
nand U7964 (N_7964,N_7027,N_7151);
xnor U7965 (N_7965,N_7140,N_7131);
or U7966 (N_7966,N_7082,N_7126);
and U7967 (N_7967,N_7344,N_7047);
and U7968 (N_7968,N_7226,N_7032);
and U7969 (N_7969,N_7300,N_7237);
and U7970 (N_7970,N_7236,N_7288);
nand U7971 (N_7971,N_7336,N_7071);
nor U7972 (N_7972,N_7063,N_7029);
nor U7973 (N_7973,N_7038,N_7080);
nor U7974 (N_7974,N_7423,N_7346);
or U7975 (N_7975,N_7377,N_7287);
or U7976 (N_7976,N_7143,N_7068);
nand U7977 (N_7977,N_7084,N_7290);
nand U7978 (N_7978,N_7204,N_7331);
or U7979 (N_7979,N_7079,N_7256);
nand U7980 (N_7980,N_7317,N_7162);
xnor U7981 (N_7981,N_7377,N_7493);
or U7982 (N_7982,N_7298,N_7449);
or U7983 (N_7983,N_7034,N_7173);
nand U7984 (N_7984,N_7233,N_7207);
nor U7985 (N_7985,N_7489,N_7272);
or U7986 (N_7986,N_7143,N_7107);
xor U7987 (N_7987,N_7269,N_7451);
or U7988 (N_7988,N_7086,N_7316);
nand U7989 (N_7989,N_7437,N_7305);
xor U7990 (N_7990,N_7300,N_7318);
nand U7991 (N_7991,N_7137,N_7120);
and U7992 (N_7992,N_7292,N_7016);
nand U7993 (N_7993,N_7040,N_7134);
nand U7994 (N_7994,N_7171,N_7060);
or U7995 (N_7995,N_7238,N_7462);
and U7996 (N_7996,N_7315,N_7077);
or U7997 (N_7997,N_7287,N_7420);
nor U7998 (N_7998,N_7237,N_7225);
or U7999 (N_7999,N_7329,N_7202);
nor U8000 (N_8000,N_7976,N_7860);
nor U8001 (N_8001,N_7908,N_7567);
nor U8002 (N_8002,N_7997,N_7564);
and U8003 (N_8003,N_7762,N_7984);
nand U8004 (N_8004,N_7663,N_7753);
or U8005 (N_8005,N_7503,N_7586);
or U8006 (N_8006,N_7689,N_7556);
nor U8007 (N_8007,N_7602,N_7927);
and U8008 (N_8008,N_7943,N_7965);
or U8009 (N_8009,N_7505,N_7871);
nand U8010 (N_8010,N_7791,N_7966);
nor U8011 (N_8011,N_7604,N_7893);
and U8012 (N_8012,N_7509,N_7831);
nor U8013 (N_8013,N_7983,N_7936);
nand U8014 (N_8014,N_7933,N_7738);
nor U8015 (N_8015,N_7818,N_7867);
nor U8016 (N_8016,N_7733,N_7882);
nand U8017 (N_8017,N_7838,N_7656);
and U8018 (N_8018,N_7999,N_7875);
nor U8019 (N_8019,N_7565,N_7916);
and U8020 (N_8020,N_7971,N_7687);
nand U8021 (N_8021,N_7819,N_7551);
or U8022 (N_8022,N_7700,N_7577);
and U8023 (N_8023,N_7562,N_7822);
nand U8024 (N_8024,N_7606,N_7519);
nor U8025 (N_8025,N_7806,N_7677);
xnor U8026 (N_8026,N_7963,N_7542);
or U8027 (N_8027,N_7845,N_7872);
nand U8028 (N_8028,N_7625,N_7920);
xnor U8029 (N_8029,N_7574,N_7977);
and U8030 (N_8030,N_7825,N_7580);
nor U8031 (N_8031,N_7731,N_7619);
nand U8032 (N_8032,N_7514,N_7967);
nor U8033 (N_8033,N_7555,N_7902);
xor U8034 (N_8034,N_7937,N_7877);
xnor U8035 (N_8035,N_7746,N_7549);
nor U8036 (N_8036,N_7608,N_7942);
or U8037 (N_8037,N_7940,N_7615);
or U8038 (N_8038,N_7830,N_7704);
nand U8039 (N_8039,N_7684,N_7850);
nand U8040 (N_8040,N_7925,N_7587);
nor U8041 (N_8041,N_7524,N_7754);
nor U8042 (N_8042,N_7705,N_7973);
nand U8043 (N_8043,N_7617,N_7773);
or U8044 (N_8044,N_7926,N_7585);
xnor U8045 (N_8045,N_7673,N_7546);
xnor U8046 (N_8046,N_7594,N_7719);
nand U8047 (N_8047,N_7905,N_7525);
and U8048 (N_8048,N_7897,N_7712);
xnor U8049 (N_8049,N_7508,N_7513);
or U8050 (N_8050,N_7647,N_7766);
or U8051 (N_8051,N_7781,N_7755);
and U8052 (N_8052,N_7785,N_7894);
nor U8053 (N_8053,N_7797,N_7723);
and U8054 (N_8054,N_7691,N_7532);
and U8055 (N_8055,N_7631,N_7708);
nand U8056 (N_8056,N_7763,N_7742);
and U8057 (N_8057,N_7868,N_7760);
or U8058 (N_8058,N_7758,N_7989);
or U8059 (N_8059,N_7857,N_7652);
xor U8060 (N_8060,N_7517,N_7750);
or U8061 (N_8061,N_7686,N_7690);
or U8062 (N_8062,N_7559,N_7826);
and U8063 (N_8063,N_7727,N_7671);
and U8064 (N_8064,N_7832,N_7840);
nand U8065 (N_8065,N_7952,N_7698);
and U8066 (N_8066,N_7887,N_7960);
or U8067 (N_8067,N_7552,N_7995);
and U8068 (N_8068,N_7911,N_7506);
nor U8069 (N_8069,N_7648,N_7804);
and U8070 (N_8070,N_7610,N_7788);
and U8071 (N_8071,N_7828,N_7855);
and U8072 (N_8072,N_7544,N_7722);
or U8073 (N_8073,N_7747,N_7575);
nand U8074 (N_8074,N_7693,N_7573);
or U8075 (N_8075,N_7789,N_7720);
and U8076 (N_8076,N_7732,N_7581);
nor U8077 (N_8077,N_7847,N_7912);
and U8078 (N_8078,N_7814,N_7557);
or U8079 (N_8079,N_7770,N_7659);
and U8080 (N_8080,N_7682,N_7834);
nand U8081 (N_8081,N_7558,N_7802);
nand U8082 (N_8082,N_7986,N_7817);
or U8083 (N_8083,N_7646,N_7523);
nor U8084 (N_8084,N_7563,N_7701);
nand U8085 (N_8085,N_7778,N_7842);
nand U8086 (N_8086,N_7672,N_7697);
or U8087 (N_8087,N_7801,N_7990);
and U8088 (N_8088,N_7643,N_7784);
nor U8089 (N_8089,N_7869,N_7991);
and U8090 (N_8090,N_7603,N_7566);
nand U8091 (N_8091,N_7721,N_7534);
nand U8092 (N_8092,N_7833,N_7675);
nand U8093 (N_8093,N_7735,N_7931);
or U8094 (N_8094,N_7730,N_7816);
nand U8095 (N_8095,N_7622,N_7707);
and U8096 (N_8096,N_7950,N_7810);
and U8097 (N_8097,N_7919,N_7741);
nand U8098 (N_8098,N_7811,N_7605);
nand U8099 (N_8099,N_7703,N_7982);
and U8100 (N_8100,N_7944,N_7512);
nor U8101 (N_8101,N_7918,N_7539);
xor U8102 (N_8102,N_7985,N_7692);
or U8103 (N_8103,N_7921,N_7772);
nor U8104 (N_8104,N_7815,N_7890);
and U8105 (N_8105,N_7764,N_7752);
nor U8106 (N_8106,N_7809,N_7792);
and U8107 (N_8107,N_7642,N_7529);
nand U8108 (N_8108,N_7666,N_7618);
nand U8109 (N_8109,N_7543,N_7669);
and U8110 (N_8110,N_7953,N_7561);
nor U8111 (N_8111,N_7545,N_7924);
xor U8112 (N_8112,N_7679,N_7592);
or U8113 (N_8113,N_7507,N_7527);
and U8114 (N_8114,N_7765,N_7694);
xnor U8115 (N_8115,N_7835,N_7824);
nand U8116 (N_8116,N_7923,N_7794);
xnor U8117 (N_8117,N_7596,N_7695);
nand U8118 (N_8118,N_7620,N_7928);
and U8119 (N_8119,N_7676,N_7530);
or U8120 (N_8120,N_7637,N_7880);
nor U8121 (N_8121,N_7862,N_7956);
or U8122 (N_8122,N_7502,N_7964);
nand U8123 (N_8123,N_7511,N_7793);
nor U8124 (N_8124,N_7548,N_7907);
nor U8125 (N_8125,N_7972,N_7888);
xor U8126 (N_8126,N_7504,N_7849);
nor U8127 (N_8127,N_7613,N_7521);
nor U8128 (N_8128,N_7678,N_7959);
nor U8129 (N_8129,N_7803,N_7807);
nand U8130 (N_8130,N_7946,N_7829);
and U8131 (N_8131,N_7598,N_7589);
nor U8132 (N_8132,N_7591,N_7994);
nor U8133 (N_8133,N_7767,N_7582);
or U8134 (N_8134,N_7533,N_7726);
nand U8135 (N_8135,N_7632,N_7630);
or U8136 (N_8136,N_7724,N_7884);
nand U8137 (N_8137,N_7651,N_7540);
and U8138 (N_8138,N_7820,N_7570);
or U8139 (N_8139,N_7547,N_7969);
and U8140 (N_8140,N_7714,N_7510);
or U8141 (N_8141,N_7629,N_7681);
nand U8142 (N_8142,N_7653,N_7590);
nand U8143 (N_8143,N_7958,N_7537);
nor U8144 (N_8144,N_7531,N_7661);
nor U8145 (N_8145,N_7866,N_7568);
or U8146 (N_8146,N_7627,N_7827);
or U8147 (N_8147,N_7650,N_7856);
and U8148 (N_8148,N_7904,N_7939);
or U8149 (N_8149,N_7914,N_7645);
and U8150 (N_8150,N_7578,N_7836);
and U8151 (N_8151,N_7846,N_7883);
xor U8152 (N_8152,N_7812,N_7736);
and U8153 (N_8153,N_7635,N_7518);
and U8154 (N_8154,N_7898,N_7528);
nand U8155 (N_8155,N_7761,N_7879);
or U8156 (N_8156,N_7680,N_7777);
or U8157 (N_8157,N_7769,N_7571);
and U8158 (N_8158,N_7706,N_7900);
nor U8159 (N_8159,N_7843,N_7639);
or U8160 (N_8160,N_7748,N_7636);
or U8161 (N_8161,N_7878,N_7938);
xnor U8162 (N_8162,N_7892,N_7696);
or U8163 (N_8163,N_7998,N_7616);
and U8164 (N_8164,N_7584,N_7853);
nand U8165 (N_8165,N_7974,N_7796);
nand U8166 (N_8166,N_7917,N_7873);
xnor U8167 (N_8167,N_7725,N_7992);
or U8168 (N_8168,N_7751,N_7716);
or U8169 (N_8169,N_7713,N_7996);
nor U8170 (N_8170,N_7955,N_7607);
or U8171 (N_8171,N_7588,N_7710);
and U8172 (N_8172,N_7699,N_7913);
or U8173 (N_8173,N_7515,N_7930);
or U8174 (N_8174,N_7711,N_7638);
or U8175 (N_8175,N_7771,N_7683);
nor U8176 (N_8176,N_7660,N_7858);
nand U8177 (N_8177,N_7805,N_7572);
or U8178 (N_8178,N_7909,N_7813);
and U8179 (N_8179,N_7979,N_7837);
nand U8180 (N_8180,N_7674,N_7612);
nand U8181 (N_8181,N_7554,N_7962);
nand U8182 (N_8182,N_7739,N_7941);
xor U8183 (N_8183,N_7729,N_7553);
or U8184 (N_8184,N_7749,N_7623);
or U8185 (N_8185,N_7945,N_7975);
or U8186 (N_8186,N_7644,N_7949);
nor U8187 (N_8187,N_7864,N_7848);
nand U8188 (N_8188,N_7621,N_7500);
or U8189 (N_8189,N_7759,N_7935);
or U8190 (N_8190,N_7968,N_7665);
and U8191 (N_8191,N_7745,N_7601);
nand U8192 (N_8192,N_7667,N_7861);
nand U8193 (N_8193,N_7609,N_7633);
or U8194 (N_8194,N_7782,N_7576);
nand U8195 (N_8195,N_7852,N_7881);
or U8196 (N_8196,N_7886,N_7839);
and U8197 (N_8197,N_7664,N_7786);
and U8198 (N_8198,N_7654,N_7717);
xnor U8199 (N_8199,N_7993,N_7611);
nand U8200 (N_8200,N_7954,N_7932);
and U8201 (N_8201,N_7655,N_7685);
nor U8202 (N_8202,N_7961,N_7541);
nor U8203 (N_8203,N_7798,N_7934);
or U8204 (N_8204,N_7628,N_7740);
nor U8205 (N_8205,N_7957,N_7970);
nand U8206 (N_8206,N_7688,N_7987);
nor U8207 (N_8207,N_7865,N_7891);
and U8208 (N_8208,N_7600,N_7841);
or U8209 (N_8209,N_7583,N_7597);
nor U8210 (N_8210,N_7768,N_7526);
and U8211 (N_8211,N_7743,N_7915);
and U8212 (N_8212,N_7657,N_7718);
nor U8213 (N_8213,N_7895,N_7981);
nor U8214 (N_8214,N_7948,N_7988);
nor U8215 (N_8215,N_7737,N_7901);
and U8216 (N_8216,N_7641,N_7595);
xor U8217 (N_8217,N_7774,N_7889);
nand U8218 (N_8218,N_7780,N_7624);
nand U8219 (N_8219,N_7538,N_7903);
nor U8220 (N_8220,N_7978,N_7980);
nor U8221 (N_8221,N_7709,N_7779);
or U8222 (N_8222,N_7787,N_7808);
nand U8223 (N_8223,N_7863,N_7910);
or U8224 (N_8224,N_7899,N_7658);
nor U8225 (N_8225,N_7614,N_7536);
xnor U8226 (N_8226,N_7634,N_7560);
nand U8227 (N_8227,N_7823,N_7756);
or U8228 (N_8228,N_7795,N_7649);
or U8229 (N_8229,N_7922,N_7896);
and U8230 (N_8230,N_7800,N_7744);
and U8231 (N_8231,N_7593,N_7640);
or U8232 (N_8232,N_7947,N_7844);
and U8233 (N_8233,N_7715,N_7516);
nand U8234 (N_8234,N_7870,N_7501);
or U8235 (N_8235,N_7859,N_7702);
and U8236 (N_8236,N_7906,N_7851);
or U8237 (N_8237,N_7626,N_7885);
and U8238 (N_8238,N_7599,N_7876);
and U8239 (N_8239,N_7757,N_7790);
nand U8240 (N_8240,N_7670,N_7821);
or U8241 (N_8241,N_7734,N_7522);
nor U8242 (N_8242,N_7520,N_7854);
or U8243 (N_8243,N_7579,N_7929);
and U8244 (N_8244,N_7535,N_7550);
and U8245 (N_8245,N_7569,N_7783);
and U8246 (N_8246,N_7951,N_7668);
and U8247 (N_8247,N_7874,N_7775);
nor U8248 (N_8248,N_7728,N_7776);
or U8249 (N_8249,N_7799,N_7662);
nor U8250 (N_8250,N_7637,N_7887);
nor U8251 (N_8251,N_7504,N_7668);
xnor U8252 (N_8252,N_7600,N_7852);
nand U8253 (N_8253,N_7594,N_7622);
nand U8254 (N_8254,N_7888,N_7600);
or U8255 (N_8255,N_7853,N_7550);
nor U8256 (N_8256,N_7703,N_7519);
xnor U8257 (N_8257,N_7646,N_7963);
nor U8258 (N_8258,N_7902,N_7588);
nor U8259 (N_8259,N_7656,N_7939);
nor U8260 (N_8260,N_7527,N_7721);
nand U8261 (N_8261,N_7524,N_7865);
nand U8262 (N_8262,N_7560,N_7713);
nand U8263 (N_8263,N_7606,N_7933);
or U8264 (N_8264,N_7683,N_7647);
and U8265 (N_8265,N_7606,N_7572);
nand U8266 (N_8266,N_7648,N_7605);
xnor U8267 (N_8267,N_7780,N_7575);
and U8268 (N_8268,N_7606,N_7795);
xnor U8269 (N_8269,N_7654,N_7831);
and U8270 (N_8270,N_7740,N_7537);
and U8271 (N_8271,N_7701,N_7626);
and U8272 (N_8272,N_7919,N_7727);
nand U8273 (N_8273,N_7839,N_7717);
nand U8274 (N_8274,N_7866,N_7880);
or U8275 (N_8275,N_7784,N_7929);
or U8276 (N_8276,N_7648,N_7998);
nand U8277 (N_8277,N_7733,N_7898);
nand U8278 (N_8278,N_7931,N_7672);
and U8279 (N_8279,N_7753,N_7632);
or U8280 (N_8280,N_7802,N_7530);
nand U8281 (N_8281,N_7585,N_7935);
and U8282 (N_8282,N_7993,N_7778);
nand U8283 (N_8283,N_7736,N_7633);
and U8284 (N_8284,N_7934,N_7834);
nand U8285 (N_8285,N_7858,N_7873);
and U8286 (N_8286,N_7583,N_7718);
or U8287 (N_8287,N_7773,N_7543);
nand U8288 (N_8288,N_7535,N_7554);
or U8289 (N_8289,N_7777,N_7623);
xor U8290 (N_8290,N_7739,N_7899);
xnor U8291 (N_8291,N_7838,N_7824);
or U8292 (N_8292,N_7828,N_7792);
nand U8293 (N_8293,N_7937,N_7820);
and U8294 (N_8294,N_7876,N_7854);
nor U8295 (N_8295,N_7973,N_7994);
nor U8296 (N_8296,N_7898,N_7980);
and U8297 (N_8297,N_7765,N_7606);
and U8298 (N_8298,N_7855,N_7763);
nand U8299 (N_8299,N_7921,N_7879);
nand U8300 (N_8300,N_7610,N_7801);
and U8301 (N_8301,N_7885,N_7935);
nor U8302 (N_8302,N_7993,N_7924);
or U8303 (N_8303,N_7958,N_7911);
and U8304 (N_8304,N_7579,N_7714);
xor U8305 (N_8305,N_7785,N_7520);
xnor U8306 (N_8306,N_7668,N_7618);
nand U8307 (N_8307,N_7871,N_7860);
and U8308 (N_8308,N_7763,N_7789);
or U8309 (N_8309,N_7854,N_7907);
nand U8310 (N_8310,N_7967,N_7789);
or U8311 (N_8311,N_7841,N_7870);
or U8312 (N_8312,N_7958,N_7503);
nand U8313 (N_8313,N_7602,N_7665);
nor U8314 (N_8314,N_7760,N_7746);
nor U8315 (N_8315,N_7864,N_7880);
nor U8316 (N_8316,N_7795,N_7893);
nor U8317 (N_8317,N_7601,N_7966);
and U8318 (N_8318,N_7928,N_7546);
and U8319 (N_8319,N_7574,N_7551);
and U8320 (N_8320,N_7584,N_7509);
or U8321 (N_8321,N_7753,N_7945);
nand U8322 (N_8322,N_7819,N_7665);
and U8323 (N_8323,N_7937,N_7940);
xor U8324 (N_8324,N_7898,N_7559);
or U8325 (N_8325,N_7712,N_7643);
nor U8326 (N_8326,N_7522,N_7872);
or U8327 (N_8327,N_7614,N_7543);
or U8328 (N_8328,N_7849,N_7729);
and U8329 (N_8329,N_7757,N_7968);
nand U8330 (N_8330,N_7517,N_7667);
and U8331 (N_8331,N_7517,N_7883);
nor U8332 (N_8332,N_7518,N_7663);
nor U8333 (N_8333,N_7711,N_7580);
nor U8334 (N_8334,N_7765,N_7729);
or U8335 (N_8335,N_7577,N_7632);
nand U8336 (N_8336,N_7878,N_7792);
nand U8337 (N_8337,N_7539,N_7710);
nand U8338 (N_8338,N_7967,N_7632);
or U8339 (N_8339,N_7966,N_7676);
and U8340 (N_8340,N_7652,N_7944);
and U8341 (N_8341,N_7756,N_7724);
or U8342 (N_8342,N_7819,N_7782);
or U8343 (N_8343,N_7855,N_7500);
and U8344 (N_8344,N_7811,N_7633);
and U8345 (N_8345,N_7759,N_7687);
and U8346 (N_8346,N_7672,N_7917);
nand U8347 (N_8347,N_7864,N_7704);
nor U8348 (N_8348,N_7939,N_7807);
and U8349 (N_8349,N_7721,N_7605);
nand U8350 (N_8350,N_7770,N_7792);
nor U8351 (N_8351,N_7823,N_7702);
xor U8352 (N_8352,N_7793,N_7590);
and U8353 (N_8353,N_7718,N_7800);
or U8354 (N_8354,N_7705,N_7832);
nand U8355 (N_8355,N_7737,N_7626);
and U8356 (N_8356,N_7850,N_7535);
nand U8357 (N_8357,N_7773,N_7534);
nand U8358 (N_8358,N_7618,N_7607);
nand U8359 (N_8359,N_7828,N_7987);
nor U8360 (N_8360,N_7697,N_7909);
nor U8361 (N_8361,N_7835,N_7915);
nand U8362 (N_8362,N_7734,N_7873);
nor U8363 (N_8363,N_7754,N_7555);
nand U8364 (N_8364,N_7923,N_7509);
and U8365 (N_8365,N_7843,N_7892);
nand U8366 (N_8366,N_7744,N_7577);
nand U8367 (N_8367,N_7647,N_7671);
xnor U8368 (N_8368,N_7520,N_7860);
nand U8369 (N_8369,N_7856,N_7873);
nor U8370 (N_8370,N_7647,N_7586);
and U8371 (N_8371,N_7640,N_7853);
and U8372 (N_8372,N_7942,N_7744);
or U8373 (N_8373,N_7891,N_7778);
and U8374 (N_8374,N_7542,N_7607);
nand U8375 (N_8375,N_7842,N_7722);
nand U8376 (N_8376,N_7704,N_7868);
xnor U8377 (N_8377,N_7945,N_7507);
nand U8378 (N_8378,N_7697,N_7832);
or U8379 (N_8379,N_7774,N_7907);
nand U8380 (N_8380,N_7768,N_7976);
nor U8381 (N_8381,N_7790,N_7759);
nand U8382 (N_8382,N_7708,N_7821);
nor U8383 (N_8383,N_7882,N_7644);
xnor U8384 (N_8384,N_7516,N_7683);
nor U8385 (N_8385,N_7618,N_7994);
nand U8386 (N_8386,N_7877,N_7791);
and U8387 (N_8387,N_7945,N_7777);
nor U8388 (N_8388,N_7996,N_7528);
and U8389 (N_8389,N_7988,N_7947);
nand U8390 (N_8390,N_7742,N_7526);
xnor U8391 (N_8391,N_7923,N_7606);
and U8392 (N_8392,N_7683,N_7746);
or U8393 (N_8393,N_7625,N_7565);
and U8394 (N_8394,N_7561,N_7906);
nand U8395 (N_8395,N_7896,N_7959);
nand U8396 (N_8396,N_7836,N_7585);
or U8397 (N_8397,N_7701,N_7811);
nand U8398 (N_8398,N_7718,N_7736);
nor U8399 (N_8399,N_7980,N_7530);
xor U8400 (N_8400,N_7556,N_7707);
or U8401 (N_8401,N_7919,N_7522);
nor U8402 (N_8402,N_7529,N_7848);
and U8403 (N_8403,N_7684,N_7864);
or U8404 (N_8404,N_7968,N_7901);
and U8405 (N_8405,N_7850,N_7906);
nand U8406 (N_8406,N_7671,N_7662);
xnor U8407 (N_8407,N_7562,N_7888);
nand U8408 (N_8408,N_7605,N_7584);
nand U8409 (N_8409,N_7614,N_7954);
xor U8410 (N_8410,N_7528,N_7676);
xor U8411 (N_8411,N_7714,N_7734);
nand U8412 (N_8412,N_7537,N_7893);
nor U8413 (N_8413,N_7654,N_7762);
nor U8414 (N_8414,N_7624,N_7529);
nand U8415 (N_8415,N_7565,N_7980);
nor U8416 (N_8416,N_7837,N_7928);
nand U8417 (N_8417,N_7622,N_7541);
nand U8418 (N_8418,N_7655,N_7601);
nand U8419 (N_8419,N_7700,N_7878);
xnor U8420 (N_8420,N_7983,N_7904);
nor U8421 (N_8421,N_7826,N_7609);
nand U8422 (N_8422,N_7710,N_7794);
nor U8423 (N_8423,N_7755,N_7953);
nor U8424 (N_8424,N_7817,N_7542);
nor U8425 (N_8425,N_7616,N_7776);
nand U8426 (N_8426,N_7664,N_7777);
and U8427 (N_8427,N_7849,N_7650);
nor U8428 (N_8428,N_7617,N_7709);
nor U8429 (N_8429,N_7535,N_7801);
nor U8430 (N_8430,N_7551,N_7559);
or U8431 (N_8431,N_7555,N_7906);
nand U8432 (N_8432,N_7714,N_7884);
or U8433 (N_8433,N_7614,N_7895);
or U8434 (N_8434,N_7849,N_7885);
nor U8435 (N_8435,N_7835,N_7791);
nand U8436 (N_8436,N_7803,N_7631);
and U8437 (N_8437,N_7909,N_7722);
nand U8438 (N_8438,N_7885,N_7735);
and U8439 (N_8439,N_7777,N_7636);
and U8440 (N_8440,N_7584,N_7585);
nand U8441 (N_8441,N_7715,N_7826);
and U8442 (N_8442,N_7857,N_7638);
xor U8443 (N_8443,N_7807,N_7779);
nor U8444 (N_8444,N_7961,N_7880);
nor U8445 (N_8445,N_7844,N_7756);
xor U8446 (N_8446,N_7575,N_7682);
or U8447 (N_8447,N_7634,N_7531);
xor U8448 (N_8448,N_7584,N_7586);
xor U8449 (N_8449,N_7705,N_7557);
xnor U8450 (N_8450,N_7718,N_7731);
xor U8451 (N_8451,N_7973,N_7874);
nand U8452 (N_8452,N_7900,N_7742);
nand U8453 (N_8453,N_7756,N_7893);
nor U8454 (N_8454,N_7992,N_7974);
nor U8455 (N_8455,N_7869,N_7844);
xor U8456 (N_8456,N_7552,N_7677);
or U8457 (N_8457,N_7728,N_7800);
or U8458 (N_8458,N_7765,N_7787);
or U8459 (N_8459,N_7899,N_7951);
and U8460 (N_8460,N_7845,N_7639);
nand U8461 (N_8461,N_7940,N_7926);
nand U8462 (N_8462,N_7869,N_7841);
nor U8463 (N_8463,N_7624,N_7756);
nor U8464 (N_8464,N_7522,N_7526);
or U8465 (N_8465,N_7740,N_7529);
nor U8466 (N_8466,N_7942,N_7847);
or U8467 (N_8467,N_7829,N_7886);
and U8468 (N_8468,N_7660,N_7806);
or U8469 (N_8469,N_7717,N_7595);
or U8470 (N_8470,N_7747,N_7833);
or U8471 (N_8471,N_7664,N_7570);
or U8472 (N_8472,N_7765,N_7665);
nor U8473 (N_8473,N_7715,N_7691);
nor U8474 (N_8474,N_7910,N_7889);
or U8475 (N_8475,N_7835,N_7733);
nor U8476 (N_8476,N_7931,N_7957);
or U8477 (N_8477,N_7753,N_7555);
and U8478 (N_8478,N_7816,N_7616);
and U8479 (N_8479,N_7813,N_7954);
and U8480 (N_8480,N_7580,N_7948);
nand U8481 (N_8481,N_7894,N_7678);
or U8482 (N_8482,N_7845,N_7909);
or U8483 (N_8483,N_7643,N_7960);
or U8484 (N_8484,N_7865,N_7911);
and U8485 (N_8485,N_7775,N_7846);
or U8486 (N_8486,N_7647,N_7871);
and U8487 (N_8487,N_7658,N_7888);
xnor U8488 (N_8488,N_7886,N_7847);
nor U8489 (N_8489,N_7905,N_7598);
or U8490 (N_8490,N_7858,N_7625);
and U8491 (N_8491,N_7598,N_7774);
nor U8492 (N_8492,N_7827,N_7783);
and U8493 (N_8493,N_7557,N_7898);
nand U8494 (N_8494,N_7643,N_7871);
nor U8495 (N_8495,N_7564,N_7908);
and U8496 (N_8496,N_7877,N_7558);
and U8497 (N_8497,N_7675,N_7965);
nor U8498 (N_8498,N_7845,N_7589);
nand U8499 (N_8499,N_7675,N_7931);
nand U8500 (N_8500,N_8323,N_8092);
nor U8501 (N_8501,N_8170,N_8411);
xor U8502 (N_8502,N_8493,N_8476);
xor U8503 (N_8503,N_8121,N_8274);
nor U8504 (N_8504,N_8388,N_8135);
nor U8505 (N_8505,N_8357,N_8262);
nand U8506 (N_8506,N_8327,N_8094);
nor U8507 (N_8507,N_8430,N_8286);
nor U8508 (N_8508,N_8478,N_8143);
nor U8509 (N_8509,N_8394,N_8372);
or U8510 (N_8510,N_8350,N_8193);
or U8511 (N_8511,N_8182,N_8043);
or U8512 (N_8512,N_8011,N_8487);
and U8513 (N_8513,N_8341,N_8335);
or U8514 (N_8514,N_8406,N_8378);
and U8515 (N_8515,N_8384,N_8112);
xnor U8516 (N_8516,N_8263,N_8412);
nor U8517 (N_8517,N_8008,N_8477);
nand U8518 (N_8518,N_8063,N_8315);
nor U8519 (N_8519,N_8024,N_8302);
and U8520 (N_8520,N_8014,N_8438);
or U8521 (N_8521,N_8303,N_8454);
nor U8522 (N_8522,N_8334,N_8171);
nor U8523 (N_8523,N_8093,N_8201);
nand U8524 (N_8524,N_8195,N_8001);
nor U8525 (N_8525,N_8108,N_8187);
or U8526 (N_8526,N_8326,N_8029);
and U8527 (N_8527,N_8453,N_8256);
xnor U8528 (N_8528,N_8047,N_8332);
nor U8529 (N_8529,N_8374,N_8348);
nor U8530 (N_8530,N_8220,N_8481);
and U8531 (N_8531,N_8206,N_8105);
and U8532 (N_8532,N_8393,N_8349);
nor U8533 (N_8533,N_8333,N_8144);
or U8534 (N_8534,N_8129,N_8319);
nor U8535 (N_8535,N_8351,N_8317);
or U8536 (N_8536,N_8181,N_8124);
and U8537 (N_8537,N_8285,N_8134);
or U8538 (N_8538,N_8486,N_8176);
nand U8539 (N_8539,N_8316,N_8455);
or U8540 (N_8540,N_8280,N_8085);
nand U8541 (N_8541,N_8208,N_8371);
or U8542 (N_8542,N_8295,N_8055);
and U8543 (N_8543,N_8346,N_8004);
or U8544 (N_8544,N_8254,N_8034);
nand U8545 (N_8545,N_8417,N_8210);
nand U8546 (N_8546,N_8272,N_8118);
xnor U8547 (N_8547,N_8185,N_8418);
nand U8548 (N_8548,N_8140,N_8373);
nor U8549 (N_8549,N_8164,N_8240);
or U8550 (N_8550,N_8192,N_8368);
and U8551 (N_8551,N_8204,N_8102);
or U8552 (N_8552,N_8083,N_8246);
xor U8553 (N_8553,N_8071,N_8475);
xor U8554 (N_8554,N_8459,N_8401);
and U8555 (N_8555,N_8050,N_8407);
or U8556 (N_8556,N_8397,N_8362);
and U8557 (N_8557,N_8474,N_8087);
nand U8558 (N_8558,N_8367,N_8441);
and U8559 (N_8559,N_8312,N_8236);
or U8560 (N_8560,N_8156,N_8032);
or U8561 (N_8561,N_8365,N_8379);
or U8562 (N_8562,N_8252,N_8157);
nor U8563 (N_8563,N_8443,N_8091);
or U8564 (N_8564,N_8084,N_8276);
nor U8565 (N_8565,N_8184,N_8101);
nor U8566 (N_8566,N_8287,N_8068);
nor U8567 (N_8567,N_8222,N_8284);
nand U8568 (N_8568,N_8098,N_8122);
nor U8569 (N_8569,N_8452,N_8211);
nor U8570 (N_8570,N_8225,N_8337);
or U8571 (N_8571,N_8313,N_8450);
nor U8572 (N_8572,N_8300,N_8456);
and U8573 (N_8573,N_8281,N_8268);
or U8574 (N_8574,N_8377,N_8429);
or U8575 (N_8575,N_8003,N_8423);
and U8576 (N_8576,N_8449,N_8433);
nand U8577 (N_8577,N_8463,N_8081);
and U8578 (N_8578,N_8392,N_8369);
nor U8579 (N_8579,N_8364,N_8307);
nor U8580 (N_8580,N_8296,N_8131);
nor U8581 (N_8581,N_8078,N_8179);
nor U8582 (N_8582,N_8328,N_8436);
xnor U8583 (N_8583,N_8126,N_8205);
nor U8584 (N_8584,N_8483,N_8191);
nand U8585 (N_8585,N_8221,N_8283);
and U8586 (N_8586,N_8239,N_8488);
nand U8587 (N_8587,N_8294,N_8103);
nand U8588 (N_8588,N_8408,N_8217);
and U8589 (N_8589,N_8036,N_8489);
nor U8590 (N_8590,N_8200,N_8203);
and U8591 (N_8591,N_8416,N_8444);
nor U8592 (N_8592,N_8405,N_8042);
xor U8593 (N_8593,N_8168,N_8067);
nand U8594 (N_8594,N_8288,N_8117);
nor U8595 (N_8595,N_8147,N_8161);
nor U8596 (N_8596,N_8304,N_8207);
or U8597 (N_8597,N_8038,N_8498);
xor U8598 (N_8598,N_8190,N_8282);
or U8599 (N_8599,N_8391,N_8451);
nor U8600 (N_8600,N_8330,N_8109);
nand U8601 (N_8601,N_8457,N_8216);
or U8602 (N_8602,N_8104,N_8089);
nor U8603 (N_8603,N_8471,N_8106);
nor U8604 (N_8604,N_8021,N_8381);
or U8605 (N_8605,N_8172,N_8426);
nand U8606 (N_8606,N_8030,N_8142);
nand U8607 (N_8607,N_8051,N_8025);
xor U8608 (N_8608,N_8226,N_8229);
nor U8609 (N_8609,N_8308,N_8037);
xnor U8610 (N_8610,N_8149,N_8027);
nand U8611 (N_8611,N_8010,N_8159);
and U8612 (N_8612,N_8301,N_8020);
nand U8613 (N_8613,N_8439,N_8244);
or U8614 (N_8614,N_8231,N_8138);
xnor U8615 (N_8615,N_8146,N_8427);
nor U8616 (N_8616,N_8228,N_8306);
nand U8617 (N_8617,N_8347,N_8005);
or U8618 (N_8618,N_8292,N_8189);
or U8619 (N_8619,N_8261,N_8044);
or U8620 (N_8620,N_8119,N_8133);
nor U8621 (N_8621,N_8165,N_8026);
xnor U8622 (N_8622,N_8458,N_8345);
and U8623 (N_8623,N_8033,N_8338);
nand U8624 (N_8624,N_8188,N_8310);
and U8625 (N_8625,N_8158,N_8479);
or U8626 (N_8626,N_8095,N_8139);
nor U8627 (N_8627,N_8052,N_8297);
or U8628 (N_8628,N_8123,N_8040);
or U8629 (N_8629,N_8311,N_8329);
xor U8630 (N_8630,N_8497,N_8363);
xor U8631 (N_8631,N_8358,N_8079);
and U8632 (N_8632,N_8445,N_8096);
nand U8633 (N_8633,N_8062,N_8414);
or U8634 (N_8634,N_8446,N_8057);
xnor U8635 (N_8635,N_8435,N_8440);
or U8636 (N_8636,N_8107,N_8464);
or U8637 (N_8637,N_8403,N_8293);
nor U8638 (N_8638,N_8421,N_8070);
or U8639 (N_8639,N_8006,N_8234);
nand U8640 (N_8640,N_8480,N_8383);
nor U8641 (N_8641,N_8413,N_8321);
nor U8642 (N_8642,N_8198,N_8279);
and U8643 (N_8643,N_8233,N_8227);
nand U8644 (N_8644,N_8495,N_8485);
or U8645 (N_8645,N_8245,N_8058);
or U8646 (N_8646,N_8342,N_8088);
nand U8647 (N_8647,N_8173,N_8237);
nor U8648 (N_8648,N_8404,N_8180);
nand U8649 (N_8649,N_8399,N_8082);
nand U8650 (N_8650,N_8097,N_8023);
and U8651 (N_8651,N_8178,N_8065);
nand U8652 (N_8652,N_8425,N_8410);
nor U8653 (N_8653,N_8484,N_8465);
xnor U8654 (N_8654,N_8039,N_8163);
and U8655 (N_8655,N_8099,N_8428);
and U8656 (N_8656,N_8309,N_8223);
and U8657 (N_8657,N_8130,N_8448);
and U8658 (N_8658,N_8437,N_8110);
and U8659 (N_8659,N_8420,N_8291);
and U8660 (N_8660,N_8253,N_8127);
nor U8661 (N_8661,N_8056,N_8271);
nor U8662 (N_8662,N_8442,N_8258);
or U8663 (N_8663,N_8366,N_8255);
nor U8664 (N_8664,N_8194,N_8270);
and U8665 (N_8665,N_8324,N_8473);
and U8666 (N_8666,N_8224,N_8382);
or U8667 (N_8667,N_8340,N_8318);
nor U8668 (N_8668,N_8015,N_8266);
nor U8669 (N_8669,N_8072,N_8431);
nor U8670 (N_8670,N_8069,N_8141);
or U8671 (N_8671,N_8202,N_8125);
or U8672 (N_8672,N_8353,N_8007);
nor U8673 (N_8673,N_8322,N_8469);
and U8674 (N_8674,N_8460,N_8273);
or U8675 (N_8675,N_8022,N_8199);
xor U8676 (N_8676,N_8048,N_8390);
or U8677 (N_8677,N_8012,N_8113);
or U8678 (N_8678,N_8213,N_8387);
xor U8679 (N_8679,N_8402,N_8235);
or U8680 (N_8680,N_8472,N_8466);
or U8681 (N_8681,N_8376,N_8230);
or U8682 (N_8682,N_8269,N_8447);
xnor U8683 (N_8683,N_8290,N_8013);
nor U8684 (N_8684,N_8061,N_8160);
nand U8685 (N_8685,N_8482,N_8242);
nand U8686 (N_8686,N_8167,N_8046);
nor U8687 (N_8687,N_8343,N_8016);
or U8688 (N_8688,N_8075,N_8064);
nand U8689 (N_8689,N_8018,N_8060);
nand U8690 (N_8690,N_8218,N_8344);
or U8691 (N_8691,N_8186,N_8002);
and U8692 (N_8692,N_8175,N_8395);
nand U8693 (N_8693,N_8074,N_8086);
xor U8694 (N_8694,N_8017,N_8137);
nor U8695 (N_8695,N_8461,N_8259);
nor U8696 (N_8696,N_8243,N_8260);
or U8697 (N_8697,N_8289,N_8132);
nor U8698 (N_8698,N_8059,N_8155);
and U8699 (N_8699,N_8257,N_8153);
or U8700 (N_8700,N_8277,N_8434);
nor U8701 (N_8701,N_8250,N_8073);
and U8702 (N_8702,N_8249,N_8152);
nand U8703 (N_8703,N_8035,N_8415);
or U8704 (N_8704,N_8177,N_8151);
nand U8705 (N_8705,N_8370,N_8183);
nand U8706 (N_8706,N_8499,N_8385);
or U8707 (N_8707,N_8009,N_8380);
nand U8708 (N_8708,N_8299,N_8494);
and U8709 (N_8709,N_8080,N_8361);
nand U8710 (N_8710,N_8215,N_8251);
nand U8711 (N_8711,N_8325,N_8145);
nor U8712 (N_8712,N_8265,N_8336);
and U8713 (N_8713,N_8264,N_8169);
or U8714 (N_8714,N_8468,N_8154);
nor U8715 (N_8715,N_8077,N_8174);
nand U8716 (N_8716,N_8400,N_8356);
nor U8717 (N_8717,N_8496,N_8424);
nor U8718 (N_8718,N_8041,N_8090);
and U8719 (N_8719,N_8120,N_8331);
and U8720 (N_8720,N_8422,N_8275);
nand U8721 (N_8721,N_8248,N_8214);
nand U8722 (N_8722,N_8491,N_8359);
and U8723 (N_8723,N_8320,N_8432);
or U8724 (N_8724,N_8467,N_8267);
and U8725 (N_8725,N_8212,N_8389);
xor U8726 (N_8726,N_8409,N_8166);
or U8727 (N_8727,N_8419,N_8111);
nor U8728 (N_8728,N_8019,N_8232);
nand U8729 (N_8729,N_8148,N_8049);
or U8730 (N_8730,N_8470,N_8219);
nor U8731 (N_8731,N_8150,N_8352);
xnor U8732 (N_8732,N_8492,N_8398);
or U8733 (N_8733,N_8462,N_8115);
nand U8734 (N_8734,N_8196,N_8000);
nor U8735 (N_8735,N_8354,N_8076);
nand U8736 (N_8736,N_8298,N_8028);
and U8737 (N_8737,N_8305,N_8128);
and U8738 (N_8738,N_8197,N_8114);
nor U8739 (N_8739,N_8355,N_8162);
and U8740 (N_8740,N_8031,N_8314);
or U8741 (N_8741,N_8360,N_8053);
or U8742 (N_8742,N_8339,N_8247);
nand U8743 (N_8743,N_8375,N_8116);
nor U8744 (N_8744,N_8100,N_8136);
or U8745 (N_8745,N_8241,N_8054);
and U8746 (N_8746,N_8278,N_8045);
nor U8747 (N_8747,N_8209,N_8490);
nand U8748 (N_8748,N_8396,N_8386);
and U8749 (N_8749,N_8066,N_8238);
xnor U8750 (N_8750,N_8101,N_8146);
or U8751 (N_8751,N_8044,N_8385);
nand U8752 (N_8752,N_8034,N_8134);
and U8753 (N_8753,N_8466,N_8062);
nor U8754 (N_8754,N_8409,N_8187);
nor U8755 (N_8755,N_8309,N_8238);
or U8756 (N_8756,N_8238,N_8190);
or U8757 (N_8757,N_8330,N_8259);
or U8758 (N_8758,N_8474,N_8440);
nand U8759 (N_8759,N_8086,N_8021);
and U8760 (N_8760,N_8276,N_8124);
and U8761 (N_8761,N_8076,N_8082);
nand U8762 (N_8762,N_8208,N_8212);
nand U8763 (N_8763,N_8014,N_8188);
or U8764 (N_8764,N_8342,N_8451);
and U8765 (N_8765,N_8421,N_8458);
and U8766 (N_8766,N_8188,N_8289);
nor U8767 (N_8767,N_8174,N_8103);
nand U8768 (N_8768,N_8171,N_8413);
nand U8769 (N_8769,N_8062,N_8376);
nand U8770 (N_8770,N_8066,N_8107);
nor U8771 (N_8771,N_8338,N_8205);
and U8772 (N_8772,N_8289,N_8396);
and U8773 (N_8773,N_8403,N_8224);
nand U8774 (N_8774,N_8035,N_8471);
xor U8775 (N_8775,N_8443,N_8440);
nor U8776 (N_8776,N_8266,N_8366);
and U8777 (N_8777,N_8272,N_8253);
nor U8778 (N_8778,N_8030,N_8063);
nand U8779 (N_8779,N_8037,N_8321);
xnor U8780 (N_8780,N_8027,N_8307);
and U8781 (N_8781,N_8177,N_8023);
nor U8782 (N_8782,N_8370,N_8477);
nand U8783 (N_8783,N_8369,N_8314);
nor U8784 (N_8784,N_8178,N_8326);
and U8785 (N_8785,N_8112,N_8329);
or U8786 (N_8786,N_8068,N_8224);
and U8787 (N_8787,N_8309,N_8217);
nand U8788 (N_8788,N_8202,N_8269);
and U8789 (N_8789,N_8171,N_8377);
nor U8790 (N_8790,N_8158,N_8082);
and U8791 (N_8791,N_8376,N_8300);
and U8792 (N_8792,N_8315,N_8162);
nand U8793 (N_8793,N_8106,N_8319);
nor U8794 (N_8794,N_8115,N_8188);
and U8795 (N_8795,N_8198,N_8463);
or U8796 (N_8796,N_8026,N_8430);
or U8797 (N_8797,N_8409,N_8178);
and U8798 (N_8798,N_8422,N_8188);
and U8799 (N_8799,N_8328,N_8217);
nand U8800 (N_8800,N_8135,N_8431);
and U8801 (N_8801,N_8061,N_8086);
nand U8802 (N_8802,N_8092,N_8386);
nor U8803 (N_8803,N_8169,N_8416);
nor U8804 (N_8804,N_8194,N_8210);
nor U8805 (N_8805,N_8067,N_8234);
nor U8806 (N_8806,N_8117,N_8322);
nand U8807 (N_8807,N_8305,N_8489);
or U8808 (N_8808,N_8462,N_8042);
and U8809 (N_8809,N_8191,N_8465);
or U8810 (N_8810,N_8207,N_8377);
and U8811 (N_8811,N_8147,N_8468);
or U8812 (N_8812,N_8425,N_8262);
nand U8813 (N_8813,N_8383,N_8278);
nand U8814 (N_8814,N_8115,N_8426);
nor U8815 (N_8815,N_8451,N_8201);
or U8816 (N_8816,N_8297,N_8028);
nand U8817 (N_8817,N_8238,N_8490);
nand U8818 (N_8818,N_8292,N_8060);
xor U8819 (N_8819,N_8372,N_8374);
or U8820 (N_8820,N_8406,N_8198);
and U8821 (N_8821,N_8123,N_8047);
nor U8822 (N_8822,N_8205,N_8327);
nor U8823 (N_8823,N_8455,N_8466);
nor U8824 (N_8824,N_8444,N_8089);
or U8825 (N_8825,N_8407,N_8295);
or U8826 (N_8826,N_8004,N_8430);
or U8827 (N_8827,N_8278,N_8292);
nor U8828 (N_8828,N_8303,N_8136);
and U8829 (N_8829,N_8204,N_8485);
and U8830 (N_8830,N_8056,N_8426);
or U8831 (N_8831,N_8324,N_8303);
and U8832 (N_8832,N_8220,N_8309);
and U8833 (N_8833,N_8079,N_8098);
nor U8834 (N_8834,N_8136,N_8011);
or U8835 (N_8835,N_8489,N_8084);
nand U8836 (N_8836,N_8173,N_8474);
xor U8837 (N_8837,N_8170,N_8302);
nor U8838 (N_8838,N_8484,N_8070);
nor U8839 (N_8839,N_8432,N_8012);
and U8840 (N_8840,N_8063,N_8359);
xnor U8841 (N_8841,N_8144,N_8421);
or U8842 (N_8842,N_8242,N_8394);
and U8843 (N_8843,N_8477,N_8177);
xor U8844 (N_8844,N_8102,N_8371);
or U8845 (N_8845,N_8193,N_8418);
or U8846 (N_8846,N_8425,N_8406);
or U8847 (N_8847,N_8329,N_8389);
nand U8848 (N_8848,N_8108,N_8129);
xor U8849 (N_8849,N_8426,N_8168);
nand U8850 (N_8850,N_8160,N_8234);
nand U8851 (N_8851,N_8231,N_8284);
and U8852 (N_8852,N_8106,N_8045);
and U8853 (N_8853,N_8274,N_8305);
nor U8854 (N_8854,N_8356,N_8054);
nor U8855 (N_8855,N_8229,N_8107);
nand U8856 (N_8856,N_8243,N_8229);
and U8857 (N_8857,N_8462,N_8239);
nand U8858 (N_8858,N_8017,N_8107);
nor U8859 (N_8859,N_8274,N_8477);
xor U8860 (N_8860,N_8028,N_8192);
nor U8861 (N_8861,N_8326,N_8153);
and U8862 (N_8862,N_8007,N_8412);
nor U8863 (N_8863,N_8439,N_8088);
and U8864 (N_8864,N_8029,N_8089);
nand U8865 (N_8865,N_8223,N_8042);
nand U8866 (N_8866,N_8194,N_8424);
nand U8867 (N_8867,N_8407,N_8076);
xnor U8868 (N_8868,N_8457,N_8031);
xor U8869 (N_8869,N_8397,N_8406);
or U8870 (N_8870,N_8136,N_8478);
and U8871 (N_8871,N_8438,N_8230);
and U8872 (N_8872,N_8274,N_8251);
and U8873 (N_8873,N_8392,N_8438);
nand U8874 (N_8874,N_8261,N_8368);
nand U8875 (N_8875,N_8007,N_8084);
or U8876 (N_8876,N_8490,N_8382);
and U8877 (N_8877,N_8420,N_8151);
xnor U8878 (N_8878,N_8275,N_8253);
or U8879 (N_8879,N_8325,N_8324);
nor U8880 (N_8880,N_8257,N_8196);
nor U8881 (N_8881,N_8200,N_8195);
nor U8882 (N_8882,N_8023,N_8406);
or U8883 (N_8883,N_8386,N_8107);
nand U8884 (N_8884,N_8117,N_8114);
and U8885 (N_8885,N_8472,N_8132);
xor U8886 (N_8886,N_8219,N_8086);
nor U8887 (N_8887,N_8441,N_8267);
and U8888 (N_8888,N_8334,N_8437);
nand U8889 (N_8889,N_8076,N_8052);
nand U8890 (N_8890,N_8359,N_8295);
nor U8891 (N_8891,N_8437,N_8189);
or U8892 (N_8892,N_8133,N_8223);
nor U8893 (N_8893,N_8203,N_8030);
nor U8894 (N_8894,N_8023,N_8234);
nand U8895 (N_8895,N_8112,N_8226);
and U8896 (N_8896,N_8237,N_8135);
and U8897 (N_8897,N_8349,N_8318);
nand U8898 (N_8898,N_8357,N_8150);
xnor U8899 (N_8899,N_8274,N_8391);
and U8900 (N_8900,N_8103,N_8098);
xor U8901 (N_8901,N_8006,N_8367);
and U8902 (N_8902,N_8126,N_8005);
nor U8903 (N_8903,N_8409,N_8176);
nand U8904 (N_8904,N_8481,N_8396);
and U8905 (N_8905,N_8151,N_8407);
and U8906 (N_8906,N_8409,N_8411);
and U8907 (N_8907,N_8085,N_8341);
or U8908 (N_8908,N_8349,N_8303);
nor U8909 (N_8909,N_8079,N_8209);
or U8910 (N_8910,N_8230,N_8272);
and U8911 (N_8911,N_8438,N_8082);
and U8912 (N_8912,N_8324,N_8381);
nand U8913 (N_8913,N_8000,N_8018);
xor U8914 (N_8914,N_8220,N_8155);
and U8915 (N_8915,N_8294,N_8171);
nand U8916 (N_8916,N_8082,N_8379);
and U8917 (N_8917,N_8213,N_8377);
and U8918 (N_8918,N_8289,N_8401);
nand U8919 (N_8919,N_8422,N_8065);
nand U8920 (N_8920,N_8472,N_8348);
or U8921 (N_8921,N_8165,N_8145);
or U8922 (N_8922,N_8083,N_8266);
or U8923 (N_8923,N_8347,N_8254);
nand U8924 (N_8924,N_8257,N_8062);
xor U8925 (N_8925,N_8083,N_8121);
nor U8926 (N_8926,N_8310,N_8435);
and U8927 (N_8927,N_8044,N_8014);
or U8928 (N_8928,N_8197,N_8291);
nand U8929 (N_8929,N_8053,N_8425);
nor U8930 (N_8930,N_8081,N_8276);
and U8931 (N_8931,N_8097,N_8205);
and U8932 (N_8932,N_8322,N_8456);
xnor U8933 (N_8933,N_8049,N_8197);
xor U8934 (N_8934,N_8430,N_8242);
xnor U8935 (N_8935,N_8274,N_8291);
nor U8936 (N_8936,N_8059,N_8355);
and U8937 (N_8937,N_8203,N_8002);
nor U8938 (N_8938,N_8423,N_8308);
or U8939 (N_8939,N_8412,N_8005);
nor U8940 (N_8940,N_8338,N_8355);
or U8941 (N_8941,N_8330,N_8413);
nor U8942 (N_8942,N_8105,N_8161);
xor U8943 (N_8943,N_8330,N_8433);
nor U8944 (N_8944,N_8159,N_8446);
or U8945 (N_8945,N_8233,N_8014);
nand U8946 (N_8946,N_8310,N_8063);
xnor U8947 (N_8947,N_8016,N_8191);
or U8948 (N_8948,N_8090,N_8452);
nor U8949 (N_8949,N_8354,N_8367);
nor U8950 (N_8950,N_8468,N_8267);
nor U8951 (N_8951,N_8288,N_8230);
nand U8952 (N_8952,N_8329,N_8492);
or U8953 (N_8953,N_8137,N_8139);
and U8954 (N_8954,N_8496,N_8108);
and U8955 (N_8955,N_8100,N_8292);
nor U8956 (N_8956,N_8266,N_8467);
or U8957 (N_8957,N_8056,N_8495);
xor U8958 (N_8958,N_8120,N_8225);
nand U8959 (N_8959,N_8260,N_8255);
and U8960 (N_8960,N_8365,N_8006);
nand U8961 (N_8961,N_8015,N_8231);
nor U8962 (N_8962,N_8286,N_8178);
xor U8963 (N_8963,N_8221,N_8019);
or U8964 (N_8964,N_8300,N_8066);
or U8965 (N_8965,N_8075,N_8489);
nor U8966 (N_8966,N_8082,N_8041);
or U8967 (N_8967,N_8024,N_8407);
nand U8968 (N_8968,N_8034,N_8315);
xnor U8969 (N_8969,N_8183,N_8022);
or U8970 (N_8970,N_8015,N_8081);
and U8971 (N_8971,N_8348,N_8073);
or U8972 (N_8972,N_8350,N_8335);
nor U8973 (N_8973,N_8205,N_8086);
nor U8974 (N_8974,N_8416,N_8278);
nand U8975 (N_8975,N_8415,N_8058);
nor U8976 (N_8976,N_8001,N_8287);
xor U8977 (N_8977,N_8023,N_8461);
nor U8978 (N_8978,N_8370,N_8482);
nand U8979 (N_8979,N_8199,N_8453);
or U8980 (N_8980,N_8357,N_8338);
nand U8981 (N_8981,N_8459,N_8223);
nor U8982 (N_8982,N_8028,N_8448);
and U8983 (N_8983,N_8469,N_8092);
or U8984 (N_8984,N_8305,N_8062);
nor U8985 (N_8985,N_8269,N_8342);
nor U8986 (N_8986,N_8404,N_8044);
or U8987 (N_8987,N_8137,N_8114);
and U8988 (N_8988,N_8040,N_8453);
xor U8989 (N_8989,N_8260,N_8264);
nor U8990 (N_8990,N_8138,N_8013);
and U8991 (N_8991,N_8014,N_8065);
nor U8992 (N_8992,N_8318,N_8460);
xor U8993 (N_8993,N_8170,N_8463);
nand U8994 (N_8994,N_8239,N_8034);
nor U8995 (N_8995,N_8439,N_8136);
nand U8996 (N_8996,N_8344,N_8009);
nand U8997 (N_8997,N_8102,N_8329);
nand U8998 (N_8998,N_8212,N_8035);
nor U8999 (N_8999,N_8251,N_8026);
nor U9000 (N_9000,N_8653,N_8710);
nand U9001 (N_9001,N_8905,N_8551);
nor U9002 (N_9002,N_8729,N_8610);
and U9003 (N_9003,N_8921,N_8867);
or U9004 (N_9004,N_8901,N_8606);
nand U9005 (N_9005,N_8812,N_8709);
nand U9006 (N_9006,N_8937,N_8603);
or U9007 (N_9007,N_8739,N_8547);
nor U9008 (N_9008,N_8839,N_8783);
and U9009 (N_9009,N_8635,N_8553);
or U9010 (N_9010,N_8652,N_8507);
nand U9011 (N_9011,N_8827,N_8963);
and U9012 (N_9012,N_8885,N_8503);
or U9013 (N_9013,N_8585,N_8773);
nand U9014 (N_9014,N_8855,N_8616);
or U9015 (N_9015,N_8985,N_8707);
nand U9016 (N_9016,N_8966,N_8968);
nor U9017 (N_9017,N_8776,N_8928);
and U9018 (N_9018,N_8557,N_8645);
and U9019 (N_9019,N_8613,N_8756);
nand U9020 (N_9020,N_8667,N_8854);
nand U9021 (N_9021,N_8987,N_8774);
or U9022 (N_9022,N_8722,N_8740);
xor U9023 (N_9023,N_8681,N_8676);
nand U9024 (N_9024,N_8835,N_8903);
or U9025 (N_9025,N_8989,N_8902);
nand U9026 (N_9026,N_8777,N_8831);
and U9027 (N_9027,N_8759,N_8699);
and U9028 (N_9028,N_8986,N_8952);
and U9029 (N_9029,N_8724,N_8510);
nand U9030 (N_9030,N_8581,N_8520);
and U9031 (N_9031,N_8723,N_8964);
nand U9032 (N_9032,N_8801,N_8809);
nand U9033 (N_9033,N_8786,N_8823);
xor U9034 (N_9034,N_8675,N_8691);
xnor U9035 (N_9035,N_8999,N_8755);
and U9036 (N_9036,N_8663,N_8982);
or U9037 (N_9037,N_8798,N_8869);
or U9038 (N_9038,N_8758,N_8925);
nand U9039 (N_9039,N_8910,N_8993);
xor U9040 (N_9040,N_8832,N_8920);
or U9041 (N_9041,N_8788,N_8545);
nand U9042 (N_9042,N_8769,N_8589);
nand U9043 (N_9043,N_8778,N_8829);
or U9044 (N_9044,N_8536,N_8518);
nor U9045 (N_9045,N_8543,N_8959);
nand U9046 (N_9046,N_8706,N_8608);
or U9047 (N_9047,N_8945,N_8612);
or U9048 (N_9048,N_8671,N_8978);
or U9049 (N_9049,N_8747,N_8844);
and U9050 (N_9050,N_8666,N_8697);
nor U9051 (N_9051,N_8750,N_8926);
xor U9052 (N_9052,N_8672,N_8833);
xnor U9053 (N_9053,N_8601,N_8524);
or U9054 (N_9054,N_8841,N_8836);
or U9055 (N_9055,N_8741,N_8872);
or U9056 (N_9056,N_8717,N_8745);
nand U9057 (N_9057,N_8818,N_8538);
and U9058 (N_9058,N_8935,N_8568);
nor U9059 (N_9059,N_8884,N_8554);
or U9060 (N_9060,N_8719,N_8701);
xnor U9061 (N_9061,N_8864,N_8771);
or U9062 (N_9062,N_8513,N_8587);
nand U9063 (N_9063,N_8757,N_8834);
nor U9064 (N_9064,N_8641,N_8782);
xnor U9065 (N_9065,N_8743,N_8787);
nor U9066 (N_9066,N_8849,N_8842);
and U9067 (N_9067,N_8916,N_8947);
nand U9068 (N_9068,N_8875,N_8821);
nor U9069 (N_9069,N_8584,N_8811);
or U9070 (N_9070,N_8772,N_8651);
and U9071 (N_9071,N_8860,N_8644);
nor U9072 (N_9072,N_8648,N_8873);
and U9073 (N_9073,N_8542,N_8992);
or U9074 (N_9074,N_8768,N_8522);
and U9075 (N_9075,N_8898,N_8752);
and U9076 (N_9076,N_8857,N_8970);
nor U9077 (N_9077,N_8558,N_8620);
nand U9078 (N_9078,N_8814,N_8725);
nor U9079 (N_9079,N_8679,N_8907);
nand U9080 (N_9080,N_8838,N_8689);
and U9081 (N_9081,N_8871,N_8617);
and U9082 (N_9082,N_8575,N_8767);
nor U9083 (N_9083,N_8586,N_8735);
xor U9084 (N_9084,N_8662,N_8677);
and U9085 (N_9085,N_8591,N_8887);
nand U9086 (N_9086,N_8983,N_8929);
xor U9087 (N_9087,N_8577,N_8944);
xnor U9088 (N_9088,N_8933,N_8540);
nand U9089 (N_9089,N_8861,N_8628);
nor U9090 (N_9090,N_8847,N_8807);
nand U9091 (N_9091,N_8618,N_8850);
nor U9092 (N_9092,N_8880,N_8523);
nand U9093 (N_9093,N_8649,N_8828);
nor U9094 (N_9094,N_8563,N_8891);
nand U9095 (N_9095,N_8664,N_8670);
nand U9096 (N_9096,N_8700,N_8981);
and U9097 (N_9097,N_8996,N_8712);
and U9098 (N_9098,N_8715,N_8537);
nor U9099 (N_9099,N_8539,N_8684);
xnor U9100 (N_9100,N_8728,N_8962);
or U9101 (N_9101,N_8848,N_8639);
nand U9102 (N_9102,N_8923,N_8549);
nor U9103 (N_9103,N_8636,N_8550);
nand U9104 (N_9104,N_8938,N_8760);
or U9105 (N_9105,N_8734,N_8846);
nor U9106 (N_9106,N_8797,N_8882);
or U9107 (N_9107,N_8804,N_8780);
nor U9108 (N_9108,N_8569,N_8504);
nor U9109 (N_9109,N_8973,N_8961);
and U9110 (N_9110,N_8535,N_8730);
and U9111 (N_9111,N_8896,N_8845);
and U9112 (N_9112,N_8599,N_8718);
nor U9113 (N_9113,N_8781,N_8856);
xnor U9114 (N_9114,N_8749,N_8622);
nor U9115 (N_9115,N_8683,N_8806);
nor U9116 (N_9116,N_8605,N_8727);
nand U9117 (N_9117,N_8704,N_8655);
nand U9118 (N_9118,N_8816,N_8579);
xnor U9119 (N_9119,N_8544,N_8826);
and U9120 (N_9120,N_8592,N_8866);
nand U9121 (N_9121,N_8531,N_8794);
nor U9122 (N_9122,N_8853,N_8934);
and U9123 (N_9123,N_8858,N_8795);
or U9124 (N_9124,N_8659,N_8556);
or U9125 (N_9125,N_8517,N_8562);
xor U9126 (N_9126,N_8576,N_8611);
xor U9127 (N_9127,N_8703,N_8874);
or U9128 (N_9128,N_8643,N_8879);
nand U9129 (N_9129,N_8984,N_8865);
nor U9130 (N_9130,N_8516,N_8694);
nor U9131 (N_9131,N_8696,N_8897);
and U9132 (N_9132,N_8682,N_8878);
and U9133 (N_9133,N_8505,N_8590);
nor U9134 (N_9134,N_8530,N_8908);
or U9135 (N_9135,N_8802,N_8762);
nand U9136 (N_9136,N_8955,N_8566);
or U9137 (N_9137,N_8693,N_8990);
nor U9138 (N_9138,N_8813,N_8702);
and U9139 (N_9139,N_8660,N_8843);
and U9140 (N_9140,N_8500,N_8790);
nor U9141 (N_9141,N_8650,N_8571);
nand U9142 (N_9142,N_8930,N_8748);
nor U9143 (N_9143,N_8669,N_8889);
or U9144 (N_9144,N_8979,N_8789);
or U9145 (N_9145,N_8936,N_8830);
nor U9146 (N_9146,N_8917,N_8570);
or U9147 (N_9147,N_8997,N_8692);
or U9148 (N_9148,N_8940,N_8764);
and U9149 (N_9149,N_8596,N_8956);
nand U9150 (N_9150,N_8942,N_8559);
nor U9151 (N_9151,N_8609,N_8588);
nor U9152 (N_9152,N_8506,N_8567);
or U9153 (N_9153,N_8892,N_8761);
and U9154 (N_9154,N_8792,N_8711);
nand U9155 (N_9155,N_8615,N_8746);
nand U9156 (N_9156,N_8852,N_8600);
or U9157 (N_9157,N_8863,N_8817);
or U9158 (N_9158,N_8883,N_8915);
or U9159 (N_9159,N_8526,N_8533);
nand U9160 (N_9160,N_8766,N_8751);
or U9161 (N_9161,N_8619,N_8661);
or U9162 (N_9162,N_8890,N_8733);
and U9163 (N_9163,N_8726,N_8647);
nor U9164 (N_9164,N_8580,N_8980);
and U9165 (N_9165,N_8509,N_8939);
and U9166 (N_9166,N_8595,N_8919);
or U9167 (N_9167,N_8674,N_8560);
nor U9168 (N_9168,N_8950,N_8627);
and U9169 (N_9169,N_8574,N_8824);
and U9170 (N_9170,N_8770,N_8582);
and U9171 (N_9171,N_8913,N_8895);
and U9172 (N_9172,N_8656,N_8573);
and U9173 (N_9173,N_8779,N_8698);
xnor U9174 (N_9174,N_8607,N_8604);
or U9175 (N_9175,N_8911,N_8529);
nand U9176 (N_9176,N_8753,N_8803);
or U9177 (N_9177,N_8521,N_8972);
nor U9178 (N_9178,N_8565,N_8991);
and U9179 (N_9179,N_8965,N_8909);
xnor U9180 (N_9180,N_8995,N_8953);
nor U9181 (N_9181,N_8501,N_8548);
or U9182 (N_9182,N_8738,N_8528);
nand U9183 (N_9183,N_8971,N_8646);
nor U9184 (N_9184,N_8881,N_8918);
nand U9185 (N_9185,N_8754,N_8893);
nor U9186 (N_9186,N_8825,N_8862);
or U9187 (N_9187,N_8927,N_8624);
and U9188 (N_9188,N_8720,N_8633);
or U9189 (N_9189,N_8578,N_8736);
nand U9190 (N_9190,N_8763,N_8638);
or U9191 (N_9191,N_8793,N_8904);
and U9192 (N_9192,N_8888,N_8931);
nor U9193 (N_9193,N_8555,N_8688);
and U9194 (N_9194,N_8631,N_8868);
or U9195 (N_9195,N_8687,N_8714);
nand U9196 (N_9196,N_8658,N_8541);
nor U9197 (N_9197,N_8532,N_8784);
nor U9198 (N_9198,N_8716,N_8886);
or U9199 (N_9199,N_8808,N_8690);
xor U9200 (N_9200,N_8791,N_8975);
nor U9201 (N_9201,N_8597,N_8899);
nand U9202 (N_9202,N_8994,N_8977);
and U9203 (N_9203,N_8906,N_8508);
or U9204 (N_9204,N_8642,N_8998);
and U9205 (N_9205,N_8870,N_8598);
and U9206 (N_9206,N_8796,N_8900);
xor U9207 (N_9207,N_8851,N_8810);
or U9208 (N_9208,N_8960,N_8625);
and U9209 (N_9209,N_8958,N_8695);
or U9210 (N_9210,N_8837,N_8922);
and U9211 (N_9211,N_8737,N_8512);
xnor U9212 (N_9212,N_8988,N_8775);
nor U9213 (N_9213,N_8534,N_8686);
nor U9214 (N_9214,N_8914,N_8621);
and U9215 (N_9215,N_8954,N_8583);
xor U9216 (N_9216,N_8614,N_8859);
and U9217 (N_9217,N_8941,N_8665);
or U9218 (N_9218,N_8502,N_8765);
and U9219 (N_9219,N_8800,N_8572);
and U9220 (N_9220,N_8546,N_8912);
or U9221 (N_9221,N_8820,N_8876);
and U9222 (N_9222,N_8630,N_8623);
nand U9223 (N_9223,N_8721,N_8974);
and U9224 (N_9224,N_8819,N_8564);
or U9225 (N_9225,N_8969,N_8976);
nand U9226 (N_9226,N_8593,N_8561);
or U9227 (N_9227,N_8822,N_8894);
nor U9228 (N_9228,N_8744,N_8680);
and U9229 (N_9229,N_8629,N_8948);
and U9230 (N_9230,N_8626,N_8668);
nor U9231 (N_9231,N_8525,N_8840);
and U9232 (N_9232,N_8949,N_8640);
and U9233 (N_9233,N_8708,N_8637);
nor U9234 (N_9234,N_8731,N_8732);
or U9235 (N_9235,N_8515,N_8946);
xor U9236 (N_9236,N_8742,N_8657);
nand U9237 (N_9237,N_8519,N_8713);
nand U9238 (N_9238,N_8967,N_8815);
nand U9239 (N_9239,N_8527,N_8785);
nand U9240 (N_9240,N_8951,N_8514);
or U9241 (N_9241,N_8632,N_8877);
or U9242 (N_9242,N_8552,N_8799);
nor U9243 (N_9243,N_8634,N_8805);
nor U9244 (N_9244,N_8943,N_8654);
or U9245 (N_9245,N_8678,N_8511);
nand U9246 (N_9246,N_8705,N_8957);
nand U9247 (N_9247,N_8932,N_8594);
or U9248 (N_9248,N_8673,N_8685);
nand U9249 (N_9249,N_8924,N_8602);
and U9250 (N_9250,N_8780,N_8664);
nor U9251 (N_9251,N_8923,N_8924);
nor U9252 (N_9252,N_8874,N_8716);
or U9253 (N_9253,N_8976,N_8955);
nand U9254 (N_9254,N_8583,N_8955);
or U9255 (N_9255,N_8869,N_8641);
and U9256 (N_9256,N_8890,N_8893);
and U9257 (N_9257,N_8952,N_8935);
nor U9258 (N_9258,N_8679,N_8602);
nand U9259 (N_9259,N_8651,N_8952);
and U9260 (N_9260,N_8927,N_8796);
nand U9261 (N_9261,N_8654,N_8861);
nor U9262 (N_9262,N_8718,N_8723);
nor U9263 (N_9263,N_8877,N_8717);
nor U9264 (N_9264,N_8736,N_8648);
or U9265 (N_9265,N_8500,N_8739);
nand U9266 (N_9266,N_8922,N_8750);
or U9267 (N_9267,N_8627,N_8974);
or U9268 (N_9268,N_8811,N_8609);
or U9269 (N_9269,N_8959,N_8761);
nor U9270 (N_9270,N_8944,N_8896);
or U9271 (N_9271,N_8953,N_8797);
nand U9272 (N_9272,N_8702,N_8918);
nand U9273 (N_9273,N_8579,N_8952);
nor U9274 (N_9274,N_8505,N_8907);
and U9275 (N_9275,N_8895,N_8659);
or U9276 (N_9276,N_8778,N_8825);
and U9277 (N_9277,N_8637,N_8999);
or U9278 (N_9278,N_8533,N_8849);
or U9279 (N_9279,N_8824,N_8914);
nor U9280 (N_9280,N_8638,N_8624);
and U9281 (N_9281,N_8904,N_8993);
nand U9282 (N_9282,N_8631,N_8675);
xnor U9283 (N_9283,N_8762,N_8892);
or U9284 (N_9284,N_8578,N_8775);
and U9285 (N_9285,N_8529,N_8839);
or U9286 (N_9286,N_8761,N_8685);
nor U9287 (N_9287,N_8849,N_8982);
nand U9288 (N_9288,N_8938,N_8543);
xnor U9289 (N_9289,N_8840,N_8951);
and U9290 (N_9290,N_8596,N_8849);
nor U9291 (N_9291,N_8781,N_8597);
or U9292 (N_9292,N_8600,N_8593);
or U9293 (N_9293,N_8935,N_8529);
nor U9294 (N_9294,N_8612,N_8532);
nand U9295 (N_9295,N_8938,N_8644);
and U9296 (N_9296,N_8811,N_8654);
xnor U9297 (N_9297,N_8901,N_8604);
or U9298 (N_9298,N_8759,N_8533);
nor U9299 (N_9299,N_8731,N_8943);
nor U9300 (N_9300,N_8598,N_8718);
nand U9301 (N_9301,N_8903,N_8682);
or U9302 (N_9302,N_8968,N_8925);
nor U9303 (N_9303,N_8830,N_8957);
xnor U9304 (N_9304,N_8992,N_8802);
xor U9305 (N_9305,N_8637,N_8633);
xnor U9306 (N_9306,N_8655,N_8793);
and U9307 (N_9307,N_8848,N_8851);
or U9308 (N_9308,N_8985,N_8732);
and U9309 (N_9309,N_8723,N_8898);
or U9310 (N_9310,N_8727,N_8980);
nor U9311 (N_9311,N_8820,N_8616);
or U9312 (N_9312,N_8815,N_8631);
or U9313 (N_9313,N_8789,N_8990);
nor U9314 (N_9314,N_8870,N_8608);
nor U9315 (N_9315,N_8799,N_8760);
or U9316 (N_9316,N_8598,N_8820);
nor U9317 (N_9317,N_8671,N_8630);
or U9318 (N_9318,N_8867,N_8725);
nand U9319 (N_9319,N_8593,N_8799);
xor U9320 (N_9320,N_8714,N_8627);
or U9321 (N_9321,N_8588,N_8885);
nand U9322 (N_9322,N_8501,N_8646);
nor U9323 (N_9323,N_8956,N_8953);
or U9324 (N_9324,N_8824,N_8561);
nor U9325 (N_9325,N_8992,N_8826);
nor U9326 (N_9326,N_8751,N_8528);
or U9327 (N_9327,N_8751,N_8671);
nand U9328 (N_9328,N_8888,N_8994);
or U9329 (N_9329,N_8620,N_8738);
nor U9330 (N_9330,N_8911,N_8919);
or U9331 (N_9331,N_8554,N_8667);
nand U9332 (N_9332,N_8915,N_8878);
nor U9333 (N_9333,N_8893,N_8978);
or U9334 (N_9334,N_8702,N_8993);
nand U9335 (N_9335,N_8834,N_8674);
and U9336 (N_9336,N_8767,N_8510);
nand U9337 (N_9337,N_8933,N_8615);
nand U9338 (N_9338,N_8934,N_8817);
nor U9339 (N_9339,N_8941,N_8885);
or U9340 (N_9340,N_8861,N_8976);
xnor U9341 (N_9341,N_8998,N_8993);
or U9342 (N_9342,N_8990,N_8950);
nand U9343 (N_9343,N_8989,N_8869);
and U9344 (N_9344,N_8841,N_8773);
nor U9345 (N_9345,N_8737,N_8666);
nor U9346 (N_9346,N_8639,N_8757);
or U9347 (N_9347,N_8616,N_8608);
or U9348 (N_9348,N_8599,N_8782);
xnor U9349 (N_9349,N_8850,N_8986);
nand U9350 (N_9350,N_8599,N_8546);
nand U9351 (N_9351,N_8890,N_8655);
nand U9352 (N_9352,N_8978,N_8628);
nor U9353 (N_9353,N_8585,N_8650);
nand U9354 (N_9354,N_8669,N_8625);
and U9355 (N_9355,N_8972,N_8533);
and U9356 (N_9356,N_8636,N_8632);
nand U9357 (N_9357,N_8667,N_8986);
nand U9358 (N_9358,N_8896,N_8633);
and U9359 (N_9359,N_8684,N_8976);
or U9360 (N_9360,N_8761,N_8543);
or U9361 (N_9361,N_8768,N_8739);
or U9362 (N_9362,N_8571,N_8530);
nand U9363 (N_9363,N_8696,N_8589);
or U9364 (N_9364,N_8692,N_8660);
nand U9365 (N_9365,N_8754,N_8519);
nand U9366 (N_9366,N_8609,N_8672);
xor U9367 (N_9367,N_8701,N_8754);
xor U9368 (N_9368,N_8742,N_8594);
nor U9369 (N_9369,N_8919,N_8529);
nor U9370 (N_9370,N_8785,N_8516);
and U9371 (N_9371,N_8809,N_8647);
or U9372 (N_9372,N_8730,N_8765);
nor U9373 (N_9373,N_8787,N_8966);
nor U9374 (N_9374,N_8623,N_8667);
and U9375 (N_9375,N_8826,N_8912);
or U9376 (N_9376,N_8870,N_8768);
and U9377 (N_9377,N_8576,N_8939);
nor U9378 (N_9378,N_8833,N_8645);
nand U9379 (N_9379,N_8894,N_8562);
and U9380 (N_9380,N_8891,N_8530);
nand U9381 (N_9381,N_8611,N_8997);
xnor U9382 (N_9382,N_8912,N_8765);
nor U9383 (N_9383,N_8953,N_8862);
nor U9384 (N_9384,N_8913,N_8789);
nor U9385 (N_9385,N_8582,N_8503);
nand U9386 (N_9386,N_8839,N_8577);
and U9387 (N_9387,N_8784,N_8824);
and U9388 (N_9388,N_8963,N_8509);
xnor U9389 (N_9389,N_8536,N_8598);
nand U9390 (N_9390,N_8846,N_8816);
nor U9391 (N_9391,N_8790,N_8738);
nand U9392 (N_9392,N_8992,N_8526);
or U9393 (N_9393,N_8679,N_8934);
nor U9394 (N_9394,N_8758,N_8837);
xnor U9395 (N_9395,N_8986,N_8605);
or U9396 (N_9396,N_8664,N_8975);
and U9397 (N_9397,N_8534,N_8829);
nor U9398 (N_9398,N_8822,N_8827);
xor U9399 (N_9399,N_8502,N_8603);
and U9400 (N_9400,N_8694,N_8542);
nor U9401 (N_9401,N_8681,N_8563);
or U9402 (N_9402,N_8981,N_8524);
and U9403 (N_9403,N_8976,N_8679);
nor U9404 (N_9404,N_8624,N_8677);
nor U9405 (N_9405,N_8636,N_8914);
nand U9406 (N_9406,N_8776,N_8851);
or U9407 (N_9407,N_8594,N_8837);
and U9408 (N_9408,N_8662,N_8881);
nand U9409 (N_9409,N_8642,N_8545);
nand U9410 (N_9410,N_8643,N_8795);
and U9411 (N_9411,N_8731,N_8955);
xor U9412 (N_9412,N_8910,N_8637);
nand U9413 (N_9413,N_8880,N_8658);
or U9414 (N_9414,N_8966,N_8833);
and U9415 (N_9415,N_8606,N_8685);
or U9416 (N_9416,N_8900,N_8960);
nand U9417 (N_9417,N_8548,N_8791);
nor U9418 (N_9418,N_8995,N_8895);
and U9419 (N_9419,N_8662,N_8684);
nor U9420 (N_9420,N_8506,N_8831);
and U9421 (N_9421,N_8852,N_8637);
or U9422 (N_9422,N_8682,N_8792);
nand U9423 (N_9423,N_8890,N_8762);
and U9424 (N_9424,N_8998,N_8767);
nand U9425 (N_9425,N_8833,N_8546);
nor U9426 (N_9426,N_8625,N_8534);
nor U9427 (N_9427,N_8883,N_8628);
nand U9428 (N_9428,N_8874,N_8685);
nand U9429 (N_9429,N_8668,N_8893);
nand U9430 (N_9430,N_8915,N_8575);
nand U9431 (N_9431,N_8899,N_8763);
nor U9432 (N_9432,N_8572,N_8552);
nor U9433 (N_9433,N_8564,N_8629);
nor U9434 (N_9434,N_8949,N_8621);
and U9435 (N_9435,N_8852,N_8684);
nor U9436 (N_9436,N_8668,N_8843);
nand U9437 (N_9437,N_8890,N_8980);
nand U9438 (N_9438,N_8948,N_8558);
nand U9439 (N_9439,N_8927,N_8993);
and U9440 (N_9440,N_8594,N_8936);
or U9441 (N_9441,N_8503,N_8720);
or U9442 (N_9442,N_8724,N_8719);
nor U9443 (N_9443,N_8756,N_8831);
or U9444 (N_9444,N_8920,N_8525);
nor U9445 (N_9445,N_8913,N_8905);
or U9446 (N_9446,N_8973,N_8782);
nor U9447 (N_9447,N_8753,N_8644);
xnor U9448 (N_9448,N_8844,N_8551);
xor U9449 (N_9449,N_8518,N_8805);
and U9450 (N_9450,N_8513,N_8961);
nor U9451 (N_9451,N_8555,N_8662);
and U9452 (N_9452,N_8540,N_8874);
or U9453 (N_9453,N_8713,N_8865);
nor U9454 (N_9454,N_8664,N_8741);
and U9455 (N_9455,N_8811,N_8540);
xor U9456 (N_9456,N_8625,N_8676);
and U9457 (N_9457,N_8509,N_8597);
nor U9458 (N_9458,N_8841,N_8732);
nand U9459 (N_9459,N_8724,N_8701);
or U9460 (N_9460,N_8893,N_8671);
nor U9461 (N_9461,N_8581,N_8941);
nand U9462 (N_9462,N_8634,N_8629);
and U9463 (N_9463,N_8850,N_8880);
xor U9464 (N_9464,N_8646,N_8685);
nand U9465 (N_9465,N_8986,N_8870);
nor U9466 (N_9466,N_8513,N_8548);
nand U9467 (N_9467,N_8976,N_8843);
and U9468 (N_9468,N_8974,N_8763);
nor U9469 (N_9469,N_8973,N_8639);
or U9470 (N_9470,N_8791,N_8820);
or U9471 (N_9471,N_8513,N_8781);
and U9472 (N_9472,N_8698,N_8781);
nor U9473 (N_9473,N_8835,N_8737);
or U9474 (N_9474,N_8677,N_8631);
or U9475 (N_9475,N_8527,N_8612);
nor U9476 (N_9476,N_8933,N_8762);
and U9477 (N_9477,N_8618,N_8605);
nor U9478 (N_9478,N_8741,N_8936);
nor U9479 (N_9479,N_8677,N_8690);
nor U9480 (N_9480,N_8964,N_8763);
and U9481 (N_9481,N_8516,N_8797);
xor U9482 (N_9482,N_8643,N_8928);
xor U9483 (N_9483,N_8970,N_8527);
or U9484 (N_9484,N_8800,N_8696);
and U9485 (N_9485,N_8550,N_8693);
nor U9486 (N_9486,N_8800,N_8901);
or U9487 (N_9487,N_8671,N_8631);
xnor U9488 (N_9488,N_8646,N_8586);
and U9489 (N_9489,N_8634,N_8771);
xnor U9490 (N_9490,N_8919,N_8741);
nor U9491 (N_9491,N_8609,N_8743);
nand U9492 (N_9492,N_8618,N_8872);
nand U9493 (N_9493,N_8677,N_8563);
nor U9494 (N_9494,N_8820,N_8715);
and U9495 (N_9495,N_8732,N_8746);
or U9496 (N_9496,N_8987,N_8507);
or U9497 (N_9497,N_8591,N_8786);
and U9498 (N_9498,N_8771,N_8957);
nand U9499 (N_9499,N_8755,N_8705);
or U9500 (N_9500,N_9043,N_9187);
xor U9501 (N_9501,N_9484,N_9070);
or U9502 (N_9502,N_9065,N_9456);
nor U9503 (N_9503,N_9454,N_9052);
and U9504 (N_9504,N_9087,N_9244);
nor U9505 (N_9505,N_9428,N_9222);
nor U9506 (N_9506,N_9108,N_9316);
and U9507 (N_9507,N_9372,N_9083);
nand U9508 (N_9508,N_9285,N_9447);
and U9509 (N_9509,N_9166,N_9129);
nand U9510 (N_9510,N_9127,N_9443);
nand U9511 (N_9511,N_9079,N_9201);
nand U9512 (N_9512,N_9377,N_9136);
nor U9513 (N_9513,N_9106,N_9220);
or U9514 (N_9514,N_9380,N_9469);
nand U9515 (N_9515,N_9286,N_9418);
nand U9516 (N_9516,N_9100,N_9496);
or U9517 (N_9517,N_9348,N_9085);
nor U9518 (N_9518,N_9210,N_9322);
or U9519 (N_9519,N_9088,N_9384);
nand U9520 (N_9520,N_9074,N_9152);
or U9521 (N_9521,N_9261,N_9373);
nand U9522 (N_9522,N_9331,N_9343);
nor U9523 (N_9523,N_9122,N_9440);
nor U9524 (N_9524,N_9059,N_9304);
nor U9525 (N_9525,N_9361,N_9207);
nand U9526 (N_9526,N_9271,N_9360);
and U9527 (N_9527,N_9481,N_9444);
or U9528 (N_9528,N_9280,N_9057);
nand U9529 (N_9529,N_9036,N_9368);
and U9530 (N_9530,N_9091,N_9296);
and U9531 (N_9531,N_9457,N_9367);
or U9532 (N_9532,N_9072,N_9090);
or U9533 (N_9533,N_9451,N_9247);
xor U9534 (N_9534,N_9149,N_9097);
nand U9535 (N_9535,N_9064,N_9270);
or U9536 (N_9536,N_9199,N_9061);
or U9537 (N_9537,N_9268,N_9459);
nor U9538 (N_9538,N_9303,N_9370);
xor U9539 (N_9539,N_9465,N_9204);
nor U9540 (N_9540,N_9463,N_9333);
nor U9541 (N_9541,N_9308,N_9223);
or U9542 (N_9542,N_9235,N_9158);
and U9543 (N_9543,N_9412,N_9144);
and U9544 (N_9544,N_9362,N_9089);
or U9545 (N_9545,N_9111,N_9030);
nor U9546 (N_9546,N_9278,N_9300);
and U9547 (N_9547,N_9497,N_9432);
and U9548 (N_9548,N_9336,N_9117);
nor U9549 (N_9549,N_9458,N_9422);
or U9550 (N_9550,N_9125,N_9265);
nor U9551 (N_9551,N_9212,N_9374);
nand U9552 (N_9552,N_9453,N_9231);
or U9553 (N_9553,N_9021,N_9234);
nand U9554 (N_9554,N_9040,N_9442);
and U9555 (N_9555,N_9340,N_9134);
nand U9556 (N_9556,N_9116,N_9033);
or U9557 (N_9557,N_9239,N_9104);
xnor U9558 (N_9558,N_9046,N_9312);
xor U9559 (N_9559,N_9275,N_9225);
or U9560 (N_9560,N_9494,N_9081);
nand U9561 (N_9561,N_9148,N_9181);
xnor U9562 (N_9562,N_9366,N_9473);
xor U9563 (N_9563,N_9172,N_9138);
and U9564 (N_9564,N_9365,N_9450);
or U9565 (N_9565,N_9405,N_9128);
xnor U9566 (N_9566,N_9363,N_9485);
or U9567 (N_9567,N_9179,N_9337);
nand U9568 (N_9568,N_9185,N_9335);
nor U9569 (N_9569,N_9154,N_9311);
xnor U9570 (N_9570,N_9407,N_9173);
nor U9571 (N_9571,N_9137,N_9119);
and U9572 (N_9572,N_9262,N_9479);
nand U9573 (N_9573,N_9398,N_9283);
and U9574 (N_9574,N_9039,N_9215);
or U9575 (N_9575,N_9486,N_9395);
and U9576 (N_9576,N_9062,N_9288);
nor U9577 (N_9577,N_9013,N_9216);
nor U9578 (N_9578,N_9324,N_9147);
nor U9579 (N_9579,N_9017,N_9411);
nor U9580 (N_9580,N_9175,N_9320);
or U9581 (N_9581,N_9048,N_9240);
nor U9582 (N_9582,N_9402,N_9047);
nand U9583 (N_9583,N_9256,N_9103);
or U9584 (N_9584,N_9291,N_9356);
and U9585 (N_9585,N_9272,N_9162);
nand U9586 (N_9586,N_9310,N_9385);
and U9587 (N_9587,N_9421,N_9430);
nand U9588 (N_9588,N_9446,N_9439);
nor U9589 (N_9589,N_9279,N_9161);
nor U9590 (N_9590,N_9050,N_9068);
or U9591 (N_9591,N_9403,N_9196);
nor U9592 (N_9592,N_9396,N_9471);
nand U9593 (N_9593,N_9435,N_9135);
nor U9594 (N_9594,N_9295,N_9153);
nand U9595 (N_9595,N_9429,N_9480);
nand U9596 (N_9596,N_9448,N_9415);
or U9597 (N_9597,N_9474,N_9198);
nor U9598 (N_9598,N_9419,N_9189);
xnor U9599 (N_9599,N_9194,N_9325);
and U9600 (N_9600,N_9101,N_9004);
and U9601 (N_9601,N_9455,N_9159);
nand U9602 (N_9602,N_9150,N_9098);
xnor U9603 (N_9603,N_9404,N_9249);
nand U9604 (N_9604,N_9109,N_9489);
and U9605 (N_9605,N_9358,N_9146);
or U9606 (N_9606,N_9264,N_9206);
nor U9607 (N_9607,N_9330,N_9160);
and U9608 (N_9608,N_9332,N_9002);
nand U9609 (N_9609,N_9130,N_9269);
and U9610 (N_9610,N_9051,N_9254);
and U9611 (N_9611,N_9390,N_9425);
and U9612 (N_9612,N_9301,N_9114);
or U9613 (N_9613,N_9092,N_9309);
xnor U9614 (N_9614,N_9099,N_9164);
nor U9615 (N_9615,N_9339,N_9277);
or U9616 (N_9616,N_9255,N_9259);
nor U9617 (N_9617,N_9214,N_9000);
nor U9618 (N_9618,N_9490,N_9260);
and U9619 (N_9619,N_9477,N_9010);
nor U9620 (N_9620,N_9078,N_9441);
or U9621 (N_9621,N_9008,N_9221);
and U9622 (N_9622,N_9349,N_9184);
nor U9623 (N_9623,N_9094,N_9230);
or U9624 (N_9624,N_9145,N_9468);
or U9625 (N_9625,N_9315,N_9382);
xor U9626 (N_9626,N_9475,N_9007);
nand U9627 (N_9627,N_9139,N_9242);
and U9628 (N_9628,N_9058,N_9218);
nor U9629 (N_9629,N_9203,N_9406);
nor U9630 (N_9630,N_9346,N_9466);
or U9631 (N_9631,N_9491,N_9341);
and U9632 (N_9632,N_9289,N_9276);
xor U9633 (N_9633,N_9393,N_9102);
nand U9634 (N_9634,N_9389,N_9282);
nor U9635 (N_9635,N_9238,N_9041);
and U9636 (N_9636,N_9193,N_9123);
and U9637 (N_9637,N_9056,N_9483);
and U9638 (N_9638,N_9096,N_9488);
and U9639 (N_9639,N_9266,N_9392);
nand U9640 (N_9640,N_9399,N_9355);
nor U9641 (N_9641,N_9375,N_9195);
or U9642 (N_9642,N_9180,N_9076);
or U9643 (N_9643,N_9328,N_9493);
or U9644 (N_9644,N_9258,N_9306);
nand U9645 (N_9645,N_9073,N_9029);
nand U9646 (N_9646,N_9387,N_9003);
nor U9647 (N_9647,N_9470,N_9174);
or U9648 (N_9648,N_9229,N_9131);
nor U9649 (N_9649,N_9274,N_9359);
xor U9650 (N_9650,N_9020,N_9209);
and U9651 (N_9651,N_9257,N_9067);
or U9652 (N_9652,N_9026,N_9250);
and U9653 (N_9653,N_9416,N_9248);
and U9654 (N_9654,N_9314,N_9191);
or U9655 (N_9655,N_9401,N_9121);
nor U9656 (N_9656,N_9434,N_9397);
nor U9657 (N_9657,N_9044,N_9287);
and U9658 (N_9658,N_9213,N_9006);
and U9659 (N_9659,N_9202,N_9351);
or U9660 (N_9660,N_9133,N_9284);
nand U9661 (N_9661,N_9253,N_9156);
or U9662 (N_9662,N_9112,N_9449);
xor U9663 (N_9663,N_9410,N_9027);
or U9664 (N_9664,N_9132,N_9294);
nand U9665 (N_9665,N_9313,N_9001);
nand U9666 (N_9666,N_9177,N_9071);
and U9667 (N_9667,N_9487,N_9298);
xnor U9668 (N_9668,N_9353,N_9031);
nor U9669 (N_9669,N_9431,N_9034);
xor U9670 (N_9670,N_9141,N_9126);
or U9671 (N_9671,N_9053,N_9305);
nand U9672 (N_9672,N_9063,N_9140);
xor U9673 (N_9673,N_9192,N_9424);
or U9674 (N_9674,N_9165,N_9120);
or U9675 (N_9675,N_9472,N_9241);
nor U9676 (N_9676,N_9009,N_9478);
nor U9677 (N_9677,N_9110,N_9438);
or U9678 (N_9678,N_9344,N_9233);
or U9679 (N_9679,N_9200,N_9226);
nor U9680 (N_9680,N_9409,N_9386);
nand U9681 (N_9681,N_9032,N_9232);
nand U9682 (N_9682,N_9095,N_9115);
nor U9683 (N_9683,N_9224,N_9476);
nor U9684 (N_9684,N_9069,N_9299);
or U9685 (N_9685,N_9077,N_9025);
or U9686 (N_9686,N_9037,N_9082);
or U9687 (N_9687,N_9236,N_9016);
nor U9688 (N_9688,N_9042,N_9022);
nand U9689 (N_9689,N_9028,N_9433);
nor U9690 (N_9690,N_9023,N_9197);
or U9691 (N_9691,N_9167,N_9329);
nor U9692 (N_9692,N_9452,N_9376);
and U9693 (N_9693,N_9292,N_9190);
and U9694 (N_9694,N_9075,N_9014);
nor U9695 (N_9695,N_9482,N_9420);
or U9696 (N_9696,N_9391,N_9080);
and U9697 (N_9697,N_9186,N_9267);
and U9698 (N_9698,N_9217,N_9228);
or U9699 (N_9699,N_9263,N_9171);
nand U9700 (N_9700,N_9290,N_9350);
nor U9701 (N_9701,N_9381,N_9105);
or U9702 (N_9702,N_9018,N_9492);
or U9703 (N_9703,N_9281,N_9086);
nor U9704 (N_9704,N_9142,N_9011);
nor U9705 (N_9705,N_9352,N_9205);
and U9706 (N_9706,N_9307,N_9252);
xnor U9707 (N_9707,N_9467,N_9499);
nor U9708 (N_9708,N_9347,N_9155);
and U9709 (N_9709,N_9163,N_9066);
and U9710 (N_9710,N_9445,N_9461);
xnor U9711 (N_9711,N_9113,N_9038);
xor U9712 (N_9712,N_9345,N_9460);
and U9713 (N_9713,N_9055,N_9378);
nand U9714 (N_9714,N_9293,N_9178);
nand U9715 (N_9715,N_9084,N_9334);
or U9716 (N_9716,N_9437,N_9243);
nor U9717 (N_9717,N_9400,N_9024);
or U9718 (N_9718,N_9093,N_9464);
or U9719 (N_9719,N_9157,N_9208);
and U9720 (N_9720,N_9369,N_9182);
or U9721 (N_9721,N_9414,N_9326);
xnor U9722 (N_9722,N_9168,N_9342);
nor U9723 (N_9723,N_9049,N_9423);
nor U9724 (N_9724,N_9327,N_9364);
nor U9725 (N_9725,N_9394,N_9436);
xor U9726 (N_9726,N_9321,N_9408);
xor U9727 (N_9727,N_9319,N_9227);
nor U9728 (N_9728,N_9237,N_9302);
or U9729 (N_9729,N_9151,N_9462);
and U9730 (N_9730,N_9118,N_9246);
nor U9731 (N_9731,N_9045,N_9054);
nor U9732 (N_9732,N_9417,N_9251);
xor U9733 (N_9733,N_9245,N_9338);
or U9734 (N_9734,N_9323,N_9035);
or U9735 (N_9735,N_9005,N_9211);
nand U9736 (N_9736,N_9124,N_9427);
nor U9737 (N_9737,N_9388,N_9357);
and U9738 (N_9738,N_9495,N_9107);
xor U9739 (N_9739,N_9015,N_9379);
and U9740 (N_9740,N_9183,N_9371);
nand U9741 (N_9741,N_9317,N_9219);
nor U9742 (N_9742,N_9297,N_9019);
or U9743 (N_9743,N_9060,N_9318);
and U9744 (N_9744,N_9169,N_9498);
nand U9745 (N_9745,N_9273,N_9176);
nor U9746 (N_9746,N_9354,N_9383);
nor U9747 (N_9747,N_9426,N_9188);
nor U9748 (N_9748,N_9170,N_9012);
or U9749 (N_9749,N_9413,N_9143);
nor U9750 (N_9750,N_9212,N_9028);
or U9751 (N_9751,N_9230,N_9172);
or U9752 (N_9752,N_9142,N_9129);
and U9753 (N_9753,N_9049,N_9086);
nand U9754 (N_9754,N_9245,N_9381);
and U9755 (N_9755,N_9378,N_9061);
xnor U9756 (N_9756,N_9129,N_9128);
or U9757 (N_9757,N_9399,N_9000);
nand U9758 (N_9758,N_9270,N_9375);
xor U9759 (N_9759,N_9201,N_9309);
nor U9760 (N_9760,N_9062,N_9325);
nand U9761 (N_9761,N_9485,N_9286);
nor U9762 (N_9762,N_9172,N_9192);
nand U9763 (N_9763,N_9285,N_9134);
nand U9764 (N_9764,N_9214,N_9313);
and U9765 (N_9765,N_9149,N_9071);
nor U9766 (N_9766,N_9090,N_9104);
or U9767 (N_9767,N_9298,N_9377);
or U9768 (N_9768,N_9421,N_9374);
nand U9769 (N_9769,N_9134,N_9215);
nand U9770 (N_9770,N_9453,N_9269);
and U9771 (N_9771,N_9011,N_9087);
or U9772 (N_9772,N_9350,N_9399);
and U9773 (N_9773,N_9423,N_9473);
nand U9774 (N_9774,N_9411,N_9484);
xnor U9775 (N_9775,N_9392,N_9013);
and U9776 (N_9776,N_9472,N_9150);
xor U9777 (N_9777,N_9370,N_9071);
nor U9778 (N_9778,N_9154,N_9236);
or U9779 (N_9779,N_9309,N_9488);
or U9780 (N_9780,N_9100,N_9260);
nor U9781 (N_9781,N_9114,N_9414);
or U9782 (N_9782,N_9306,N_9377);
nand U9783 (N_9783,N_9338,N_9306);
nand U9784 (N_9784,N_9187,N_9317);
nor U9785 (N_9785,N_9202,N_9226);
and U9786 (N_9786,N_9282,N_9109);
nor U9787 (N_9787,N_9484,N_9474);
and U9788 (N_9788,N_9251,N_9496);
nand U9789 (N_9789,N_9327,N_9281);
and U9790 (N_9790,N_9026,N_9145);
or U9791 (N_9791,N_9384,N_9222);
nor U9792 (N_9792,N_9112,N_9187);
or U9793 (N_9793,N_9248,N_9369);
nand U9794 (N_9794,N_9143,N_9475);
nand U9795 (N_9795,N_9420,N_9004);
and U9796 (N_9796,N_9134,N_9275);
nor U9797 (N_9797,N_9207,N_9274);
and U9798 (N_9798,N_9261,N_9470);
and U9799 (N_9799,N_9197,N_9293);
xor U9800 (N_9800,N_9445,N_9131);
nor U9801 (N_9801,N_9315,N_9073);
nor U9802 (N_9802,N_9425,N_9244);
and U9803 (N_9803,N_9371,N_9442);
or U9804 (N_9804,N_9403,N_9320);
and U9805 (N_9805,N_9320,N_9140);
nand U9806 (N_9806,N_9233,N_9415);
and U9807 (N_9807,N_9026,N_9006);
nand U9808 (N_9808,N_9151,N_9481);
nor U9809 (N_9809,N_9432,N_9196);
nand U9810 (N_9810,N_9238,N_9468);
nand U9811 (N_9811,N_9160,N_9169);
or U9812 (N_9812,N_9219,N_9493);
nor U9813 (N_9813,N_9294,N_9260);
or U9814 (N_9814,N_9247,N_9020);
nor U9815 (N_9815,N_9147,N_9304);
or U9816 (N_9816,N_9327,N_9367);
or U9817 (N_9817,N_9155,N_9129);
nand U9818 (N_9818,N_9036,N_9129);
and U9819 (N_9819,N_9059,N_9013);
or U9820 (N_9820,N_9049,N_9051);
nand U9821 (N_9821,N_9020,N_9477);
or U9822 (N_9822,N_9027,N_9491);
nor U9823 (N_9823,N_9139,N_9271);
nor U9824 (N_9824,N_9002,N_9314);
nand U9825 (N_9825,N_9124,N_9168);
nand U9826 (N_9826,N_9481,N_9115);
nand U9827 (N_9827,N_9412,N_9323);
or U9828 (N_9828,N_9068,N_9492);
and U9829 (N_9829,N_9014,N_9047);
nor U9830 (N_9830,N_9153,N_9111);
or U9831 (N_9831,N_9443,N_9032);
nor U9832 (N_9832,N_9116,N_9284);
or U9833 (N_9833,N_9146,N_9004);
nand U9834 (N_9834,N_9278,N_9337);
xnor U9835 (N_9835,N_9060,N_9480);
or U9836 (N_9836,N_9352,N_9107);
and U9837 (N_9837,N_9244,N_9313);
and U9838 (N_9838,N_9063,N_9055);
or U9839 (N_9839,N_9089,N_9353);
nor U9840 (N_9840,N_9083,N_9299);
nand U9841 (N_9841,N_9266,N_9077);
and U9842 (N_9842,N_9373,N_9054);
or U9843 (N_9843,N_9487,N_9326);
nor U9844 (N_9844,N_9191,N_9092);
or U9845 (N_9845,N_9305,N_9339);
and U9846 (N_9846,N_9324,N_9059);
nor U9847 (N_9847,N_9371,N_9283);
nor U9848 (N_9848,N_9023,N_9420);
xnor U9849 (N_9849,N_9387,N_9365);
nand U9850 (N_9850,N_9365,N_9259);
and U9851 (N_9851,N_9340,N_9235);
or U9852 (N_9852,N_9179,N_9449);
and U9853 (N_9853,N_9458,N_9069);
and U9854 (N_9854,N_9050,N_9205);
nand U9855 (N_9855,N_9321,N_9193);
and U9856 (N_9856,N_9309,N_9364);
nand U9857 (N_9857,N_9408,N_9040);
or U9858 (N_9858,N_9055,N_9368);
or U9859 (N_9859,N_9185,N_9478);
xnor U9860 (N_9860,N_9017,N_9409);
xor U9861 (N_9861,N_9217,N_9299);
or U9862 (N_9862,N_9474,N_9189);
xnor U9863 (N_9863,N_9244,N_9442);
nor U9864 (N_9864,N_9333,N_9151);
and U9865 (N_9865,N_9080,N_9187);
nand U9866 (N_9866,N_9372,N_9019);
or U9867 (N_9867,N_9358,N_9118);
or U9868 (N_9868,N_9139,N_9367);
nand U9869 (N_9869,N_9369,N_9241);
or U9870 (N_9870,N_9240,N_9418);
nand U9871 (N_9871,N_9028,N_9211);
and U9872 (N_9872,N_9435,N_9234);
nor U9873 (N_9873,N_9291,N_9305);
xnor U9874 (N_9874,N_9223,N_9402);
or U9875 (N_9875,N_9260,N_9309);
nand U9876 (N_9876,N_9352,N_9088);
or U9877 (N_9877,N_9427,N_9058);
or U9878 (N_9878,N_9252,N_9270);
nor U9879 (N_9879,N_9476,N_9453);
nor U9880 (N_9880,N_9167,N_9241);
nand U9881 (N_9881,N_9223,N_9125);
nand U9882 (N_9882,N_9345,N_9339);
nor U9883 (N_9883,N_9409,N_9313);
nor U9884 (N_9884,N_9050,N_9416);
nand U9885 (N_9885,N_9058,N_9333);
or U9886 (N_9886,N_9261,N_9440);
or U9887 (N_9887,N_9121,N_9328);
xor U9888 (N_9888,N_9087,N_9139);
xor U9889 (N_9889,N_9323,N_9276);
nand U9890 (N_9890,N_9382,N_9125);
or U9891 (N_9891,N_9181,N_9103);
and U9892 (N_9892,N_9225,N_9043);
and U9893 (N_9893,N_9253,N_9281);
nor U9894 (N_9894,N_9114,N_9305);
or U9895 (N_9895,N_9276,N_9303);
or U9896 (N_9896,N_9010,N_9439);
or U9897 (N_9897,N_9086,N_9358);
xor U9898 (N_9898,N_9313,N_9326);
nor U9899 (N_9899,N_9052,N_9279);
or U9900 (N_9900,N_9254,N_9345);
xor U9901 (N_9901,N_9427,N_9147);
xor U9902 (N_9902,N_9214,N_9065);
and U9903 (N_9903,N_9034,N_9156);
xor U9904 (N_9904,N_9361,N_9411);
or U9905 (N_9905,N_9193,N_9184);
xnor U9906 (N_9906,N_9029,N_9002);
and U9907 (N_9907,N_9257,N_9116);
and U9908 (N_9908,N_9188,N_9149);
and U9909 (N_9909,N_9306,N_9070);
nor U9910 (N_9910,N_9122,N_9485);
nor U9911 (N_9911,N_9058,N_9357);
and U9912 (N_9912,N_9347,N_9488);
xnor U9913 (N_9913,N_9058,N_9377);
or U9914 (N_9914,N_9346,N_9268);
nand U9915 (N_9915,N_9262,N_9270);
xnor U9916 (N_9916,N_9332,N_9115);
xnor U9917 (N_9917,N_9314,N_9481);
nor U9918 (N_9918,N_9385,N_9376);
nand U9919 (N_9919,N_9478,N_9482);
nor U9920 (N_9920,N_9280,N_9059);
or U9921 (N_9921,N_9005,N_9207);
or U9922 (N_9922,N_9317,N_9412);
nand U9923 (N_9923,N_9134,N_9197);
nand U9924 (N_9924,N_9044,N_9102);
nand U9925 (N_9925,N_9241,N_9429);
and U9926 (N_9926,N_9433,N_9388);
nor U9927 (N_9927,N_9317,N_9086);
nand U9928 (N_9928,N_9387,N_9290);
nand U9929 (N_9929,N_9279,N_9343);
and U9930 (N_9930,N_9183,N_9333);
or U9931 (N_9931,N_9025,N_9303);
or U9932 (N_9932,N_9155,N_9362);
or U9933 (N_9933,N_9178,N_9252);
nor U9934 (N_9934,N_9041,N_9089);
and U9935 (N_9935,N_9410,N_9057);
nand U9936 (N_9936,N_9089,N_9477);
nand U9937 (N_9937,N_9034,N_9209);
xor U9938 (N_9938,N_9315,N_9155);
nand U9939 (N_9939,N_9347,N_9292);
and U9940 (N_9940,N_9409,N_9322);
nor U9941 (N_9941,N_9150,N_9366);
or U9942 (N_9942,N_9005,N_9034);
nand U9943 (N_9943,N_9197,N_9271);
xor U9944 (N_9944,N_9062,N_9425);
nand U9945 (N_9945,N_9437,N_9400);
xor U9946 (N_9946,N_9364,N_9322);
or U9947 (N_9947,N_9105,N_9428);
nor U9948 (N_9948,N_9276,N_9066);
and U9949 (N_9949,N_9290,N_9145);
and U9950 (N_9950,N_9028,N_9344);
nor U9951 (N_9951,N_9108,N_9286);
nor U9952 (N_9952,N_9337,N_9223);
and U9953 (N_9953,N_9083,N_9243);
nor U9954 (N_9954,N_9321,N_9458);
nor U9955 (N_9955,N_9104,N_9340);
nor U9956 (N_9956,N_9144,N_9194);
and U9957 (N_9957,N_9216,N_9201);
xor U9958 (N_9958,N_9394,N_9282);
nor U9959 (N_9959,N_9381,N_9314);
xnor U9960 (N_9960,N_9334,N_9163);
or U9961 (N_9961,N_9396,N_9385);
nor U9962 (N_9962,N_9266,N_9064);
and U9963 (N_9963,N_9022,N_9327);
nand U9964 (N_9964,N_9479,N_9105);
and U9965 (N_9965,N_9020,N_9319);
nand U9966 (N_9966,N_9092,N_9038);
nand U9967 (N_9967,N_9247,N_9316);
xnor U9968 (N_9968,N_9396,N_9118);
nor U9969 (N_9969,N_9148,N_9279);
nand U9970 (N_9970,N_9207,N_9161);
nor U9971 (N_9971,N_9032,N_9053);
or U9972 (N_9972,N_9118,N_9200);
nor U9973 (N_9973,N_9428,N_9406);
nor U9974 (N_9974,N_9150,N_9463);
or U9975 (N_9975,N_9059,N_9292);
or U9976 (N_9976,N_9047,N_9124);
or U9977 (N_9977,N_9147,N_9077);
nor U9978 (N_9978,N_9181,N_9220);
nor U9979 (N_9979,N_9384,N_9004);
or U9980 (N_9980,N_9006,N_9132);
nor U9981 (N_9981,N_9448,N_9106);
or U9982 (N_9982,N_9211,N_9300);
and U9983 (N_9983,N_9182,N_9305);
nor U9984 (N_9984,N_9165,N_9043);
or U9985 (N_9985,N_9482,N_9097);
xnor U9986 (N_9986,N_9009,N_9162);
nand U9987 (N_9987,N_9110,N_9452);
and U9988 (N_9988,N_9282,N_9397);
xor U9989 (N_9989,N_9476,N_9427);
nor U9990 (N_9990,N_9042,N_9046);
and U9991 (N_9991,N_9376,N_9119);
and U9992 (N_9992,N_9259,N_9271);
nor U9993 (N_9993,N_9107,N_9177);
nor U9994 (N_9994,N_9178,N_9417);
or U9995 (N_9995,N_9393,N_9359);
and U9996 (N_9996,N_9286,N_9229);
nand U9997 (N_9997,N_9255,N_9422);
or U9998 (N_9998,N_9164,N_9317);
nor U9999 (N_9999,N_9398,N_9151);
or UO_0 (O_0,N_9581,N_9711);
or UO_1 (O_1,N_9716,N_9720);
and UO_2 (O_2,N_9831,N_9806);
nor UO_3 (O_3,N_9650,N_9507);
nand UO_4 (O_4,N_9566,N_9722);
or UO_5 (O_5,N_9809,N_9953);
and UO_6 (O_6,N_9896,N_9772);
and UO_7 (O_7,N_9934,N_9580);
nor UO_8 (O_8,N_9647,N_9593);
nor UO_9 (O_9,N_9827,N_9639);
nand UO_10 (O_10,N_9980,N_9890);
and UO_11 (O_11,N_9741,N_9565);
or UO_12 (O_12,N_9958,N_9626);
nor UO_13 (O_13,N_9978,N_9868);
nor UO_14 (O_14,N_9740,N_9582);
and UO_15 (O_15,N_9805,N_9757);
nand UO_16 (O_16,N_9972,N_9508);
or UO_17 (O_17,N_9574,N_9898);
nor UO_18 (O_18,N_9587,N_9993);
nor UO_19 (O_19,N_9552,N_9586);
and UO_20 (O_20,N_9847,N_9705);
nand UO_21 (O_21,N_9967,N_9707);
or UO_22 (O_22,N_9816,N_9951);
nand UO_23 (O_23,N_9556,N_9825);
nand UO_24 (O_24,N_9840,N_9889);
nor UO_25 (O_25,N_9937,N_9697);
or UO_26 (O_26,N_9532,N_9622);
nor UO_27 (O_27,N_9842,N_9683);
nor UO_28 (O_28,N_9925,N_9742);
nand UO_29 (O_29,N_9504,N_9519);
and UO_30 (O_30,N_9863,N_9845);
or UO_31 (O_31,N_9962,N_9916);
nor UO_32 (O_32,N_9744,N_9878);
or UO_33 (O_33,N_9685,N_9866);
or UO_34 (O_34,N_9540,N_9834);
nor UO_35 (O_35,N_9558,N_9724);
nor UO_36 (O_36,N_9652,N_9846);
nor UO_37 (O_37,N_9636,N_9909);
or UO_38 (O_38,N_9715,N_9555);
nand UO_39 (O_39,N_9512,N_9858);
and UO_40 (O_40,N_9598,N_9968);
xnor UO_41 (O_41,N_9952,N_9538);
and UO_42 (O_42,N_9543,N_9838);
or UO_43 (O_43,N_9928,N_9974);
nor UO_44 (O_44,N_9982,N_9762);
nand UO_45 (O_45,N_9698,N_9988);
or UO_46 (O_46,N_9960,N_9571);
nor UO_47 (O_47,N_9785,N_9750);
or UO_48 (O_48,N_9500,N_9549);
nand UO_49 (O_49,N_9600,N_9634);
xnor UO_50 (O_50,N_9933,N_9595);
and UO_51 (O_51,N_9906,N_9651);
nand UO_52 (O_52,N_9841,N_9696);
nor UO_53 (O_53,N_9665,N_9568);
nor UO_54 (O_54,N_9624,N_9601);
nand UO_55 (O_55,N_9609,N_9536);
nand UO_56 (O_56,N_9644,N_9918);
nor UO_57 (O_57,N_9915,N_9527);
nor UO_58 (O_58,N_9767,N_9525);
xnor UO_59 (O_59,N_9637,N_9688);
and UO_60 (O_60,N_9701,N_9623);
nand UO_61 (O_61,N_9812,N_9931);
or UO_62 (O_62,N_9784,N_9681);
and UO_63 (O_63,N_9513,N_9761);
nor UO_64 (O_64,N_9714,N_9717);
or UO_65 (O_65,N_9760,N_9964);
xor UO_66 (O_66,N_9794,N_9506);
or UO_67 (O_67,N_9535,N_9975);
and UO_68 (O_68,N_9655,N_9584);
or UO_69 (O_69,N_9718,N_9577);
or UO_70 (O_70,N_9611,N_9853);
nor UO_71 (O_71,N_9766,N_9779);
nor UO_72 (O_72,N_9596,N_9563);
and UO_73 (O_73,N_9514,N_9541);
nor UO_74 (O_74,N_9755,N_9894);
nor UO_75 (O_75,N_9654,N_9804);
and UO_76 (O_76,N_9857,N_9808);
or UO_77 (O_77,N_9927,N_9682);
and UO_78 (O_78,N_9979,N_9664);
or UO_79 (O_79,N_9815,N_9656);
and UO_80 (O_80,N_9738,N_9795);
and UO_81 (O_81,N_9613,N_9899);
or UO_82 (O_82,N_9771,N_9893);
or UO_83 (O_83,N_9822,N_9924);
nand UO_84 (O_84,N_9989,N_9884);
or UO_85 (O_85,N_9604,N_9678);
nand UO_86 (O_86,N_9887,N_9542);
or UO_87 (O_87,N_9510,N_9502);
nand UO_88 (O_88,N_9932,N_9904);
nand UO_89 (O_89,N_9920,N_9559);
nand UO_90 (O_90,N_9686,N_9533);
xnor UO_91 (O_91,N_9873,N_9632);
nand UO_92 (O_92,N_9914,N_9780);
nand UO_93 (O_93,N_9680,N_9672);
xnor UO_94 (O_94,N_9796,N_9905);
and UO_95 (O_95,N_9522,N_9912);
or UO_96 (O_96,N_9712,N_9941);
or UO_97 (O_97,N_9590,N_9743);
or UO_98 (O_98,N_9764,N_9801);
or UO_99 (O_99,N_9782,N_9814);
or UO_100 (O_100,N_9800,N_9709);
nand UO_101 (O_101,N_9999,N_9923);
or UO_102 (O_102,N_9769,N_9629);
or UO_103 (O_103,N_9560,N_9944);
nand UO_104 (O_104,N_9728,N_9876);
nand UO_105 (O_105,N_9903,N_9936);
nand UO_106 (O_106,N_9957,N_9839);
nand UO_107 (O_107,N_9830,N_9684);
nor UO_108 (O_108,N_9710,N_9702);
nor UO_109 (O_109,N_9687,N_9669);
and UO_110 (O_110,N_9546,N_9950);
and UO_111 (O_111,N_9592,N_9947);
nand UO_112 (O_112,N_9786,N_9956);
or UO_113 (O_113,N_9792,N_9589);
nor UO_114 (O_114,N_9921,N_9737);
and UO_115 (O_115,N_9976,N_9564);
or UO_116 (O_116,N_9658,N_9554);
or UO_117 (O_117,N_9612,N_9700);
nand UO_118 (O_118,N_9864,N_9640);
and UO_119 (O_119,N_9691,N_9511);
nor UO_120 (O_120,N_9872,N_9783);
nor UO_121 (O_121,N_9692,N_9505);
or UO_122 (O_122,N_9575,N_9843);
and UO_123 (O_123,N_9745,N_9770);
and UO_124 (O_124,N_9620,N_9938);
nor UO_125 (O_125,N_9917,N_9746);
or UO_126 (O_126,N_9539,N_9621);
nor UO_127 (O_127,N_9567,N_9673);
nor UO_128 (O_128,N_9668,N_9942);
and UO_129 (O_129,N_9959,N_9667);
nor UO_130 (O_130,N_9823,N_9985);
and UO_131 (O_131,N_9641,N_9579);
and UO_132 (O_132,N_9523,N_9562);
nor UO_133 (O_133,N_9662,N_9693);
nor UO_134 (O_134,N_9790,N_9824);
nor UO_135 (O_135,N_9895,N_9799);
xor UO_136 (O_136,N_9869,N_9836);
or UO_137 (O_137,N_9572,N_9984);
nand UO_138 (O_138,N_9851,N_9892);
nand UO_139 (O_139,N_9930,N_9754);
nand UO_140 (O_140,N_9594,N_9676);
nand UO_141 (O_141,N_9550,N_9987);
and UO_142 (O_142,N_9605,N_9671);
and UO_143 (O_143,N_9802,N_9759);
nand UO_144 (O_144,N_9534,N_9588);
and UO_145 (O_145,N_9585,N_9674);
or UO_146 (O_146,N_9633,N_9977);
or UO_147 (O_147,N_9602,N_9570);
nand UO_148 (O_148,N_9775,N_9619);
and UO_149 (O_149,N_9614,N_9756);
nor UO_150 (O_150,N_9530,N_9578);
and UO_151 (O_151,N_9569,N_9954);
and UO_152 (O_152,N_9807,N_9996);
or UO_153 (O_153,N_9850,N_9990);
nor UO_154 (O_154,N_9791,N_9854);
or UO_155 (O_155,N_9627,N_9888);
nor UO_156 (O_156,N_9798,N_9897);
nor UO_157 (O_157,N_9926,N_9518);
and UO_158 (O_158,N_9865,N_9666);
nor UO_159 (O_159,N_9970,N_9739);
nor UO_160 (O_160,N_9945,N_9994);
and UO_161 (O_161,N_9529,N_9969);
or UO_162 (O_162,N_9777,N_9955);
nor UO_163 (O_163,N_9591,N_9638);
or UO_164 (O_164,N_9885,N_9544);
or UO_165 (O_165,N_9811,N_9768);
nor UO_166 (O_166,N_9731,N_9880);
xnor UO_167 (O_167,N_9723,N_9875);
and UO_168 (O_168,N_9788,N_9599);
or UO_169 (O_169,N_9521,N_9732);
nand UO_170 (O_170,N_9597,N_9660);
and UO_171 (O_171,N_9689,N_9736);
xnor UO_172 (O_172,N_9793,N_9703);
or UO_173 (O_173,N_9520,N_9528);
and UO_174 (O_174,N_9751,N_9747);
nand UO_175 (O_175,N_9910,N_9733);
and UO_176 (O_176,N_9835,N_9630);
and UO_177 (O_177,N_9818,N_9643);
nor UO_178 (O_178,N_9606,N_9503);
nand UO_179 (O_179,N_9729,N_9870);
nor UO_180 (O_180,N_9922,N_9734);
nand UO_181 (O_181,N_9603,N_9860);
nor UO_182 (O_182,N_9855,N_9907);
and UO_183 (O_183,N_9810,N_9908);
nand UO_184 (O_184,N_9803,N_9561);
nand UO_185 (O_185,N_9774,N_9981);
or UO_186 (O_186,N_9642,N_9879);
nor UO_187 (O_187,N_9670,N_9752);
nor UO_188 (O_188,N_9832,N_9617);
xor UO_189 (O_189,N_9911,N_9929);
nand UO_190 (O_190,N_9826,N_9776);
and UO_191 (O_191,N_9919,N_9852);
nand UO_192 (O_192,N_9758,N_9699);
nor UO_193 (O_193,N_9615,N_9719);
or UO_194 (O_194,N_9961,N_9874);
nor UO_195 (O_195,N_9573,N_9861);
xor UO_196 (O_196,N_9787,N_9725);
nor UO_197 (O_197,N_9935,N_9986);
xor UO_198 (O_198,N_9721,N_9881);
or UO_199 (O_199,N_9995,N_9648);
or UO_200 (O_200,N_9649,N_9653);
and UO_201 (O_201,N_9773,N_9713);
xor UO_202 (O_202,N_9867,N_9677);
and UO_203 (O_203,N_9829,N_9659);
or UO_204 (O_204,N_9663,N_9516);
and UO_205 (O_205,N_9859,N_9797);
nand UO_206 (O_206,N_9628,N_9781);
nor UO_207 (O_207,N_9833,N_9973);
nand UO_208 (O_208,N_9849,N_9509);
nand UO_209 (O_209,N_9545,N_9862);
nor UO_210 (O_210,N_9661,N_9675);
nand UO_211 (O_211,N_9548,N_9608);
nand UO_212 (O_212,N_9837,N_9871);
and UO_213 (O_213,N_9690,N_9616);
nand UO_214 (O_214,N_9631,N_9813);
or UO_215 (O_215,N_9856,N_9943);
nor UO_216 (O_216,N_9991,N_9891);
and UO_217 (O_217,N_9635,N_9902);
nor UO_218 (O_218,N_9547,N_9646);
nand UO_219 (O_219,N_9576,N_9694);
or UO_220 (O_220,N_9966,N_9983);
nand UO_221 (O_221,N_9553,N_9848);
nand UO_222 (O_222,N_9517,N_9763);
or UO_223 (O_223,N_9963,N_9735);
or UO_224 (O_224,N_9515,N_9992);
and UO_225 (O_225,N_9765,N_9583);
xor UO_226 (O_226,N_9708,N_9940);
nand UO_227 (O_227,N_9749,N_9501);
and UO_228 (O_228,N_9730,N_9820);
and UO_229 (O_229,N_9551,N_9883);
and UO_230 (O_230,N_9971,N_9997);
nor UO_231 (O_231,N_9531,N_9704);
or UO_232 (O_232,N_9607,N_9695);
nand UO_233 (O_233,N_9789,N_9657);
and UO_234 (O_234,N_9948,N_9965);
and UO_235 (O_235,N_9524,N_9753);
nand UO_236 (O_236,N_9625,N_9778);
or UO_237 (O_237,N_9828,N_9877);
nor UO_238 (O_238,N_9882,N_9886);
nand UO_239 (O_239,N_9998,N_9706);
and UO_240 (O_240,N_9913,N_9610);
and UO_241 (O_241,N_9946,N_9817);
or UO_242 (O_242,N_9679,N_9844);
nand UO_243 (O_243,N_9726,N_9821);
and UO_244 (O_244,N_9939,N_9949);
nand UO_245 (O_245,N_9537,N_9900);
or UO_246 (O_246,N_9901,N_9727);
nand UO_247 (O_247,N_9645,N_9526);
or UO_248 (O_248,N_9748,N_9819);
or UO_249 (O_249,N_9557,N_9618);
or UO_250 (O_250,N_9793,N_9598);
nand UO_251 (O_251,N_9739,N_9707);
nor UO_252 (O_252,N_9903,N_9746);
nand UO_253 (O_253,N_9713,N_9703);
nor UO_254 (O_254,N_9575,N_9635);
nor UO_255 (O_255,N_9832,N_9620);
or UO_256 (O_256,N_9709,N_9525);
or UO_257 (O_257,N_9883,N_9910);
nand UO_258 (O_258,N_9665,N_9900);
nand UO_259 (O_259,N_9832,N_9740);
xnor UO_260 (O_260,N_9938,N_9595);
and UO_261 (O_261,N_9678,N_9875);
or UO_262 (O_262,N_9998,N_9860);
nand UO_263 (O_263,N_9626,N_9719);
nor UO_264 (O_264,N_9758,N_9915);
nand UO_265 (O_265,N_9863,N_9731);
nor UO_266 (O_266,N_9609,N_9845);
or UO_267 (O_267,N_9982,N_9561);
nor UO_268 (O_268,N_9508,N_9783);
xor UO_269 (O_269,N_9959,N_9966);
nor UO_270 (O_270,N_9982,N_9970);
and UO_271 (O_271,N_9542,N_9961);
and UO_272 (O_272,N_9716,N_9882);
or UO_273 (O_273,N_9981,N_9814);
nor UO_274 (O_274,N_9547,N_9604);
nor UO_275 (O_275,N_9574,N_9522);
or UO_276 (O_276,N_9610,N_9807);
nand UO_277 (O_277,N_9561,N_9546);
nand UO_278 (O_278,N_9646,N_9822);
and UO_279 (O_279,N_9748,N_9942);
nand UO_280 (O_280,N_9535,N_9839);
nand UO_281 (O_281,N_9530,N_9790);
nor UO_282 (O_282,N_9918,N_9777);
nand UO_283 (O_283,N_9850,N_9719);
xnor UO_284 (O_284,N_9993,N_9585);
nor UO_285 (O_285,N_9958,N_9967);
nor UO_286 (O_286,N_9733,N_9602);
or UO_287 (O_287,N_9623,N_9606);
or UO_288 (O_288,N_9503,N_9530);
and UO_289 (O_289,N_9613,N_9996);
or UO_290 (O_290,N_9781,N_9961);
and UO_291 (O_291,N_9896,N_9821);
and UO_292 (O_292,N_9662,N_9941);
xnor UO_293 (O_293,N_9793,N_9796);
nor UO_294 (O_294,N_9750,N_9529);
xor UO_295 (O_295,N_9932,N_9990);
and UO_296 (O_296,N_9639,N_9814);
xnor UO_297 (O_297,N_9853,N_9617);
and UO_298 (O_298,N_9807,N_9918);
and UO_299 (O_299,N_9511,N_9745);
nand UO_300 (O_300,N_9598,N_9720);
and UO_301 (O_301,N_9508,N_9926);
nand UO_302 (O_302,N_9821,N_9546);
nor UO_303 (O_303,N_9888,N_9686);
or UO_304 (O_304,N_9889,N_9557);
xnor UO_305 (O_305,N_9821,N_9717);
and UO_306 (O_306,N_9882,N_9979);
nand UO_307 (O_307,N_9838,N_9825);
or UO_308 (O_308,N_9860,N_9967);
nand UO_309 (O_309,N_9590,N_9852);
nand UO_310 (O_310,N_9712,N_9686);
and UO_311 (O_311,N_9638,N_9846);
or UO_312 (O_312,N_9974,N_9513);
nand UO_313 (O_313,N_9832,N_9697);
nand UO_314 (O_314,N_9756,N_9969);
nand UO_315 (O_315,N_9674,N_9540);
nor UO_316 (O_316,N_9808,N_9604);
and UO_317 (O_317,N_9739,N_9677);
or UO_318 (O_318,N_9870,N_9536);
nand UO_319 (O_319,N_9729,N_9908);
or UO_320 (O_320,N_9730,N_9583);
or UO_321 (O_321,N_9584,N_9637);
and UO_322 (O_322,N_9922,N_9867);
or UO_323 (O_323,N_9817,N_9919);
or UO_324 (O_324,N_9634,N_9973);
nor UO_325 (O_325,N_9536,N_9996);
nor UO_326 (O_326,N_9551,N_9597);
or UO_327 (O_327,N_9601,N_9796);
and UO_328 (O_328,N_9814,N_9832);
nand UO_329 (O_329,N_9582,N_9638);
nor UO_330 (O_330,N_9776,N_9967);
and UO_331 (O_331,N_9729,N_9840);
nand UO_332 (O_332,N_9624,N_9616);
or UO_333 (O_333,N_9935,N_9573);
xnor UO_334 (O_334,N_9866,N_9706);
nor UO_335 (O_335,N_9921,N_9857);
nand UO_336 (O_336,N_9853,N_9733);
and UO_337 (O_337,N_9710,N_9740);
nor UO_338 (O_338,N_9625,N_9645);
nand UO_339 (O_339,N_9979,N_9989);
and UO_340 (O_340,N_9844,N_9994);
nor UO_341 (O_341,N_9836,N_9643);
xor UO_342 (O_342,N_9730,N_9788);
nand UO_343 (O_343,N_9889,N_9948);
and UO_344 (O_344,N_9863,N_9738);
nor UO_345 (O_345,N_9597,N_9626);
nand UO_346 (O_346,N_9811,N_9550);
nand UO_347 (O_347,N_9572,N_9903);
nand UO_348 (O_348,N_9606,N_9980);
and UO_349 (O_349,N_9875,N_9671);
or UO_350 (O_350,N_9579,N_9834);
nor UO_351 (O_351,N_9864,N_9958);
or UO_352 (O_352,N_9753,N_9519);
nand UO_353 (O_353,N_9739,N_9546);
and UO_354 (O_354,N_9723,N_9677);
nor UO_355 (O_355,N_9938,N_9743);
nor UO_356 (O_356,N_9619,N_9560);
and UO_357 (O_357,N_9613,N_9625);
or UO_358 (O_358,N_9840,N_9862);
nand UO_359 (O_359,N_9690,N_9937);
or UO_360 (O_360,N_9979,N_9751);
and UO_361 (O_361,N_9792,N_9722);
nor UO_362 (O_362,N_9762,N_9573);
or UO_363 (O_363,N_9811,N_9877);
nor UO_364 (O_364,N_9975,N_9719);
or UO_365 (O_365,N_9651,N_9844);
nor UO_366 (O_366,N_9651,N_9843);
or UO_367 (O_367,N_9882,N_9599);
or UO_368 (O_368,N_9743,N_9768);
nor UO_369 (O_369,N_9509,N_9983);
and UO_370 (O_370,N_9525,N_9649);
nand UO_371 (O_371,N_9735,N_9803);
or UO_372 (O_372,N_9831,N_9960);
and UO_373 (O_373,N_9789,N_9600);
xor UO_374 (O_374,N_9780,N_9899);
nor UO_375 (O_375,N_9944,N_9888);
or UO_376 (O_376,N_9923,N_9621);
nor UO_377 (O_377,N_9934,N_9870);
nand UO_378 (O_378,N_9847,N_9605);
nand UO_379 (O_379,N_9618,N_9825);
and UO_380 (O_380,N_9790,N_9740);
xor UO_381 (O_381,N_9686,N_9670);
nand UO_382 (O_382,N_9779,N_9770);
and UO_383 (O_383,N_9990,N_9825);
xor UO_384 (O_384,N_9813,N_9636);
and UO_385 (O_385,N_9914,N_9583);
and UO_386 (O_386,N_9895,N_9605);
and UO_387 (O_387,N_9694,N_9922);
or UO_388 (O_388,N_9895,N_9914);
xor UO_389 (O_389,N_9735,N_9521);
and UO_390 (O_390,N_9712,N_9999);
nor UO_391 (O_391,N_9999,N_9919);
nand UO_392 (O_392,N_9567,N_9979);
nand UO_393 (O_393,N_9713,N_9629);
or UO_394 (O_394,N_9571,N_9792);
xnor UO_395 (O_395,N_9640,N_9593);
and UO_396 (O_396,N_9523,N_9522);
nor UO_397 (O_397,N_9960,N_9842);
nor UO_398 (O_398,N_9700,N_9735);
nand UO_399 (O_399,N_9600,N_9831);
or UO_400 (O_400,N_9757,N_9941);
nor UO_401 (O_401,N_9976,N_9715);
or UO_402 (O_402,N_9796,N_9859);
nor UO_403 (O_403,N_9652,N_9796);
nor UO_404 (O_404,N_9944,N_9842);
nand UO_405 (O_405,N_9698,N_9996);
or UO_406 (O_406,N_9820,N_9663);
nand UO_407 (O_407,N_9550,N_9805);
or UO_408 (O_408,N_9960,N_9753);
nand UO_409 (O_409,N_9765,N_9533);
or UO_410 (O_410,N_9673,N_9933);
or UO_411 (O_411,N_9822,N_9605);
or UO_412 (O_412,N_9674,N_9933);
xnor UO_413 (O_413,N_9744,N_9628);
xor UO_414 (O_414,N_9936,N_9774);
xor UO_415 (O_415,N_9940,N_9550);
nand UO_416 (O_416,N_9555,N_9579);
nor UO_417 (O_417,N_9540,N_9955);
nor UO_418 (O_418,N_9970,N_9641);
or UO_419 (O_419,N_9997,N_9709);
xnor UO_420 (O_420,N_9816,N_9994);
nand UO_421 (O_421,N_9511,N_9810);
and UO_422 (O_422,N_9614,N_9838);
nand UO_423 (O_423,N_9935,N_9726);
or UO_424 (O_424,N_9746,N_9638);
and UO_425 (O_425,N_9578,N_9815);
or UO_426 (O_426,N_9860,N_9612);
nor UO_427 (O_427,N_9770,N_9748);
nor UO_428 (O_428,N_9682,N_9734);
nor UO_429 (O_429,N_9744,N_9777);
or UO_430 (O_430,N_9508,N_9776);
xnor UO_431 (O_431,N_9953,N_9501);
nor UO_432 (O_432,N_9864,N_9849);
and UO_433 (O_433,N_9553,N_9707);
nor UO_434 (O_434,N_9657,N_9864);
or UO_435 (O_435,N_9958,N_9706);
nor UO_436 (O_436,N_9586,N_9604);
nor UO_437 (O_437,N_9824,N_9537);
nand UO_438 (O_438,N_9715,N_9556);
nor UO_439 (O_439,N_9808,N_9954);
nand UO_440 (O_440,N_9780,N_9992);
or UO_441 (O_441,N_9587,N_9793);
or UO_442 (O_442,N_9985,N_9848);
and UO_443 (O_443,N_9698,N_9937);
nor UO_444 (O_444,N_9735,N_9603);
xor UO_445 (O_445,N_9907,N_9542);
or UO_446 (O_446,N_9586,N_9769);
nand UO_447 (O_447,N_9630,N_9897);
and UO_448 (O_448,N_9795,N_9584);
nand UO_449 (O_449,N_9834,N_9989);
nor UO_450 (O_450,N_9813,N_9906);
or UO_451 (O_451,N_9650,N_9620);
nor UO_452 (O_452,N_9656,N_9580);
and UO_453 (O_453,N_9634,N_9607);
nor UO_454 (O_454,N_9869,N_9685);
or UO_455 (O_455,N_9942,N_9605);
or UO_456 (O_456,N_9547,N_9573);
nand UO_457 (O_457,N_9990,N_9552);
or UO_458 (O_458,N_9633,N_9802);
nor UO_459 (O_459,N_9986,N_9968);
nor UO_460 (O_460,N_9506,N_9863);
nand UO_461 (O_461,N_9838,N_9818);
and UO_462 (O_462,N_9746,N_9641);
nand UO_463 (O_463,N_9693,N_9503);
and UO_464 (O_464,N_9793,N_9848);
or UO_465 (O_465,N_9688,N_9661);
and UO_466 (O_466,N_9949,N_9522);
nor UO_467 (O_467,N_9607,N_9793);
or UO_468 (O_468,N_9882,N_9617);
and UO_469 (O_469,N_9818,N_9727);
nand UO_470 (O_470,N_9682,N_9739);
or UO_471 (O_471,N_9814,N_9699);
or UO_472 (O_472,N_9866,N_9729);
nor UO_473 (O_473,N_9763,N_9571);
nor UO_474 (O_474,N_9629,N_9845);
or UO_475 (O_475,N_9921,N_9877);
or UO_476 (O_476,N_9782,N_9623);
nor UO_477 (O_477,N_9915,N_9920);
and UO_478 (O_478,N_9872,N_9695);
nor UO_479 (O_479,N_9777,N_9880);
or UO_480 (O_480,N_9694,N_9962);
or UO_481 (O_481,N_9951,N_9682);
nand UO_482 (O_482,N_9786,N_9561);
nand UO_483 (O_483,N_9509,N_9719);
or UO_484 (O_484,N_9911,N_9899);
and UO_485 (O_485,N_9762,N_9991);
and UO_486 (O_486,N_9738,N_9942);
and UO_487 (O_487,N_9540,N_9650);
nor UO_488 (O_488,N_9861,N_9584);
or UO_489 (O_489,N_9963,N_9975);
or UO_490 (O_490,N_9637,N_9914);
nand UO_491 (O_491,N_9927,N_9841);
and UO_492 (O_492,N_9928,N_9653);
and UO_493 (O_493,N_9868,N_9957);
xor UO_494 (O_494,N_9816,N_9796);
and UO_495 (O_495,N_9907,N_9957);
nand UO_496 (O_496,N_9984,N_9974);
xnor UO_497 (O_497,N_9939,N_9919);
xnor UO_498 (O_498,N_9724,N_9693);
or UO_499 (O_499,N_9703,N_9639);
or UO_500 (O_500,N_9856,N_9522);
xnor UO_501 (O_501,N_9525,N_9785);
nor UO_502 (O_502,N_9535,N_9922);
nand UO_503 (O_503,N_9882,N_9597);
or UO_504 (O_504,N_9695,N_9741);
or UO_505 (O_505,N_9697,N_9645);
or UO_506 (O_506,N_9776,N_9852);
xnor UO_507 (O_507,N_9732,N_9907);
nand UO_508 (O_508,N_9837,N_9629);
or UO_509 (O_509,N_9999,N_9546);
nand UO_510 (O_510,N_9932,N_9771);
and UO_511 (O_511,N_9560,N_9599);
nor UO_512 (O_512,N_9503,N_9917);
nor UO_513 (O_513,N_9979,N_9973);
nor UO_514 (O_514,N_9788,N_9949);
and UO_515 (O_515,N_9578,N_9548);
or UO_516 (O_516,N_9754,N_9855);
or UO_517 (O_517,N_9708,N_9790);
nor UO_518 (O_518,N_9941,N_9810);
xor UO_519 (O_519,N_9988,N_9608);
nor UO_520 (O_520,N_9830,N_9622);
nand UO_521 (O_521,N_9524,N_9542);
or UO_522 (O_522,N_9986,N_9521);
and UO_523 (O_523,N_9646,N_9827);
or UO_524 (O_524,N_9937,N_9936);
nand UO_525 (O_525,N_9852,N_9908);
and UO_526 (O_526,N_9762,N_9900);
and UO_527 (O_527,N_9549,N_9761);
or UO_528 (O_528,N_9928,N_9607);
and UO_529 (O_529,N_9542,N_9790);
or UO_530 (O_530,N_9882,N_9680);
xor UO_531 (O_531,N_9994,N_9553);
and UO_532 (O_532,N_9977,N_9520);
nor UO_533 (O_533,N_9790,N_9737);
nor UO_534 (O_534,N_9570,N_9974);
and UO_535 (O_535,N_9709,N_9868);
nor UO_536 (O_536,N_9505,N_9532);
and UO_537 (O_537,N_9623,N_9737);
nand UO_538 (O_538,N_9672,N_9798);
nor UO_539 (O_539,N_9507,N_9866);
nand UO_540 (O_540,N_9510,N_9562);
nand UO_541 (O_541,N_9649,N_9609);
nand UO_542 (O_542,N_9760,N_9996);
or UO_543 (O_543,N_9560,N_9992);
or UO_544 (O_544,N_9516,N_9762);
xor UO_545 (O_545,N_9958,N_9754);
and UO_546 (O_546,N_9619,N_9795);
nand UO_547 (O_547,N_9942,N_9588);
and UO_548 (O_548,N_9872,N_9874);
or UO_549 (O_549,N_9530,N_9717);
or UO_550 (O_550,N_9532,N_9524);
or UO_551 (O_551,N_9728,N_9830);
and UO_552 (O_552,N_9944,N_9723);
or UO_553 (O_553,N_9797,N_9545);
or UO_554 (O_554,N_9668,N_9976);
nor UO_555 (O_555,N_9941,N_9917);
nand UO_556 (O_556,N_9708,N_9770);
or UO_557 (O_557,N_9738,N_9640);
nand UO_558 (O_558,N_9521,N_9970);
nor UO_559 (O_559,N_9838,N_9947);
nor UO_560 (O_560,N_9977,N_9954);
or UO_561 (O_561,N_9686,N_9862);
or UO_562 (O_562,N_9681,N_9694);
nand UO_563 (O_563,N_9928,N_9834);
nor UO_564 (O_564,N_9878,N_9804);
nor UO_565 (O_565,N_9649,N_9775);
nor UO_566 (O_566,N_9729,N_9720);
nand UO_567 (O_567,N_9576,N_9744);
and UO_568 (O_568,N_9977,N_9777);
and UO_569 (O_569,N_9805,N_9934);
or UO_570 (O_570,N_9805,N_9652);
nand UO_571 (O_571,N_9912,N_9632);
and UO_572 (O_572,N_9824,N_9709);
nand UO_573 (O_573,N_9627,N_9880);
nor UO_574 (O_574,N_9793,N_9898);
and UO_575 (O_575,N_9963,N_9730);
nor UO_576 (O_576,N_9673,N_9819);
and UO_577 (O_577,N_9890,N_9949);
nand UO_578 (O_578,N_9973,N_9937);
and UO_579 (O_579,N_9855,N_9535);
and UO_580 (O_580,N_9598,N_9605);
nand UO_581 (O_581,N_9811,N_9868);
nand UO_582 (O_582,N_9953,N_9817);
nor UO_583 (O_583,N_9866,N_9760);
xnor UO_584 (O_584,N_9873,N_9918);
or UO_585 (O_585,N_9969,N_9913);
nand UO_586 (O_586,N_9524,N_9971);
xor UO_587 (O_587,N_9959,N_9680);
nor UO_588 (O_588,N_9554,N_9504);
and UO_589 (O_589,N_9811,N_9883);
nor UO_590 (O_590,N_9944,N_9714);
nor UO_591 (O_591,N_9673,N_9703);
or UO_592 (O_592,N_9927,N_9749);
nand UO_593 (O_593,N_9706,N_9599);
nor UO_594 (O_594,N_9831,N_9842);
or UO_595 (O_595,N_9825,N_9551);
and UO_596 (O_596,N_9568,N_9781);
and UO_597 (O_597,N_9707,N_9862);
nor UO_598 (O_598,N_9681,N_9749);
xor UO_599 (O_599,N_9812,N_9513);
nor UO_600 (O_600,N_9634,N_9936);
and UO_601 (O_601,N_9857,N_9608);
nand UO_602 (O_602,N_9570,N_9868);
nand UO_603 (O_603,N_9631,N_9683);
nor UO_604 (O_604,N_9709,N_9834);
or UO_605 (O_605,N_9555,N_9732);
nand UO_606 (O_606,N_9771,N_9860);
and UO_607 (O_607,N_9596,N_9656);
nand UO_608 (O_608,N_9750,N_9515);
and UO_609 (O_609,N_9657,N_9886);
and UO_610 (O_610,N_9825,N_9972);
or UO_611 (O_611,N_9795,N_9739);
nor UO_612 (O_612,N_9562,N_9964);
nor UO_613 (O_613,N_9942,N_9691);
xor UO_614 (O_614,N_9881,N_9646);
nand UO_615 (O_615,N_9809,N_9534);
nor UO_616 (O_616,N_9635,N_9777);
nor UO_617 (O_617,N_9572,N_9929);
nand UO_618 (O_618,N_9578,N_9869);
and UO_619 (O_619,N_9704,N_9944);
nand UO_620 (O_620,N_9519,N_9730);
and UO_621 (O_621,N_9993,N_9507);
nor UO_622 (O_622,N_9516,N_9766);
or UO_623 (O_623,N_9830,N_9911);
and UO_624 (O_624,N_9854,N_9610);
and UO_625 (O_625,N_9662,N_9767);
or UO_626 (O_626,N_9989,N_9723);
and UO_627 (O_627,N_9759,N_9972);
xnor UO_628 (O_628,N_9611,N_9642);
nor UO_629 (O_629,N_9868,N_9764);
or UO_630 (O_630,N_9913,N_9713);
nor UO_631 (O_631,N_9613,N_9597);
nor UO_632 (O_632,N_9819,N_9618);
or UO_633 (O_633,N_9871,N_9755);
nor UO_634 (O_634,N_9742,N_9541);
nor UO_635 (O_635,N_9712,N_9698);
nor UO_636 (O_636,N_9839,N_9880);
nor UO_637 (O_637,N_9736,N_9725);
and UO_638 (O_638,N_9936,N_9866);
nor UO_639 (O_639,N_9972,N_9620);
or UO_640 (O_640,N_9859,N_9773);
nor UO_641 (O_641,N_9828,N_9712);
nor UO_642 (O_642,N_9789,N_9656);
nand UO_643 (O_643,N_9831,N_9698);
nor UO_644 (O_644,N_9802,N_9626);
or UO_645 (O_645,N_9529,N_9792);
xor UO_646 (O_646,N_9959,N_9682);
or UO_647 (O_647,N_9537,N_9555);
or UO_648 (O_648,N_9724,N_9835);
and UO_649 (O_649,N_9981,N_9729);
nand UO_650 (O_650,N_9563,N_9932);
or UO_651 (O_651,N_9544,N_9592);
or UO_652 (O_652,N_9568,N_9879);
nor UO_653 (O_653,N_9601,N_9668);
and UO_654 (O_654,N_9927,N_9505);
or UO_655 (O_655,N_9583,N_9985);
nor UO_656 (O_656,N_9561,N_9575);
or UO_657 (O_657,N_9705,N_9756);
or UO_658 (O_658,N_9841,N_9561);
and UO_659 (O_659,N_9954,N_9804);
or UO_660 (O_660,N_9842,N_9929);
or UO_661 (O_661,N_9692,N_9729);
nor UO_662 (O_662,N_9590,N_9679);
nand UO_663 (O_663,N_9869,N_9737);
nor UO_664 (O_664,N_9510,N_9519);
or UO_665 (O_665,N_9885,N_9964);
or UO_666 (O_666,N_9671,N_9952);
or UO_667 (O_667,N_9632,N_9812);
nand UO_668 (O_668,N_9723,N_9658);
or UO_669 (O_669,N_9818,N_9555);
nor UO_670 (O_670,N_9560,N_9855);
xnor UO_671 (O_671,N_9918,N_9944);
and UO_672 (O_672,N_9891,N_9555);
nand UO_673 (O_673,N_9729,N_9815);
or UO_674 (O_674,N_9993,N_9836);
nor UO_675 (O_675,N_9986,N_9547);
nand UO_676 (O_676,N_9600,N_9935);
nor UO_677 (O_677,N_9708,N_9845);
and UO_678 (O_678,N_9677,N_9974);
nand UO_679 (O_679,N_9736,N_9571);
or UO_680 (O_680,N_9977,N_9951);
nor UO_681 (O_681,N_9854,N_9762);
nor UO_682 (O_682,N_9997,N_9981);
nand UO_683 (O_683,N_9717,N_9594);
and UO_684 (O_684,N_9996,N_9663);
or UO_685 (O_685,N_9760,N_9865);
and UO_686 (O_686,N_9671,N_9596);
or UO_687 (O_687,N_9563,N_9826);
nor UO_688 (O_688,N_9929,N_9755);
nand UO_689 (O_689,N_9887,N_9932);
and UO_690 (O_690,N_9979,N_9892);
xor UO_691 (O_691,N_9825,N_9794);
nand UO_692 (O_692,N_9832,N_9938);
or UO_693 (O_693,N_9651,N_9963);
or UO_694 (O_694,N_9756,N_9862);
nor UO_695 (O_695,N_9771,N_9912);
and UO_696 (O_696,N_9853,N_9559);
and UO_697 (O_697,N_9761,N_9978);
nor UO_698 (O_698,N_9901,N_9932);
and UO_699 (O_699,N_9561,N_9591);
and UO_700 (O_700,N_9886,N_9822);
nor UO_701 (O_701,N_9968,N_9991);
and UO_702 (O_702,N_9898,N_9980);
nand UO_703 (O_703,N_9587,N_9571);
nand UO_704 (O_704,N_9662,N_9977);
and UO_705 (O_705,N_9960,N_9642);
nand UO_706 (O_706,N_9686,N_9997);
or UO_707 (O_707,N_9765,N_9791);
nand UO_708 (O_708,N_9695,N_9714);
nor UO_709 (O_709,N_9572,N_9883);
nand UO_710 (O_710,N_9582,N_9710);
nand UO_711 (O_711,N_9665,N_9679);
and UO_712 (O_712,N_9741,N_9865);
nor UO_713 (O_713,N_9867,N_9989);
xnor UO_714 (O_714,N_9665,N_9861);
nor UO_715 (O_715,N_9577,N_9813);
and UO_716 (O_716,N_9702,N_9807);
or UO_717 (O_717,N_9751,N_9788);
or UO_718 (O_718,N_9861,N_9812);
or UO_719 (O_719,N_9715,N_9518);
nand UO_720 (O_720,N_9566,N_9574);
xor UO_721 (O_721,N_9956,N_9818);
nor UO_722 (O_722,N_9741,N_9708);
and UO_723 (O_723,N_9695,N_9804);
or UO_724 (O_724,N_9704,N_9503);
or UO_725 (O_725,N_9913,N_9662);
nor UO_726 (O_726,N_9966,N_9578);
or UO_727 (O_727,N_9561,N_9745);
and UO_728 (O_728,N_9910,N_9690);
or UO_729 (O_729,N_9684,N_9952);
xor UO_730 (O_730,N_9993,N_9615);
nand UO_731 (O_731,N_9942,N_9832);
and UO_732 (O_732,N_9688,N_9966);
and UO_733 (O_733,N_9894,N_9966);
nand UO_734 (O_734,N_9881,N_9966);
nor UO_735 (O_735,N_9893,N_9684);
nand UO_736 (O_736,N_9937,N_9577);
or UO_737 (O_737,N_9754,N_9542);
nand UO_738 (O_738,N_9658,N_9515);
xor UO_739 (O_739,N_9978,N_9662);
nand UO_740 (O_740,N_9778,N_9548);
or UO_741 (O_741,N_9544,N_9556);
or UO_742 (O_742,N_9790,N_9825);
nor UO_743 (O_743,N_9912,N_9836);
nand UO_744 (O_744,N_9615,N_9731);
and UO_745 (O_745,N_9942,N_9737);
and UO_746 (O_746,N_9802,N_9679);
and UO_747 (O_747,N_9915,N_9940);
and UO_748 (O_748,N_9921,N_9853);
nor UO_749 (O_749,N_9984,N_9858);
nand UO_750 (O_750,N_9514,N_9502);
nand UO_751 (O_751,N_9957,N_9697);
nand UO_752 (O_752,N_9625,N_9987);
nor UO_753 (O_753,N_9554,N_9797);
nor UO_754 (O_754,N_9698,N_9856);
nor UO_755 (O_755,N_9917,N_9888);
or UO_756 (O_756,N_9558,N_9523);
xnor UO_757 (O_757,N_9902,N_9607);
nand UO_758 (O_758,N_9615,N_9983);
or UO_759 (O_759,N_9973,N_9790);
nor UO_760 (O_760,N_9596,N_9629);
or UO_761 (O_761,N_9698,N_9968);
or UO_762 (O_762,N_9719,N_9800);
and UO_763 (O_763,N_9745,N_9944);
nand UO_764 (O_764,N_9968,N_9629);
nand UO_765 (O_765,N_9744,N_9855);
xor UO_766 (O_766,N_9898,N_9870);
or UO_767 (O_767,N_9595,N_9630);
nand UO_768 (O_768,N_9745,N_9710);
or UO_769 (O_769,N_9774,N_9613);
nor UO_770 (O_770,N_9882,N_9732);
nor UO_771 (O_771,N_9731,N_9976);
xor UO_772 (O_772,N_9599,N_9977);
nand UO_773 (O_773,N_9501,N_9764);
or UO_774 (O_774,N_9639,N_9501);
nand UO_775 (O_775,N_9642,N_9591);
or UO_776 (O_776,N_9597,N_9530);
and UO_777 (O_777,N_9592,N_9999);
nor UO_778 (O_778,N_9796,N_9803);
nand UO_779 (O_779,N_9844,N_9652);
xor UO_780 (O_780,N_9694,N_9936);
and UO_781 (O_781,N_9926,N_9819);
nor UO_782 (O_782,N_9951,N_9587);
nor UO_783 (O_783,N_9576,N_9837);
nor UO_784 (O_784,N_9946,N_9573);
nand UO_785 (O_785,N_9578,N_9757);
and UO_786 (O_786,N_9799,N_9640);
and UO_787 (O_787,N_9518,N_9533);
nand UO_788 (O_788,N_9930,N_9969);
and UO_789 (O_789,N_9765,N_9761);
and UO_790 (O_790,N_9983,N_9752);
and UO_791 (O_791,N_9959,N_9742);
and UO_792 (O_792,N_9638,N_9549);
xnor UO_793 (O_793,N_9995,N_9963);
and UO_794 (O_794,N_9665,N_9595);
nand UO_795 (O_795,N_9966,N_9531);
nor UO_796 (O_796,N_9540,N_9531);
nor UO_797 (O_797,N_9703,N_9745);
nor UO_798 (O_798,N_9557,N_9527);
or UO_799 (O_799,N_9743,N_9986);
xnor UO_800 (O_800,N_9775,N_9892);
and UO_801 (O_801,N_9818,N_9714);
nand UO_802 (O_802,N_9571,N_9540);
and UO_803 (O_803,N_9643,N_9649);
nand UO_804 (O_804,N_9760,N_9637);
nor UO_805 (O_805,N_9798,N_9836);
xor UO_806 (O_806,N_9534,N_9988);
and UO_807 (O_807,N_9817,N_9518);
nand UO_808 (O_808,N_9656,N_9911);
or UO_809 (O_809,N_9728,N_9864);
nand UO_810 (O_810,N_9640,N_9905);
or UO_811 (O_811,N_9650,N_9996);
or UO_812 (O_812,N_9805,N_9779);
nor UO_813 (O_813,N_9674,N_9511);
nand UO_814 (O_814,N_9500,N_9867);
or UO_815 (O_815,N_9969,N_9799);
and UO_816 (O_816,N_9971,N_9778);
nor UO_817 (O_817,N_9712,N_9551);
or UO_818 (O_818,N_9592,N_9670);
nand UO_819 (O_819,N_9740,N_9879);
nor UO_820 (O_820,N_9761,N_9855);
nor UO_821 (O_821,N_9946,N_9884);
and UO_822 (O_822,N_9853,N_9944);
nand UO_823 (O_823,N_9930,N_9759);
nand UO_824 (O_824,N_9500,N_9817);
or UO_825 (O_825,N_9832,N_9525);
and UO_826 (O_826,N_9925,N_9824);
or UO_827 (O_827,N_9927,N_9536);
and UO_828 (O_828,N_9731,N_9710);
or UO_829 (O_829,N_9991,N_9538);
xnor UO_830 (O_830,N_9538,N_9620);
xnor UO_831 (O_831,N_9697,N_9583);
or UO_832 (O_832,N_9821,N_9548);
nand UO_833 (O_833,N_9651,N_9691);
or UO_834 (O_834,N_9578,N_9787);
and UO_835 (O_835,N_9788,N_9666);
xnor UO_836 (O_836,N_9560,N_9709);
nand UO_837 (O_837,N_9807,N_9707);
and UO_838 (O_838,N_9591,N_9666);
and UO_839 (O_839,N_9589,N_9968);
or UO_840 (O_840,N_9706,N_9707);
and UO_841 (O_841,N_9753,N_9617);
nand UO_842 (O_842,N_9980,N_9860);
and UO_843 (O_843,N_9548,N_9925);
xnor UO_844 (O_844,N_9736,N_9894);
nor UO_845 (O_845,N_9977,N_9764);
or UO_846 (O_846,N_9591,N_9709);
nand UO_847 (O_847,N_9615,N_9623);
nand UO_848 (O_848,N_9887,N_9927);
and UO_849 (O_849,N_9988,N_9564);
or UO_850 (O_850,N_9869,N_9529);
nand UO_851 (O_851,N_9615,N_9827);
nand UO_852 (O_852,N_9707,N_9916);
or UO_853 (O_853,N_9913,N_9925);
xor UO_854 (O_854,N_9583,N_9835);
nor UO_855 (O_855,N_9855,N_9555);
and UO_856 (O_856,N_9724,N_9603);
and UO_857 (O_857,N_9598,N_9922);
nand UO_858 (O_858,N_9580,N_9971);
nand UO_859 (O_859,N_9938,N_9593);
or UO_860 (O_860,N_9651,N_9532);
nand UO_861 (O_861,N_9695,N_9823);
nor UO_862 (O_862,N_9939,N_9556);
or UO_863 (O_863,N_9634,N_9926);
nor UO_864 (O_864,N_9903,N_9608);
xor UO_865 (O_865,N_9647,N_9840);
or UO_866 (O_866,N_9974,N_9771);
nand UO_867 (O_867,N_9943,N_9883);
nor UO_868 (O_868,N_9622,N_9786);
nor UO_869 (O_869,N_9759,N_9558);
and UO_870 (O_870,N_9994,N_9520);
or UO_871 (O_871,N_9598,N_9561);
or UO_872 (O_872,N_9804,N_9643);
or UO_873 (O_873,N_9934,N_9630);
nor UO_874 (O_874,N_9684,N_9781);
and UO_875 (O_875,N_9526,N_9517);
nand UO_876 (O_876,N_9611,N_9607);
nor UO_877 (O_877,N_9762,N_9796);
nand UO_878 (O_878,N_9929,N_9683);
nand UO_879 (O_879,N_9946,N_9680);
nand UO_880 (O_880,N_9880,N_9861);
nor UO_881 (O_881,N_9633,N_9910);
or UO_882 (O_882,N_9695,N_9647);
nand UO_883 (O_883,N_9928,N_9567);
and UO_884 (O_884,N_9639,N_9635);
and UO_885 (O_885,N_9657,N_9739);
nor UO_886 (O_886,N_9609,N_9926);
and UO_887 (O_887,N_9955,N_9950);
nand UO_888 (O_888,N_9728,N_9608);
and UO_889 (O_889,N_9907,N_9789);
and UO_890 (O_890,N_9566,N_9696);
xor UO_891 (O_891,N_9965,N_9854);
and UO_892 (O_892,N_9756,N_9811);
nand UO_893 (O_893,N_9782,N_9680);
and UO_894 (O_894,N_9944,N_9987);
or UO_895 (O_895,N_9519,N_9507);
nor UO_896 (O_896,N_9555,N_9788);
xnor UO_897 (O_897,N_9651,N_9693);
nor UO_898 (O_898,N_9709,N_9693);
xor UO_899 (O_899,N_9961,N_9681);
xnor UO_900 (O_900,N_9585,N_9947);
or UO_901 (O_901,N_9687,N_9683);
or UO_902 (O_902,N_9797,N_9674);
or UO_903 (O_903,N_9735,N_9505);
nor UO_904 (O_904,N_9641,N_9930);
nand UO_905 (O_905,N_9665,N_9687);
and UO_906 (O_906,N_9812,N_9672);
or UO_907 (O_907,N_9693,N_9716);
nor UO_908 (O_908,N_9940,N_9852);
and UO_909 (O_909,N_9567,N_9623);
or UO_910 (O_910,N_9679,N_9757);
and UO_911 (O_911,N_9586,N_9577);
and UO_912 (O_912,N_9532,N_9590);
or UO_913 (O_913,N_9700,N_9959);
and UO_914 (O_914,N_9778,N_9957);
or UO_915 (O_915,N_9553,N_9657);
nor UO_916 (O_916,N_9845,N_9976);
xor UO_917 (O_917,N_9692,N_9696);
nor UO_918 (O_918,N_9691,N_9503);
nand UO_919 (O_919,N_9504,N_9995);
or UO_920 (O_920,N_9943,N_9621);
nor UO_921 (O_921,N_9513,N_9652);
nor UO_922 (O_922,N_9819,N_9808);
and UO_923 (O_923,N_9623,N_9647);
nor UO_924 (O_924,N_9680,N_9516);
nor UO_925 (O_925,N_9815,N_9804);
and UO_926 (O_926,N_9727,N_9558);
or UO_927 (O_927,N_9682,N_9565);
and UO_928 (O_928,N_9780,N_9525);
nand UO_929 (O_929,N_9682,N_9719);
and UO_930 (O_930,N_9852,N_9766);
and UO_931 (O_931,N_9724,N_9879);
nand UO_932 (O_932,N_9894,N_9646);
nand UO_933 (O_933,N_9761,N_9533);
or UO_934 (O_934,N_9955,N_9813);
and UO_935 (O_935,N_9746,N_9989);
or UO_936 (O_936,N_9574,N_9835);
or UO_937 (O_937,N_9810,N_9915);
and UO_938 (O_938,N_9853,N_9779);
nor UO_939 (O_939,N_9574,N_9623);
and UO_940 (O_940,N_9912,N_9514);
and UO_941 (O_941,N_9986,N_9853);
nor UO_942 (O_942,N_9671,N_9609);
nand UO_943 (O_943,N_9645,N_9596);
and UO_944 (O_944,N_9623,N_9992);
or UO_945 (O_945,N_9976,N_9893);
nand UO_946 (O_946,N_9643,N_9767);
and UO_947 (O_947,N_9866,N_9779);
and UO_948 (O_948,N_9618,N_9846);
and UO_949 (O_949,N_9522,N_9573);
or UO_950 (O_950,N_9780,N_9795);
nand UO_951 (O_951,N_9755,N_9970);
xnor UO_952 (O_952,N_9861,N_9813);
and UO_953 (O_953,N_9717,N_9685);
and UO_954 (O_954,N_9889,N_9912);
or UO_955 (O_955,N_9936,N_9553);
and UO_956 (O_956,N_9788,N_9950);
and UO_957 (O_957,N_9926,N_9611);
nand UO_958 (O_958,N_9505,N_9925);
nand UO_959 (O_959,N_9663,N_9808);
nor UO_960 (O_960,N_9768,N_9517);
and UO_961 (O_961,N_9564,N_9806);
nand UO_962 (O_962,N_9755,N_9959);
or UO_963 (O_963,N_9713,N_9724);
and UO_964 (O_964,N_9988,N_9664);
or UO_965 (O_965,N_9689,N_9991);
nand UO_966 (O_966,N_9760,N_9658);
or UO_967 (O_967,N_9787,N_9970);
or UO_968 (O_968,N_9660,N_9703);
and UO_969 (O_969,N_9743,N_9844);
or UO_970 (O_970,N_9641,N_9677);
nor UO_971 (O_971,N_9699,N_9762);
xor UO_972 (O_972,N_9622,N_9744);
nand UO_973 (O_973,N_9554,N_9682);
nor UO_974 (O_974,N_9904,N_9662);
nand UO_975 (O_975,N_9762,N_9648);
nor UO_976 (O_976,N_9880,N_9802);
or UO_977 (O_977,N_9879,N_9628);
nor UO_978 (O_978,N_9594,N_9593);
nand UO_979 (O_979,N_9971,N_9954);
xnor UO_980 (O_980,N_9653,N_9589);
and UO_981 (O_981,N_9537,N_9642);
nand UO_982 (O_982,N_9501,N_9660);
nor UO_983 (O_983,N_9823,N_9525);
and UO_984 (O_984,N_9511,N_9937);
and UO_985 (O_985,N_9691,N_9569);
xor UO_986 (O_986,N_9822,N_9593);
nor UO_987 (O_987,N_9641,N_9578);
nor UO_988 (O_988,N_9991,N_9894);
and UO_989 (O_989,N_9658,N_9597);
or UO_990 (O_990,N_9978,N_9807);
and UO_991 (O_991,N_9874,N_9771);
or UO_992 (O_992,N_9625,N_9585);
nand UO_993 (O_993,N_9962,N_9682);
or UO_994 (O_994,N_9553,N_9614);
or UO_995 (O_995,N_9823,N_9749);
and UO_996 (O_996,N_9651,N_9717);
and UO_997 (O_997,N_9897,N_9860);
nand UO_998 (O_998,N_9632,N_9829);
and UO_999 (O_999,N_9685,N_9855);
nand UO_1000 (O_1000,N_9718,N_9559);
and UO_1001 (O_1001,N_9738,N_9554);
or UO_1002 (O_1002,N_9813,N_9705);
nor UO_1003 (O_1003,N_9979,N_9752);
nor UO_1004 (O_1004,N_9752,N_9900);
or UO_1005 (O_1005,N_9604,N_9504);
nand UO_1006 (O_1006,N_9860,N_9607);
and UO_1007 (O_1007,N_9525,N_9659);
nor UO_1008 (O_1008,N_9527,N_9581);
nor UO_1009 (O_1009,N_9813,N_9698);
and UO_1010 (O_1010,N_9735,N_9508);
nor UO_1011 (O_1011,N_9684,N_9615);
and UO_1012 (O_1012,N_9584,N_9572);
nand UO_1013 (O_1013,N_9997,N_9838);
xor UO_1014 (O_1014,N_9561,N_9734);
or UO_1015 (O_1015,N_9583,N_9825);
and UO_1016 (O_1016,N_9502,N_9958);
nand UO_1017 (O_1017,N_9775,N_9760);
nor UO_1018 (O_1018,N_9858,N_9605);
nor UO_1019 (O_1019,N_9816,N_9643);
nand UO_1020 (O_1020,N_9897,N_9535);
nand UO_1021 (O_1021,N_9703,N_9667);
and UO_1022 (O_1022,N_9603,N_9629);
or UO_1023 (O_1023,N_9677,N_9826);
xor UO_1024 (O_1024,N_9740,N_9581);
xor UO_1025 (O_1025,N_9653,N_9706);
nand UO_1026 (O_1026,N_9907,N_9562);
nor UO_1027 (O_1027,N_9557,N_9947);
and UO_1028 (O_1028,N_9669,N_9619);
xor UO_1029 (O_1029,N_9821,N_9989);
and UO_1030 (O_1030,N_9515,N_9872);
and UO_1031 (O_1031,N_9687,N_9981);
and UO_1032 (O_1032,N_9697,N_9565);
and UO_1033 (O_1033,N_9580,N_9724);
nand UO_1034 (O_1034,N_9593,N_9531);
and UO_1035 (O_1035,N_9606,N_9612);
nand UO_1036 (O_1036,N_9720,N_9664);
nand UO_1037 (O_1037,N_9605,N_9670);
nand UO_1038 (O_1038,N_9685,N_9652);
xnor UO_1039 (O_1039,N_9911,N_9978);
or UO_1040 (O_1040,N_9925,N_9708);
and UO_1041 (O_1041,N_9713,N_9745);
nand UO_1042 (O_1042,N_9888,N_9928);
nand UO_1043 (O_1043,N_9651,N_9791);
nor UO_1044 (O_1044,N_9900,N_9835);
nor UO_1045 (O_1045,N_9676,N_9861);
and UO_1046 (O_1046,N_9785,N_9935);
or UO_1047 (O_1047,N_9940,N_9826);
nor UO_1048 (O_1048,N_9604,N_9869);
or UO_1049 (O_1049,N_9526,N_9989);
nand UO_1050 (O_1050,N_9639,N_9627);
nor UO_1051 (O_1051,N_9862,N_9951);
or UO_1052 (O_1052,N_9741,N_9791);
or UO_1053 (O_1053,N_9822,N_9563);
or UO_1054 (O_1054,N_9551,N_9688);
and UO_1055 (O_1055,N_9713,N_9982);
nor UO_1056 (O_1056,N_9772,N_9882);
nor UO_1057 (O_1057,N_9621,N_9678);
nand UO_1058 (O_1058,N_9981,N_9669);
or UO_1059 (O_1059,N_9821,N_9827);
nand UO_1060 (O_1060,N_9904,N_9681);
and UO_1061 (O_1061,N_9878,N_9928);
nor UO_1062 (O_1062,N_9659,N_9790);
xnor UO_1063 (O_1063,N_9695,N_9772);
nand UO_1064 (O_1064,N_9774,N_9893);
xnor UO_1065 (O_1065,N_9745,N_9657);
or UO_1066 (O_1066,N_9738,N_9849);
nand UO_1067 (O_1067,N_9836,N_9574);
and UO_1068 (O_1068,N_9748,N_9537);
and UO_1069 (O_1069,N_9821,N_9851);
or UO_1070 (O_1070,N_9546,N_9883);
and UO_1071 (O_1071,N_9980,N_9642);
nor UO_1072 (O_1072,N_9935,N_9875);
nand UO_1073 (O_1073,N_9879,N_9826);
xnor UO_1074 (O_1074,N_9890,N_9677);
nor UO_1075 (O_1075,N_9778,N_9763);
or UO_1076 (O_1076,N_9514,N_9523);
nand UO_1077 (O_1077,N_9756,N_9775);
nor UO_1078 (O_1078,N_9850,N_9906);
or UO_1079 (O_1079,N_9569,N_9897);
or UO_1080 (O_1080,N_9767,N_9584);
and UO_1081 (O_1081,N_9874,N_9858);
nor UO_1082 (O_1082,N_9527,N_9787);
and UO_1083 (O_1083,N_9872,N_9992);
or UO_1084 (O_1084,N_9508,N_9803);
or UO_1085 (O_1085,N_9581,N_9833);
and UO_1086 (O_1086,N_9628,N_9919);
nor UO_1087 (O_1087,N_9513,N_9729);
xor UO_1088 (O_1088,N_9632,N_9619);
or UO_1089 (O_1089,N_9800,N_9782);
and UO_1090 (O_1090,N_9700,N_9721);
nand UO_1091 (O_1091,N_9943,N_9558);
or UO_1092 (O_1092,N_9659,N_9916);
or UO_1093 (O_1093,N_9796,N_9783);
or UO_1094 (O_1094,N_9959,N_9587);
nand UO_1095 (O_1095,N_9708,N_9661);
and UO_1096 (O_1096,N_9529,N_9897);
nor UO_1097 (O_1097,N_9635,N_9790);
nor UO_1098 (O_1098,N_9504,N_9970);
or UO_1099 (O_1099,N_9631,N_9867);
and UO_1100 (O_1100,N_9568,N_9707);
nand UO_1101 (O_1101,N_9608,N_9604);
and UO_1102 (O_1102,N_9720,N_9932);
or UO_1103 (O_1103,N_9610,N_9531);
xor UO_1104 (O_1104,N_9641,N_9816);
xnor UO_1105 (O_1105,N_9932,N_9853);
or UO_1106 (O_1106,N_9565,N_9901);
and UO_1107 (O_1107,N_9938,N_9594);
nand UO_1108 (O_1108,N_9606,N_9994);
nor UO_1109 (O_1109,N_9520,N_9688);
nand UO_1110 (O_1110,N_9995,N_9983);
and UO_1111 (O_1111,N_9553,N_9952);
or UO_1112 (O_1112,N_9871,N_9804);
xnor UO_1113 (O_1113,N_9522,N_9646);
nor UO_1114 (O_1114,N_9740,N_9607);
or UO_1115 (O_1115,N_9533,N_9573);
nor UO_1116 (O_1116,N_9587,N_9545);
nand UO_1117 (O_1117,N_9936,N_9605);
and UO_1118 (O_1118,N_9744,N_9912);
and UO_1119 (O_1119,N_9778,N_9668);
and UO_1120 (O_1120,N_9850,N_9665);
or UO_1121 (O_1121,N_9600,N_9747);
and UO_1122 (O_1122,N_9995,N_9772);
nor UO_1123 (O_1123,N_9513,N_9639);
and UO_1124 (O_1124,N_9662,N_9801);
and UO_1125 (O_1125,N_9533,N_9981);
and UO_1126 (O_1126,N_9975,N_9704);
and UO_1127 (O_1127,N_9642,N_9996);
xor UO_1128 (O_1128,N_9689,N_9679);
xor UO_1129 (O_1129,N_9554,N_9703);
and UO_1130 (O_1130,N_9676,N_9786);
and UO_1131 (O_1131,N_9686,N_9841);
or UO_1132 (O_1132,N_9859,N_9655);
and UO_1133 (O_1133,N_9997,N_9677);
or UO_1134 (O_1134,N_9891,N_9723);
nor UO_1135 (O_1135,N_9698,N_9547);
nand UO_1136 (O_1136,N_9992,N_9896);
and UO_1137 (O_1137,N_9920,N_9691);
xor UO_1138 (O_1138,N_9570,N_9926);
xor UO_1139 (O_1139,N_9982,N_9622);
or UO_1140 (O_1140,N_9992,N_9853);
nand UO_1141 (O_1141,N_9693,N_9854);
nor UO_1142 (O_1142,N_9871,N_9728);
and UO_1143 (O_1143,N_9868,N_9864);
nand UO_1144 (O_1144,N_9833,N_9519);
nor UO_1145 (O_1145,N_9871,N_9918);
or UO_1146 (O_1146,N_9716,N_9822);
xnor UO_1147 (O_1147,N_9912,N_9647);
or UO_1148 (O_1148,N_9568,N_9567);
nor UO_1149 (O_1149,N_9918,N_9943);
nand UO_1150 (O_1150,N_9773,N_9541);
nor UO_1151 (O_1151,N_9750,N_9749);
nor UO_1152 (O_1152,N_9968,N_9507);
and UO_1153 (O_1153,N_9942,N_9604);
nand UO_1154 (O_1154,N_9610,N_9694);
and UO_1155 (O_1155,N_9941,N_9610);
and UO_1156 (O_1156,N_9966,N_9570);
nand UO_1157 (O_1157,N_9806,N_9677);
and UO_1158 (O_1158,N_9664,N_9620);
and UO_1159 (O_1159,N_9820,N_9671);
xor UO_1160 (O_1160,N_9747,N_9604);
or UO_1161 (O_1161,N_9505,N_9993);
and UO_1162 (O_1162,N_9701,N_9800);
or UO_1163 (O_1163,N_9872,N_9789);
nor UO_1164 (O_1164,N_9757,N_9571);
nand UO_1165 (O_1165,N_9765,N_9694);
and UO_1166 (O_1166,N_9769,N_9778);
xnor UO_1167 (O_1167,N_9745,N_9631);
and UO_1168 (O_1168,N_9877,N_9583);
and UO_1169 (O_1169,N_9635,N_9522);
or UO_1170 (O_1170,N_9712,N_9514);
or UO_1171 (O_1171,N_9750,N_9706);
xnor UO_1172 (O_1172,N_9797,N_9583);
or UO_1173 (O_1173,N_9584,N_9658);
or UO_1174 (O_1174,N_9745,N_9651);
nand UO_1175 (O_1175,N_9641,N_9588);
or UO_1176 (O_1176,N_9658,N_9844);
and UO_1177 (O_1177,N_9574,N_9614);
xnor UO_1178 (O_1178,N_9866,N_9999);
nor UO_1179 (O_1179,N_9780,N_9515);
or UO_1180 (O_1180,N_9953,N_9674);
xor UO_1181 (O_1181,N_9791,N_9889);
nand UO_1182 (O_1182,N_9864,N_9977);
nand UO_1183 (O_1183,N_9714,N_9744);
xnor UO_1184 (O_1184,N_9624,N_9774);
nor UO_1185 (O_1185,N_9876,N_9999);
xor UO_1186 (O_1186,N_9626,N_9701);
nand UO_1187 (O_1187,N_9561,N_9942);
nor UO_1188 (O_1188,N_9636,N_9740);
nand UO_1189 (O_1189,N_9975,N_9886);
xor UO_1190 (O_1190,N_9633,N_9678);
nand UO_1191 (O_1191,N_9785,N_9694);
nor UO_1192 (O_1192,N_9773,N_9620);
nand UO_1193 (O_1193,N_9903,N_9731);
nor UO_1194 (O_1194,N_9642,N_9991);
nor UO_1195 (O_1195,N_9745,N_9562);
or UO_1196 (O_1196,N_9850,N_9689);
nor UO_1197 (O_1197,N_9578,N_9570);
or UO_1198 (O_1198,N_9965,N_9864);
or UO_1199 (O_1199,N_9813,N_9674);
or UO_1200 (O_1200,N_9853,N_9570);
and UO_1201 (O_1201,N_9933,N_9642);
nor UO_1202 (O_1202,N_9996,N_9636);
nor UO_1203 (O_1203,N_9518,N_9655);
nand UO_1204 (O_1204,N_9971,N_9881);
or UO_1205 (O_1205,N_9514,N_9744);
or UO_1206 (O_1206,N_9797,N_9798);
nand UO_1207 (O_1207,N_9932,N_9601);
nor UO_1208 (O_1208,N_9548,N_9924);
nand UO_1209 (O_1209,N_9686,N_9730);
nand UO_1210 (O_1210,N_9512,N_9958);
or UO_1211 (O_1211,N_9526,N_9531);
nor UO_1212 (O_1212,N_9931,N_9829);
nand UO_1213 (O_1213,N_9835,N_9764);
xnor UO_1214 (O_1214,N_9674,N_9852);
nor UO_1215 (O_1215,N_9514,N_9977);
and UO_1216 (O_1216,N_9745,N_9625);
or UO_1217 (O_1217,N_9995,N_9572);
nor UO_1218 (O_1218,N_9655,N_9605);
nand UO_1219 (O_1219,N_9784,N_9894);
and UO_1220 (O_1220,N_9703,N_9586);
and UO_1221 (O_1221,N_9739,N_9506);
nor UO_1222 (O_1222,N_9906,N_9879);
and UO_1223 (O_1223,N_9979,N_9971);
nor UO_1224 (O_1224,N_9824,N_9565);
or UO_1225 (O_1225,N_9597,N_9896);
xnor UO_1226 (O_1226,N_9746,N_9534);
nor UO_1227 (O_1227,N_9932,N_9699);
nand UO_1228 (O_1228,N_9588,N_9573);
or UO_1229 (O_1229,N_9615,N_9525);
nor UO_1230 (O_1230,N_9857,N_9757);
nand UO_1231 (O_1231,N_9777,N_9989);
nand UO_1232 (O_1232,N_9760,N_9927);
and UO_1233 (O_1233,N_9934,N_9896);
nor UO_1234 (O_1234,N_9573,N_9876);
nor UO_1235 (O_1235,N_9504,N_9892);
and UO_1236 (O_1236,N_9711,N_9693);
nor UO_1237 (O_1237,N_9687,N_9551);
and UO_1238 (O_1238,N_9772,N_9991);
and UO_1239 (O_1239,N_9647,N_9640);
nand UO_1240 (O_1240,N_9843,N_9556);
xnor UO_1241 (O_1241,N_9794,N_9650);
nand UO_1242 (O_1242,N_9599,N_9782);
or UO_1243 (O_1243,N_9566,N_9534);
nor UO_1244 (O_1244,N_9981,N_9975);
nor UO_1245 (O_1245,N_9853,N_9972);
xnor UO_1246 (O_1246,N_9687,N_9782);
nor UO_1247 (O_1247,N_9817,N_9758);
nor UO_1248 (O_1248,N_9918,N_9767);
nor UO_1249 (O_1249,N_9547,N_9918);
and UO_1250 (O_1250,N_9985,N_9718);
nand UO_1251 (O_1251,N_9523,N_9935);
and UO_1252 (O_1252,N_9930,N_9611);
nor UO_1253 (O_1253,N_9659,N_9717);
xor UO_1254 (O_1254,N_9608,N_9582);
or UO_1255 (O_1255,N_9863,N_9928);
and UO_1256 (O_1256,N_9560,N_9819);
or UO_1257 (O_1257,N_9572,N_9735);
nor UO_1258 (O_1258,N_9800,N_9840);
nand UO_1259 (O_1259,N_9562,N_9819);
nand UO_1260 (O_1260,N_9606,N_9689);
nand UO_1261 (O_1261,N_9861,N_9799);
nand UO_1262 (O_1262,N_9829,N_9575);
or UO_1263 (O_1263,N_9598,N_9581);
nor UO_1264 (O_1264,N_9703,N_9893);
and UO_1265 (O_1265,N_9725,N_9869);
and UO_1266 (O_1266,N_9927,N_9837);
nor UO_1267 (O_1267,N_9746,N_9700);
and UO_1268 (O_1268,N_9774,N_9653);
or UO_1269 (O_1269,N_9570,N_9999);
and UO_1270 (O_1270,N_9951,N_9501);
or UO_1271 (O_1271,N_9950,N_9852);
and UO_1272 (O_1272,N_9745,N_9836);
and UO_1273 (O_1273,N_9690,N_9740);
and UO_1274 (O_1274,N_9995,N_9915);
or UO_1275 (O_1275,N_9631,N_9554);
and UO_1276 (O_1276,N_9822,N_9624);
or UO_1277 (O_1277,N_9903,N_9941);
nand UO_1278 (O_1278,N_9652,N_9773);
xor UO_1279 (O_1279,N_9989,N_9952);
or UO_1280 (O_1280,N_9675,N_9617);
xnor UO_1281 (O_1281,N_9554,N_9717);
or UO_1282 (O_1282,N_9653,N_9800);
nand UO_1283 (O_1283,N_9785,N_9985);
or UO_1284 (O_1284,N_9756,N_9849);
nor UO_1285 (O_1285,N_9932,N_9742);
and UO_1286 (O_1286,N_9541,N_9741);
nor UO_1287 (O_1287,N_9632,N_9916);
xor UO_1288 (O_1288,N_9510,N_9767);
and UO_1289 (O_1289,N_9596,N_9545);
xor UO_1290 (O_1290,N_9762,N_9987);
or UO_1291 (O_1291,N_9787,N_9997);
nand UO_1292 (O_1292,N_9585,N_9690);
nand UO_1293 (O_1293,N_9705,N_9990);
or UO_1294 (O_1294,N_9635,N_9700);
nand UO_1295 (O_1295,N_9920,N_9578);
nor UO_1296 (O_1296,N_9696,N_9864);
nor UO_1297 (O_1297,N_9950,N_9634);
and UO_1298 (O_1298,N_9943,N_9871);
and UO_1299 (O_1299,N_9852,N_9945);
and UO_1300 (O_1300,N_9579,N_9611);
or UO_1301 (O_1301,N_9505,N_9817);
nand UO_1302 (O_1302,N_9825,N_9540);
xnor UO_1303 (O_1303,N_9600,N_9820);
and UO_1304 (O_1304,N_9910,N_9596);
and UO_1305 (O_1305,N_9564,N_9577);
and UO_1306 (O_1306,N_9782,N_9878);
nor UO_1307 (O_1307,N_9620,N_9934);
xor UO_1308 (O_1308,N_9820,N_9659);
or UO_1309 (O_1309,N_9652,N_9868);
xor UO_1310 (O_1310,N_9782,N_9633);
and UO_1311 (O_1311,N_9559,N_9524);
nor UO_1312 (O_1312,N_9658,N_9560);
nand UO_1313 (O_1313,N_9706,N_9528);
xnor UO_1314 (O_1314,N_9895,N_9858);
and UO_1315 (O_1315,N_9650,N_9745);
nor UO_1316 (O_1316,N_9675,N_9961);
or UO_1317 (O_1317,N_9672,N_9652);
nor UO_1318 (O_1318,N_9845,N_9630);
nand UO_1319 (O_1319,N_9567,N_9817);
and UO_1320 (O_1320,N_9764,N_9520);
or UO_1321 (O_1321,N_9775,N_9833);
nand UO_1322 (O_1322,N_9772,N_9574);
nand UO_1323 (O_1323,N_9702,N_9717);
or UO_1324 (O_1324,N_9681,N_9717);
or UO_1325 (O_1325,N_9571,N_9750);
xor UO_1326 (O_1326,N_9643,N_9923);
or UO_1327 (O_1327,N_9645,N_9505);
and UO_1328 (O_1328,N_9795,N_9629);
and UO_1329 (O_1329,N_9752,N_9741);
and UO_1330 (O_1330,N_9741,N_9947);
and UO_1331 (O_1331,N_9771,N_9816);
nor UO_1332 (O_1332,N_9793,N_9993);
and UO_1333 (O_1333,N_9876,N_9705);
and UO_1334 (O_1334,N_9925,N_9962);
nand UO_1335 (O_1335,N_9802,N_9675);
or UO_1336 (O_1336,N_9500,N_9984);
or UO_1337 (O_1337,N_9814,N_9522);
xnor UO_1338 (O_1338,N_9598,N_9818);
or UO_1339 (O_1339,N_9873,N_9548);
xor UO_1340 (O_1340,N_9798,N_9906);
nor UO_1341 (O_1341,N_9679,N_9557);
xor UO_1342 (O_1342,N_9898,N_9995);
and UO_1343 (O_1343,N_9807,N_9746);
and UO_1344 (O_1344,N_9610,N_9627);
and UO_1345 (O_1345,N_9872,N_9743);
nand UO_1346 (O_1346,N_9524,N_9829);
nand UO_1347 (O_1347,N_9794,N_9822);
nor UO_1348 (O_1348,N_9873,N_9894);
nand UO_1349 (O_1349,N_9605,N_9616);
nand UO_1350 (O_1350,N_9633,N_9651);
nand UO_1351 (O_1351,N_9849,N_9852);
and UO_1352 (O_1352,N_9917,N_9690);
xor UO_1353 (O_1353,N_9553,N_9959);
or UO_1354 (O_1354,N_9669,N_9610);
nand UO_1355 (O_1355,N_9585,N_9971);
nor UO_1356 (O_1356,N_9861,N_9992);
nor UO_1357 (O_1357,N_9560,N_9987);
and UO_1358 (O_1358,N_9700,N_9758);
and UO_1359 (O_1359,N_9649,N_9770);
nand UO_1360 (O_1360,N_9986,N_9913);
or UO_1361 (O_1361,N_9554,N_9920);
and UO_1362 (O_1362,N_9696,N_9926);
xor UO_1363 (O_1363,N_9849,N_9645);
or UO_1364 (O_1364,N_9688,N_9671);
xnor UO_1365 (O_1365,N_9923,N_9765);
nand UO_1366 (O_1366,N_9525,N_9805);
or UO_1367 (O_1367,N_9504,N_9624);
nor UO_1368 (O_1368,N_9627,N_9843);
nor UO_1369 (O_1369,N_9593,N_9949);
and UO_1370 (O_1370,N_9726,N_9759);
or UO_1371 (O_1371,N_9564,N_9905);
and UO_1372 (O_1372,N_9972,N_9580);
xnor UO_1373 (O_1373,N_9621,N_9684);
or UO_1374 (O_1374,N_9605,N_9931);
nand UO_1375 (O_1375,N_9810,N_9762);
and UO_1376 (O_1376,N_9934,N_9956);
nand UO_1377 (O_1377,N_9587,N_9681);
and UO_1378 (O_1378,N_9606,N_9598);
nor UO_1379 (O_1379,N_9559,N_9898);
and UO_1380 (O_1380,N_9936,N_9606);
and UO_1381 (O_1381,N_9883,N_9719);
or UO_1382 (O_1382,N_9526,N_9770);
nand UO_1383 (O_1383,N_9606,N_9674);
nand UO_1384 (O_1384,N_9991,N_9658);
xnor UO_1385 (O_1385,N_9664,N_9776);
and UO_1386 (O_1386,N_9629,N_9752);
or UO_1387 (O_1387,N_9670,N_9984);
xor UO_1388 (O_1388,N_9552,N_9958);
or UO_1389 (O_1389,N_9635,N_9543);
or UO_1390 (O_1390,N_9842,N_9676);
nor UO_1391 (O_1391,N_9701,N_9678);
nand UO_1392 (O_1392,N_9692,N_9632);
or UO_1393 (O_1393,N_9805,N_9972);
or UO_1394 (O_1394,N_9565,N_9717);
nor UO_1395 (O_1395,N_9971,N_9505);
nor UO_1396 (O_1396,N_9557,N_9934);
xnor UO_1397 (O_1397,N_9585,N_9734);
and UO_1398 (O_1398,N_9697,N_9623);
xor UO_1399 (O_1399,N_9997,N_9527);
nand UO_1400 (O_1400,N_9562,N_9706);
or UO_1401 (O_1401,N_9788,N_9567);
or UO_1402 (O_1402,N_9658,N_9565);
or UO_1403 (O_1403,N_9786,N_9862);
and UO_1404 (O_1404,N_9944,N_9534);
nand UO_1405 (O_1405,N_9897,N_9921);
nor UO_1406 (O_1406,N_9594,N_9626);
xor UO_1407 (O_1407,N_9656,N_9681);
xnor UO_1408 (O_1408,N_9796,N_9638);
nand UO_1409 (O_1409,N_9801,N_9524);
xnor UO_1410 (O_1410,N_9996,N_9867);
nor UO_1411 (O_1411,N_9818,N_9853);
nand UO_1412 (O_1412,N_9631,N_9852);
and UO_1413 (O_1413,N_9588,N_9804);
nor UO_1414 (O_1414,N_9635,N_9677);
nor UO_1415 (O_1415,N_9527,N_9688);
xor UO_1416 (O_1416,N_9823,N_9885);
and UO_1417 (O_1417,N_9593,N_9895);
nor UO_1418 (O_1418,N_9524,N_9880);
or UO_1419 (O_1419,N_9745,N_9826);
and UO_1420 (O_1420,N_9803,N_9783);
nand UO_1421 (O_1421,N_9858,N_9869);
nor UO_1422 (O_1422,N_9813,N_9515);
nor UO_1423 (O_1423,N_9680,N_9768);
or UO_1424 (O_1424,N_9720,N_9769);
or UO_1425 (O_1425,N_9904,N_9525);
or UO_1426 (O_1426,N_9545,N_9868);
nor UO_1427 (O_1427,N_9810,N_9795);
or UO_1428 (O_1428,N_9826,N_9667);
xor UO_1429 (O_1429,N_9852,N_9938);
nor UO_1430 (O_1430,N_9720,N_9576);
or UO_1431 (O_1431,N_9683,N_9872);
nor UO_1432 (O_1432,N_9665,N_9755);
nand UO_1433 (O_1433,N_9688,N_9840);
xor UO_1434 (O_1434,N_9660,N_9533);
nand UO_1435 (O_1435,N_9695,N_9687);
xnor UO_1436 (O_1436,N_9888,N_9593);
nand UO_1437 (O_1437,N_9588,N_9734);
nand UO_1438 (O_1438,N_9662,N_9923);
nor UO_1439 (O_1439,N_9887,N_9968);
and UO_1440 (O_1440,N_9995,N_9873);
nand UO_1441 (O_1441,N_9708,N_9856);
nand UO_1442 (O_1442,N_9643,N_9685);
nor UO_1443 (O_1443,N_9878,N_9909);
nand UO_1444 (O_1444,N_9992,N_9733);
nor UO_1445 (O_1445,N_9977,N_9664);
and UO_1446 (O_1446,N_9763,N_9586);
and UO_1447 (O_1447,N_9712,N_9693);
and UO_1448 (O_1448,N_9888,N_9586);
and UO_1449 (O_1449,N_9758,N_9702);
xor UO_1450 (O_1450,N_9775,N_9998);
nor UO_1451 (O_1451,N_9637,N_9956);
xnor UO_1452 (O_1452,N_9932,N_9722);
or UO_1453 (O_1453,N_9717,N_9830);
nand UO_1454 (O_1454,N_9686,N_9787);
or UO_1455 (O_1455,N_9975,N_9608);
and UO_1456 (O_1456,N_9916,N_9611);
xor UO_1457 (O_1457,N_9978,N_9878);
nor UO_1458 (O_1458,N_9994,N_9800);
and UO_1459 (O_1459,N_9900,N_9673);
or UO_1460 (O_1460,N_9517,N_9643);
and UO_1461 (O_1461,N_9825,N_9653);
or UO_1462 (O_1462,N_9629,N_9899);
xor UO_1463 (O_1463,N_9555,N_9923);
nor UO_1464 (O_1464,N_9739,N_9556);
nor UO_1465 (O_1465,N_9704,N_9913);
xnor UO_1466 (O_1466,N_9959,N_9600);
nand UO_1467 (O_1467,N_9946,N_9725);
nor UO_1468 (O_1468,N_9567,N_9641);
or UO_1469 (O_1469,N_9891,N_9623);
xnor UO_1470 (O_1470,N_9903,N_9629);
or UO_1471 (O_1471,N_9880,N_9828);
or UO_1472 (O_1472,N_9973,N_9907);
or UO_1473 (O_1473,N_9576,N_9668);
and UO_1474 (O_1474,N_9547,N_9733);
and UO_1475 (O_1475,N_9520,N_9875);
and UO_1476 (O_1476,N_9617,N_9732);
and UO_1477 (O_1477,N_9800,N_9567);
and UO_1478 (O_1478,N_9778,N_9722);
nor UO_1479 (O_1479,N_9634,N_9865);
and UO_1480 (O_1480,N_9737,N_9583);
or UO_1481 (O_1481,N_9819,N_9998);
nand UO_1482 (O_1482,N_9841,N_9807);
nand UO_1483 (O_1483,N_9593,N_9555);
or UO_1484 (O_1484,N_9684,N_9542);
nor UO_1485 (O_1485,N_9872,N_9875);
nor UO_1486 (O_1486,N_9932,N_9745);
nor UO_1487 (O_1487,N_9600,N_9858);
xor UO_1488 (O_1488,N_9872,N_9758);
and UO_1489 (O_1489,N_9517,N_9620);
and UO_1490 (O_1490,N_9831,N_9783);
or UO_1491 (O_1491,N_9903,N_9811);
nor UO_1492 (O_1492,N_9813,N_9541);
nor UO_1493 (O_1493,N_9719,N_9587);
or UO_1494 (O_1494,N_9665,N_9940);
nor UO_1495 (O_1495,N_9760,N_9948);
xor UO_1496 (O_1496,N_9600,N_9641);
nand UO_1497 (O_1497,N_9958,N_9652);
or UO_1498 (O_1498,N_9897,N_9614);
or UO_1499 (O_1499,N_9583,N_9853);
endmodule