module basic_500_3000_500_6_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_335,In_122);
nor U1 (N_1,In_334,In_473);
xor U2 (N_2,In_248,In_109);
nand U3 (N_3,In_485,In_167);
nand U4 (N_4,In_216,In_209);
nand U5 (N_5,In_2,In_117);
and U6 (N_6,In_446,In_38);
or U7 (N_7,In_25,In_19);
nand U8 (N_8,In_72,In_3);
nor U9 (N_9,In_361,In_272);
xnor U10 (N_10,In_83,In_244);
or U11 (N_11,In_47,In_342);
and U12 (N_12,In_292,In_429);
nand U13 (N_13,In_252,In_291);
xor U14 (N_14,In_424,In_145);
or U15 (N_15,In_368,In_389);
nand U16 (N_16,In_377,In_360);
nand U17 (N_17,In_298,In_385);
nor U18 (N_18,In_493,In_12);
or U19 (N_19,In_285,In_181);
xor U20 (N_20,In_128,In_137);
nand U21 (N_21,In_226,In_266);
nand U22 (N_22,In_449,In_198);
nand U23 (N_23,In_238,In_401);
or U24 (N_24,In_444,In_460);
nand U25 (N_25,In_75,In_118);
or U26 (N_26,In_228,In_270);
nand U27 (N_27,In_210,In_410);
nor U28 (N_28,In_315,In_139);
and U29 (N_29,In_462,In_231);
or U30 (N_30,In_400,In_195);
or U31 (N_31,In_146,In_409);
nand U32 (N_32,In_77,In_290);
and U33 (N_33,In_459,In_352);
or U34 (N_34,In_476,In_204);
or U35 (N_35,In_61,In_15);
and U36 (N_36,In_14,In_323);
nand U37 (N_37,In_324,In_229);
xor U38 (N_38,In_1,In_156);
xor U39 (N_39,In_293,In_168);
or U40 (N_40,In_218,In_163);
nor U41 (N_41,In_397,In_84);
or U42 (N_42,In_375,In_121);
and U43 (N_43,In_354,In_297);
and U44 (N_44,In_472,In_454);
xnor U45 (N_45,In_470,In_332);
nor U46 (N_46,In_382,In_431);
nor U47 (N_47,In_379,In_349);
nand U48 (N_48,In_126,In_65);
xor U49 (N_49,In_144,In_249);
xnor U50 (N_50,In_213,In_246);
xor U51 (N_51,In_456,In_461);
and U52 (N_52,In_189,In_8);
nor U53 (N_53,In_46,In_414);
nor U54 (N_54,In_458,In_316);
nor U55 (N_55,In_164,In_225);
xor U56 (N_56,In_135,In_176);
nor U57 (N_57,In_363,In_366);
xnor U58 (N_58,In_419,In_495);
nor U59 (N_59,In_96,In_173);
xnor U60 (N_60,In_11,In_346);
or U61 (N_61,In_388,In_378);
and U62 (N_62,In_203,In_27);
nor U63 (N_63,In_471,In_196);
nand U64 (N_64,In_275,In_74);
and U65 (N_65,In_4,In_70);
or U66 (N_66,In_24,In_237);
nor U67 (N_67,In_170,In_442);
xor U68 (N_68,In_387,In_104);
nor U69 (N_69,In_386,In_212);
xor U70 (N_70,In_234,In_50);
or U71 (N_71,In_450,In_439);
nor U72 (N_72,In_69,In_49);
xor U73 (N_73,In_344,In_131);
nand U74 (N_74,In_314,In_256);
and U75 (N_75,In_134,In_29);
and U76 (N_76,In_404,In_222);
nand U77 (N_77,In_488,In_205);
and U78 (N_78,In_66,In_331);
or U79 (N_79,In_60,In_464);
xnor U80 (N_80,In_261,In_182);
or U81 (N_81,In_0,In_381);
xnor U82 (N_82,In_183,In_311);
nor U83 (N_83,In_97,In_367);
nor U84 (N_84,In_100,In_227);
and U85 (N_85,In_423,In_408);
and U86 (N_86,In_34,In_341);
and U87 (N_87,In_465,In_257);
and U88 (N_88,In_482,In_294);
nor U89 (N_89,In_492,In_251);
and U90 (N_90,In_80,In_466);
or U91 (N_91,In_9,In_59);
and U92 (N_92,In_398,In_330);
xor U93 (N_93,In_197,In_158);
nor U94 (N_94,In_175,In_174);
and U95 (N_95,In_171,In_313);
xor U96 (N_96,In_265,In_347);
and U97 (N_97,In_299,In_87);
nand U98 (N_98,In_373,In_396);
or U99 (N_99,In_223,In_374);
or U100 (N_100,In_17,In_303);
nand U101 (N_101,In_108,In_151);
xor U102 (N_102,In_358,In_201);
and U103 (N_103,In_40,In_202);
and U104 (N_104,In_486,In_54);
and U105 (N_105,In_271,In_440);
and U106 (N_106,In_154,In_68);
xnor U107 (N_107,In_23,In_428);
nand U108 (N_108,In_190,In_242);
xnor U109 (N_109,In_160,In_129);
and U110 (N_110,In_76,In_165);
nor U111 (N_111,In_35,In_362);
and U112 (N_112,In_452,In_477);
nor U113 (N_113,In_399,In_498);
nor U114 (N_114,In_407,In_57);
and U115 (N_115,In_287,In_186);
nand U116 (N_116,In_430,In_411);
and U117 (N_117,In_451,In_425);
nor U118 (N_118,In_64,In_119);
nor U119 (N_119,In_309,In_112);
nand U120 (N_120,In_22,In_63);
nor U121 (N_121,In_107,In_105);
nand U122 (N_122,In_127,In_73);
and U123 (N_123,In_45,In_16);
nor U124 (N_124,In_353,In_130);
nor U125 (N_125,In_260,In_79);
xor U126 (N_126,In_21,In_269);
and U127 (N_127,In_113,In_274);
or U128 (N_128,In_51,In_81);
nand U129 (N_129,In_82,In_178);
nor U130 (N_130,In_253,In_336);
xnor U131 (N_131,In_364,In_337);
nor U132 (N_132,In_235,In_372);
nor U133 (N_133,In_71,In_243);
and U134 (N_134,In_282,In_427);
nand U135 (N_135,In_180,In_296);
or U136 (N_136,In_94,In_365);
nor U137 (N_137,In_95,In_172);
and U138 (N_138,In_191,In_88);
and U139 (N_139,In_207,In_489);
and U140 (N_140,In_217,In_371);
nor U141 (N_141,In_93,In_494);
xnor U142 (N_142,In_405,In_312);
xor U143 (N_143,In_255,In_115);
nand U144 (N_144,In_31,In_420);
and U145 (N_145,In_98,In_343);
nor U146 (N_146,In_125,In_41);
or U147 (N_147,In_149,In_447);
and U148 (N_148,In_491,In_267);
and U149 (N_149,In_280,In_13);
nor U150 (N_150,In_99,In_369);
or U151 (N_151,In_37,In_468);
or U152 (N_152,In_390,In_351);
xor U153 (N_153,In_141,In_478);
nor U154 (N_154,In_32,In_329);
xor U155 (N_155,In_62,In_91);
xor U156 (N_156,In_42,In_453);
or U157 (N_157,In_200,In_230);
or U158 (N_158,In_6,In_161);
and U159 (N_159,In_56,In_20);
nand U160 (N_160,In_469,In_277);
nand U161 (N_161,In_264,In_273);
or U162 (N_162,In_239,In_276);
nor U163 (N_163,In_421,In_10);
nor U164 (N_164,In_422,In_232);
and U165 (N_165,In_438,In_259);
nand U166 (N_166,In_480,In_263);
nor U167 (N_167,In_33,In_380);
and U168 (N_168,In_262,In_92);
or U169 (N_169,In_350,In_284);
nand U170 (N_170,In_184,In_30);
nor U171 (N_171,In_395,In_43);
nand U172 (N_172,In_339,In_384);
xor U173 (N_173,In_150,In_310);
or U174 (N_174,In_250,In_433);
nor U175 (N_175,In_124,In_67);
or U176 (N_176,In_441,In_245);
nand U177 (N_177,In_394,In_258);
or U178 (N_178,In_463,In_177);
xor U179 (N_179,In_221,In_357);
or U180 (N_180,In_110,In_162);
xnor U181 (N_181,In_53,In_123);
nand U182 (N_182,In_159,In_283);
nor U183 (N_183,In_153,In_355);
nand U184 (N_184,In_348,In_448);
xor U185 (N_185,In_187,In_481);
xnor U186 (N_186,In_338,In_236);
nor U187 (N_187,In_327,In_194);
nor U188 (N_188,In_215,In_157);
or U189 (N_189,In_320,In_148);
nor U190 (N_190,In_356,In_417);
or U191 (N_191,In_306,In_443);
nand U192 (N_192,In_208,In_457);
nand U193 (N_193,In_147,In_132);
nand U194 (N_194,In_326,In_90);
or U195 (N_195,In_305,In_302);
nand U196 (N_196,In_487,In_307);
and U197 (N_197,In_321,In_308);
and U198 (N_198,In_304,In_497);
nand U199 (N_199,In_211,In_152);
or U200 (N_200,In_418,In_188);
and U201 (N_201,In_426,In_142);
and U202 (N_202,In_78,In_55);
nor U203 (N_203,In_359,In_206);
or U204 (N_204,In_402,In_254);
nor U205 (N_205,In_467,In_328);
or U206 (N_206,In_474,In_301);
and U207 (N_207,In_101,In_415);
or U208 (N_208,In_490,In_475);
nand U209 (N_209,In_286,In_102);
nand U210 (N_210,In_289,In_383);
nand U211 (N_211,In_89,In_143);
nand U212 (N_212,In_241,In_240);
nor U213 (N_213,In_416,In_318);
and U214 (N_214,In_317,In_52);
nor U215 (N_215,In_28,In_333);
and U216 (N_216,In_295,In_484);
and U217 (N_217,In_39,In_412);
nor U218 (N_218,In_140,In_18);
or U219 (N_219,In_233,In_319);
or U220 (N_220,In_403,In_499);
xnor U221 (N_221,In_58,In_133);
nor U222 (N_222,In_413,In_278);
xor U223 (N_223,In_5,In_44);
or U224 (N_224,In_214,In_111);
xnor U225 (N_225,In_26,In_445);
nand U226 (N_226,In_220,In_483);
or U227 (N_227,In_85,In_391);
or U228 (N_228,In_322,In_36);
and U229 (N_229,In_392,In_86);
nand U230 (N_230,In_288,In_199);
nand U231 (N_231,In_166,In_432);
nand U232 (N_232,In_393,In_48);
nor U233 (N_233,In_437,In_455);
or U234 (N_234,In_345,In_370);
xnor U235 (N_235,In_192,In_179);
nand U236 (N_236,In_434,In_138);
nand U237 (N_237,In_155,In_479);
or U238 (N_238,In_268,In_7);
nand U239 (N_239,In_376,In_136);
nor U240 (N_240,In_496,In_340);
nand U241 (N_241,In_436,In_169);
and U242 (N_242,In_185,In_300);
xor U243 (N_243,In_219,In_435);
and U244 (N_244,In_406,In_193);
xnor U245 (N_245,In_103,In_325);
nor U246 (N_246,In_106,In_247);
nand U247 (N_247,In_116,In_114);
or U248 (N_248,In_279,In_281);
xnor U249 (N_249,In_224,In_120);
and U250 (N_250,In_382,In_407);
xor U251 (N_251,In_199,In_3);
xnor U252 (N_252,In_470,In_394);
and U253 (N_253,In_302,In_34);
nor U254 (N_254,In_302,In_164);
and U255 (N_255,In_308,In_150);
xor U256 (N_256,In_84,In_297);
or U257 (N_257,In_270,In_410);
xnor U258 (N_258,In_274,In_263);
and U259 (N_259,In_245,In_66);
nor U260 (N_260,In_493,In_377);
and U261 (N_261,In_237,In_25);
xnor U262 (N_262,In_399,In_248);
xnor U263 (N_263,In_50,In_403);
nand U264 (N_264,In_54,In_401);
xnor U265 (N_265,In_203,In_269);
nand U266 (N_266,In_291,In_236);
or U267 (N_267,In_19,In_358);
nand U268 (N_268,In_177,In_46);
nand U269 (N_269,In_281,In_388);
nand U270 (N_270,In_95,In_102);
xor U271 (N_271,In_441,In_124);
or U272 (N_272,In_405,In_331);
nor U273 (N_273,In_123,In_38);
xnor U274 (N_274,In_397,In_410);
nand U275 (N_275,In_312,In_204);
nand U276 (N_276,In_226,In_140);
xor U277 (N_277,In_117,In_453);
and U278 (N_278,In_476,In_151);
or U279 (N_279,In_490,In_282);
or U280 (N_280,In_1,In_409);
nor U281 (N_281,In_83,In_125);
nand U282 (N_282,In_109,In_299);
or U283 (N_283,In_13,In_355);
and U284 (N_284,In_170,In_291);
nor U285 (N_285,In_91,In_96);
nand U286 (N_286,In_128,In_488);
nand U287 (N_287,In_211,In_445);
nor U288 (N_288,In_225,In_148);
or U289 (N_289,In_365,In_194);
or U290 (N_290,In_43,In_401);
and U291 (N_291,In_377,In_389);
and U292 (N_292,In_79,In_432);
and U293 (N_293,In_223,In_127);
nand U294 (N_294,In_44,In_127);
xor U295 (N_295,In_106,In_374);
xor U296 (N_296,In_10,In_487);
or U297 (N_297,In_143,In_13);
or U298 (N_298,In_314,In_87);
and U299 (N_299,In_400,In_130);
and U300 (N_300,In_432,In_61);
nand U301 (N_301,In_353,In_160);
and U302 (N_302,In_318,In_12);
nand U303 (N_303,In_120,In_45);
and U304 (N_304,In_267,In_495);
xnor U305 (N_305,In_334,In_32);
nand U306 (N_306,In_494,In_392);
xnor U307 (N_307,In_220,In_210);
nor U308 (N_308,In_438,In_155);
nor U309 (N_309,In_57,In_296);
nand U310 (N_310,In_65,In_481);
or U311 (N_311,In_24,In_59);
or U312 (N_312,In_237,In_313);
nand U313 (N_313,In_429,In_381);
xnor U314 (N_314,In_159,In_237);
nand U315 (N_315,In_42,In_367);
or U316 (N_316,In_98,In_368);
nand U317 (N_317,In_412,In_282);
nor U318 (N_318,In_496,In_359);
xnor U319 (N_319,In_44,In_292);
nor U320 (N_320,In_253,In_291);
or U321 (N_321,In_409,In_376);
nand U322 (N_322,In_18,In_175);
xnor U323 (N_323,In_240,In_280);
nor U324 (N_324,In_404,In_469);
xor U325 (N_325,In_109,In_216);
xnor U326 (N_326,In_327,In_165);
nor U327 (N_327,In_401,In_153);
xor U328 (N_328,In_313,In_177);
nand U329 (N_329,In_169,In_285);
nand U330 (N_330,In_440,In_484);
xor U331 (N_331,In_453,In_212);
or U332 (N_332,In_496,In_188);
or U333 (N_333,In_198,In_303);
xor U334 (N_334,In_491,In_403);
nand U335 (N_335,In_180,In_215);
nand U336 (N_336,In_468,In_381);
and U337 (N_337,In_160,In_292);
xor U338 (N_338,In_279,In_299);
and U339 (N_339,In_399,In_56);
nand U340 (N_340,In_373,In_235);
nand U341 (N_341,In_138,In_199);
and U342 (N_342,In_227,In_215);
xor U343 (N_343,In_74,In_498);
and U344 (N_344,In_351,In_276);
nor U345 (N_345,In_62,In_297);
nor U346 (N_346,In_164,In_233);
or U347 (N_347,In_418,In_310);
xor U348 (N_348,In_265,In_340);
and U349 (N_349,In_207,In_365);
nand U350 (N_350,In_253,In_128);
or U351 (N_351,In_469,In_379);
nand U352 (N_352,In_100,In_61);
nor U353 (N_353,In_375,In_295);
nor U354 (N_354,In_452,In_472);
and U355 (N_355,In_438,In_32);
or U356 (N_356,In_105,In_441);
nand U357 (N_357,In_339,In_250);
or U358 (N_358,In_136,In_293);
or U359 (N_359,In_151,In_491);
and U360 (N_360,In_492,In_464);
xnor U361 (N_361,In_276,In_399);
nor U362 (N_362,In_254,In_183);
and U363 (N_363,In_440,In_214);
or U364 (N_364,In_37,In_393);
nor U365 (N_365,In_260,In_366);
xnor U366 (N_366,In_263,In_262);
or U367 (N_367,In_112,In_9);
or U368 (N_368,In_99,In_29);
nor U369 (N_369,In_146,In_230);
nor U370 (N_370,In_24,In_321);
nand U371 (N_371,In_161,In_0);
nor U372 (N_372,In_296,In_366);
nand U373 (N_373,In_279,In_223);
nand U374 (N_374,In_365,In_18);
or U375 (N_375,In_318,In_54);
xor U376 (N_376,In_475,In_236);
or U377 (N_377,In_96,In_81);
xnor U378 (N_378,In_26,In_304);
nor U379 (N_379,In_58,In_430);
nor U380 (N_380,In_125,In_315);
xor U381 (N_381,In_81,In_364);
or U382 (N_382,In_152,In_66);
and U383 (N_383,In_178,In_213);
nor U384 (N_384,In_116,In_261);
and U385 (N_385,In_12,In_42);
nor U386 (N_386,In_472,In_338);
and U387 (N_387,In_305,In_193);
nor U388 (N_388,In_31,In_216);
xor U389 (N_389,In_452,In_285);
nor U390 (N_390,In_215,In_241);
nor U391 (N_391,In_248,In_400);
or U392 (N_392,In_223,In_59);
nand U393 (N_393,In_359,In_219);
xnor U394 (N_394,In_205,In_80);
xnor U395 (N_395,In_446,In_476);
nand U396 (N_396,In_201,In_259);
and U397 (N_397,In_378,In_70);
or U398 (N_398,In_392,In_490);
or U399 (N_399,In_496,In_229);
nor U400 (N_400,In_254,In_415);
and U401 (N_401,In_368,In_93);
or U402 (N_402,In_151,In_242);
xnor U403 (N_403,In_128,In_104);
nor U404 (N_404,In_454,In_4);
xnor U405 (N_405,In_490,In_313);
xnor U406 (N_406,In_363,In_156);
and U407 (N_407,In_122,In_38);
or U408 (N_408,In_445,In_333);
or U409 (N_409,In_387,In_444);
or U410 (N_410,In_459,In_392);
and U411 (N_411,In_130,In_279);
or U412 (N_412,In_130,In_216);
nor U413 (N_413,In_315,In_229);
and U414 (N_414,In_235,In_498);
or U415 (N_415,In_498,In_298);
or U416 (N_416,In_79,In_207);
nand U417 (N_417,In_72,In_347);
and U418 (N_418,In_97,In_25);
xor U419 (N_419,In_266,In_260);
and U420 (N_420,In_249,In_498);
nand U421 (N_421,In_476,In_62);
or U422 (N_422,In_377,In_239);
xnor U423 (N_423,In_417,In_14);
and U424 (N_424,In_95,In_275);
or U425 (N_425,In_396,In_61);
or U426 (N_426,In_28,In_195);
and U427 (N_427,In_119,In_24);
or U428 (N_428,In_407,In_203);
nand U429 (N_429,In_228,In_72);
nand U430 (N_430,In_461,In_362);
nand U431 (N_431,In_171,In_464);
and U432 (N_432,In_284,In_358);
nand U433 (N_433,In_496,In_391);
nand U434 (N_434,In_449,In_487);
nand U435 (N_435,In_26,In_395);
nor U436 (N_436,In_253,In_148);
nor U437 (N_437,In_409,In_242);
or U438 (N_438,In_14,In_135);
xnor U439 (N_439,In_390,In_218);
nor U440 (N_440,In_473,In_272);
or U441 (N_441,In_277,In_30);
or U442 (N_442,In_362,In_277);
xor U443 (N_443,In_219,In_70);
nand U444 (N_444,In_58,In_282);
nor U445 (N_445,In_100,In_196);
or U446 (N_446,In_490,In_315);
nand U447 (N_447,In_14,In_358);
nor U448 (N_448,In_244,In_394);
or U449 (N_449,In_250,In_212);
and U450 (N_450,In_152,In_61);
and U451 (N_451,In_225,In_235);
nor U452 (N_452,In_132,In_178);
nor U453 (N_453,In_269,In_123);
xor U454 (N_454,In_220,In_411);
and U455 (N_455,In_368,In_135);
and U456 (N_456,In_327,In_310);
and U457 (N_457,In_14,In_258);
or U458 (N_458,In_496,In_140);
or U459 (N_459,In_194,In_34);
nand U460 (N_460,In_54,In_273);
xor U461 (N_461,In_186,In_57);
xor U462 (N_462,In_121,In_9);
xor U463 (N_463,In_108,In_156);
nand U464 (N_464,In_206,In_424);
and U465 (N_465,In_327,In_288);
nand U466 (N_466,In_324,In_18);
nand U467 (N_467,In_408,In_139);
nand U468 (N_468,In_380,In_394);
nor U469 (N_469,In_457,In_187);
nor U470 (N_470,In_46,In_174);
nor U471 (N_471,In_6,In_58);
xor U472 (N_472,In_456,In_408);
or U473 (N_473,In_391,In_389);
nor U474 (N_474,In_165,In_277);
and U475 (N_475,In_453,In_483);
or U476 (N_476,In_354,In_136);
or U477 (N_477,In_341,In_247);
nand U478 (N_478,In_430,In_120);
and U479 (N_479,In_0,In_212);
or U480 (N_480,In_268,In_291);
and U481 (N_481,In_62,In_36);
xnor U482 (N_482,In_252,In_277);
and U483 (N_483,In_94,In_434);
and U484 (N_484,In_247,In_46);
nor U485 (N_485,In_361,In_60);
or U486 (N_486,In_29,In_261);
nand U487 (N_487,In_387,In_459);
nand U488 (N_488,In_244,In_298);
or U489 (N_489,In_445,In_359);
nor U490 (N_490,In_0,In_493);
xnor U491 (N_491,In_472,In_449);
and U492 (N_492,In_60,In_132);
nand U493 (N_493,In_23,In_222);
nor U494 (N_494,In_498,In_269);
nand U495 (N_495,In_326,In_299);
and U496 (N_496,In_134,In_330);
nand U497 (N_497,In_265,In_271);
xnor U498 (N_498,In_135,In_382);
nor U499 (N_499,In_77,In_365);
nor U500 (N_500,N_152,N_201);
and U501 (N_501,N_359,N_316);
nand U502 (N_502,N_397,N_75);
nor U503 (N_503,N_449,N_144);
or U504 (N_504,N_17,N_289);
nand U505 (N_505,N_265,N_391);
nand U506 (N_506,N_320,N_68);
and U507 (N_507,N_103,N_81);
nand U508 (N_508,N_481,N_107);
xor U509 (N_509,N_198,N_196);
or U510 (N_510,N_21,N_483);
xnor U511 (N_511,N_156,N_175);
nand U512 (N_512,N_204,N_452);
nor U513 (N_513,N_244,N_199);
or U514 (N_514,N_381,N_86);
and U515 (N_515,N_277,N_146);
xnor U516 (N_516,N_362,N_132);
and U517 (N_517,N_141,N_271);
xor U518 (N_518,N_84,N_45);
or U519 (N_519,N_470,N_28);
and U520 (N_520,N_484,N_65);
xnor U521 (N_521,N_208,N_380);
xor U522 (N_522,N_233,N_499);
nor U523 (N_523,N_465,N_280);
nand U524 (N_524,N_50,N_370);
or U525 (N_525,N_210,N_411);
xnor U526 (N_526,N_177,N_49);
nand U527 (N_527,N_474,N_150);
and U528 (N_528,N_477,N_267);
and U529 (N_529,N_352,N_47);
or U530 (N_530,N_339,N_323);
xnor U531 (N_531,N_281,N_133);
xor U532 (N_532,N_379,N_264);
xor U533 (N_533,N_384,N_363);
nand U534 (N_534,N_46,N_443);
nor U535 (N_535,N_192,N_155);
xor U536 (N_536,N_371,N_3);
and U537 (N_537,N_270,N_344);
and U538 (N_538,N_451,N_285);
xor U539 (N_539,N_429,N_420);
or U540 (N_540,N_182,N_416);
or U541 (N_541,N_194,N_274);
or U542 (N_542,N_482,N_467);
nand U543 (N_543,N_473,N_64);
nand U544 (N_544,N_367,N_180);
and U545 (N_545,N_406,N_229);
xnor U546 (N_546,N_297,N_444);
xor U547 (N_547,N_471,N_168);
xor U548 (N_548,N_216,N_385);
and U549 (N_549,N_403,N_25);
or U550 (N_550,N_450,N_448);
xor U551 (N_551,N_43,N_400);
or U552 (N_552,N_129,N_459);
nand U553 (N_553,N_157,N_213);
and U554 (N_554,N_402,N_159);
nand U555 (N_555,N_190,N_44);
or U556 (N_556,N_125,N_410);
xnor U557 (N_557,N_153,N_237);
or U558 (N_558,N_200,N_166);
xnor U559 (N_559,N_181,N_307);
or U560 (N_560,N_395,N_26);
nor U561 (N_561,N_135,N_239);
nand U562 (N_562,N_305,N_67);
and U563 (N_563,N_327,N_424);
and U564 (N_564,N_487,N_418);
and U565 (N_565,N_268,N_492);
or U566 (N_566,N_51,N_350);
xnor U567 (N_567,N_24,N_456);
and U568 (N_568,N_209,N_295);
or U569 (N_569,N_214,N_337);
and U570 (N_570,N_372,N_80);
nor U571 (N_571,N_234,N_472);
nand U572 (N_572,N_187,N_476);
nor U573 (N_573,N_290,N_15);
nand U574 (N_574,N_292,N_419);
or U575 (N_575,N_161,N_435);
or U576 (N_576,N_167,N_253);
or U577 (N_577,N_478,N_334);
nand U578 (N_578,N_225,N_230);
xnor U579 (N_579,N_446,N_173);
nor U580 (N_580,N_324,N_108);
nand U581 (N_581,N_77,N_238);
nor U582 (N_582,N_296,N_61);
nor U583 (N_583,N_396,N_147);
xor U584 (N_584,N_52,N_109);
nand U585 (N_585,N_215,N_205);
xor U586 (N_586,N_257,N_99);
or U587 (N_587,N_138,N_343);
nor U588 (N_588,N_171,N_34);
and U589 (N_589,N_489,N_131);
xor U590 (N_590,N_258,N_145);
nand U591 (N_591,N_54,N_221);
and U592 (N_592,N_259,N_408);
xnor U593 (N_593,N_462,N_83);
nor U594 (N_594,N_48,N_70);
or U595 (N_595,N_154,N_136);
nor U596 (N_596,N_461,N_386);
nor U597 (N_597,N_466,N_57);
or U598 (N_598,N_63,N_341);
or U599 (N_599,N_357,N_358);
or U600 (N_600,N_162,N_498);
xnor U601 (N_601,N_6,N_468);
nand U602 (N_602,N_338,N_226);
nand U603 (N_603,N_114,N_364);
nand U604 (N_604,N_189,N_373);
nor U605 (N_605,N_7,N_5);
or U606 (N_606,N_92,N_22);
xnor U607 (N_607,N_104,N_299);
nor U608 (N_608,N_250,N_405);
nor U609 (N_609,N_486,N_184);
xnor U610 (N_610,N_310,N_261);
and U611 (N_611,N_365,N_88);
nor U612 (N_612,N_101,N_245);
nand U613 (N_613,N_283,N_366);
and U614 (N_614,N_491,N_480);
and U615 (N_615,N_356,N_211);
xor U616 (N_616,N_72,N_148);
and U617 (N_617,N_100,N_224);
nand U618 (N_618,N_98,N_304);
xnor U619 (N_619,N_306,N_407);
or U620 (N_620,N_41,N_431);
and U621 (N_621,N_421,N_422);
nor U622 (N_622,N_35,N_164);
nand U623 (N_623,N_329,N_56);
xnor U624 (N_624,N_353,N_97);
nor U625 (N_625,N_325,N_309);
xnor U626 (N_626,N_117,N_497);
xnor U627 (N_627,N_207,N_376);
nand U628 (N_628,N_94,N_252);
and U629 (N_629,N_149,N_219);
or U630 (N_630,N_140,N_4);
or U631 (N_631,N_163,N_423);
nor U632 (N_632,N_151,N_123);
and U633 (N_633,N_59,N_413);
or U634 (N_634,N_33,N_31);
and U635 (N_635,N_298,N_42);
nor U636 (N_636,N_255,N_433);
and U637 (N_637,N_58,N_269);
xor U638 (N_638,N_236,N_232);
nand U639 (N_639,N_401,N_312);
nor U640 (N_640,N_340,N_282);
and U641 (N_641,N_14,N_23);
and U642 (N_642,N_203,N_479);
or U643 (N_643,N_399,N_328);
nor U644 (N_644,N_398,N_293);
nand U645 (N_645,N_315,N_39);
nand U646 (N_646,N_89,N_263);
and U647 (N_647,N_197,N_87);
or U648 (N_648,N_186,N_249);
and U649 (N_649,N_102,N_354);
nand U650 (N_650,N_112,N_458);
and U651 (N_651,N_447,N_311);
nand U652 (N_652,N_319,N_178);
nand U653 (N_653,N_95,N_392);
or U654 (N_654,N_30,N_393);
nor U655 (N_655,N_348,N_463);
nor U656 (N_656,N_8,N_128);
xnor U657 (N_657,N_383,N_273);
and U658 (N_658,N_12,N_439);
and U659 (N_659,N_251,N_287);
xnor U660 (N_660,N_368,N_248);
nand U661 (N_661,N_10,N_347);
nor U662 (N_662,N_493,N_260);
or U663 (N_663,N_317,N_32);
or U664 (N_664,N_242,N_330);
and U665 (N_665,N_442,N_460);
nor U666 (N_666,N_279,N_457);
xnor U667 (N_667,N_124,N_389);
and U668 (N_668,N_276,N_342);
xnor U669 (N_669,N_172,N_169);
xor U670 (N_670,N_69,N_16);
and U671 (N_671,N_119,N_432);
nand U672 (N_672,N_142,N_485);
xnor U673 (N_673,N_336,N_286);
and U674 (N_674,N_294,N_53);
nand U675 (N_675,N_235,N_110);
nand U676 (N_676,N_469,N_183);
xnor U677 (N_677,N_223,N_212);
xor U678 (N_678,N_90,N_262);
nor U679 (N_679,N_243,N_160);
and U680 (N_680,N_332,N_404);
and U681 (N_681,N_300,N_415);
nor U682 (N_682,N_228,N_496);
xor U683 (N_683,N_79,N_165);
or U684 (N_684,N_360,N_227);
nor U685 (N_685,N_382,N_222);
nor U686 (N_686,N_220,N_488);
or U687 (N_687,N_247,N_137);
nand U688 (N_688,N_193,N_9);
and U689 (N_689,N_333,N_445);
nand U690 (N_690,N_428,N_272);
nor U691 (N_691,N_375,N_143);
and U692 (N_692,N_85,N_369);
nand U693 (N_693,N_37,N_240);
nor U694 (N_694,N_394,N_134);
or U695 (N_695,N_38,N_76);
or U696 (N_696,N_349,N_390);
nor U697 (N_697,N_351,N_122);
nand U698 (N_698,N_361,N_27);
nor U699 (N_699,N_116,N_437);
nor U700 (N_700,N_454,N_206);
nor U701 (N_701,N_326,N_0);
nand U702 (N_702,N_118,N_455);
nor U703 (N_703,N_331,N_409);
and U704 (N_704,N_71,N_174);
nor U705 (N_705,N_256,N_321);
nand U706 (N_706,N_170,N_464);
xor U707 (N_707,N_231,N_78);
and U708 (N_708,N_127,N_73);
and U709 (N_709,N_241,N_106);
nor U710 (N_710,N_288,N_278);
or U711 (N_711,N_91,N_275);
or U712 (N_712,N_427,N_388);
nor U713 (N_713,N_303,N_414);
or U714 (N_714,N_195,N_490);
and U715 (N_715,N_29,N_2);
nor U716 (N_716,N_335,N_434);
or U717 (N_717,N_176,N_453);
or U718 (N_718,N_1,N_387);
xnor U719 (N_719,N_246,N_62);
nor U720 (N_720,N_121,N_301);
and U721 (N_721,N_139,N_74);
nand U722 (N_722,N_113,N_19);
xnor U723 (N_723,N_93,N_291);
nor U724 (N_724,N_11,N_374);
nor U725 (N_725,N_440,N_36);
or U726 (N_726,N_266,N_111);
nand U727 (N_727,N_346,N_126);
xor U728 (N_728,N_20,N_284);
and U729 (N_729,N_308,N_218);
nor U730 (N_730,N_494,N_355);
xnor U731 (N_731,N_430,N_202);
or U732 (N_732,N_254,N_438);
or U733 (N_733,N_185,N_426);
and U734 (N_734,N_378,N_425);
nor U735 (N_735,N_115,N_436);
and U736 (N_736,N_322,N_217);
nor U737 (N_737,N_82,N_314);
or U738 (N_738,N_13,N_18);
nand U739 (N_739,N_412,N_377);
and U740 (N_740,N_495,N_179);
and U741 (N_741,N_475,N_158);
nand U742 (N_742,N_441,N_60);
nand U743 (N_743,N_318,N_96);
or U744 (N_744,N_66,N_130);
nor U745 (N_745,N_417,N_345);
xnor U746 (N_746,N_55,N_188);
nand U747 (N_747,N_313,N_302);
and U748 (N_748,N_105,N_191);
or U749 (N_749,N_120,N_40);
nor U750 (N_750,N_144,N_41);
or U751 (N_751,N_395,N_20);
and U752 (N_752,N_433,N_214);
and U753 (N_753,N_74,N_366);
nand U754 (N_754,N_456,N_37);
nand U755 (N_755,N_184,N_438);
nand U756 (N_756,N_160,N_267);
nor U757 (N_757,N_21,N_130);
and U758 (N_758,N_415,N_384);
and U759 (N_759,N_36,N_432);
nor U760 (N_760,N_102,N_79);
and U761 (N_761,N_144,N_82);
and U762 (N_762,N_6,N_291);
and U763 (N_763,N_482,N_192);
nand U764 (N_764,N_291,N_190);
and U765 (N_765,N_282,N_431);
nor U766 (N_766,N_51,N_282);
xor U767 (N_767,N_189,N_381);
and U768 (N_768,N_116,N_478);
nor U769 (N_769,N_354,N_239);
nor U770 (N_770,N_219,N_221);
nand U771 (N_771,N_235,N_266);
and U772 (N_772,N_493,N_450);
and U773 (N_773,N_289,N_426);
xor U774 (N_774,N_113,N_305);
or U775 (N_775,N_97,N_66);
xor U776 (N_776,N_262,N_226);
xnor U777 (N_777,N_413,N_103);
nor U778 (N_778,N_493,N_247);
nor U779 (N_779,N_38,N_99);
nand U780 (N_780,N_44,N_386);
xor U781 (N_781,N_124,N_5);
or U782 (N_782,N_444,N_289);
nor U783 (N_783,N_81,N_410);
nand U784 (N_784,N_391,N_269);
xor U785 (N_785,N_356,N_226);
and U786 (N_786,N_317,N_72);
nand U787 (N_787,N_399,N_54);
xnor U788 (N_788,N_460,N_167);
xnor U789 (N_789,N_278,N_279);
xnor U790 (N_790,N_97,N_455);
and U791 (N_791,N_337,N_277);
nand U792 (N_792,N_49,N_372);
and U793 (N_793,N_297,N_110);
or U794 (N_794,N_71,N_55);
nor U795 (N_795,N_124,N_190);
xnor U796 (N_796,N_441,N_115);
nor U797 (N_797,N_305,N_127);
and U798 (N_798,N_459,N_193);
nor U799 (N_799,N_284,N_208);
or U800 (N_800,N_486,N_398);
nor U801 (N_801,N_63,N_114);
and U802 (N_802,N_119,N_242);
nor U803 (N_803,N_238,N_223);
nand U804 (N_804,N_23,N_56);
xnor U805 (N_805,N_60,N_206);
nand U806 (N_806,N_64,N_155);
nor U807 (N_807,N_319,N_403);
xnor U808 (N_808,N_415,N_480);
and U809 (N_809,N_144,N_438);
nor U810 (N_810,N_78,N_127);
or U811 (N_811,N_81,N_162);
or U812 (N_812,N_257,N_436);
xnor U813 (N_813,N_310,N_420);
and U814 (N_814,N_391,N_267);
xnor U815 (N_815,N_438,N_45);
or U816 (N_816,N_93,N_79);
and U817 (N_817,N_461,N_456);
nand U818 (N_818,N_356,N_224);
nand U819 (N_819,N_70,N_379);
and U820 (N_820,N_413,N_16);
nand U821 (N_821,N_485,N_286);
and U822 (N_822,N_325,N_360);
xnor U823 (N_823,N_465,N_58);
nand U824 (N_824,N_224,N_45);
nor U825 (N_825,N_231,N_201);
or U826 (N_826,N_157,N_212);
and U827 (N_827,N_410,N_307);
nor U828 (N_828,N_470,N_230);
xnor U829 (N_829,N_161,N_396);
and U830 (N_830,N_73,N_287);
and U831 (N_831,N_248,N_267);
xor U832 (N_832,N_202,N_442);
nor U833 (N_833,N_294,N_223);
or U834 (N_834,N_392,N_469);
xor U835 (N_835,N_328,N_3);
nor U836 (N_836,N_42,N_316);
nor U837 (N_837,N_16,N_320);
nor U838 (N_838,N_96,N_146);
nand U839 (N_839,N_261,N_472);
nor U840 (N_840,N_94,N_87);
nor U841 (N_841,N_355,N_481);
or U842 (N_842,N_225,N_87);
nor U843 (N_843,N_137,N_244);
xnor U844 (N_844,N_352,N_75);
xor U845 (N_845,N_299,N_363);
xnor U846 (N_846,N_223,N_196);
or U847 (N_847,N_138,N_374);
nand U848 (N_848,N_357,N_82);
and U849 (N_849,N_80,N_428);
nand U850 (N_850,N_63,N_471);
nor U851 (N_851,N_42,N_174);
or U852 (N_852,N_26,N_316);
nand U853 (N_853,N_104,N_438);
xor U854 (N_854,N_91,N_218);
and U855 (N_855,N_490,N_166);
nor U856 (N_856,N_117,N_307);
or U857 (N_857,N_445,N_281);
and U858 (N_858,N_120,N_80);
nor U859 (N_859,N_218,N_460);
xnor U860 (N_860,N_153,N_336);
and U861 (N_861,N_130,N_267);
or U862 (N_862,N_382,N_242);
nor U863 (N_863,N_479,N_57);
or U864 (N_864,N_43,N_284);
or U865 (N_865,N_152,N_96);
nand U866 (N_866,N_314,N_320);
nand U867 (N_867,N_406,N_143);
nor U868 (N_868,N_97,N_220);
nand U869 (N_869,N_344,N_323);
or U870 (N_870,N_55,N_334);
xnor U871 (N_871,N_422,N_49);
xor U872 (N_872,N_198,N_357);
and U873 (N_873,N_126,N_269);
nand U874 (N_874,N_132,N_79);
nand U875 (N_875,N_261,N_103);
xnor U876 (N_876,N_154,N_348);
and U877 (N_877,N_293,N_446);
nand U878 (N_878,N_48,N_42);
nand U879 (N_879,N_352,N_102);
nor U880 (N_880,N_375,N_225);
xnor U881 (N_881,N_207,N_95);
nor U882 (N_882,N_164,N_10);
xor U883 (N_883,N_178,N_109);
and U884 (N_884,N_270,N_195);
xnor U885 (N_885,N_59,N_309);
nor U886 (N_886,N_79,N_69);
nor U887 (N_887,N_435,N_134);
nand U888 (N_888,N_200,N_233);
and U889 (N_889,N_465,N_189);
nor U890 (N_890,N_398,N_430);
nand U891 (N_891,N_172,N_139);
xnor U892 (N_892,N_252,N_100);
nand U893 (N_893,N_365,N_488);
nor U894 (N_894,N_4,N_244);
and U895 (N_895,N_261,N_322);
xor U896 (N_896,N_216,N_99);
or U897 (N_897,N_295,N_357);
or U898 (N_898,N_230,N_336);
xnor U899 (N_899,N_310,N_51);
xor U900 (N_900,N_284,N_300);
nor U901 (N_901,N_270,N_92);
nor U902 (N_902,N_157,N_21);
nor U903 (N_903,N_456,N_404);
xnor U904 (N_904,N_181,N_344);
and U905 (N_905,N_256,N_364);
xnor U906 (N_906,N_182,N_28);
or U907 (N_907,N_193,N_256);
nand U908 (N_908,N_190,N_184);
nand U909 (N_909,N_55,N_480);
xnor U910 (N_910,N_496,N_268);
xnor U911 (N_911,N_70,N_170);
or U912 (N_912,N_139,N_239);
nor U913 (N_913,N_123,N_304);
and U914 (N_914,N_238,N_123);
nand U915 (N_915,N_200,N_381);
and U916 (N_916,N_490,N_190);
nand U917 (N_917,N_222,N_460);
or U918 (N_918,N_277,N_103);
xnor U919 (N_919,N_138,N_386);
or U920 (N_920,N_446,N_31);
nand U921 (N_921,N_479,N_272);
nor U922 (N_922,N_270,N_33);
or U923 (N_923,N_450,N_290);
nand U924 (N_924,N_351,N_381);
nand U925 (N_925,N_314,N_254);
or U926 (N_926,N_57,N_317);
or U927 (N_927,N_203,N_122);
xnor U928 (N_928,N_96,N_458);
or U929 (N_929,N_470,N_258);
or U930 (N_930,N_337,N_278);
nor U931 (N_931,N_266,N_452);
xor U932 (N_932,N_76,N_235);
and U933 (N_933,N_398,N_279);
nor U934 (N_934,N_397,N_235);
nand U935 (N_935,N_233,N_348);
nor U936 (N_936,N_460,N_350);
xnor U937 (N_937,N_318,N_435);
nor U938 (N_938,N_126,N_107);
xnor U939 (N_939,N_432,N_490);
nor U940 (N_940,N_117,N_136);
xnor U941 (N_941,N_263,N_308);
nand U942 (N_942,N_8,N_390);
and U943 (N_943,N_118,N_272);
nor U944 (N_944,N_459,N_256);
and U945 (N_945,N_395,N_160);
nand U946 (N_946,N_350,N_452);
nor U947 (N_947,N_353,N_25);
or U948 (N_948,N_209,N_27);
nand U949 (N_949,N_267,N_216);
nand U950 (N_950,N_333,N_254);
xor U951 (N_951,N_122,N_295);
xor U952 (N_952,N_209,N_238);
nor U953 (N_953,N_49,N_221);
or U954 (N_954,N_219,N_22);
xnor U955 (N_955,N_485,N_332);
nand U956 (N_956,N_161,N_468);
or U957 (N_957,N_393,N_360);
and U958 (N_958,N_306,N_292);
and U959 (N_959,N_231,N_335);
xnor U960 (N_960,N_5,N_315);
or U961 (N_961,N_51,N_386);
nor U962 (N_962,N_213,N_194);
or U963 (N_963,N_63,N_198);
xnor U964 (N_964,N_259,N_296);
nor U965 (N_965,N_312,N_222);
and U966 (N_966,N_12,N_450);
xor U967 (N_967,N_154,N_1);
nand U968 (N_968,N_54,N_351);
and U969 (N_969,N_31,N_375);
xnor U970 (N_970,N_338,N_130);
or U971 (N_971,N_49,N_259);
nand U972 (N_972,N_97,N_370);
or U973 (N_973,N_388,N_14);
and U974 (N_974,N_252,N_89);
xnor U975 (N_975,N_241,N_74);
nor U976 (N_976,N_75,N_46);
xnor U977 (N_977,N_127,N_7);
nor U978 (N_978,N_248,N_389);
nand U979 (N_979,N_293,N_341);
nand U980 (N_980,N_92,N_422);
or U981 (N_981,N_441,N_207);
and U982 (N_982,N_21,N_435);
nor U983 (N_983,N_48,N_474);
and U984 (N_984,N_183,N_427);
nor U985 (N_985,N_354,N_6);
nor U986 (N_986,N_11,N_406);
and U987 (N_987,N_94,N_268);
or U988 (N_988,N_90,N_181);
nor U989 (N_989,N_386,N_340);
xor U990 (N_990,N_255,N_443);
nand U991 (N_991,N_268,N_384);
and U992 (N_992,N_119,N_86);
or U993 (N_993,N_190,N_368);
or U994 (N_994,N_373,N_194);
nand U995 (N_995,N_408,N_441);
xnor U996 (N_996,N_227,N_7);
or U997 (N_997,N_432,N_323);
nand U998 (N_998,N_307,N_211);
xnor U999 (N_999,N_67,N_352);
nand U1000 (N_1000,N_841,N_635);
xnor U1001 (N_1001,N_738,N_881);
or U1002 (N_1002,N_566,N_505);
xnor U1003 (N_1003,N_741,N_705);
or U1004 (N_1004,N_551,N_682);
or U1005 (N_1005,N_941,N_863);
and U1006 (N_1006,N_812,N_930);
and U1007 (N_1007,N_886,N_686);
nand U1008 (N_1008,N_593,N_585);
and U1009 (N_1009,N_791,N_595);
and U1010 (N_1010,N_772,N_872);
nor U1011 (N_1011,N_656,N_898);
and U1012 (N_1012,N_858,N_644);
xnor U1013 (N_1013,N_890,N_565);
nor U1014 (N_1014,N_664,N_807);
nor U1015 (N_1015,N_878,N_591);
nand U1016 (N_1016,N_727,N_750);
nor U1017 (N_1017,N_717,N_776);
nor U1018 (N_1018,N_833,N_651);
and U1019 (N_1019,N_934,N_891);
or U1020 (N_1020,N_852,N_979);
or U1021 (N_1021,N_980,N_603);
xor U1022 (N_1022,N_574,N_536);
xnor U1023 (N_1023,N_785,N_676);
and U1024 (N_1024,N_967,N_987);
nor U1025 (N_1025,N_530,N_758);
nor U1026 (N_1026,N_757,N_828);
or U1027 (N_1027,N_628,N_547);
xor U1028 (N_1028,N_670,N_517);
xor U1029 (N_1029,N_838,N_846);
nand U1030 (N_1030,N_808,N_775);
nor U1031 (N_1031,N_689,N_883);
and U1032 (N_1032,N_630,N_924);
xor U1033 (N_1033,N_617,N_866);
nor U1034 (N_1034,N_760,N_926);
xnor U1035 (N_1035,N_780,N_744);
nor U1036 (N_1036,N_929,N_935);
nor U1037 (N_1037,N_901,N_570);
nor U1038 (N_1038,N_857,N_687);
or U1039 (N_1039,N_995,N_711);
nand U1040 (N_1040,N_948,N_539);
and U1041 (N_1041,N_618,N_779);
nor U1042 (N_1042,N_634,N_994);
nor U1043 (N_1043,N_888,N_722);
or U1044 (N_1044,N_625,N_751);
nand U1045 (N_1045,N_562,N_700);
and U1046 (N_1046,N_900,N_733);
nor U1047 (N_1047,N_940,N_734);
and U1048 (N_1048,N_704,N_746);
or U1049 (N_1049,N_867,N_993);
and U1050 (N_1050,N_699,N_516);
nand U1051 (N_1051,N_899,N_633);
xor U1052 (N_1052,N_729,N_554);
or U1053 (N_1053,N_507,N_894);
nand U1054 (N_1054,N_798,N_567);
and U1055 (N_1055,N_902,N_963);
or U1056 (N_1056,N_865,N_600);
or U1057 (N_1057,N_928,N_690);
and U1058 (N_1058,N_815,N_725);
and U1059 (N_1059,N_859,N_860);
nand U1060 (N_1060,N_893,N_832);
nand U1061 (N_1061,N_715,N_939);
and U1062 (N_1062,N_895,N_827);
nand U1063 (N_1063,N_589,N_549);
and U1064 (N_1064,N_970,N_641);
and U1065 (N_1065,N_788,N_560);
nand U1066 (N_1066,N_792,N_569);
xor U1067 (N_1067,N_923,N_611);
and U1068 (N_1068,N_956,N_916);
and U1069 (N_1069,N_578,N_802);
nand U1070 (N_1070,N_583,N_801);
and U1071 (N_1071,N_519,N_564);
or U1072 (N_1072,N_876,N_936);
or U1073 (N_1073,N_666,N_974);
nor U1074 (N_1074,N_647,N_680);
or U1075 (N_1075,N_679,N_524);
nand U1076 (N_1076,N_982,N_669);
nor U1077 (N_1077,N_931,N_909);
nor U1078 (N_1078,N_981,N_712);
xor U1079 (N_1079,N_730,N_971);
nand U1080 (N_1080,N_826,N_906);
xnor U1081 (N_1081,N_740,N_553);
nor U1082 (N_1082,N_825,N_868);
nand U1083 (N_1083,N_642,N_783);
xor U1084 (N_1084,N_984,N_607);
or U1085 (N_1085,N_576,N_702);
nand U1086 (N_1086,N_912,N_584);
xor U1087 (N_1087,N_768,N_694);
nand U1088 (N_1088,N_806,N_723);
xnor U1089 (N_1089,N_770,N_763);
nor U1090 (N_1090,N_586,N_731);
nor U1091 (N_1091,N_639,N_718);
nor U1092 (N_1092,N_648,N_778);
and U1093 (N_1093,N_847,N_631);
nand U1094 (N_1094,N_752,N_532);
nor U1095 (N_1095,N_977,N_691);
or U1096 (N_1096,N_668,N_880);
or U1097 (N_1097,N_552,N_657);
nand U1098 (N_1098,N_575,N_513);
xnor U1099 (N_1099,N_864,N_765);
and U1100 (N_1100,N_945,N_875);
and U1101 (N_1101,N_514,N_663);
and U1102 (N_1102,N_716,N_834);
nor U1103 (N_1103,N_571,N_706);
or U1104 (N_1104,N_774,N_612);
or U1105 (N_1105,N_511,N_811);
xnor U1106 (N_1106,N_673,N_597);
xnor U1107 (N_1107,N_590,N_955);
or U1108 (N_1108,N_685,N_962);
nand U1109 (N_1109,N_879,N_887);
xor U1110 (N_1110,N_708,N_777);
and U1111 (N_1111,N_787,N_973);
nor U1112 (N_1112,N_696,N_526);
nand U1113 (N_1113,N_545,N_721);
nor U1114 (N_1114,N_767,N_515);
xor U1115 (N_1115,N_509,N_755);
and U1116 (N_1116,N_698,N_855);
and U1117 (N_1117,N_605,N_810);
nor U1118 (N_1118,N_816,N_558);
and U1119 (N_1119,N_596,N_947);
nor U1120 (N_1120,N_546,N_794);
or U1121 (N_1121,N_804,N_919);
nand U1122 (N_1122,N_813,N_869);
nand U1123 (N_1123,N_527,N_822);
xnor U1124 (N_1124,N_998,N_897);
xor U1125 (N_1125,N_573,N_732);
nand U1126 (N_1126,N_528,N_692);
or U1127 (N_1127,N_502,N_925);
xnor U1128 (N_1128,N_658,N_922);
nor U1129 (N_1129,N_580,N_819);
or U1130 (N_1130,N_501,N_749);
xor U1131 (N_1131,N_942,N_960);
or U1132 (N_1132,N_983,N_623);
and U1133 (N_1133,N_622,N_835);
and U1134 (N_1134,N_874,N_914);
nand U1135 (N_1135,N_823,N_609);
or U1136 (N_1136,N_862,N_885);
xor U1137 (N_1137,N_938,N_559);
xnor U1138 (N_1138,N_557,N_769);
or U1139 (N_1139,N_614,N_743);
xor U1140 (N_1140,N_572,N_969);
and U1141 (N_1141,N_845,N_720);
or U1142 (N_1142,N_683,N_681);
nor U1143 (N_1143,N_753,N_976);
and U1144 (N_1144,N_952,N_991);
and U1145 (N_1145,N_512,N_677);
and U1146 (N_1146,N_629,N_660);
nor U1147 (N_1147,N_742,N_793);
or U1148 (N_1148,N_745,N_620);
and U1149 (N_1149,N_621,N_703);
xnor U1150 (N_1150,N_824,N_882);
nand U1151 (N_1151,N_908,N_563);
and U1152 (N_1152,N_643,N_964);
xor U1153 (N_1153,N_637,N_649);
nor U1154 (N_1154,N_771,N_951);
xnor U1155 (N_1155,N_905,N_548);
nand U1156 (N_1156,N_661,N_544);
xnor U1157 (N_1157,N_726,N_920);
xor U1158 (N_1158,N_958,N_937);
nand U1159 (N_1159,N_638,N_829);
or U1160 (N_1160,N_653,N_608);
xnor U1161 (N_1161,N_766,N_896);
or U1162 (N_1162,N_599,N_587);
and U1163 (N_1163,N_839,N_795);
xor U1164 (N_1164,N_541,N_781);
nor U1165 (N_1165,N_606,N_821);
nand U1166 (N_1166,N_943,N_662);
nand U1167 (N_1167,N_619,N_695);
nor U1168 (N_1168,N_739,N_582);
and U1169 (N_1169,N_830,N_650);
and U1170 (N_1170,N_535,N_884);
or U1171 (N_1171,N_627,N_904);
nor U1172 (N_1172,N_959,N_616);
xor U1173 (N_1173,N_927,N_594);
nand U1174 (N_1174,N_799,N_784);
nand U1175 (N_1175,N_665,N_533);
xor U1176 (N_1176,N_871,N_697);
and U1177 (N_1177,N_975,N_921);
and U1178 (N_1178,N_508,N_719);
or U1179 (N_1179,N_978,N_932);
or U1180 (N_1180,N_579,N_645);
xnor U1181 (N_1181,N_988,N_675);
nor U1182 (N_1182,N_844,N_534);
or U1183 (N_1183,N_803,N_856);
nor U1184 (N_1184,N_748,N_790);
or U1185 (N_1185,N_735,N_877);
xor U1186 (N_1186,N_550,N_761);
nand U1187 (N_1187,N_626,N_672);
nand U1188 (N_1188,N_688,N_701);
xor U1189 (N_1189,N_809,N_671);
and U1190 (N_1190,N_840,N_949);
nor U1191 (N_1191,N_820,N_849);
nor U1192 (N_1192,N_624,N_518);
nand U1193 (N_1193,N_503,N_933);
and U1194 (N_1194,N_854,N_654);
nor U1195 (N_1195,N_773,N_831);
nor U1196 (N_1196,N_917,N_556);
nand U1197 (N_1197,N_610,N_525);
nor U1198 (N_1198,N_889,N_613);
and U1199 (N_1199,N_997,N_543);
or U1200 (N_1200,N_965,N_713);
xnor U1201 (N_1201,N_667,N_789);
nand U1202 (N_1202,N_674,N_693);
and U1203 (N_1203,N_850,N_818);
nor U1204 (N_1204,N_842,N_837);
nand U1205 (N_1205,N_907,N_851);
or U1206 (N_1206,N_954,N_989);
nand U1207 (N_1207,N_747,N_996);
nand U1208 (N_1208,N_555,N_523);
nor U1209 (N_1209,N_966,N_782);
and U1210 (N_1210,N_796,N_800);
nand U1211 (N_1211,N_754,N_646);
nand U1212 (N_1212,N_615,N_870);
xor U1213 (N_1213,N_853,N_836);
nor U1214 (N_1214,N_805,N_944);
xnor U1215 (N_1215,N_506,N_588);
nor U1216 (N_1216,N_848,N_957);
nand U1217 (N_1217,N_521,N_985);
and U1218 (N_1218,N_762,N_710);
or U1219 (N_1219,N_986,N_972);
nand U1220 (N_1220,N_659,N_540);
xor U1221 (N_1221,N_709,N_764);
and U1222 (N_1222,N_542,N_520);
nand U1223 (N_1223,N_592,N_737);
and U1224 (N_1224,N_861,N_707);
nand U1225 (N_1225,N_918,N_814);
nand U1226 (N_1226,N_684,N_601);
or U1227 (N_1227,N_602,N_568);
and U1228 (N_1228,N_843,N_728);
nor U1229 (N_1229,N_678,N_946);
or U1230 (N_1230,N_636,N_913);
xnor U1231 (N_1231,N_640,N_786);
and U1232 (N_1232,N_652,N_537);
nand U1233 (N_1233,N_992,N_950);
xnor U1234 (N_1234,N_873,N_577);
and U1235 (N_1235,N_892,N_724);
nand U1236 (N_1236,N_510,N_911);
nor U1237 (N_1237,N_915,N_817);
nor U1238 (N_1238,N_632,N_968);
and U1239 (N_1239,N_714,N_500);
xnor U1240 (N_1240,N_961,N_522);
and U1241 (N_1241,N_598,N_736);
and U1242 (N_1242,N_999,N_759);
or U1243 (N_1243,N_504,N_990);
xnor U1244 (N_1244,N_604,N_903);
or U1245 (N_1245,N_910,N_756);
nand U1246 (N_1246,N_953,N_538);
nor U1247 (N_1247,N_561,N_581);
or U1248 (N_1248,N_655,N_531);
and U1249 (N_1249,N_529,N_797);
nor U1250 (N_1250,N_640,N_608);
xnor U1251 (N_1251,N_541,N_546);
nor U1252 (N_1252,N_593,N_589);
nor U1253 (N_1253,N_512,N_570);
nand U1254 (N_1254,N_503,N_851);
xor U1255 (N_1255,N_862,N_533);
nor U1256 (N_1256,N_674,N_832);
xor U1257 (N_1257,N_972,N_932);
or U1258 (N_1258,N_925,N_579);
or U1259 (N_1259,N_874,N_781);
xnor U1260 (N_1260,N_842,N_963);
or U1261 (N_1261,N_507,N_836);
xor U1262 (N_1262,N_919,N_525);
nor U1263 (N_1263,N_644,N_565);
xnor U1264 (N_1264,N_932,N_924);
xnor U1265 (N_1265,N_608,N_505);
or U1266 (N_1266,N_701,N_696);
nor U1267 (N_1267,N_784,N_837);
nor U1268 (N_1268,N_503,N_854);
or U1269 (N_1269,N_996,N_797);
and U1270 (N_1270,N_997,N_516);
xor U1271 (N_1271,N_965,N_863);
and U1272 (N_1272,N_786,N_798);
and U1273 (N_1273,N_839,N_976);
and U1274 (N_1274,N_723,N_988);
xor U1275 (N_1275,N_551,N_933);
or U1276 (N_1276,N_677,N_870);
nor U1277 (N_1277,N_578,N_793);
or U1278 (N_1278,N_989,N_578);
and U1279 (N_1279,N_751,N_543);
or U1280 (N_1280,N_973,N_999);
or U1281 (N_1281,N_884,N_865);
and U1282 (N_1282,N_703,N_692);
nor U1283 (N_1283,N_707,N_946);
xor U1284 (N_1284,N_684,N_859);
nand U1285 (N_1285,N_859,N_780);
nand U1286 (N_1286,N_907,N_523);
nor U1287 (N_1287,N_571,N_760);
xor U1288 (N_1288,N_990,N_537);
or U1289 (N_1289,N_963,N_557);
nor U1290 (N_1290,N_676,N_553);
xor U1291 (N_1291,N_652,N_947);
or U1292 (N_1292,N_976,N_961);
or U1293 (N_1293,N_878,N_825);
nor U1294 (N_1294,N_639,N_799);
or U1295 (N_1295,N_922,N_960);
nor U1296 (N_1296,N_875,N_974);
nand U1297 (N_1297,N_919,N_844);
xnor U1298 (N_1298,N_667,N_718);
nor U1299 (N_1299,N_984,N_762);
xnor U1300 (N_1300,N_978,N_517);
and U1301 (N_1301,N_565,N_744);
or U1302 (N_1302,N_950,N_741);
or U1303 (N_1303,N_631,N_979);
or U1304 (N_1304,N_553,N_801);
xnor U1305 (N_1305,N_677,N_782);
nand U1306 (N_1306,N_834,N_662);
and U1307 (N_1307,N_973,N_545);
nand U1308 (N_1308,N_939,N_598);
or U1309 (N_1309,N_799,N_821);
xor U1310 (N_1310,N_690,N_848);
or U1311 (N_1311,N_672,N_562);
nand U1312 (N_1312,N_916,N_648);
nand U1313 (N_1313,N_546,N_564);
and U1314 (N_1314,N_507,N_573);
and U1315 (N_1315,N_517,N_642);
nand U1316 (N_1316,N_730,N_699);
nor U1317 (N_1317,N_939,N_663);
nor U1318 (N_1318,N_747,N_697);
nand U1319 (N_1319,N_571,N_798);
and U1320 (N_1320,N_979,N_977);
xnor U1321 (N_1321,N_674,N_639);
nand U1322 (N_1322,N_989,N_786);
xnor U1323 (N_1323,N_714,N_846);
nand U1324 (N_1324,N_537,N_974);
nor U1325 (N_1325,N_512,N_975);
nor U1326 (N_1326,N_610,N_568);
nand U1327 (N_1327,N_871,N_707);
or U1328 (N_1328,N_662,N_857);
nor U1329 (N_1329,N_772,N_700);
and U1330 (N_1330,N_706,N_715);
or U1331 (N_1331,N_781,N_701);
xor U1332 (N_1332,N_867,N_824);
or U1333 (N_1333,N_770,N_938);
xor U1334 (N_1334,N_589,N_939);
nand U1335 (N_1335,N_948,N_787);
nand U1336 (N_1336,N_970,N_532);
or U1337 (N_1337,N_601,N_602);
nand U1338 (N_1338,N_971,N_974);
or U1339 (N_1339,N_687,N_738);
or U1340 (N_1340,N_994,N_534);
nor U1341 (N_1341,N_545,N_901);
nand U1342 (N_1342,N_761,N_854);
nor U1343 (N_1343,N_963,N_749);
and U1344 (N_1344,N_940,N_817);
xnor U1345 (N_1345,N_646,N_772);
and U1346 (N_1346,N_910,N_621);
nor U1347 (N_1347,N_606,N_704);
and U1348 (N_1348,N_839,N_895);
nand U1349 (N_1349,N_581,N_893);
and U1350 (N_1350,N_801,N_989);
xnor U1351 (N_1351,N_736,N_504);
nand U1352 (N_1352,N_952,N_559);
or U1353 (N_1353,N_761,N_775);
nor U1354 (N_1354,N_835,N_601);
nand U1355 (N_1355,N_708,N_634);
xor U1356 (N_1356,N_965,N_522);
nand U1357 (N_1357,N_797,N_876);
or U1358 (N_1358,N_774,N_989);
nand U1359 (N_1359,N_676,N_889);
nor U1360 (N_1360,N_778,N_553);
xnor U1361 (N_1361,N_938,N_767);
nor U1362 (N_1362,N_879,N_747);
xnor U1363 (N_1363,N_674,N_547);
or U1364 (N_1364,N_828,N_690);
nor U1365 (N_1365,N_578,N_837);
nor U1366 (N_1366,N_771,N_945);
or U1367 (N_1367,N_775,N_736);
nand U1368 (N_1368,N_722,N_542);
nand U1369 (N_1369,N_885,N_695);
or U1370 (N_1370,N_869,N_921);
and U1371 (N_1371,N_595,N_883);
or U1372 (N_1372,N_731,N_668);
nor U1373 (N_1373,N_703,N_672);
xnor U1374 (N_1374,N_775,N_636);
xnor U1375 (N_1375,N_627,N_737);
and U1376 (N_1376,N_974,N_741);
xnor U1377 (N_1377,N_659,N_691);
nand U1378 (N_1378,N_634,N_761);
or U1379 (N_1379,N_879,N_986);
and U1380 (N_1380,N_739,N_831);
and U1381 (N_1381,N_650,N_620);
nand U1382 (N_1382,N_588,N_531);
nand U1383 (N_1383,N_917,N_863);
nand U1384 (N_1384,N_558,N_943);
nor U1385 (N_1385,N_735,N_940);
nor U1386 (N_1386,N_992,N_758);
nor U1387 (N_1387,N_852,N_631);
xnor U1388 (N_1388,N_972,N_966);
or U1389 (N_1389,N_866,N_703);
nand U1390 (N_1390,N_849,N_823);
xnor U1391 (N_1391,N_764,N_786);
nor U1392 (N_1392,N_926,N_556);
or U1393 (N_1393,N_984,N_514);
nand U1394 (N_1394,N_626,N_788);
xor U1395 (N_1395,N_537,N_825);
nor U1396 (N_1396,N_966,N_659);
xnor U1397 (N_1397,N_683,N_751);
or U1398 (N_1398,N_852,N_709);
xor U1399 (N_1399,N_749,N_962);
or U1400 (N_1400,N_582,N_899);
xor U1401 (N_1401,N_596,N_657);
nor U1402 (N_1402,N_808,N_758);
nand U1403 (N_1403,N_557,N_538);
xnor U1404 (N_1404,N_546,N_792);
or U1405 (N_1405,N_678,N_880);
xor U1406 (N_1406,N_545,N_551);
xnor U1407 (N_1407,N_694,N_700);
or U1408 (N_1408,N_814,N_564);
nand U1409 (N_1409,N_938,N_645);
nand U1410 (N_1410,N_654,N_807);
and U1411 (N_1411,N_827,N_661);
nor U1412 (N_1412,N_579,N_845);
nand U1413 (N_1413,N_982,N_873);
and U1414 (N_1414,N_764,N_939);
nand U1415 (N_1415,N_861,N_562);
nor U1416 (N_1416,N_559,N_504);
or U1417 (N_1417,N_525,N_854);
or U1418 (N_1418,N_884,N_782);
or U1419 (N_1419,N_580,N_559);
nor U1420 (N_1420,N_696,N_871);
xnor U1421 (N_1421,N_570,N_842);
or U1422 (N_1422,N_785,N_646);
nor U1423 (N_1423,N_740,N_508);
xnor U1424 (N_1424,N_629,N_903);
or U1425 (N_1425,N_715,N_574);
or U1426 (N_1426,N_550,N_630);
or U1427 (N_1427,N_845,N_574);
nand U1428 (N_1428,N_760,N_718);
xor U1429 (N_1429,N_719,N_743);
or U1430 (N_1430,N_892,N_756);
nand U1431 (N_1431,N_663,N_623);
xnor U1432 (N_1432,N_816,N_915);
xor U1433 (N_1433,N_635,N_756);
or U1434 (N_1434,N_703,N_997);
and U1435 (N_1435,N_703,N_968);
nor U1436 (N_1436,N_949,N_715);
and U1437 (N_1437,N_932,N_685);
xor U1438 (N_1438,N_871,N_516);
and U1439 (N_1439,N_938,N_795);
nor U1440 (N_1440,N_591,N_626);
xnor U1441 (N_1441,N_993,N_579);
nand U1442 (N_1442,N_836,N_758);
nand U1443 (N_1443,N_763,N_717);
nand U1444 (N_1444,N_765,N_729);
nor U1445 (N_1445,N_666,N_864);
and U1446 (N_1446,N_612,N_935);
nor U1447 (N_1447,N_739,N_574);
nor U1448 (N_1448,N_910,N_752);
nand U1449 (N_1449,N_622,N_963);
or U1450 (N_1450,N_560,N_629);
nor U1451 (N_1451,N_806,N_767);
nand U1452 (N_1452,N_785,N_760);
and U1453 (N_1453,N_975,N_721);
nor U1454 (N_1454,N_758,N_618);
nand U1455 (N_1455,N_856,N_762);
nand U1456 (N_1456,N_877,N_557);
or U1457 (N_1457,N_953,N_821);
nor U1458 (N_1458,N_721,N_831);
xor U1459 (N_1459,N_907,N_563);
xnor U1460 (N_1460,N_940,N_538);
nand U1461 (N_1461,N_984,N_756);
or U1462 (N_1462,N_619,N_584);
nor U1463 (N_1463,N_838,N_946);
nor U1464 (N_1464,N_868,N_838);
nand U1465 (N_1465,N_913,N_971);
or U1466 (N_1466,N_897,N_740);
or U1467 (N_1467,N_777,N_619);
nor U1468 (N_1468,N_757,N_758);
nor U1469 (N_1469,N_837,N_952);
or U1470 (N_1470,N_625,N_580);
and U1471 (N_1471,N_526,N_728);
xnor U1472 (N_1472,N_917,N_561);
nor U1473 (N_1473,N_606,N_770);
xor U1474 (N_1474,N_982,N_790);
or U1475 (N_1475,N_859,N_739);
or U1476 (N_1476,N_914,N_533);
nor U1477 (N_1477,N_958,N_848);
nor U1478 (N_1478,N_989,N_835);
or U1479 (N_1479,N_506,N_653);
nand U1480 (N_1480,N_583,N_838);
xnor U1481 (N_1481,N_836,N_963);
xor U1482 (N_1482,N_555,N_645);
or U1483 (N_1483,N_670,N_946);
xnor U1484 (N_1484,N_717,N_670);
nor U1485 (N_1485,N_766,N_947);
and U1486 (N_1486,N_553,N_996);
nand U1487 (N_1487,N_547,N_848);
and U1488 (N_1488,N_784,N_891);
and U1489 (N_1489,N_550,N_773);
and U1490 (N_1490,N_772,N_512);
and U1491 (N_1491,N_884,N_941);
and U1492 (N_1492,N_990,N_632);
nand U1493 (N_1493,N_553,N_578);
nand U1494 (N_1494,N_955,N_697);
xor U1495 (N_1495,N_869,N_929);
xor U1496 (N_1496,N_814,N_902);
xor U1497 (N_1497,N_967,N_574);
or U1498 (N_1498,N_969,N_877);
or U1499 (N_1499,N_846,N_939);
or U1500 (N_1500,N_1276,N_1497);
and U1501 (N_1501,N_1306,N_1304);
xor U1502 (N_1502,N_1287,N_1153);
or U1503 (N_1503,N_1208,N_1060);
or U1504 (N_1504,N_1041,N_1318);
nand U1505 (N_1505,N_1009,N_1038);
nand U1506 (N_1506,N_1417,N_1131);
or U1507 (N_1507,N_1434,N_1213);
and U1508 (N_1508,N_1335,N_1339);
and U1509 (N_1509,N_1371,N_1337);
xnor U1510 (N_1510,N_1274,N_1112);
nand U1511 (N_1511,N_1286,N_1082);
or U1512 (N_1512,N_1118,N_1151);
nand U1513 (N_1513,N_1178,N_1152);
and U1514 (N_1514,N_1261,N_1415);
nor U1515 (N_1515,N_1249,N_1048);
or U1516 (N_1516,N_1404,N_1350);
nor U1517 (N_1517,N_1332,N_1169);
or U1518 (N_1518,N_1227,N_1210);
and U1519 (N_1519,N_1228,N_1262);
nor U1520 (N_1520,N_1466,N_1224);
and U1521 (N_1521,N_1174,N_1381);
nand U1522 (N_1522,N_1327,N_1014);
nand U1523 (N_1523,N_1285,N_1264);
xor U1524 (N_1524,N_1126,N_1421);
nor U1525 (N_1525,N_1006,N_1030);
xor U1526 (N_1526,N_1297,N_1344);
xor U1527 (N_1527,N_1023,N_1348);
nand U1528 (N_1528,N_1076,N_1099);
or U1529 (N_1529,N_1267,N_1439);
nor U1530 (N_1530,N_1104,N_1320);
nand U1531 (N_1531,N_1314,N_1062);
nand U1532 (N_1532,N_1345,N_1427);
nor U1533 (N_1533,N_1061,N_1295);
and U1534 (N_1534,N_1369,N_1103);
xor U1535 (N_1535,N_1486,N_1219);
xnor U1536 (N_1536,N_1065,N_1007);
nand U1537 (N_1537,N_1107,N_1479);
nor U1538 (N_1538,N_1447,N_1383);
xor U1539 (N_1539,N_1201,N_1209);
nor U1540 (N_1540,N_1498,N_1311);
nor U1541 (N_1541,N_1307,N_1167);
xor U1542 (N_1542,N_1142,N_1423);
nand U1543 (N_1543,N_1111,N_1260);
xnor U1544 (N_1544,N_1438,N_1275);
xnor U1545 (N_1545,N_1263,N_1199);
nor U1546 (N_1546,N_1172,N_1257);
nand U1547 (N_1547,N_1347,N_1252);
or U1548 (N_1548,N_1412,N_1380);
nand U1549 (N_1549,N_1265,N_1308);
xnor U1550 (N_1550,N_1487,N_1455);
and U1551 (N_1551,N_1122,N_1458);
nand U1552 (N_1552,N_1204,N_1217);
or U1553 (N_1553,N_1385,N_1341);
and U1554 (N_1554,N_1467,N_1315);
xor U1555 (N_1555,N_1042,N_1231);
nor U1556 (N_1556,N_1351,N_1493);
nand U1557 (N_1557,N_1402,N_1273);
and U1558 (N_1558,N_1135,N_1093);
nor U1559 (N_1559,N_1134,N_1205);
nand U1560 (N_1560,N_1336,N_1294);
xnor U1561 (N_1561,N_1250,N_1226);
nor U1562 (N_1562,N_1125,N_1079);
nor U1563 (N_1563,N_1182,N_1472);
nand U1564 (N_1564,N_1074,N_1046);
xor U1565 (N_1565,N_1435,N_1324);
nand U1566 (N_1566,N_1051,N_1272);
xor U1567 (N_1567,N_1194,N_1155);
xnor U1568 (N_1568,N_1407,N_1058);
or U1569 (N_1569,N_1496,N_1021);
xnor U1570 (N_1570,N_1084,N_1181);
and U1571 (N_1571,N_1379,N_1358);
and U1572 (N_1572,N_1083,N_1049);
nor U1573 (N_1573,N_1214,N_1095);
nor U1574 (N_1574,N_1384,N_1138);
xnor U1575 (N_1575,N_1397,N_1368);
or U1576 (N_1576,N_1270,N_1491);
or U1577 (N_1577,N_1080,N_1396);
or U1578 (N_1578,N_1037,N_1357);
and U1579 (N_1579,N_1203,N_1206);
xnor U1580 (N_1580,N_1137,N_1161);
nand U1581 (N_1581,N_1393,N_1490);
nor U1582 (N_1582,N_1476,N_1441);
nand U1583 (N_1583,N_1445,N_1164);
and U1584 (N_1584,N_1313,N_1352);
or U1585 (N_1585,N_1431,N_1400);
and U1586 (N_1586,N_1334,N_1179);
or U1587 (N_1587,N_1081,N_1303);
nand U1588 (N_1588,N_1443,N_1026);
or U1589 (N_1589,N_1477,N_1321);
nor U1590 (N_1590,N_1386,N_1216);
xor U1591 (N_1591,N_1063,N_1086);
nor U1592 (N_1592,N_1359,N_1378);
xnor U1593 (N_1593,N_1360,N_1162);
xor U1594 (N_1594,N_1188,N_1448);
nor U1595 (N_1595,N_1140,N_1193);
and U1596 (N_1596,N_1150,N_1364);
and U1597 (N_1597,N_1132,N_1073);
and U1598 (N_1598,N_1373,N_1293);
xnor U1599 (N_1599,N_1408,N_1464);
nand U1600 (N_1600,N_1144,N_1059);
xor U1601 (N_1601,N_1392,N_1401);
nor U1602 (N_1602,N_1003,N_1409);
and U1603 (N_1603,N_1141,N_1077);
and U1604 (N_1604,N_1291,N_1354);
and U1605 (N_1605,N_1361,N_1362);
and U1606 (N_1606,N_1159,N_1094);
or U1607 (N_1607,N_1485,N_1449);
or U1608 (N_1608,N_1461,N_1154);
xnor U1609 (N_1609,N_1075,N_1020);
xor U1610 (N_1610,N_1316,N_1090);
nand U1611 (N_1611,N_1478,N_1489);
nor U1612 (N_1612,N_1376,N_1419);
xor U1613 (N_1613,N_1370,N_1196);
nand U1614 (N_1614,N_1015,N_1105);
and U1615 (N_1615,N_1230,N_1266);
nor U1616 (N_1616,N_1184,N_1148);
xnor U1617 (N_1617,N_1403,N_1156);
nor U1618 (N_1618,N_1028,N_1004);
xor U1619 (N_1619,N_1200,N_1413);
and U1620 (N_1620,N_1067,N_1317);
nor U1621 (N_1621,N_1319,N_1469);
and U1622 (N_1622,N_1165,N_1171);
or U1623 (N_1623,N_1106,N_1254);
and U1624 (N_1624,N_1124,N_1198);
xor U1625 (N_1625,N_1070,N_1390);
nand U1626 (N_1626,N_1387,N_1101);
and U1627 (N_1627,N_1012,N_1475);
xnor U1628 (N_1628,N_1177,N_1452);
xor U1629 (N_1629,N_1289,N_1168);
nand U1630 (N_1630,N_1047,N_1459);
or U1631 (N_1631,N_1221,N_1157);
xor U1632 (N_1632,N_1225,N_1146);
or U1633 (N_1633,N_1256,N_1139);
nand U1634 (N_1634,N_1398,N_1096);
and U1635 (N_1635,N_1282,N_1278);
and U1636 (N_1636,N_1245,N_1000);
or U1637 (N_1637,N_1300,N_1430);
and U1638 (N_1638,N_1338,N_1192);
nand U1639 (N_1639,N_1055,N_1202);
nor U1640 (N_1640,N_1440,N_1022);
or U1641 (N_1641,N_1032,N_1495);
and U1642 (N_1642,N_1251,N_1108);
or U1643 (N_1643,N_1087,N_1343);
or U1644 (N_1644,N_1024,N_1328);
or U1645 (N_1645,N_1323,N_1040);
and U1646 (N_1646,N_1480,N_1484);
nor U1647 (N_1647,N_1411,N_1259);
xor U1648 (N_1648,N_1388,N_1422);
xnor U1649 (N_1649,N_1160,N_1457);
or U1650 (N_1650,N_1456,N_1190);
nor U1651 (N_1651,N_1414,N_1248);
and U1652 (N_1652,N_1091,N_1223);
nor U1653 (N_1653,N_1143,N_1322);
xnor U1654 (N_1654,N_1483,N_1002);
or U1655 (N_1655,N_1068,N_1005);
xnor U1656 (N_1656,N_1450,N_1340);
and U1657 (N_1657,N_1391,N_1429);
xor U1658 (N_1658,N_1468,N_1033);
and U1659 (N_1659,N_1416,N_1482);
or U1660 (N_1660,N_1292,N_1097);
nor U1661 (N_1661,N_1284,N_1454);
nand U1662 (N_1662,N_1191,N_1240);
nor U1663 (N_1663,N_1418,N_1269);
or U1664 (N_1664,N_1098,N_1246);
nand U1665 (N_1665,N_1029,N_1136);
nor U1666 (N_1666,N_1089,N_1277);
nand U1667 (N_1667,N_1211,N_1355);
xor U1668 (N_1668,N_1129,N_1039);
nor U1669 (N_1669,N_1045,N_1365);
and U1670 (N_1670,N_1050,N_1149);
nor U1671 (N_1671,N_1460,N_1442);
or U1672 (N_1672,N_1071,N_1183);
nor U1673 (N_1673,N_1053,N_1302);
xor U1674 (N_1674,N_1372,N_1013);
and U1675 (N_1675,N_1333,N_1235);
and U1676 (N_1676,N_1399,N_1356);
or U1677 (N_1677,N_1481,N_1187);
or U1678 (N_1678,N_1078,N_1301);
and U1679 (N_1679,N_1255,N_1446);
xor U1680 (N_1680,N_1465,N_1025);
or U1681 (N_1681,N_1166,N_1044);
nand U1682 (N_1682,N_1389,N_1019);
and U1683 (N_1683,N_1236,N_1375);
nand U1684 (N_1684,N_1218,N_1405);
nor U1685 (N_1685,N_1253,N_1027);
xor U1686 (N_1686,N_1410,N_1451);
or U1687 (N_1687,N_1170,N_1102);
nand U1688 (N_1688,N_1054,N_1064);
and U1689 (N_1689,N_1433,N_1242);
xnor U1690 (N_1690,N_1463,N_1471);
xor U1691 (N_1691,N_1377,N_1367);
nor U1692 (N_1692,N_1117,N_1426);
or U1693 (N_1693,N_1305,N_1492);
or U1694 (N_1694,N_1395,N_1428);
nor U1695 (N_1695,N_1353,N_1494);
nand U1696 (N_1696,N_1215,N_1330);
and U1697 (N_1697,N_1069,N_1420);
nand U1698 (N_1698,N_1127,N_1279);
and U1699 (N_1699,N_1057,N_1100);
and U1700 (N_1700,N_1299,N_1232);
nand U1701 (N_1701,N_1271,N_1298);
and U1702 (N_1702,N_1290,N_1382);
xor U1703 (N_1703,N_1229,N_1220);
nor U1704 (N_1704,N_1189,N_1346);
nand U1705 (N_1705,N_1116,N_1173);
nor U1706 (N_1706,N_1043,N_1052);
and U1707 (N_1707,N_1238,N_1056);
or U1708 (N_1708,N_1268,N_1366);
xor U1709 (N_1709,N_1121,N_1437);
nand U1710 (N_1710,N_1241,N_1234);
xnor U1711 (N_1711,N_1444,N_1186);
nand U1712 (N_1712,N_1309,N_1394);
and U1713 (N_1713,N_1010,N_1243);
nand U1714 (N_1714,N_1473,N_1329);
or U1715 (N_1715,N_1034,N_1488);
nand U1716 (N_1716,N_1175,N_1436);
nand U1717 (N_1717,N_1147,N_1072);
nand U1718 (N_1718,N_1197,N_1180);
xor U1719 (N_1719,N_1212,N_1247);
xnor U1720 (N_1720,N_1130,N_1283);
nand U1721 (N_1721,N_1331,N_1066);
and U1722 (N_1722,N_1119,N_1239);
xor U1723 (N_1723,N_1462,N_1296);
or U1724 (N_1724,N_1374,N_1031);
nor U1725 (N_1725,N_1123,N_1280);
or U1726 (N_1726,N_1244,N_1085);
nand U1727 (N_1727,N_1092,N_1453);
and U1728 (N_1728,N_1258,N_1088);
nor U1729 (N_1729,N_1474,N_1110);
nor U1730 (N_1730,N_1128,N_1349);
or U1731 (N_1731,N_1158,N_1018);
and U1732 (N_1732,N_1133,N_1017);
and U1733 (N_1733,N_1310,N_1176);
and U1734 (N_1734,N_1424,N_1432);
and U1735 (N_1735,N_1185,N_1222);
or U1736 (N_1736,N_1342,N_1326);
or U1737 (N_1737,N_1325,N_1499);
nand U1738 (N_1738,N_1163,N_1312);
and U1739 (N_1739,N_1114,N_1036);
nand U1740 (N_1740,N_1035,N_1281);
xor U1741 (N_1741,N_1113,N_1288);
xnor U1742 (N_1742,N_1363,N_1001);
nor U1743 (N_1743,N_1237,N_1120);
or U1744 (N_1744,N_1425,N_1207);
nor U1745 (N_1745,N_1011,N_1233);
or U1746 (N_1746,N_1008,N_1195);
nand U1747 (N_1747,N_1145,N_1016);
xnor U1748 (N_1748,N_1109,N_1115);
or U1749 (N_1749,N_1470,N_1406);
or U1750 (N_1750,N_1020,N_1331);
and U1751 (N_1751,N_1104,N_1150);
nor U1752 (N_1752,N_1209,N_1080);
xor U1753 (N_1753,N_1319,N_1006);
nor U1754 (N_1754,N_1247,N_1138);
nor U1755 (N_1755,N_1417,N_1050);
and U1756 (N_1756,N_1217,N_1375);
xor U1757 (N_1757,N_1258,N_1045);
xor U1758 (N_1758,N_1041,N_1408);
xor U1759 (N_1759,N_1366,N_1023);
nand U1760 (N_1760,N_1149,N_1028);
xor U1761 (N_1761,N_1299,N_1379);
nand U1762 (N_1762,N_1237,N_1016);
or U1763 (N_1763,N_1083,N_1048);
nand U1764 (N_1764,N_1403,N_1052);
nand U1765 (N_1765,N_1112,N_1130);
and U1766 (N_1766,N_1196,N_1469);
and U1767 (N_1767,N_1127,N_1364);
and U1768 (N_1768,N_1154,N_1382);
or U1769 (N_1769,N_1087,N_1441);
nor U1770 (N_1770,N_1019,N_1237);
xor U1771 (N_1771,N_1267,N_1049);
nand U1772 (N_1772,N_1487,N_1152);
or U1773 (N_1773,N_1194,N_1032);
or U1774 (N_1774,N_1368,N_1450);
and U1775 (N_1775,N_1218,N_1372);
or U1776 (N_1776,N_1087,N_1351);
nor U1777 (N_1777,N_1232,N_1115);
nor U1778 (N_1778,N_1003,N_1343);
or U1779 (N_1779,N_1412,N_1131);
nand U1780 (N_1780,N_1469,N_1399);
nor U1781 (N_1781,N_1121,N_1305);
and U1782 (N_1782,N_1300,N_1111);
or U1783 (N_1783,N_1228,N_1054);
or U1784 (N_1784,N_1340,N_1455);
and U1785 (N_1785,N_1397,N_1358);
nand U1786 (N_1786,N_1478,N_1196);
and U1787 (N_1787,N_1270,N_1010);
and U1788 (N_1788,N_1276,N_1414);
and U1789 (N_1789,N_1167,N_1408);
or U1790 (N_1790,N_1442,N_1462);
nor U1791 (N_1791,N_1156,N_1371);
and U1792 (N_1792,N_1357,N_1319);
nor U1793 (N_1793,N_1385,N_1376);
and U1794 (N_1794,N_1401,N_1217);
nor U1795 (N_1795,N_1194,N_1024);
and U1796 (N_1796,N_1362,N_1319);
or U1797 (N_1797,N_1450,N_1145);
or U1798 (N_1798,N_1112,N_1450);
nor U1799 (N_1799,N_1373,N_1235);
and U1800 (N_1800,N_1402,N_1431);
or U1801 (N_1801,N_1437,N_1232);
or U1802 (N_1802,N_1282,N_1389);
nor U1803 (N_1803,N_1008,N_1051);
nand U1804 (N_1804,N_1277,N_1201);
and U1805 (N_1805,N_1456,N_1122);
nor U1806 (N_1806,N_1100,N_1429);
nand U1807 (N_1807,N_1422,N_1447);
nor U1808 (N_1808,N_1429,N_1366);
nor U1809 (N_1809,N_1493,N_1290);
xnor U1810 (N_1810,N_1013,N_1130);
or U1811 (N_1811,N_1306,N_1369);
or U1812 (N_1812,N_1453,N_1039);
or U1813 (N_1813,N_1431,N_1278);
and U1814 (N_1814,N_1424,N_1153);
nor U1815 (N_1815,N_1396,N_1207);
nor U1816 (N_1816,N_1253,N_1406);
and U1817 (N_1817,N_1154,N_1165);
nand U1818 (N_1818,N_1472,N_1129);
and U1819 (N_1819,N_1253,N_1184);
nand U1820 (N_1820,N_1498,N_1419);
nor U1821 (N_1821,N_1004,N_1074);
xnor U1822 (N_1822,N_1169,N_1053);
nand U1823 (N_1823,N_1131,N_1193);
and U1824 (N_1824,N_1063,N_1273);
and U1825 (N_1825,N_1304,N_1486);
and U1826 (N_1826,N_1367,N_1228);
xor U1827 (N_1827,N_1163,N_1244);
and U1828 (N_1828,N_1218,N_1153);
nor U1829 (N_1829,N_1327,N_1190);
or U1830 (N_1830,N_1223,N_1468);
and U1831 (N_1831,N_1342,N_1218);
nor U1832 (N_1832,N_1117,N_1403);
or U1833 (N_1833,N_1484,N_1369);
nor U1834 (N_1834,N_1030,N_1178);
xnor U1835 (N_1835,N_1157,N_1401);
nor U1836 (N_1836,N_1244,N_1207);
and U1837 (N_1837,N_1476,N_1200);
xnor U1838 (N_1838,N_1454,N_1205);
and U1839 (N_1839,N_1118,N_1190);
or U1840 (N_1840,N_1106,N_1246);
or U1841 (N_1841,N_1364,N_1190);
xnor U1842 (N_1842,N_1420,N_1436);
xor U1843 (N_1843,N_1334,N_1019);
nand U1844 (N_1844,N_1235,N_1467);
xnor U1845 (N_1845,N_1233,N_1198);
xor U1846 (N_1846,N_1083,N_1463);
and U1847 (N_1847,N_1484,N_1034);
nand U1848 (N_1848,N_1389,N_1453);
nor U1849 (N_1849,N_1120,N_1063);
xor U1850 (N_1850,N_1177,N_1164);
and U1851 (N_1851,N_1188,N_1197);
and U1852 (N_1852,N_1292,N_1412);
nand U1853 (N_1853,N_1028,N_1052);
nand U1854 (N_1854,N_1096,N_1468);
or U1855 (N_1855,N_1317,N_1063);
and U1856 (N_1856,N_1084,N_1006);
xor U1857 (N_1857,N_1196,N_1294);
and U1858 (N_1858,N_1307,N_1235);
and U1859 (N_1859,N_1296,N_1088);
or U1860 (N_1860,N_1383,N_1387);
nand U1861 (N_1861,N_1019,N_1463);
or U1862 (N_1862,N_1499,N_1158);
nand U1863 (N_1863,N_1464,N_1070);
nand U1864 (N_1864,N_1129,N_1227);
or U1865 (N_1865,N_1134,N_1037);
and U1866 (N_1866,N_1198,N_1043);
and U1867 (N_1867,N_1324,N_1484);
nor U1868 (N_1868,N_1138,N_1117);
xor U1869 (N_1869,N_1000,N_1236);
and U1870 (N_1870,N_1393,N_1033);
nand U1871 (N_1871,N_1411,N_1253);
and U1872 (N_1872,N_1419,N_1418);
and U1873 (N_1873,N_1046,N_1204);
xor U1874 (N_1874,N_1377,N_1095);
nor U1875 (N_1875,N_1112,N_1080);
and U1876 (N_1876,N_1103,N_1038);
xnor U1877 (N_1877,N_1242,N_1153);
nand U1878 (N_1878,N_1109,N_1004);
or U1879 (N_1879,N_1058,N_1072);
and U1880 (N_1880,N_1052,N_1074);
nor U1881 (N_1881,N_1186,N_1157);
and U1882 (N_1882,N_1197,N_1404);
xor U1883 (N_1883,N_1106,N_1187);
and U1884 (N_1884,N_1328,N_1402);
or U1885 (N_1885,N_1197,N_1201);
nor U1886 (N_1886,N_1375,N_1298);
or U1887 (N_1887,N_1348,N_1152);
xnor U1888 (N_1888,N_1290,N_1225);
nor U1889 (N_1889,N_1230,N_1299);
nor U1890 (N_1890,N_1170,N_1348);
nand U1891 (N_1891,N_1338,N_1015);
xnor U1892 (N_1892,N_1415,N_1316);
xor U1893 (N_1893,N_1197,N_1030);
nand U1894 (N_1894,N_1262,N_1056);
nor U1895 (N_1895,N_1474,N_1419);
or U1896 (N_1896,N_1397,N_1139);
or U1897 (N_1897,N_1265,N_1222);
nand U1898 (N_1898,N_1110,N_1385);
nor U1899 (N_1899,N_1046,N_1117);
and U1900 (N_1900,N_1286,N_1303);
nor U1901 (N_1901,N_1332,N_1310);
nand U1902 (N_1902,N_1154,N_1410);
nand U1903 (N_1903,N_1220,N_1164);
nor U1904 (N_1904,N_1072,N_1412);
or U1905 (N_1905,N_1269,N_1161);
nand U1906 (N_1906,N_1012,N_1114);
nor U1907 (N_1907,N_1066,N_1214);
or U1908 (N_1908,N_1061,N_1333);
nor U1909 (N_1909,N_1466,N_1305);
nand U1910 (N_1910,N_1318,N_1136);
xnor U1911 (N_1911,N_1054,N_1070);
nand U1912 (N_1912,N_1220,N_1074);
or U1913 (N_1913,N_1318,N_1261);
nor U1914 (N_1914,N_1481,N_1294);
xor U1915 (N_1915,N_1177,N_1134);
or U1916 (N_1916,N_1188,N_1090);
and U1917 (N_1917,N_1039,N_1300);
or U1918 (N_1918,N_1187,N_1387);
and U1919 (N_1919,N_1190,N_1484);
and U1920 (N_1920,N_1163,N_1081);
nand U1921 (N_1921,N_1119,N_1019);
and U1922 (N_1922,N_1104,N_1374);
or U1923 (N_1923,N_1261,N_1009);
nor U1924 (N_1924,N_1012,N_1295);
or U1925 (N_1925,N_1227,N_1452);
nor U1926 (N_1926,N_1492,N_1053);
nor U1927 (N_1927,N_1465,N_1067);
nor U1928 (N_1928,N_1052,N_1201);
xnor U1929 (N_1929,N_1101,N_1263);
xor U1930 (N_1930,N_1387,N_1208);
or U1931 (N_1931,N_1372,N_1440);
xnor U1932 (N_1932,N_1419,N_1189);
xnor U1933 (N_1933,N_1266,N_1208);
and U1934 (N_1934,N_1290,N_1231);
and U1935 (N_1935,N_1295,N_1458);
nor U1936 (N_1936,N_1132,N_1207);
or U1937 (N_1937,N_1245,N_1010);
xnor U1938 (N_1938,N_1122,N_1125);
nand U1939 (N_1939,N_1002,N_1289);
nor U1940 (N_1940,N_1251,N_1393);
and U1941 (N_1941,N_1062,N_1433);
nand U1942 (N_1942,N_1291,N_1244);
xor U1943 (N_1943,N_1471,N_1239);
and U1944 (N_1944,N_1301,N_1095);
nand U1945 (N_1945,N_1029,N_1032);
nor U1946 (N_1946,N_1171,N_1499);
xnor U1947 (N_1947,N_1226,N_1042);
or U1948 (N_1948,N_1481,N_1486);
nand U1949 (N_1949,N_1090,N_1285);
or U1950 (N_1950,N_1063,N_1196);
and U1951 (N_1951,N_1406,N_1189);
nand U1952 (N_1952,N_1062,N_1037);
or U1953 (N_1953,N_1136,N_1491);
nor U1954 (N_1954,N_1056,N_1305);
nand U1955 (N_1955,N_1100,N_1493);
and U1956 (N_1956,N_1203,N_1452);
or U1957 (N_1957,N_1339,N_1011);
nor U1958 (N_1958,N_1364,N_1237);
nand U1959 (N_1959,N_1071,N_1358);
or U1960 (N_1960,N_1189,N_1040);
xnor U1961 (N_1961,N_1379,N_1234);
nand U1962 (N_1962,N_1494,N_1305);
or U1963 (N_1963,N_1457,N_1235);
xor U1964 (N_1964,N_1079,N_1287);
and U1965 (N_1965,N_1098,N_1464);
and U1966 (N_1966,N_1319,N_1444);
nor U1967 (N_1967,N_1161,N_1363);
xnor U1968 (N_1968,N_1367,N_1347);
xnor U1969 (N_1969,N_1083,N_1230);
nor U1970 (N_1970,N_1128,N_1118);
xnor U1971 (N_1971,N_1058,N_1204);
nand U1972 (N_1972,N_1181,N_1482);
xor U1973 (N_1973,N_1223,N_1229);
or U1974 (N_1974,N_1150,N_1043);
xor U1975 (N_1975,N_1342,N_1362);
xnor U1976 (N_1976,N_1079,N_1261);
xor U1977 (N_1977,N_1010,N_1347);
or U1978 (N_1978,N_1454,N_1091);
nand U1979 (N_1979,N_1423,N_1149);
xor U1980 (N_1980,N_1489,N_1069);
and U1981 (N_1981,N_1380,N_1154);
nand U1982 (N_1982,N_1476,N_1112);
or U1983 (N_1983,N_1360,N_1412);
nand U1984 (N_1984,N_1076,N_1470);
nor U1985 (N_1985,N_1060,N_1024);
nor U1986 (N_1986,N_1111,N_1060);
nor U1987 (N_1987,N_1142,N_1309);
xor U1988 (N_1988,N_1218,N_1418);
nand U1989 (N_1989,N_1099,N_1219);
nand U1990 (N_1990,N_1217,N_1281);
nand U1991 (N_1991,N_1106,N_1478);
xor U1992 (N_1992,N_1216,N_1259);
and U1993 (N_1993,N_1471,N_1260);
nand U1994 (N_1994,N_1412,N_1248);
and U1995 (N_1995,N_1028,N_1097);
xnor U1996 (N_1996,N_1150,N_1236);
and U1997 (N_1997,N_1222,N_1427);
or U1998 (N_1998,N_1487,N_1314);
or U1999 (N_1999,N_1410,N_1184);
nand U2000 (N_2000,N_1793,N_1850);
and U2001 (N_2001,N_1831,N_1991);
nor U2002 (N_2002,N_1860,N_1971);
and U2003 (N_2003,N_1821,N_1804);
xnor U2004 (N_2004,N_1689,N_1788);
nor U2005 (N_2005,N_1958,N_1923);
and U2006 (N_2006,N_1506,N_1531);
xor U2007 (N_2007,N_1735,N_1976);
or U2008 (N_2008,N_1630,N_1586);
nand U2009 (N_2009,N_1818,N_1786);
xnor U2010 (N_2010,N_1704,N_1887);
nand U2011 (N_2011,N_1798,N_1867);
xnor U2012 (N_2012,N_1766,N_1619);
xor U2013 (N_2013,N_1799,N_1683);
xnor U2014 (N_2014,N_1679,N_1741);
or U2015 (N_2015,N_1845,N_1714);
nor U2016 (N_2016,N_1589,N_1925);
xnor U2017 (N_2017,N_1864,N_1903);
xor U2018 (N_2018,N_1542,N_1848);
and U2019 (N_2019,N_1566,N_1885);
and U2020 (N_2020,N_1708,N_1994);
xor U2021 (N_2021,N_1792,N_1772);
or U2022 (N_2022,N_1745,N_1549);
nand U2023 (N_2023,N_1904,N_1762);
or U2024 (N_2024,N_1871,N_1776);
xor U2025 (N_2025,N_1604,N_1596);
nor U2026 (N_2026,N_1629,N_1802);
nor U2027 (N_2027,N_1832,N_1633);
or U2028 (N_2028,N_1677,N_1547);
nor U2029 (N_2029,N_1754,N_1657);
or U2030 (N_2030,N_1613,N_1882);
nand U2031 (N_2031,N_1599,N_1699);
nand U2032 (N_2032,N_1623,N_1628);
and U2033 (N_2033,N_1846,N_1855);
xnor U2034 (N_2034,N_1739,N_1526);
xnor U2035 (N_2035,N_1931,N_1934);
xnor U2036 (N_2036,N_1724,N_1866);
nand U2037 (N_2037,N_1890,N_1517);
nand U2038 (N_2038,N_1666,N_1511);
or U2039 (N_2039,N_1625,N_1889);
and U2040 (N_2040,N_1642,N_1954);
nand U2041 (N_2041,N_1686,N_1997);
nor U2042 (N_2042,N_1952,N_1847);
or U2043 (N_2043,N_1999,N_1896);
xor U2044 (N_2044,N_1988,N_1508);
nand U2045 (N_2045,N_1669,N_1600);
nand U2046 (N_2046,N_1513,N_1986);
and U2047 (N_2047,N_1873,N_1612);
nor U2048 (N_2048,N_1833,N_1587);
xor U2049 (N_2049,N_1869,N_1639);
and U2050 (N_2050,N_1715,N_1995);
or U2051 (N_2051,N_1702,N_1656);
nand U2052 (N_2052,N_1938,N_1554);
nor U2053 (N_2053,N_1909,N_1729);
xor U2054 (N_2054,N_1897,N_1533);
and U2055 (N_2055,N_1933,N_1945);
or U2056 (N_2056,N_1783,N_1912);
nor U2057 (N_2057,N_1543,N_1774);
and U2058 (N_2058,N_1911,N_1528);
and U2059 (N_2059,N_1981,N_1921);
and U2060 (N_2060,N_1602,N_1555);
and U2061 (N_2061,N_1725,N_1539);
xor U2062 (N_2062,N_1615,N_1658);
nand U2063 (N_2063,N_1722,N_1881);
xnor U2064 (N_2064,N_1789,N_1915);
and U2065 (N_2065,N_1919,N_1693);
nor U2066 (N_2066,N_1521,N_1744);
and U2067 (N_2067,N_1757,N_1536);
nand U2068 (N_2068,N_1721,N_1593);
nand U2069 (N_2069,N_1849,N_1730);
or U2070 (N_2070,N_1734,N_1634);
or U2071 (N_2071,N_1537,N_1863);
and U2072 (N_2072,N_1961,N_1578);
xor U2073 (N_2073,N_1910,N_1718);
nor U2074 (N_2074,N_1501,N_1719);
nand U2075 (N_2075,N_1514,N_1857);
xnor U2076 (N_2076,N_1892,N_1582);
xor U2077 (N_2077,N_1532,N_1842);
nand U2078 (N_2078,N_1862,N_1756);
or U2079 (N_2079,N_1812,N_1510);
nor U2080 (N_2080,N_1970,N_1703);
or U2081 (N_2081,N_1787,N_1894);
and U2082 (N_2082,N_1993,N_1740);
or U2083 (N_2083,N_1579,N_1837);
and U2084 (N_2084,N_1784,N_1825);
nand U2085 (N_2085,N_1843,N_1667);
nor U2086 (N_2086,N_1879,N_1975);
or U2087 (N_2087,N_1810,N_1559);
nand U2088 (N_2088,N_1968,N_1632);
and U2089 (N_2089,N_1983,N_1678);
and U2090 (N_2090,N_1760,N_1636);
and U2091 (N_2091,N_1583,N_1764);
nand U2092 (N_2092,N_1808,N_1935);
nand U2093 (N_2093,N_1717,N_1965);
xor U2094 (N_2094,N_1705,N_1814);
or U2095 (N_2095,N_1541,N_1820);
xnor U2096 (N_2096,N_1569,N_1858);
xor U2097 (N_2097,N_1564,N_1753);
or U2098 (N_2098,N_1824,N_1626);
and U2099 (N_2099,N_1813,N_1861);
xor U2100 (N_2100,N_1989,N_1829);
xnor U2101 (N_2101,N_1967,N_1807);
nor U2102 (N_2102,N_1617,N_1936);
nor U2103 (N_2103,N_1771,N_1560);
xor U2104 (N_2104,N_1643,N_1969);
nor U2105 (N_2105,N_1763,N_1709);
and U2106 (N_2106,N_1877,N_1777);
nor U2107 (N_2107,N_1844,N_1665);
nand U2108 (N_2108,N_1811,N_1752);
nor U2109 (N_2109,N_1778,N_1738);
or U2110 (N_2110,N_1584,N_1562);
and U2111 (N_2111,N_1621,N_1716);
or U2112 (N_2112,N_1926,N_1782);
nor U2113 (N_2113,N_1822,N_1962);
xor U2114 (N_2114,N_1751,N_1640);
xor U2115 (N_2115,N_1817,N_1594);
nor U2116 (N_2116,N_1690,N_1980);
nand U2117 (N_2117,N_1797,N_1960);
and U2118 (N_2118,N_1876,N_1875);
nand U2119 (N_2119,N_1736,N_1966);
nand U2120 (N_2120,N_1785,N_1920);
nand U2121 (N_2121,N_1803,N_1561);
or U2122 (N_2122,N_1567,N_1828);
nand U2123 (N_2123,N_1801,N_1504);
xor U2124 (N_2124,N_1950,N_1978);
xor U2125 (N_2125,N_1611,N_1840);
and U2126 (N_2126,N_1609,N_1556);
xnor U2127 (N_2127,N_1916,N_1512);
nand U2128 (N_2128,N_1701,N_1868);
nor U2129 (N_2129,N_1758,N_1688);
or U2130 (N_2130,N_1949,N_1522);
nor U2131 (N_2131,N_1550,N_1509);
xnor U2132 (N_2132,N_1670,N_1598);
and U2133 (N_2133,N_1838,N_1823);
nand U2134 (N_2134,N_1710,N_1700);
xor U2135 (N_2135,N_1947,N_1618);
and U2136 (N_2136,N_1859,N_1548);
xnor U2137 (N_2137,N_1518,N_1647);
nand U2138 (N_2138,N_1992,N_1796);
or U2139 (N_2139,N_1886,N_1750);
nand U2140 (N_2140,N_1930,N_1530);
nor U2141 (N_2141,N_1963,N_1726);
and U2142 (N_2142,N_1515,N_1595);
and U2143 (N_2143,N_1565,N_1905);
nor U2144 (N_2144,N_1806,N_1856);
nand U2145 (N_2145,N_1768,N_1918);
xor U2146 (N_2146,N_1637,N_1638);
and U2147 (N_2147,N_1507,N_1898);
or U2148 (N_2148,N_1749,N_1676);
or U2149 (N_2149,N_1500,N_1675);
nor U2150 (N_2150,N_1695,N_1607);
xor U2151 (N_2151,N_1941,N_1544);
or U2152 (N_2152,N_1851,N_1523);
nor U2153 (N_2153,N_1815,N_1557);
or U2154 (N_2154,N_1672,N_1723);
xor U2155 (N_2155,N_1652,N_1805);
nor U2156 (N_2156,N_1767,N_1570);
nand U2157 (N_2157,N_1924,N_1895);
nand U2158 (N_2158,N_1552,N_1616);
and U2159 (N_2159,N_1940,N_1592);
and U2160 (N_2160,N_1891,N_1917);
and U2161 (N_2161,N_1932,N_1697);
nor U2162 (N_2162,N_1728,N_1694);
xnor U2163 (N_2163,N_1692,N_1955);
or U2164 (N_2164,N_1827,N_1835);
nand U2165 (N_2165,N_1977,N_1819);
and U2166 (N_2166,N_1527,N_1575);
xnor U2167 (N_2167,N_1780,N_1631);
xnor U2168 (N_2168,N_1576,N_1707);
xor U2169 (N_2169,N_1538,N_1770);
nor U2170 (N_2170,N_1671,N_1928);
and U2171 (N_2171,N_1635,N_1908);
and U2172 (N_2172,N_1650,N_1839);
xor U2173 (N_2173,N_1899,N_1922);
and U2174 (N_2174,N_1585,N_1742);
nor U2175 (N_2175,N_1668,N_1577);
and U2176 (N_2176,N_1588,N_1684);
and U2177 (N_2177,N_1534,N_1563);
or U2178 (N_2178,N_1505,N_1608);
nand U2179 (N_2179,N_1959,N_1568);
nor U2180 (N_2180,N_1591,N_1956);
xor U2181 (N_2181,N_1791,N_1893);
nor U2182 (N_2182,N_1957,N_1880);
or U2183 (N_2183,N_1914,N_1525);
xnor U2184 (N_2184,N_1622,N_1545);
nor U2185 (N_2185,N_1964,N_1651);
xnor U2186 (N_2186,N_1900,N_1743);
nor U2187 (N_2187,N_1929,N_1990);
nand U2188 (N_2188,N_1951,N_1878);
nand U2189 (N_2189,N_1946,N_1907);
xnor U2190 (N_2190,N_1759,N_1737);
nand U2191 (N_2191,N_1673,N_1769);
and U2192 (N_2192,N_1502,N_1661);
and U2193 (N_2193,N_1888,N_1836);
nor U2194 (N_2194,N_1746,N_1901);
nand U2195 (N_2195,N_1503,N_1641);
nor U2196 (N_2196,N_1727,N_1685);
or U2197 (N_2197,N_1996,N_1597);
nor U2198 (N_2198,N_1681,N_1646);
nand U2199 (N_2199,N_1800,N_1590);
or U2200 (N_2200,N_1558,N_1942);
and U2201 (N_2201,N_1551,N_1606);
and U2202 (N_2202,N_1655,N_1627);
nor U2203 (N_2203,N_1654,N_1906);
and U2204 (N_2204,N_1872,N_1733);
nand U2205 (N_2205,N_1937,N_1540);
or U2206 (N_2206,N_1614,N_1865);
xnor U2207 (N_2207,N_1573,N_1982);
xor U2208 (N_2208,N_1790,N_1645);
nand U2209 (N_2209,N_1553,N_1546);
nor U2210 (N_2210,N_1748,N_1696);
nor U2211 (N_2211,N_1826,N_1712);
or U2212 (N_2212,N_1765,N_1747);
xnor U2213 (N_2213,N_1610,N_1662);
nand U2214 (N_2214,N_1974,N_1659);
and U2215 (N_2215,N_1620,N_1535);
nand U2216 (N_2216,N_1841,N_1948);
xnor U2217 (N_2217,N_1581,N_1816);
and U2218 (N_2218,N_1713,N_1674);
nand U2219 (N_2219,N_1572,N_1939);
or U2220 (N_2220,N_1720,N_1687);
and U2221 (N_2221,N_1682,N_1884);
nand U2222 (N_2222,N_1998,N_1601);
or U2223 (N_2223,N_1516,N_1603);
nand U2224 (N_2224,N_1698,N_1660);
nand U2225 (N_2225,N_1571,N_1644);
and U2226 (N_2226,N_1913,N_1985);
nor U2227 (N_2227,N_1711,N_1809);
and U2228 (N_2228,N_1834,N_1927);
nand U2229 (N_2229,N_1520,N_1902);
or U2230 (N_2230,N_1732,N_1574);
xnor U2231 (N_2231,N_1649,N_1987);
nand U2232 (N_2232,N_1779,N_1663);
and U2233 (N_2233,N_1852,N_1605);
or U2234 (N_2234,N_1883,N_1624);
nand U2235 (N_2235,N_1524,N_1984);
or U2236 (N_2236,N_1664,N_1870);
or U2237 (N_2237,N_1944,N_1706);
nand U2238 (N_2238,N_1755,N_1781);
and U2239 (N_2239,N_1653,N_1794);
xnor U2240 (N_2240,N_1691,N_1761);
and U2241 (N_2241,N_1972,N_1854);
and U2242 (N_2242,N_1648,N_1795);
nor U2243 (N_2243,N_1773,N_1973);
nor U2244 (N_2244,N_1519,N_1580);
nand U2245 (N_2245,N_1731,N_1943);
nor U2246 (N_2246,N_1874,N_1680);
or U2247 (N_2247,N_1979,N_1529);
nand U2248 (N_2248,N_1830,N_1853);
nand U2249 (N_2249,N_1775,N_1953);
nand U2250 (N_2250,N_1645,N_1555);
and U2251 (N_2251,N_1590,N_1722);
or U2252 (N_2252,N_1737,N_1968);
or U2253 (N_2253,N_1767,N_1647);
nor U2254 (N_2254,N_1867,N_1628);
nor U2255 (N_2255,N_1623,N_1546);
nor U2256 (N_2256,N_1600,N_1707);
and U2257 (N_2257,N_1574,N_1716);
and U2258 (N_2258,N_1579,N_1685);
nand U2259 (N_2259,N_1585,N_1526);
nor U2260 (N_2260,N_1597,N_1946);
and U2261 (N_2261,N_1554,N_1538);
nand U2262 (N_2262,N_1781,N_1599);
xnor U2263 (N_2263,N_1580,N_1757);
nand U2264 (N_2264,N_1698,N_1935);
and U2265 (N_2265,N_1633,N_1954);
and U2266 (N_2266,N_1558,N_1582);
or U2267 (N_2267,N_1869,N_1823);
xor U2268 (N_2268,N_1587,N_1719);
nand U2269 (N_2269,N_1763,N_1989);
nor U2270 (N_2270,N_1979,N_1804);
nor U2271 (N_2271,N_1622,N_1921);
and U2272 (N_2272,N_1959,N_1864);
or U2273 (N_2273,N_1718,N_1960);
xor U2274 (N_2274,N_1739,N_1765);
and U2275 (N_2275,N_1658,N_1594);
or U2276 (N_2276,N_1798,N_1584);
and U2277 (N_2277,N_1582,N_1806);
nand U2278 (N_2278,N_1593,N_1881);
and U2279 (N_2279,N_1694,N_1845);
xnor U2280 (N_2280,N_1754,N_1711);
or U2281 (N_2281,N_1673,N_1997);
xor U2282 (N_2282,N_1836,N_1842);
nor U2283 (N_2283,N_1878,N_1912);
xnor U2284 (N_2284,N_1568,N_1744);
nor U2285 (N_2285,N_1874,N_1990);
nor U2286 (N_2286,N_1739,N_1563);
nor U2287 (N_2287,N_1667,N_1771);
and U2288 (N_2288,N_1632,N_1824);
nand U2289 (N_2289,N_1994,N_1636);
nand U2290 (N_2290,N_1645,N_1600);
nor U2291 (N_2291,N_1975,N_1704);
nor U2292 (N_2292,N_1599,N_1765);
and U2293 (N_2293,N_1943,N_1772);
nor U2294 (N_2294,N_1999,N_1555);
nand U2295 (N_2295,N_1906,N_1819);
nand U2296 (N_2296,N_1855,N_1561);
or U2297 (N_2297,N_1530,N_1619);
nor U2298 (N_2298,N_1735,N_1669);
xnor U2299 (N_2299,N_1711,N_1538);
and U2300 (N_2300,N_1533,N_1855);
xor U2301 (N_2301,N_1830,N_1615);
nand U2302 (N_2302,N_1707,N_1930);
or U2303 (N_2303,N_1766,N_1675);
and U2304 (N_2304,N_1652,N_1740);
nand U2305 (N_2305,N_1796,N_1533);
xnor U2306 (N_2306,N_1818,N_1830);
xnor U2307 (N_2307,N_1628,N_1992);
xor U2308 (N_2308,N_1782,N_1723);
or U2309 (N_2309,N_1689,N_1598);
nand U2310 (N_2310,N_1751,N_1670);
or U2311 (N_2311,N_1544,N_1536);
or U2312 (N_2312,N_1502,N_1664);
or U2313 (N_2313,N_1734,N_1864);
xnor U2314 (N_2314,N_1774,N_1854);
nand U2315 (N_2315,N_1614,N_1916);
nand U2316 (N_2316,N_1641,N_1515);
and U2317 (N_2317,N_1819,N_1871);
nand U2318 (N_2318,N_1588,N_1806);
and U2319 (N_2319,N_1619,N_1621);
and U2320 (N_2320,N_1621,N_1999);
and U2321 (N_2321,N_1946,N_1761);
nand U2322 (N_2322,N_1678,N_1985);
or U2323 (N_2323,N_1546,N_1947);
or U2324 (N_2324,N_1713,N_1709);
xor U2325 (N_2325,N_1966,N_1583);
nand U2326 (N_2326,N_1700,N_1919);
xor U2327 (N_2327,N_1994,N_1661);
xnor U2328 (N_2328,N_1964,N_1869);
nand U2329 (N_2329,N_1928,N_1935);
nor U2330 (N_2330,N_1588,N_1587);
nand U2331 (N_2331,N_1757,N_1702);
nor U2332 (N_2332,N_1721,N_1564);
nor U2333 (N_2333,N_1747,N_1996);
nand U2334 (N_2334,N_1806,N_1818);
or U2335 (N_2335,N_1841,N_1748);
xnor U2336 (N_2336,N_1581,N_1874);
nor U2337 (N_2337,N_1581,N_1623);
nor U2338 (N_2338,N_1715,N_1575);
and U2339 (N_2339,N_1717,N_1792);
and U2340 (N_2340,N_1501,N_1534);
and U2341 (N_2341,N_1928,N_1911);
and U2342 (N_2342,N_1787,N_1663);
xnor U2343 (N_2343,N_1661,N_1549);
xnor U2344 (N_2344,N_1956,N_1564);
nor U2345 (N_2345,N_1778,N_1685);
nor U2346 (N_2346,N_1611,N_1602);
and U2347 (N_2347,N_1573,N_1662);
xnor U2348 (N_2348,N_1867,N_1719);
or U2349 (N_2349,N_1890,N_1713);
nand U2350 (N_2350,N_1997,N_1684);
nor U2351 (N_2351,N_1559,N_1707);
nand U2352 (N_2352,N_1915,N_1768);
or U2353 (N_2353,N_1565,N_1825);
and U2354 (N_2354,N_1684,N_1539);
xor U2355 (N_2355,N_1839,N_1974);
or U2356 (N_2356,N_1512,N_1907);
nor U2357 (N_2357,N_1872,N_1725);
or U2358 (N_2358,N_1576,N_1982);
or U2359 (N_2359,N_1515,N_1854);
or U2360 (N_2360,N_1682,N_1762);
or U2361 (N_2361,N_1829,N_1879);
nand U2362 (N_2362,N_1584,N_1800);
or U2363 (N_2363,N_1853,N_1763);
or U2364 (N_2364,N_1804,N_1654);
nor U2365 (N_2365,N_1888,N_1534);
and U2366 (N_2366,N_1668,N_1595);
and U2367 (N_2367,N_1779,N_1861);
nand U2368 (N_2368,N_1972,N_1879);
xnor U2369 (N_2369,N_1720,N_1516);
nand U2370 (N_2370,N_1906,N_1714);
xor U2371 (N_2371,N_1966,N_1546);
and U2372 (N_2372,N_1879,N_1720);
xnor U2373 (N_2373,N_1823,N_1814);
nor U2374 (N_2374,N_1820,N_1957);
and U2375 (N_2375,N_1676,N_1648);
nor U2376 (N_2376,N_1594,N_1640);
xor U2377 (N_2377,N_1874,N_1667);
or U2378 (N_2378,N_1901,N_1978);
nand U2379 (N_2379,N_1895,N_1592);
or U2380 (N_2380,N_1756,N_1929);
nand U2381 (N_2381,N_1913,N_1772);
or U2382 (N_2382,N_1519,N_1672);
or U2383 (N_2383,N_1755,N_1545);
nor U2384 (N_2384,N_1576,N_1951);
nand U2385 (N_2385,N_1986,N_1747);
nand U2386 (N_2386,N_1503,N_1695);
nand U2387 (N_2387,N_1719,N_1931);
nor U2388 (N_2388,N_1751,N_1655);
and U2389 (N_2389,N_1886,N_1773);
xor U2390 (N_2390,N_1992,N_1611);
or U2391 (N_2391,N_1740,N_1863);
nand U2392 (N_2392,N_1713,N_1624);
or U2393 (N_2393,N_1890,N_1977);
and U2394 (N_2394,N_1645,N_1902);
nand U2395 (N_2395,N_1518,N_1958);
xor U2396 (N_2396,N_1518,N_1981);
and U2397 (N_2397,N_1570,N_1754);
xnor U2398 (N_2398,N_1744,N_1613);
xor U2399 (N_2399,N_1666,N_1567);
and U2400 (N_2400,N_1616,N_1648);
nor U2401 (N_2401,N_1592,N_1682);
xnor U2402 (N_2402,N_1643,N_1757);
and U2403 (N_2403,N_1830,N_1598);
xnor U2404 (N_2404,N_1647,N_1918);
nand U2405 (N_2405,N_1612,N_1540);
or U2406 (N_2406,N_1786,N_1522);
or U2407 (N_2407,N_1777,N_1978);
and U2408 (N_2408,N_1568,N_1882);
nor U2409 (N_2409,N_1746,N_1641);
xnor U2410 (N_2410,N_1642,N_1892);
nor U2411 (N_2411,N_1553,N_1694);
and U2412 (N_2412,N_1604,N_1670);
xor U2413 (N_2413,N_1598,N_1805);
xor U2414 (N_2414,N_1729,N_1886);
nand U2415 (N_2415,N_1952,N_1638);
nand U2416 (N_2416,N_1986,N_1566);
and U2417 (N_2417,N_1500,N_1700);
or U2418 (N_2418,N_1532,N_1764);
nor U2419 (N_2419,N_1509,N_1560);
xnor U2420 (N_2420,N_1811,N_1813);
xor U2421 (N_2421,N_1706,N_1605);
or U2422 (N_2422,N_1610,N_1896);
or U2423 (N_2423,N_1663,N_1783);
xnor U2424 (N_2424,N_1735,N_1662);
xor U2425 (N_2425,N_1564,N_1701);
nand U2426 (N_2426,N_1851,N_1989);
or U2427 (N_2427,N_1590,N_1967);
nor U2428 (N_2428,N_1757,N_1504);
xnor U2429 (N_2429,N_1848,N_1997);
and U2430 (N_2430,N_1815,N_1785);
or U2431 (N_2431,N_1844,N_1767);
or U2432 (N_2432,N_1836,N_1633);
xnor U2433 (N_2433,N_1984,N_1555);
nor U2434 (N_2434,N_1786,N_1529);
or U2435 (N_2435,N_1720,N_1864);
nor U2436 (N_2436,N_1761,N_1885);
and U2437 (N_2437,N_1951,N_1870);
or U2438 (N_2438,N_1894,N_1640);
and U2439 (N_2439,N_1807,N_1725);
and U2440 (N_2440,N_1613,N_1524);
xnor U2441 (N_2441,N_1721,N_1892);
and U2442 (N_2442,N_1957,N_1696);
and U2443 (N_2443,N_1594,N_1964);
nor U2444 (N_2444,N_1537,N_1737);
xnor U2445 (N_2445,N_1504,N_1574);
and U2446 (N_2446,N_1923,N_1763);
nor U2447 (N_2447,N_1875,N_1903);
and U2448 (N_2448,N_1673,N_1585);
nand U2449 (N_2449,N_1507,N_1727);
and U2450 (N_2450,N_1736,N_1559);
nand U2451 (N_2451,N_1574,N_1953);
xor U2452 (N_2452,N_1523,N_1741);
nand U2453 (N_2453,N_1976,N_1897);
xnor U2454 (N_2454,N_1910,N_1890);
nor U2455 (N_2455,N_1856,N_1522);
and U2456 (N_2456,N_1673,N_1621);
and U2457 (N_2457,N_1520,N_1828);
nor U2458 (N_2458,N_1703,N_1597);
and U2459 (N_2459,N_1625,N_1552);
or U2460 (N_2460,N_1667,N_1867);
nand U2461 (N_2461,N_1753,N_1546);
nor U2462 (N_2462,N_1552,N_1907);
nand U2463 (N_2463,N_1579,N_1648);
xnor U2464 (N_2464,N_1811,N_1658);
or U2465 (N_2465,N_1687,N_1620);
nand U2466 (N_2466,N_1795,N_1843);
and U2467 (N_2467,N_1828,N_1710);
nand U2468 (N_2468,N_1731,N_1846);
and U2469 (N_2469,N_1695,N_1561);
nor U2470 (N_2470,N_1650,N_1913);
nor U2471 (N_2471,N_1888,N_1819);
or U2472 (N_2472,N_1830,N_1807);
and U2473 (N_2473,N_1988,N_1997);
xnor U2474 (N_2474,N_1724,N_1940);
xnor U2475 (N_2475,N_1686,N_1850);
xnor U2476 (N_2476,N_1745,N_1767);
nand U2477 (N_2477,N_1951,N_1729);
nor U2478 (N_2478,N_1659,N_1784);
or U2479 (N_2479,N_1965,N_1691);
or U2480 (N_2480,N_1850,N_1791);
and U2481 (N_2481,N_1673,N_1876);
and U2482 (N_2482,N_1916,N_1847);
and U2483 (N_2483,N_1702,N_1668);
or U2484 (N_2484,N_1866,N_1531);
or U2485 (N_2485,N_1747,N_1583);
nand U2486 (N_2486,N_1657,N_1973);
nand U2487 (N_2487,N_1793,N_1753);
nand U2488 (N_2488,N_1736,N_1663);
and U2489 (N_2489,N_1900,N_1678);
xnor U2490 (N_2490,N_1737,N_1803);
and U2491 (N_2491,N_1783,N_1722);
xnor U2492 (N_2492,N_1583,N_1846);
nor U2493 (N_2493,N_1977,N_1573);
xnor U2494 (N_2494,N_1893,N_1745);
and U2495 (N_2495,N_1615,N_1650);
xor U2496 (N_2496,N_1948,N_1781);
nor U2497 (N_2497,N_1787,N_1982);
nor U2498 (N_2498,N_1629,N_1804);
and U2499 (N_2499,N_1850,N_1595);
xnor U2500 (N_2500,N_2330,N_2002);
xor U2501 (N_2501,N_2094,N_2498);
nor U2502 (N_2502,N_2285,N_2365);
nand U2503 (N_2503,N_2339,N_2407);
nand U2504 (N_2504,N_2359,N_2165);
nor U2505 (N_2505,N_2401,N_2026);
or U2506 (N_2506,N_2448,N_2430);
or U2507 (N_2507,N_2280,N_2218);
and U2508 (N_2508,N_2289,N_2173);
and U2509 (N_2509,N_2308,N_2356);
or U2510 (N_2510,N_2471,N_2248);
and U2511 (N_2511,N_2244,N_2364);
or U2512 (N_2512,N_2159,N_2467);
nand U2513 (N_2513,N_2425,N_2465);
or U2514 (N_2514,N_2001,N_2306);
xor U2515 (N_2515,N_2117,N_2442);
xnor U2516 (N_2516,N_2437,N_2399);
nand U2517 (N_2517,N_2362,N_2441);
xor U2518 (N_2518,N_2347,N_2294);
xnor U2519 (N_2519,N_2110,N_2046);
and U2520 (N_2520,N_2403,N_2411);
xnor U2521 (N_2521,N_2491,N_2469);
and U2522 (N_2522,N_2231,N_2319);
and U2523 (N_2523,N_2355,N_2346);
or U2524 (N_2524,N_2220,N_2102);
or U2525 (N_2525,N_2088,N_2238);
xor U2526 (N_2526,N_2418,N_2071);
nand U2527 (N_2527,N_2064,N_2291);
nand U2528 (N_2528,N_2039,N_2196);
xnor U2529 (N_2529,N_2156,N_2379);
or U2530 (N_2530,N_2472,N_2006);
or U2531 (N_2531,N_2348,N_2481);
or U2532 (N_2532,N_2149,N_2367);
and U2533 (N_2533,N_2022,N_2462);
nor U2534 (N_2534,N_2052,N_2181);
xor U2535 (N_2535,N_2300,N_2482);
nor U2536 (N_2536,N_2353,N_2409);
nor U2537 (N_2537,N_2487,N_2408);
nor U2538 (N_2538,N_2322,N_2390);
and U2539 (N_2539,N_2394,N_2420);
or U2540 (N_2540,N_2233,N_2416);
nor U2541 (N_2541,N_2301,N_2092);
nand U2542 (N_2542,N_2323,N_2192);
and U2543 (N_2543,N_2259,N_2205);
and U2544 (N_2544,N_2337,N_2386);
or U2545 (N_2545,N_2107,N_2007);
nand U2546 (N_2546,N_2009,N_2225);
nor U2547 (N_2547,N_2402,N_2393);
xnor U2548 (N_2548,N_2254,N_2184);
or U2549 (N_2549,N_2056,N_2211);
nand U2550 (N_2550,N_2243,N_2201);
xor U2551 (N_2551,N_2179,N_2320);
and U2552 (N_2552,N_2455,N_2397);
nand U2553 (N_2553,N_2119,N_2313);
or U2554 (N_2554,N_2068,N_2219);
nor U2555 (N_2555,N_2395,N_2368);
and U2556 (N_2556,N_2299,N_2032);
xor U2557 (N_2557,N_2494,N_2097);
or U2558 (N_2558,N_2154,N_2457);
or U2559 (N_2559,N_2050,N_2011);
xor U2560 (N_2560,N_2069,N_2459);
and U2561 (N_2561,N_2072,N_2264);
xor U2562 (N_2562,N_2153,N_2090);
nand U2563 (N_2563,N_2261,N_2336);
nand U2564 (N_2564,N_2369,N_2172);
nor U2565 (N_2565,N_2163,N_2311);
xnor U2566 (N_2566,N_2164,N_2490);
nor U2567 (N_2567,N_2054,N_2429);
nand U2568 (N_2568,N_2450,N_2398);
nand U2569 (N_2569,N_2496,N_2096);
xor U2570 (N_2570,N_2489,N_2332);
nor U2571 (N_2571,N_2152,N_2255);
nand U2572 (N_2572,N_2229,N_2035);
xnor U2573 (N_2573,N_2423,N_2115);
xnor U2574 (N_2574,N_2295,N_2005);
xnor U2575 (N_2575,N_2384,N_2488);
nand U2576 (N_2576,N_2282,N_2155);
nand U2577 (N_2577,N_2334,N_2449);
and U2578 (N_2578,N_2131,N_2422);
xnor U2579 (N_2579,N_2093,N_2008);
nand U2580 (N_2580,N_2185,N_2036);
nor U2581 (N_2581,N_2486,N_2215);
xor U2582 (N_2582,N_2475,N_2098);
and U2583 (N_2583,N_2373,N_2105);
nor U2584 (N_2584,N_2053,N_2345);
or U2585 (N_2585,N_2175,N_2250);
and U2586 (N_2586,N_2171,N_2344);
nor U2587 (N_2587,N_2112,N_2023);
and U2588 (N_2588,N_2309,N_2141);
or U2589 (N_2589,N_2195,N_2410);
nor U2590 (N_2590,N_2451,N_2197);
or U2591 (N_2591,N_2101,N_2366);
nand U2592 (N_2592,N_2066,N_2456);
xnor U2593 (N_2593,N_2142,N_2081);
nor U2594 (N_2594,N_2341,N_2061);
nor U2595 (N_2595,N_2342,N_2360);
or U2596 (N_2596,N_2321,N_2147);
or U2597 (N_2597,N_2439,N_2024);
nand U2598 (N_2598,N_2000,N_2380);
nor U2599 (N_2599,N_2166,N_2004);
and U2600 (N_2600,N_2424,N_2129);
nor U2601 (N_2601,N_2303,N_2431);
and U2602 (N_2602,N_2060,N_2378);
nor U2603 (N_2603,N_2350,N_2202);
xor U2604 (N_2604,N_2241,N_2038);
nor U2605 (N_2605,N_2176,N_2417);
and U2606 (N_2606,N_2003,N_2329);
nor U2607 (N_2607,N_2432,N_2389);
xor U2608 (N_2608,N_2239,N_2076);
or U2609 (N_2609,N_2468,N_2249);
nor U2610 (N_2610,N_2351,N_2130);
or U2611 (N_2611,N_2288,N_2314);
and U2612 (N_2612,N_2278,N_2221);
nor U2613 (N_2613,N_2144,N_2213);
nor U2614 (N_2614,N_2100,N_2349);
and U2615 (N_2615,N_2017,N_2287);
or U2616 (N_2616,N_2392,N_2376);
nand U2617 (N_2617,N_2284,N_2232);
xor U2618 (N_2618,N_2271,N_2041);
or U2619 (N_2619,N_2474,N_2157);
nand U2620 (N_2620,N_2020,N_2025);
nand U2621 (N_2621,N_2048,N_2018);
nor U2622 (N_2622,N_2116,N_2310);
nand U2623 (N_2623,N_2082,N_2492);
xnor U2624 (N_2624,N_2143,N_2358);
and U2625 (N_2625,N_2019,N_2325);
nand U2626 (N_2626,N_2135,N_2391);
xnor U2627 (N_2627,N_2252,N_2274);
or U2628 (N_2628,N_2224,N_2139);
nor U2629 (N_2629,N_2150,N_2447);
or U2630 (N_2630,N_2208,N_2027);
xor U2631 (N_2631,N_2145,N_2466);
nand U2632 (N_2632,N_2108,N_2083);
or U2633 (N_2633,N_2304,N_2037);
or U2634 (N_2634,N_2148,N_2340);
and U2635 (N_2635,N_2222,N_2089);
nand U2636 (N_2636,N_2260,N_2227);
nand U2637 (N_2637,N_2123,N_2435);
or U2638 (N_2638,N_2206,N_2381);
xnor U2639 (N_2639,N_2216,N_2134);
nand U2640 (N_2640,N_2279,N_2104);
xor U2641 (N_2641,N_2015,N_2335);
nand U2642 (N_2642,N_2086,N_2461);
xnor U2643 (N_2643,N_2385,N_2114);
and U2644 (N_2644,N_2151,N_2272);
nor U2645 (N_2645,N_2016,N_2078);
and U2646 (N_2646,N_2257,N_2405);
nor U2647 (N_2647,N_2290,N_2180);
nand U2648 (N_2648,N_2217,N_2055);
nor U2649 (N_2649,N_2497,N_2338);
nand U2650 (N_2650,N_2012,N_2434);
or U2651 (N_2651,N_2415,N_2464);
nand U2652 (N_2652,N_2352,N_2140);
or U2653 (N_2653,N_2188,N_2286);
or U2654 (N_2654,N_2388,N_2267);
xnor U2655 (N_2655,N_2236,N_2273);
or U2656 (N_2656,N_2269,N_2182);
or U2657 (N_2657,N_2463,N_2333);
and U2658 (N_2658,N_2194,N_2132);
or U2659 (N_2659,N_2209,N_2324);
and U2660 (N_2660,N_2230,N_2028);
and U2661 (N_2661,N_2204,N_2212);
and U2662 (N_2662,N_2029,N_2298);
xnor U2663 (N_2663,N_2453,N_2283);
nor U2664 (N_2664,N_2479,N_2074);
nor U2665 (N_2665,N_2328,N_2057);
nand U2666 (N_2666,N_2458,N_2327);
nand U2667 (N_2667,N_2404,N_2161);
nand U2668 (N_2668,N_2034,N_2480);
xor U2669 (N_2669,N_2127,N_2443);
xor U2670 (N_2670,N_2421,N_2318);
nand U2671 (N_2671,N_2296,N_2124);
or U2672 (N_2672,N_2275,N_2021);
nor U2673 (N_2673,N_2013,N_2315);
or U2674 (N_2674,N_2357,N_2276);
nand U2675 (N_2675,N_2113,N_2103);
nor U2676 (N_2676,N_2162,N_2210);
and U2677 (N_2677,N_2044,N_2374);
xnor U2678 (N_2678,N_2075,N_2067);
nand U2679 (N_2679,N_2136,N_2400);
xnor U2680 (N_2680,N_2138,N_2436);
nand U2681 (N_2681,N_2049,N_2292);
nand U2682 (N_2682,N_2109,N_2207);
nand U2683 (N_2683,N_2033,N_2361);
and U2684 (N_2684,N_2189,N_2106);
and U2685 (N_2685,N_2199,N_2237);
xnor U2686 (N_2686,N_2406,N_2228);
or U2687 (N_2687,N_2091,N_2235);
nand U2688 (N_2688,N_2412,N_2031);
nand U2689 (N_2689,N_2268,N_2087);
and U2690 (N_2690,N_2499,N_2169);
nor U2691 (N_2691,N_2263,N_2484);
nor U2692 (N_2692,N_2079,N_2121);
nor U2693 (N_2693,N_2178,N_2387);
xor U2694 (N_2694,N_2226,N_2478);
nand U2695 (N_2695,N_2133,N_2307);
xnor U2696 (N_2696,N_2059,N_2234);
and U2697 (N_2697,N_2190,N_2168);
nand U2698 (N_2698,N_2158,N_2354);
and U2699 (N_2699,N_2383,N_2187);
and U2700 (N_2700,N_2118,N_2242);
and U2701 (N_2701,N_2363,N_2495);
nor U2702 (N_2702,N_2170,N_2160);
xor U2703 (N_2703,N_2146,N_2122);
xor U2704 (N_2704,N_2191,N_2485);
xnor U2705 (N_2705,N_2312,N_2281);
and U2706 (N_2706,N_2473,N_2293);
or U2707 (N_2707,N_2177,N_2183);
and U2708 (N_2708,N_2452,N_2099);
nor U2709 (N_2709,N_2266,N_2198);
nor U2710 (N_2710,N_2063,N_2270);
and U2711 (N_2711,N_2265,N_2256);
nand U2712 (N_2712,N_2030,N_2070);
or U2713 (N_2713,N_2111,N_2277);
xnor U2714 (N_2714,N_2317,N_2302);
nor U2715 (N_2715,N_2065,N_2371);
or U2716 (N_2716,N_2440,N_2095);
and U2717 (N_2717,N_2240,N_2316);
xnor U2718 (N_2718,N_2446,N_2246);
and U2719 (N_2719,N_2331,N_2433);
or U2720 (N_2720,N_2203,N_2444);
xor U2721 (N_2721,N_2253,N_2326);
xor U2722 (N_2722,N_2047,N_2454);
nor U2723 (N_2723,N_2062,N_2058);
and U2724 (N_2724,N_2120,N_2040);
or U2725 (N_2725,N_2382,N_2186);
or U2726 (N_2726,N_2460,N_2128);
nor U2727 (N_2727,N_2426,N_2085);
and U2728 (N_2728,N_2438,N_2077);
xnor U2729 (N_2729,N_2084,N_2043);
xnor U2730 (N_2730,N_2045,N_2193);
or U2731 (N_2731,N_2223,N_2414);
and U2732 (N_2732,N_2427,N_2014);
nor U2733 (N_2733,N_2305,N_2377);
and U2734 (N_2734,N_2080,N_2493);
nor U2735 (N_2735,N_2419,N_2167);
nor U2736 (N_2736,N_2375,N_2372);
nor U2737 (N_2737,N_2174,N_2483);
or U2738 (N_2738,N_2476,N_2214);
or U2739 (N_2739,N_2042,N_2413);
nand U2740 (N_2740,N_2470,N_2258);
nand U2741 (N_2741,N_2396,N_2247);
nand U2742 (N_2742,N_2200,N_2428);
xor U2743 (N_2743,N_2125,N_2051);
or U2744 (N_2744,N_2010,N_2262);
nand U2745 (N_2745,N_2251,N_2245);
nor U2746 (N_2746,N_2343,N_2297);
and U2747 (N_2747,N_2445,N_2370);
or U2748 (N_2748,N_2073,N_2477);
nand U2749 (N_2749,N_2137,N_2126);
and U2750 (N_2750,N_2411,N_2336);
xnor U2751 (N_2751,N_2135,N_2386);
xnor U2752 (N_2752,N_2257,N_2054);
and U2753 (N_2753,N_2228,N_2096);
and U2754 (N_2754,N_2100,N_2485);
and U2755 (N_2755,N_2284,N_2156);
nor U2756 (N_2756,N_2370,N_2425);
xor U2757 (N_2757,N_2200,N_2236);
nand U2758 (N_2758,N_2333,N_2239);
nand U2759 (N_2759,N_2060,N_2196);
and U2760 (N_2760,N_2431,N_2466);
nor U2761 (N_2761,N_2277,N_2050);
nand U2762 (N_2762,N_2338,N_2170);
nor U2763 (N_2763,N_2415,N_2495);
nand U2764 (N_2764,N_2148,N_2392);
xor U2765 (N_2765,N_2140,N_2439);
xnor U2766 (N_2766,N_2339,N_2478);
xnor U2767 (N_2767,N_2256,N_2309);
and U2768 (N_2768,N_2489,N_2396);
nand U2769 (N_2769,N_2048,N_2024);
nand U2770 (N_2770,N_2099,N_2389);
nor U2771 (N_2771,N_2359,N_2044);
nor U2772 (N_2772,N_2318,N_2429);
or U2773 (N_2773,N_2463,N_2487);
or U2774 (N_2774,N_2253,N_2246);
and U2775 (N_2775,N_2010,N_2232);
and U2776 (N_2776,N_2429,N_2194);
nor U2777 (N_2777,N_2014,N_2258);
nor U2778 (N_2778,N_2138,N_2333);
and U2779 (N_2779,N_2492,N_2308);
and U2780 (N_2780,N_2481,N_2182);
nand U2781 (N_2781,N_2229,N_2160);
or U2782 (N_2782,N_2321,N_2398);
or U2783 (N_2783,N_2217,N_2443);
and U2784 (N_2784,N_2200,N_2414);
nand U2785 (N_2785,N_2297,N_2352);
or U2786 (N_2786,N_2096,N_2350);
and U2787 (N_2787,N_2441,N_2209);
or U2788 (N_2788,N_2348,N_2231);
and U2789 (N_2789,N_2437,N_2388);
or U2790 (N_2790,N_2433,N_2241);
nor U2791 (N_2791,N_2423,N_2156);
nand U2792 (N_2792,N_2359,N_2488);
nand U2793 (N_2793,N_2116,N_2093);
nor U2794 (N_2794,N_2105,N_2311);
nand U2795 (N_2795,N_2044,N_2445);
or U2796 (N_2796,N_2148,N_2227);
nor U2797 (N_2797,N_2391,N_2293);
and U2798 (N_2798,N_2324,N_2364);
nor U2799 (N_2799,N_2062,N_2066);
nor U2800 (N_2800,N_2216,N_2202);
or U2801 (N_2801,N_2414,N_2285);
xor U2802 (N_2802,N_2203,N_2358);
or U2803 (N_2803,N_2318,N_2333);
xnor U2804 (N_2804,N_2467,N_2472);
nand U2805 (N_2805,N_2215,N_2233);
and U2806 (N_2806,N_2328,N_2218);
nand U2807 (N_2807,N_2148,N_2330);
or U2808 (N_2808,N_2086,N_2282);
or U2809 (N_2809,N_2262,N_2207);
or U2810 (N_2810,N_2216,N_2080);
or U2811 (N_2811,N_2182,N_2409);
nand U2812 (N_2812,N_2077,N_2313);
and U2813 (N_2813,N_2237,N_2314);
nor U2814 (N_2814,N_2213,N_2289);
and U2815 (N_2815,N_2163,N_2317);
nand U2816 (N_2816,N_2321,N_2360);
nor U2817 (N_2817,N_2467,N_2421);
nand U2818 (N_2818,N_2464,N_2109);
nand U2819 (N_2819,N_2088,N_2367);
xnor U2820 (N_2820,N_2391,N_2495);
nand U2821 (N_2821,N_2298,N_2433);
xor U2822 (N_2822,N_2376,N_2331);
nor U2823 (N_2823,N_2350,N_2421);
nand U2824 (N_2824,N_2400,N_2175);
xnor U2825 (N_2825,N_2239,N_2413);
nand U2826 (N_2826,N_2146,N_2227);
xnor U2827 (N_2827,N_2199,N_2064);
and U2828 (N_2828,N_2299,N_2137);
and U2829 (N_2829,N_2471,N_2259);
or U2830 (N_2830,N_2497,N_2133);
xor U2831 (N_2831,N_2462,N_2319);
xor U2832 (N_2832,N_2025,N_2295);
nor U2833 (N_2833,N_2140,N_2052);
nor U2834 (N_2834,N_2167,N_2431);
nand U2835 (N_2835,N_2462,N_2424);
and U2836 (N_2836,N_2032,N_2213);
and U2837 (N_2837,N_2149,N_2313);
and U2838 (N_2838,N_2346,N_2352);
nand U2839 (N_2839,N_2005,N_2002);
xor U2840 (N_2840,N_2383,N_2023);
xor U2841 (N_2841,N_2003,N_2428);
xnor U2842 (N_2842,N_2185,N_2191);
and U2843 (N_2843,N_2140,N_2274);
or U2844 (N_2844,N_2143,N_2437);
and U2845 (N_2845,N_2317,N_2344);
nor U2846 (N_2846,N_2365,N_2083);
nand U2847 (N_2847,N_2319,N_2498);
or U2848 (N_2848,N_2477,N_2052);
nand U2849 (N_2849,N_2193,N_2267);
or U2850 (N_2850,N_2315,N_2355);
xnor U2851 (N_2851,N_2038,N_2050);
or U2852 (N_2852,N_2164,N_2097);
and U2853 (N_2853,N_2193,N_2014);
nand U2854 (N_2854,N_2128,N_2206);
xor U2855 (N_2855,N_2433,N_2200);
or U2856 (N_2856,N_2264,N_2236);
xnor U2857 (N_2857,N_2258,N_2493);
nor U2858 (N_2858,N_2188,N_2104);
and U2859 (N_2859,N_2035,N_2376);
xnor U2860 (N_2860,N_2076,N_2446);
or U2861 (N_2861,N_2388,N_2222);
xor U2862 (N_2862,N_2264,N_2344);
nand U2863 (N_2863,N_2382,N_2184);
nand U2864 (N_2864,N_2117,N_2094);
nand U2865 (N_2865,N_2035,N_2493);
nand U2866 (N_2866,N_2278,N_2453);
and U2867 (N_2867,N_2300,N_2158);
nor U2868 (N_2868,N_2185,N_2498);
xor U2869 (N_2869,N_2168,N_2053);
xor U2870 (N_2870,N_2276,N_2154);
xor U2871 (N_2871,N_2179,N_2085);
nand U2872 (N_2872,N_2461,N_2323);
or U2873 (N_2873,N_2470,N_2181);
or U2874 (N_2874,N_2457,N_2367);
xor U2875 (N_2875,N_2262,N_2069);
nand U2876 (N_2876,N_2463,N_2438);
and U2877 (N_2877,N_2302,N_2061);
nor U2878 (N_2878,N_2354,N_2465);
nand U2879 (N_2879,N_2390,N_2102);
nand U2880 (N_2880,N_2188,N_2402);
or U2881 (N_2881,N_2025,N_2410);
nor U2882 (N_2882,N_2159,N_2033);
xnor U2883 (N_2883,N_2176,N_2020);
nand U2884 (N_2884,N_2192,N_2372);
nand U2885 (N_2885,N_2123,N_2491);
nand U2886 (N_2886,N_2225,N_2275);
nand U2887 (N_2887,N_2074,N_2336);
or U2888 (N_2888,N_2386,N_2249);
or U2889 (N_2889,N_2190,N_2031);
and U2890 (N_2890,N_2484,N_2050);
and U2891 (N_2891,N_2276,N_2403);
and U2892 (N_2892,N_2302,N_2205);
or U2893 (N_2893,N_2435,N_2491);
and U2894 (N_2894,N_2082,N_2441);
xor U2895 (N_2895,N_2041,N_2127);
xor U2896 (N_2896,N_2169,N_2124);
or U2897 (N_2897,N_2437,N_2255);
or U2898 (N_2898,N_2373,N_2478);
nor U2899 (N_2899,N_2272,N_2487);
and U2900 (N_2900,N_2428,N_2024);
and U2901 (N_2901,N_2120,N_2235);
nor U2902 (N_2902,N_2252,N_2271);
and U2903 (N_2903,N_2300,N_2123);
and U2904 (N_2904,N_2353,N_2319);
xor U2905 (N_2905,N_2018,N_2192);
xnor U2906 (N_2906,N_2038,N_2185);
xor U2907 (N_2907,N_2364,N_2382);
nor U2908 (N_2908,N_2412,N_2049);
and U2909 (N_2909,N_2365,N_2416);
or U2910 (N_2910,N_2008,N_2479);
and U2911 (N_2911,N_2156,N_2415);
xnor U2912 (N_2912,N_2269,N_2413);
nand U2913 (N_2913,N_2434,N_2288);
nand U2914 (N_2914,N_2333,N_2116);
or U2915 (N_2915,N_2341,N_2423);
and U2916 (N_2916,N_2021,N_2180);
and U2917 (N_2917,N_2278,N_2368);
and U2918 (N_2918,N_2021,N_2273);
and U2919 (N_2919,N_2018,N_2305);
or U2920 (N_2920,N_2037,N_2404);
or U2921 (N_2921,N_2302,N_2110);
nor U2922 (N_2922,N_2253,N_2232);
nor U2923 (N_2923,N_2191,N_2467);
or U2924 (N_2924,N_2216,N_2289);
nand U2925 (N_2925,N_2148,N_2237);
nor U2926 (N_2926,N_2092,N_2397);
nor U2927 (N_2927,N_2228,N_2229);
nand U2928 (N_2928,N_2026,N_2467);
xor U2929 (N_2929,N_2061,N_2091);
and U2930 (N_2930,N_2177,N_2096);
or U2931 (N_2931,N_2307,N_2054);
and U2932 (N_2932,N_2495,N_2113);
nand U2933 (N_2933,N_2462,N_2097);
xnor U2934 (N_2934,N_2312,N_2167);
and U2935 (N_2935,N_2188,N_2187);
or U2936 (N_2936,N_2353,N_2130);
xnor U2937 (N_2937,N_2374,N_2029);
nand U2938 (N_2938,N_2395,N_2367);
and U2939 (N_2939,N_2285,N_2119);
nand U2940 (N_2940,N_2459,N_2460);
nand U2941 (N_2941,N_2107,N_2464);
xnor U2942 (N_2942,N_2067,N_2487);
xor U2943 (N_2943,N_2490,N_2380);
and U2944 (N_2944,N_2328,N_2022);
xor U2945 (N_2945,N_2278,N_2129);
xor U2946 (N_2946,N_2106,N_2070);
nand U2947 (N_2947,N_2024,N_2430);
nor U2948 (N_2948,N_2239,N_2326);
nor U2949 (N_2949,N_2042,N_2010);
nor U2950 (N_2950,N_2053,N_2145);
nand U2951 (N_2951,N_2364,N_2077);
xor U2952 (N_2952,N_2179,N_2200);
nor U2953 (N_2953,N_2021,N_2190);
nor U2954 (N_2954,N_2313,N_2014);
nand U2955 (N_2955,N_2219,N_2264);
nor U2956 (N_2956,N_2069,N_2395);
nand U2957 (N_2957,N_2222,N_2356);
or U2958 (N_2958,N_2391,N_2336);
xor U2959 (N_2959,N_2229,N_2344);
or U2960 (N_2960,N_2274,N_2036);
nand U2961 (N_2961,N_2294,N_2422);
xor U2962 (N_2962,N_2408,N_2422);
nor U2963 (N_2963,N_2281,N_2085);
and U2964 (N_2964,N_2354,N_2433);
or U2965 (N_2965,N_2215,N_2371);
or U2966 (N_2966,N_2279,N_2184);
xnor U2967 (N_2967,N_2157,N_2049);
nand U2968 (N_2968,N_2365,N_2097);
xor U2969 (N_2969,N_2492,N_2305);
or U2970 (N_2970,N_2263,N_2367);
nor U2971 (N_2971,N_2224,N_2338);
or U2972 (N_2972,N_2073,N_2284);
or U2973 (N_2973,N_2456,N_2262);
or U2974 (N_2974,N_2123,N_2306);
and U2975 (N_2975,N_2249,N_2058);
nor U2976 (N_2976,N_2245,N_2101);
nand U2977 (N_2977,N_2349,N_2381);
nand U2978 (N_2978,N_2179,N_2036);
or U2979 (N_2979,N_2157,N_2016);
nand U2980 (N_2980,N_2290,N_2441);
nor U2981 (N_2981,N_2213,N_2209);
xor U2982 (N_2982,N_2210,N_2130);
nand U2983 (N_2983,N_2060,N_2207);
nand U2984 (N_2984,N_2394,N_2266);
nor U2985 (N_2985,N_2141,N_2390);
or U2986 (N_2986,N_2426,N_2081);
nand U2987 (N_2987,N_2000,N_2390);
nor U2988 (N_2988,N_2313,N_2406);
nand U2989 (N_2989,N_2028,N_2253);
nand U2990 (N_2990,N_2076,N_2303);
nand U2991 (N_2991,N_2478,N_2082);
or U2992 (N_2992,N_2099,N_2026);
xnor U2993 (N_2993,N_2000,N_2101);
nor U2994 (N_2994,N_2420,N_2494);
or U2995 (N_2995,N_2127,N_2067);
nand U2996 (N_2996,N_2455,N_2179);
nand U2997 (N_2997,N_2205,N_2420);
xor U2998 (N_2998,N_2006,N_2146);
xnor U2999 (N_2999,N_2142,N_2169);
or UO_0 (O_0,N_2705,N_2981);
or UO_1 (O_1,N_2666,N_2583);
xor UO_2 (O_2,N_2584,N_2727);
nor UO_3 (O_3,N_2910,N_2648);
nand UO_4 (O_4,N_2655,N_2553);
nor UO_5 (O_5,N_2808,N_2963);
nor UO_6 (O_6,N_2735,N_2762);
xor UO_7 (O_7,N_2987,N_2608);
nand UO_8 (O_8,N_2976,N_2721);
or UO_9 (O_9,N_2603,N_2884);
xnor UO_10 (O_10,N_2786,N_2813);
nor UO_11 (O_11,N_2975,N_2552);
nor UO_12 (O_12,N_2689,N_2869);
or UO_13 (O_13,N_2513,N_2969);
or UO_14 (O_14,N_2596,N_2709);
nor UO_15 (O_15,N_2960,N_2802);
or UO_16 (O_16,N_2807,N_2548);
or UO_17 (O_17,N_2887,N_2746);
nor UO_18 (O_18,N_2863,N_2895);
nor UO_19 (O_19,N_2586,N_2780);
and UO_20 (O_20,N_2794,N_2631);
xnor UO_21 (O_21,N_2977,N_2741);
nor UO_22 (O_22,N_2628,N_2751);
and UO_23 (O_23,N_2955,N_2509);
nor UO_24 (O_24,N_2771,N_2728);
nor UO_25 (O_25,N_2602,N_2950);
nand UO_26 (O_26,N_2770,N_2874);
nor UO_27 (O_27,N_2616,N_2962);
xnor UO_28 (O_28,N_2953,N_2979);
or UO_29 (O_29,N_2902,N_2997);
xor UO_30 (O_30,N_2637,N_2672);
xor UO_31 (O_31,N_2778,N_2833);
nand UO_32 (O_32,N_2738,N_2879);
nor UO_33 (O_33,N_2761,N_2825);
nor UO_34 (O_34,N_2551,N_2888);
or UO_35 (O_35,N_2543,N_2734);
xnor UO_36 (O_36,N_2704,N_2768);
nor UO_37 (O_37,N_2624,N_2809);
xnor UO_38 (O_38,N_2795,N_2886);
nand UO_39 (O_39,N_2922,N_2806);
nor UO_40 (O_40,N_2816,N_2772);
xor UO_41 (O_41,N_2933,N_2562);
nand UO_42 (O_42,N_2827,N_2555);
or UO_43 (O_43,N_2822,N_2831);
or UO_44 (O_44,N_2604,N_2645);
or UO_45 (O_45,N_2821,N_2711);
nand UO_46 (O_46,N_2701,N_2924);
xnor UO_47 (O_47,N_2859,N_2622);
nor UO_48 (O_48,N_2832,N_2841);
or UO_49 (O_49,N_2714,N_2935);
or UO_50 (O_50,N_2578,N_2871);
or UO_51 (O_51,N_2872,N_2718);
nor UO_52 (O_52,N_2911,N_2812);
xor UO_53 (O_53,N_2629,N_2725);
or UO_54 (O_54,N_2860,N_2691);
nor UO_55 (O_55,N_2627,N_2759);
xor UO_56 (O_56,N_2653,N_2625);
nand UO_57 (O_57,N_2995,N_2908);
and UO_58 (O_58,N_2528,N_2820);
and UO_59 (O_59,N_2817,N_2563);
nand UO_60 (O_60,N_2729,N_2906);
or UO_61 (O_61,N_2654,N_2531);
and UO_62 (O_62,N_2894,N_2830);
or UO_63 (O_63,N_2643,N_2524);
or UO_64 (O_64,N_2564,N_2712);
nand UO_65 (O_65,N_2865,N_2743);
nand UO_66 (O_66,N_2905,N_2919);
nand UO_67 (O_67,N_2686,N_2515);
nor UO_68 (O_68,N_2992,N_2796);
xnor UO_69 (O_69,N_2588,N_2681);
or UO_70 (O_70,N_2517,N_2749);
nor UO_71 (O_71,N_2511,N_2967);
xnor UO_72 (O_72,N_2527,N_2736);
or UO_73 (O_73,N_2670,N_2610);
and UO_74 (O_74,N_2909,N_2638);
or UO_75 (O_75,N_2695,N_2939);
xnor UO_76 (O_76,N_2642,N_2788);
or UO_77 (O_77,N_2811,N_2618);
nor UO_78 (O_78,N_2640,N_2641);
and UO_79 (O_79,N_2623,N_2556);
nand UO_80 (O_80,N_2614,N_2918);
or UO_81 (O_81,N_2932,N_2684);
and UO_82 (O_82,N_2839,N_2876);
xor UO_83 (O_83,N_2696,N_2844);
or UO_84 (O_84,N_2934,N_2514);
nand UO_85 (O_85,N_2769,N_2713);
nand UO_86 (O_86,N_2507,N_2706);
and UO_87 (O_87,N_2582,N_2739);
or UO_88 (O_88,N_2723,N_2561);
nor UO_89 (O_89,N_2698,N_2677);
and UO_90 (O_90,N_2708,N_2612);
xor UO_91 (O_91,N_2877,N_2752);
and UO_92 (O_92,N_2605,N_2609);
and UO_93 (O_93,N_2800,N_2592);
or UO_94 (O_94,N_2500,N_2998);
xnor UO_95 (O_95,N_2882,N_2569);
nand UO_96 (O_96,N_2855,N_2972);
nor UO_97 (O_97,N_2798,N_2927);
nor UO_98 (O_98,N_2545,N_2547);
or UO_99 (O_99,N_2898,N_2510);
xnor UO_100 (O_100,N_2529,N_2667);
nor UO_101 (O_101,N_2946,N_2595);
nor UO_102 (O_102,N_2707,N_2502);
or UO_103 (O_103,N_2923,N_2740);
or UO_104 (O_104,N_2779,N_2617);
nand UO_105 (O_105,N_2546,N_2916);
nand UO_106 (O_106,N_2693,N_2699);
xnor UO_107 (O_107,N_2757,N_2947);
nand UO_108 (O_108,N_2733,N_2819);
nand UO_109 (O_109,N_2890,N_2636);
xor UO_110 (O_110,N_2716,N_2959);
xnor UO_111 (O_111,N_2626,N_2787);
or UO_112 (O_112,N_2845,N_2828);
nor UO_113 (O_113,N_2717,N_2781);
or UO_114 (O_114,N_2744,N_2942);
or UO_115 (O_115,N_2760,N_2957);
xnor UO_116 (O_116,N_2773,N_2889);
nor UO_117 (O_117,N_2917,N_2538);
and UO_118 (O_118,N_2748,N_2753);
nor UO_119 (O_119,N_2742,N_2526);
nand UO_120 (O_120,N_2615,N_2697);
nand UO_121 (O_121,N_2837,N_2797);
or UO_122 (O_122,N_2776,N_2580);
xor UO_123 (O_123,N_2758,N_2914);
and UO_124 (O_124,N_2680,N_2973);
xnor UO_125 (O_125,N_2941,N_2767);
xnor UO_126 (O_126,N_2523,N_2980);
xnor UO_127 (O_127,N_2926,N_2650);
xnor UO_128 (O_128,N_2991,N_2519);
and UO_129 (O_129,N_2936,N_2850);
and UO_130 (O_130,N_2810,N_2613);
xor UO_131 (O_131,N_2694,N_2745);
and UO_132 (O_132,N_2647,N_2961);
and UO_133 (O_133,N_2804,N_2594);
xnor UO_134 (O_134,N_2883,N_2585);
nand UO_135 (O_135,N_2662,N_2852);
or UO_136 (O_136,N_2750,N_2956);
nand UO_137 (O_137,N_2783,N_2838);
and UO_138 (O_138,N_2799,N_2568);
nor UO_139 (O_139,N_2685,N_2814);
xnor UO_140 (O_140,N_2921,N_2574);
or UO_141 (O_141,N_2669,N_2756);
nand UO_142 (O_142,N_2836,N_2668);
xnor UO_143 (O_143,N_2826,N_2703);
or UO_144 (O_144,N_2673,N_2943);
nor UO_145 (O_145,N_2525,N_2840);
or UO_146 (O_146,N_2864,N_2520);
xor UO_147 (O_147,N_2853,N_2978);
or UO_148 (O_148,N_2620,N_2782);
xor UO_149 (O_149,N_2516,N_2829);
xor UO_150 (O_150,N_2854,N_2530);
xor UO_151 (O_151,N_2937,N_2966);
or UO_152 (O_152,N_2931,N_2903);
and UO_153 (O_153,N_2897,N_2983);
and UO_154 (O_154,N_2536,N_2710);
nand UO_155 (O_155,N_2777,N_2533);
or UO_156 (O_156,N_2875,N_2644);
nand UO_157 (O_157,N_2593,N_2896);
or UO_158 (O_158,N_2732,N_2868);
nor UO_159 (O_159,N_2632,N_2607);
nand UO_160 (O_160,N_2971,N_2823);
and UO_161 (O_161,N_2534,N_2521);
or UO_162 (O_162,N_2503,N_2576);
nor UO_163 (O_163,N_2656,N_2660);
and UO_164 (O_164,N_2652,N_2571);
nand UO_165 (O_165,N_2873,N_2848);
xor UO_166 (O_166,N_2968,N_2784);
xnor UO_167 (O_167,N_2982,N_2881);
nor UO_168 (O_168,N_2692,N_2554);
nand UO_169 (O_169,N_2633,N_2646);
nor UO_170 (O_170,N_2630,N_2891);
xnor UO_171 (O_171,N_2557,N_2549);
nand UO_172 (O_172,N_2687,N_2948);
nand UO_173 (O_173,N_2700,N_2904);
and UO_174 (O_174,N_2920,N_2913);
xor UO_175 (O_175,N_2754,N_2715);
and UO_176 (O_176,N_2591,N_2512);
and UO_177 (O_177,N_2532,N_2683);
nand UO_178 (O_178,N_2843,N_2985);
and UO_179 (O_179,N_2504,N_2658);
nand UO_180 (O_180,N_2567,N_2550);
nand UO_181 (O_181,N_2522,N_2835);
and UO_182 (O_182,N_2559,N_2834);
nor UO_183 (O_183,N_2880,N_2634);
xor UO_184 (O_184,N_2726,N_2506);
nor UO_185 (O_185,N_2993,N_2952);
xnor UO_186 (O_186,N_2970,N_2930);
nor UO_187 (O_187,N_2951,N_2907);
nor UO_188 (O_188,N_2679,N_2566);
xnor UO_189 (O_189,N_2665,N_2996);
nand UO_190 (O_190,N_2899,N_2621);
and UO_191 (O_191,N_2944,N_2535);
and UO_192 (O_192,N_2597,N_2893);
xor UO_193 (O_193,N_2581,N_2537);
nand UO_194 (O_194,N_2501,N_2573);
and UO_195 (O_195,N_2824,N_2540);
nor UO_196 (O_196,N_2682,N_2565);
xnor UO_197 (O_197,N_2851,N_2539);
xor UO_198 (O_198,N_2803,N_2846);
and UO_199 (O_199,N_2518,N_2579);
or UO_200 (O_200,N_2587,N_2929);
or UO_201 (O_201,N_2719,N_2671);
xor UO_202 (O_202,N_2702,N_2847);
and UO_203 (O_203,N_2600,N_2954);
nand UO_204 (O_204,N_2747,N_2805);
nor UO_205 (O_205,N_2558,N_2599);
xor UO_206 (O_206,N_2639,N_2663);
and UO_207 (O_207,N_2928,N_2590);
nor UO_208 (O_208,N_2755,N_2589);
xnor UO_209 (O_209,N_2878,N_2775);
and UO_210 (O_210,N_2945,N_2986);
nand UO_211 (O_211,N_2570,N_2988);
or UO_212 (O_212,N_2737,N_2676);
nand UO_213 (O_213,N_2764,N_2858);
and UO_214 (O_214,N_2999,N_2792);
xor UO_215 (O_215,N_2940,N_2601);
nor UO_216 (O_216,N_2958,N_2938);
and UO_217 (O_217,N_2842,N_2785);
nand UO_218 (O_218,N_2560,N_2611);
and UO_219 (O_219,N_2661,N_2870);
or UO_220 (O_220,N_2678,N_2790);
nor UO_221 (O_221,N_2577,N_2965);
nor UO_222 (O_222,N_2866,N_2818);
nand UO_223 (O_223,N_2815,N_2505);
xor UO_224 (O_224,N_2763,N_2664);
and UO_225 (O_225,N_2949,N_2659);
or UO_226 (O_226,N_2856,N_2724);
nor UO_227 (O_227,N_2849,N_2862);
and UO_228 (O_228,N_2789,N_2575);
xnor UO_229 (O_229,N_2635,N_2994);
or UO_230 (O_230,N_2974,N_2861);
nand UO_231 (O_231,N_2675,N_2619);
or UO_232 (O_232,N_2649,N_2572);
and UO_233 (O_233,N_2731,N_2722);
nor UO_234 (O_234,N_2984,N_2765);
xor UO_235 (O_235,N_2885,N_2542);
xor UO_236 (O_236,N_2793,N_2900);
xor UO_237 (O_237,N_2892,N_2674);
or UO_238 (O_238,N_2720,N_2801);
or UO_239 (O_239,N_2774,N_2867);
or UO_240 (O_240,N_2989,N_2791);
and UO_241 (O_241,N_2925,N_2901);
nand UO_242 (O_242,N_2657,N_2730);
or UO_243 (O_243,N_2857,N_2766);
or UO_244 (O_244,N_2544,N_2688);
xnor UO_245 (O_245,N_2508,N_2690);
xnor UO_246 (O_246,N_2606,N_2651);
nand UO_247 (O_247,N_2598,N_2990);
xor UO_248 (O_248,N_2964,N_2541);
and UO_249 (O_249,N_2915,N_2912);
nand UO_250 (O_250,N_2670,N_2913);
nand UO_251 (O_251,N_2906,N_2990);
and UO_252 (O_252,N_2565,N_2543);
nor UO_253 (O_253,N_2659,N_2952);
or UO_254 (O_254,N_2547,N_2867);
nand UO_255 (O_255,N_2622,N_2631);
xor UO_256 (O_256,N_2931,N_2550);
nor UO_257 (O_257,N_2871,N_2820);
and UO_258 (O_258,N_2663,N_2840);
nor UO_259 (O_259,N_2673,N_2997);
xnor UO_260 (O_260,N_2711,N_2674);
nand UO_261 (O_261,N_2610,N_2562);
nor UO_262 (O_262,N_2880,N_2763);
nand UO_263 (O_263,N_2946,N_2927);
nand UO_264 (O_264,N_2850,N_2750);
nand UO_265 (O_265,N_2838,N_2500);
nor UO_266 (O_266,N_2661,N_2968);
nand UO_267 (O_267,N_2821,N_2866);
nand UO_268 (O_268,N_2759,N_2711);
nand UO_269 (O_269,N_2761,N_2693);
or UO_270 (O_270,N_2518,N_2673);
or UO_271 (O_271,N_2769,N_2647);
nor UO_272 (O_272,N_2992,N_2587);
nor UO_273 (O_273,N_2577,N_2818);
nand UO_274 (O_274,N_2662,N_2578);
xnor UO_275 (O_275,N_2719,N_2689);
xor UO_276 (O_276,N_2837,N_2709);
xor UO_277 (O_277,N_2797,N_2938);
nand UO_278 (O_278,N_2885,N_2970);
xor UO_279 (O_279,N_2899,N_2750);
and UO_280 (O_280,N_2779,N_2516);
xor UO_281 (O_281,N_2608,N_2618);
nand UO_282 (O_282,N_2727,N_2814);
or UO_283 (O_283,N_2777,N_2645);
or UO_284 (O_284,N_2591,N_2520);
and UO_285 (O_285,N_2925,N_2777);
xnor UO_286 (O_286,N_2769,N_2960);
or UO_287 (O_287,N_2882,N_2818);
nand UO_288 (O_288,N_2624,N_2867);
nand UO_289 (O_289,N_2860,N_2598);
nand UO_290 (O_290,N_2627,N_2897);
nor UO_291 (O_291,N_2818,N_2974);
and UO_292 (O_292,N_2705,N_2885);
xnor UO_293 (O_293,N_2535,N_2662);
and UO_294 (O_294,N_2655,N_2880);
nor UO_295 (O_295,N_2725,N_2507);
or UO_296 (O_296,N_2847,N_2795);
xor UO_297 (O_297,N_2897,N_2755);
nand UO_298 (O_298,N_2779,N_2934);
xnor UO_299 (O_299,N_2964,N_2580);
and UO_300 (O_300,N_2903,N_2988);
nor UO_301 (O_301,N_2756,N_2726);
nor UO_302 (O_302,N_2998,N_2928);
or UO_303 (O_303,N_2646,N_2729);
nand UO_304 (O_304,N_2700,N_2655);
or UO_305 (O_305,N_2847,N_2584);
or UO_306 (O_306,N_2775,N_2536);
xnor UO_307 (O_307,N_2684,N_2825);
and UO_308 (O_308,N_2729,N_2551);
or UO_309 (O_309,N_2944,N_2811);
xor UO_310 (O_310,N_2990,N_2607);
or UO_311 (O_311,N_2907,N_2917);
xnor UO_312 (O_312,N_2512,N_2545);
and UO_313 (O_313,N_2757,N_2535);
xnor UO_314 (O_314,N_2995,N_2853);
nor UO_315 (O_315,N_2728,N_2703);
nor UO_316 (O_316,N_2858,N_2793);
or UO_317 (O_317,N_2550,N_2674);
nand UO_318 (O_318,N_2528,N_2828);
or UO_319 (O_319,N_2640,N_2730);
nor UO_320 (O_320,N_2935,N_2704);
nand UO_321 (O_321,N_2830,N_2596);
nor UO_322 (O_322,N_2544,N_2625);
nor UO_323 (O_323,N_2611,N_2757);
nand UO_324 (O_324,N_2757,N_2929);
and UO_325 (O_325,N_2670,N_2503);
and UO_326 (O_326,N_2906,N_2761);
or UO_327 (O_327,N_2857,N_2991);
xor UO_328 (O_328,N_2692,N_2544);
nor UO_329 (O_329,N_2569,N_2724);
or UO_330 (O_330,N_2532,N_2806);
and UO_331 (O_331,N_2956,N_2594);
and UO_332 (O_332,N_2876,N_2706);
nor UO_333 (O_333,N_2535,N_2858);
xor UO_334 (O_334,N_2805,N_2829);
and UO_335 (O_335,N_2936,N_2637);
and UO_336 (O_336,N_2832,N_2787);
or UO_337 (O_337,N_2952,N_2536);
and UO_338 (O_338,N_2875,N_2626);
nor UO_339 (O_339,N_2557,N_2885);
or UO_340 (O_340,N_2502,N_2633);
nand UO_341 (O_341,N_2865,N_2834);
and UO_342 (O_342,N_2637,N_2750);
nand UO_343 (O_343,N_2918,N_2754);
or UO_344 (O_344,N_2899,N_2580);
nand UO_345 (O_345,N_2841,N_2758);
nor UO_346 (O_346,N_2562,N_2957);
and UO_347 (O_347,N_2674,N_2846);
nor UO_348 (O_348,N_2764,N_2937);
nand UO_349 (O_349,N_2957,N_2644);
or UO_350 (O_350,N_2825,N_2549);
nand UO_351 (O_351,N_2797,N_2749);
or UO_352 (O_352,N_2759,N_2603);
xnor UO_353 (O_353,N_2636,N_2840);
or UO_354 (O_354,N_2518,N_2721);
xnor UO_355 (O_355,N_2952,N_2566);
xor UO_356 (O_356,N_2960,N_2983);
or UO_357 (O_357,N_2745,N_2866);
nand UO_358 (O_358,N_2637,N_2894);
xor UO_359 (O_359,N_2953,N_2880);
nor UO_360 (O_360,N_2902,N_2992);
nor UO_361 (O_361,N_2748,N_2889);
nor UO_362 (O_362,N_2585,N_2938);
nand UO_363 (O_363,N_2515,N_2565);
xor UO_364 (O_364,N_2613,N_2582);
xor UO_365 (O_365,N_2571,N_2656);
or UO_366 (O_366,N_2737,N_2516);
or UO_367 (O_367,N_2761,N_2674);
and UO_368 (O_368,N_2570,N_2744);
xor UO_369 (O_369,N_2962,N_2806);
and UO_370 (O_370,N_2580,N_2903);
nor UO_371 (O_371,N_2680,N_2516);
nand UO_372 (O_372,N_2956,N_2801);
and UO_373 (O_373,N_2780,N_2706);
xnor UO_374 (O_374,N_2624,N_2540);
xor UO_375 (O_375,N_2635,N_2822);
xnor UO_376 (O_376,N_2770,N_2541);
nand UO_377 (O_377,N_2925,N_2721);
nand UO_378 (O_378,N_2780,N_2583);
xnor UO_379 (O_379,N_2713,N_2549);
or UO_380 (O_380,N_2605,N_2582);
nor UO_381 (O_381,N_2580,N_2558);
or UO_382 (O_382,N_2795,N_2627);
and UO_383 (O_383,N_2530,N_2841);
nor UO_384 (O_384,N_2701,N_2929);
or UO_385 (O_385,N_2525,N_2867);
nor UO_386 (O_386,N_2529,N_2737);
nor UO_387 (O_387,N_2647,N_2774);
or UO_388 (O_388,N_2523,N_2993);
and UO_389 (O_389,N_2562,N_2885);
and UO_390 (O_390,N_2517,N_2874);
or UO_391 (O_391,N_2967,N_2811);
nor UO_392 (O_392,N_2689,N_2555);
xnor UO_393 (O_393,N_2608,N_2879);
nand UO_394 (O_394,N_2553,N_2722);
xor UO_395 (O_395,N_2752,N_2813);
xnor UO_396 (O_396,N_2943,N_2732);
nand UO_397 (O_397,N_2578,N_2845);
nor UO_398 (O_398,N_2888,N_2580);
or UO_399 (O_399,N_2883,N_2967);
xor UO_400 (O_400,N_2638,N_2954);
xor UO_401 (O_401,N_2523,N_2845);
nor UO_402 (O_402,N_2622,N_2512);
nor UO_403 (O_403,N_2777,N_2990);
nand UO_404 (O_404,N_2629,N_2581);
xor UO_405 (O_405,N_2511,N_2778);
xor UO_406 (O_406,N_2866,N_2738);
nor UO_407 (O_407,N_2613,N_2733);
or UO_408 (O_408,N_2628,N_2890);
or UO_409 (O_409,N_2995,N_2833);
or UO_410 (O_410,N_2520,N_2953);
and UO_411 (O_411,N_2707,N_2716);
and UO_412 (O_412,N_2704,N_2612);
nand UO_413 (O_413,N_2718,N_2611);
nand UO_414 (O_414,N_2748,N_2932);
and UO_415 (O_415,N_2547,N_2890);
nor UO_416 (O_416,N_2777,N_2854);
xor UO_417 (O_417,N_2521,N_2677);
or UO_418 (O_418,N_2944,N_2759);
xnor UO_419 (O_419,N_2664,N_2658);
and UO_420 (O_420,N_2894,N_2962);
nand UO_421 (O_421,N_2645,N_2565);
and UO_422 (O_422,N_2513,N_2855);
or UO_423 (O_423,N_2880,N_2931);
and UO_424 (O_424,N_2987,N_2743);
and UO_425 (O_425,N_2752,N_2843);
or UO_426 (O_426,N_2519,N_2956);
and UO_427 (O_427,N_2880,N_2526);
nand UO_428 (O_428,N_2624,N_2791);
and UO_429 (O_429,N_2605,N_2514);
xnor UO_430 (O_430,N_2676,N_2534);
nor UO_431 (O_431,N_2847,N_2849);
or UO_432 (O_432,N_2551,N_2950);
nand UO_433 (O_433,N_2708,N_2536);
xor UO_434 (O_434,N_2796,N_2625);
nor UO_435 (O_435,N_2516,N_2983);
or UO_436 (O_436,N_2577,N_2547);
nor UO_437 (O_437,N_2526,N_2653);
and UO_438 (O_438,N_2780,N_2713);
or UO_439 (O_439,N_2632,N_2924);
nand UO_440 (O_440,N_2835,N_2788);
or UO_441 (O_441,N_2863,N_2847);
nand UO_442 (O_442,N_2924,N_2568);
xnor UO_443 (O_443,N_2957,N_2968);
nor UO_444 (O_444,N_2775,N_2962);
nand UO_445 (O_445,N_2710,N_2685);
or UO_446 (O_446,N_2540,N_2864);
nor UO_447 (O_447,N_2605,N_2781);
or UO_448 (O_448,N_2680,N_2989);
nor UO_449 (O_449,N_2874,N_2712);
nand UO_450 (O_450,N_2504,N_2805);
or UO_451 (O_451,N_2682,N_2535);
or UO_452 (O_452,N_2695,N_2716);
or UO_453 (O_453,N_2849,N_2767);
xnor UO_454 (O_454,N_2904,N_2687);
or UO_455 (O_455,N_2629,N_2935);
or UO_456 (O_456,N_2820,N_2558);
xnor UO_457 (O_457,N_2848,N_2962);
or UO_458 (O_458,N_2645,N_2561);
and UO_459 (O_459,N_2698,N_2993);
and UO_460 (O_460,N_2761,N_2855);
nor UO_461 (O_461,N_2888,N_2843);
nor UO_462 (O_462,N_2851,N_2615);
nor UO_463 (O_463,N_2640,N_2731);
xnor UO_464 (O_464,N_2618,N_2836);
nand UO_465 (O_465,N_2647,N_2506);
and UO_466 (O_466,N_2614,N_2909);
xnor UO_467 (O_467,N_2722,N_2889);
nor UO_468 (O_468,N_2545,N_2852);
nor UO_469 (O_469,N_2951,N_2686);
xor UO_470 (O_470,N_2772,N_2836);
or UO_471 (O_471,N_2677,N_2533);
nand UO_472 (O_472,N_2969,N_2635);
nand UO_473 (O_473,N_2857,N_2909);
nor UO_474 (O_474,N_2542,N_2627);
and UO_475 (O_475,N_2568,N_2888);
nand UO_476 (O_476,N_2859,N_2676);
and UO_477 (O_477,N_2866,N_2877);
and UO_478 (O_478,N_2990,N_2921);
or UO_479 (O_479,N_2792,N_2570);
and UO_480 (O_480,N_2692,N_2872);
and UO_481 (O_481,N_2828,N_2692);
and UO_482 (O_482,N_2813,N_2651);
xnor UO_483 (O_483,N_2764,N_2932);
nand UO_484 (O_484,N_2742,N_2554);
nand UO_485 (O_485,N_2524,N_2585);
or UO_486 (O_486,N_2611,N_2836);
and UO_487 (O_487,N_2967,N_2973);
nor UO_488 (O_488,N_2895,N_2711);
nor UO_489 (O_489,N_2558,N_2989);
and UO_490 (O_490,N_2517,N_2935);
xnor UO_491 (O_491,N_2641,N_2764);
nor UO_492 (O_492,N_2933,N_2811);
nor UO_493 (O_493,N_2959,N_2792);
xor UO_494 (O_494,N_2882,N_2711);
xor UO_495 (O_495,N_2879,N_2776);
nand UO_496 (O_496,N_2644,N_2586);
nand UO_497 (O_497,N_2908,N_2674);
xnor UO_498 (O_498,N_2553,N_2502);
nand UO_499 (O_499,N_2997,N_2852);
endmodule