module basic_1500_15000_2000_5_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_490,In_30);
nor U1 (N_1,In_1223,In_1242);
and U2 (N_2,In_1082,In_950);
nor U3 (N_3,In_40,In_1463);
nand U4 (N_4,In_85,In_68);
and U5 (N_5,In_293,In_1419);
nand U6 (N_6,In_735,In_836);
nand U7 (N_7,In_731,In_325);
nand U8 (N_8,In_182,In_23);
and U9 (N_9,In_673,In_1368);
or U10 (N_10,In_807,In_1052);
and U11 (N_11,In_782,In_1323);
or U12 (N_12,In_1011,In_801);
nand U13 (N_13,In_174,In_1343);
and U14 (N_14,In_18,In_1133);
nand U15 (N_15,In_592,In_1248);
and U16 (N_16,In_932,In_1355);
xor U17 (N_17,In_1428,In_1267);
nand U18 (N_18,In_944,In_9);
nand U19 (N_19,In_196,In_1288);
and U20 (N_20,In_522,In_415);
and U21 (N_21,In_388,In_759);
or U22 (N_22,In_63,In_506);
and U23 (N_23,In_997,In_686);
and U24 (N_24,In_840,In_202);
and U25 (N_25,In_267,In_960);
nor U26 (N_26,In_626,In_1426);
or U27 (N_27,In_965,In_1353);
nor U28 (N_28,In_134,In_546);
and U29 (N_29,In_1348,In_283);
xor U30 (N_30,In_1453,In_1497);
nor U31 (N_31,In_1452,In_683);
nand U32 (N_32,In_426,In_273);
nor U33 (N_33,In_321,In_631);
nand U34 (N_34,In_778,In_480);
and U35 (N_35,In_757,In_1277);
or U36 (N_36,In_353,In_1179);
nand U37 (N_37,In_1423,In_269);
or U38 (N_38,In_622,In_1016);
and U39 (N_39,In_292,In_27);
and U40 (N_40,In_959,In_514);
or U41 (N_41,In_372,In_691);
or U42 (N_42,In_1313,In_1163);
and U43 (N_43,In_240,In_1151);
nand U44 (N_44,In_1382,In_334);
nand U45 (N_45,In_1220,In_1410);
nand U46 (N_46,In_632,In_983);
nand U47 (N_47,In_1192,In_1101);
nor U48 (N_48,In_98,In_880);
nor U49 (N_49,In_695,In_105);
nand U50 (N_50,In_1122,In_311);
or U51 (N_51,In_1448,In_1204);
and U52 (N_52,In_164,In_1456);
or U53 (N_53,In_1252,In_796);
nand U54 (N_54,In_1404,In_760);
nor U55 (N_55,In_655,In_275);
nor U56 (N_56,In_579,In_837);
nand U57 (N_57,In_200,In_727);
nand U58 (N_58,In_1218,In_1467);
nand U59 (N_59,In_1222,In_570);
nor U60 (N_60,In_847,In_675);
or U61 (N_61,In_1216,In_447);
and U62 (N_62,In_995,In_423);
or U63 (N_63,In_1339,In_729);
and U64 (N_64,In_1200,In_912);
and U65 (N_65,In_985,In_52);
or U66 (N_66,In_1257,In_254);
or U67 (N_67,In_694,In_397);
nand U68 (N_68,In_216,In_1137);
and U69 (N_69,In_584,In_750);
nand U70 (N_70,In_463,In_1292);
nand U71 (N_71,In_690,In_1077);
nor U72 (N_72,In_1271,In_804);
nor U73 (N_73,In_156,In_820);
nand U74 (N_74,In_851,In_1202);
and U75 (N_75,In_1173,In_1031);
nand U76 (N_76,In_488,In_1033);
nand U77 (N_77,In_385,In_43);
nand U78 (N_78,In_1268,In_331);
nand U79 (N_79,In_365,In_1004);
and U80 (N_80,In_1334,In_633);
or U81 (N_81,In_509,In_671);
nor U82 (N_82,In_253,In_556);
and U83 (N_83,In_888,In_79);
nor U84 (N_84,In_747,In_351);
or U85 (N_85,In_13,In_1363);
or U86 (N_86,In_223,In_1241);
nand U87 (N_87,In_537,In_493);
nor U88 (N_88,In_14,In_176);
and U89 (N_89,In_19,In_641);
nor U90 (N_90,In_974,In_1296);
and U91 (N_91,In_1272,In_420);
nand U92 (N_92,In_827,In_235);
or U93 (N_93,In_868,In_1225);
or U94 (N_94,In_154,In_472);
nand U95 (N_95,In_896,In_724);
or U96 (N_96,In_878,In_162);
nor U97 (N_97,In_986,In_175);
nand U98 (N_98,In_1000,In_924);
or U99 (N_99,In_966,In_354);
or U100 (N_100,In_1067,In_891);
nand U101 (N_101,In_1307,In_1025);
nand U102 (N_102,In_203,In_369);
or U103 (N_103,In_71,In_566);
and U104 (N_104,In_455,In_258);
or U105 (N_105,In_1215,In_39);
nor U106 (N_106,In_76,In_94);
nand U107 (N_107,In_722,In_437);
or U108 (N_108,In_91,In_305);
nor U109 (N_109,In_511,In_232);
or U110 (N_110,In_497,In_850);
nand U111 (N_111,In_728,In_679);
nand U112 (N_112,In_245,In_1312);
or U113 (N_113,In_1152,In_120);
and U114 (N_114,In_194,In_770);
and U115 (N_115,In_875,In_557);
and U116 (N_116,In_1354,In_865);
and U117 (N_117,In_356,In_835);
nor U118 (N_118,In_1008,In_1273);
and U119 (N_119,In_863,In_650);
or U120 (N_120,In_862,In_771);
or U121 (N_121,In_719,In_1325);
and U122 (N_122,In_743,In_853);
nor U123 (N_123,In_20,In_589);
nand U124 (N_124,In_26,In_541);
nor U125 (N_125,In_1338,In_1182);
nand U126 (N_126,In_512,In_1145);
and U127 (N_127,In_1364,In_1141);
nor U128 (N_128,In_1086,In_439);
nor U129 (N_129,In_227,In_1177);
or U130 (N_130,In_1037,In_768);
nor U131 (N_131,In_1347,In_1205);
and U132 (N_132,In_1349,In_1367);
or U133 (N_133,In_859,In_1214);
nand U134 (N_134,In_125,In_1116);
nand U135 (N_135,In_158,In_143);
nand U136 (N_136,In_921,In_848);
and U137 (N_137,In_1121,In_296);
nor U138 (N_138,In_1442,In_487);
and U139 (N_139,In_1158,In_975);
and U140 (N_140,In_976,In_559);
or U141 (N_141,In_565,In_773);
nor U142 (N_142,In_979,In_1262);
nand U143 (N_143,In_1130,In_380);
nor U144 (N_144,In_842,In_212);
nor U145 (N_145,In_234,In_1118);
nand U146 (N_146,In_282,In_1405);
or U147 (N_147,In_1079,In_247);
and U148 (N_148,In_568,In_454);
or U149 (N_149,In_1491,In_1386);
and U150 (N_150,In_360,In_218);
nand U151 (N_151,In_871,In_133);
nand U152 (N_152,In_1139,In_621);
nor U153 (N_153,In_821,In_1026);
nand U154 (N_154,In_1134,In_1490);
nor U155 (N_155,In_1302,In_1253);
or U156 (N_156,In_682,In_0);
nand U157 (N_157,In_517,In_484);
xor U158 (N_158,In_295,In_357);
and U159 (N_159,In_744,In_1281);
or U160 (N_160,In_1260,In_337);
or U161 (N_161,In_117,In_1068);
and U162 (N_162,In_1468,In_1);
and U163 (N_163,In_665,In_1258);
or U164 (N_164,In_841,In_935);
nand U165 (N_165,In_536,In_1366);
or U166 (N_166,In_1032,In_65);
and U167 (N_167,In_1473,In_1084);
or U168 (N_168,In_126,In_301);
and U169 (N_169,In_1399,In_149);
and U170 (N_170,In_704,In_1434);
or U171 (N_171,In_1249,In_160);
nand U172 (N_172,In_988,In_712);
or U173 (N_173,In_338,In_1286);
and U174 (N_174,In_1411,In_663);
nand U175 (N_175,In_115,In_816);
nand U176 (N_176,In_786,In_696);
or U177 (N_177,In_806,In_41);
nand U178 (N_178,In_51,In_1425);
and U179 (N_179,In_1328,In_659);
and U180 (N_180,In_1290,In_425);
nand U181 (N_181,In_407,In_900);
nor U182 (N_182,In_70,In_424);
or U183 (N_183,In_767,In_687);
and U184 (N_184,In_329,In_623);
nand U185 (N_185,In_1065,In_739);
nor U186 (N_186,In_297,In_142);
nand U187 (N_187,In_774,In_1400);
and U188 (N_188,In_37,In_737);
nand U189 (N_189,In_917,In_317);
or U190 (N_190,In_595,In_714);
nand U191 (N_191,In_102,In_401);
or U192 (N_192,In_1007,In_766);
nor U193 (N_193,In_812,In_1309);
or U194 (N_194,In_281,In_1345);
and U195 (N_195,In_503,In_1104);
nor U196 (N_196,In_95,In_499);
and U197 (N_197,In_1298,In_779);
nor U198 (N_198,In_649,In_1458);
or U199 (N_199,In_1185,In_1306);
or U200 (N_200,In_756,In_593);
xor U201 (N_201,In_89,In_127);
nand U202 (N_202,In_1264,In_1237);
nand U203 (N_203,In_1254,In_1380);
and U204 (N_204,In_874,In_918);
or U205 (N_205,In_408,In_998);
nand U206 (N_206,In_1318,In_1107);
or U207 (N_207,In_1293,In_942);
nand U208 (N_208,In_251,In_962);
nor U209 (N_209,In_1112,In_1147);
or U210 (N_210,In_231,In_318);
or U211 (N_211,In_617,In_518);
or U212 (N_212,In_416,In_280);
and U213 (N_213,In_1002,In_1224);
nor U214 (N_214,In_1213,In_791);
or U215 (N_215,In_452,In_1431);
or U216 (N_216,In_1009,In_1369);
nand U217 (N_217,In_936,In_899);
or U218 (N_218,In_1395,In_1209);
and U219 (N_219,In_530,In_1211);
nand U220 (N_220,In_605,In_99);
and U221 (N_221,In_754,In_226);
and U222 (N_222,In_474,In_1146);
nor U223 (N_223,In_954,In_738);
or U224 (N_224,In_560,In_562);
or U225 (N_225,In_945,In_558);
and U226 (N_226,In_758,In_846);
and U227 (N_227,In_1094,In_1229);
nor U228 (N_228,In_179,In_97);
or U229 (N_229,In_1384,In_1403);
nand U230 (N_230,In_478,In_1184);
and U231 (N_231,In_475,In_186);
nand U232 (N_232,In_916,In_931);
and U233 (N_233,In_140,In_1427);
nand U234 (N_234,In_968,In_1437);
or U235 (N_235,In_101,In_438);
or U236 (N_236,In_667,In_1350);
nor U237 (N_237,In_528,In_531);
or U238 (N_238,In_930,In_1370);
nand U239 (N_239,In_1378,In_630);
and U240 (N_240,In_1415,In_1451);
nor U241 (N_241,In_765,In_845);
and U242 (N_242,In_529,In_831);
and U243 (N_243,In_1362,In_306);
or U244 (N_244,In_926,In_440);
nand U245 (N_245,In_1206,In_892);
and U246 (N_246,In_343,In_172);
or U247 (N_247,In_393,In_996);
nor U248 (N_248,In_249,In_469);
and U249 (N_249,In_272,In_199);
nor U250 (N_250,In_1232,In_898);
nand U251 (N_251,In_165,In_795);
and U252 (N_252,In_973,In_1465);
and U253 (N_253,In_31,In_1441);
and U254 (N_254,In_138,In_550);
nand U255 (N_255,In_1059,In_443);
nand U256 (N_256,In_711,In_384);
xor U257 (N_257,In_64,In_681);
or U258 (N_258,In_316,In_590);
and U259 (N_259,In_48,In_1233);
nand U260 (N_260,In_1476,In_1398);
nor U261 (N_261,In_951,In_603);
nor U262 (N_262,In_1110,In_628);
and U263 (N_263,In_1055,In_1183);
nor U264 (N_264,In_1157,In_1475);
nor U265 (N_265,In_312,In_920);
nor U266 (N_266,In_1289,In_1351);
or U267 (N_267,In_349,In_1436);
and U268 (N_268,In_905,In_168);
nor U269 (N_269,In_1221,In_77);
nor U270 (N_270,In_647,In_145);
nor U271 (N_271,In_533,In_1484);
nor U272 (N_272,In_585,In_150);
or U273 (N_273,In_243,In_672);
nor U274 (N_274,In_370,In_1247);
nand U275 (N_275,In_109,In_1054);
nor U276 (N_276,In_67,In_587);
nand U277 (N_277,In_225,In_341);
nand U278 (N_278,In_940,In_328);
or U279 (N_279,In_725,In_800);
and U280 (N_280,In_1064,In_1250);
nor U281 (N_281,In_525,In_1056);
nand U282 (N_282,In_978,In_594);
nand U283 (N_283,In_471,In_575);
and U284 (N_284,In_1044,In_551);
and U285 (N_285,In_1303,In_886);
nand U286 (N_286,In_468,In_326);
or U287 (N_287,In_394,In_1015);
nand U288 (N_288,In_265,In_404);
and U289 (N_289,In_923,In_433);
nor U290 (N_290,In_830,In_347);
nand U291 (N_291,In_524,In_1352);
or U292 (N_292,In_1418,In_1461);
or U293 (N_293,In_428,In_664);
or U294 (N_294,In_709,In_609);
nand U295 (N_295,In_1159,In_10);
or U296 (N_296,In_1308,In_266);
nand U297 (N_297,In_364,In_646);
or U298 (N_298,In_1043,In_1492);
xor U299 (N_299,In_289,In_763);
nand U300 (N_300,In_308,In_780);
nor U301 (N_301,In_1375,In_1049);
or U302 (N_302,In_173,In_1329);
nand U303 (N_303,In_654,In_144);
xnor U304 (N_304,In_335,In_399);
and U305 (N_305,In_799,In_832);
and U306 (N_306,In_611,In_470);
or U307 (N_307,In_1337,In_718);
nand U308 (N_308,In_599,In_1024);
or U309 (N_309,In_1317,In_824);
and U310 (N_310,In_939,In_166);
nand U311 (N_311,In_462,In_66);
and U312 (N_312,In_262,In_178);
and U313 (N_313,In_17,In_1193);
or U314 (N_314,In_359,In_54);
and U315 (N_315,In_1278,In_1063);
and U316 (N_316,In_432,In_1344);
and U317 (N_317,In_1361,In_1447);
or U318 (N_318,In_1488,In_1171);
nor U319 (N_319,In_139,In_124);
nor U320 (N_320,In_1228,In_502);
or U321 (N_321,In_598,In_467);
nor U322 (N_322,In_1156,In_706);
and U323 (N_323,In_35,In_481);
nor U324 (N_324,In_1150,In_1439);
and U325 (N_325,In_540,In_882);
xnor U326 (N_326,In_1335,In_999);
nand U327 (N_327,In_57,In_1078);
nand U328 (N_328,In_1172,In_860);
nor U329 (N_329,In_844,In_319);
and U330 (N_330,In_58,In_1495);
and U331 (N_331,In_277,In_521);
and U332 (N_332,In_406,In_928);
nor U333 (N_333,In_793,In_376);
nor U334 (N_334,In_181,In_1489);
nand U335 (N_335,In_1165,In_368);
nand U336 (N_336,In_1036,In_702);
and U337 (N_337,In_1301,In_1187);
nor U338 (N_338,In_442,In_866);
and U339 (N_339,In_285,In_1305);
or U340 (N_340,In_1095,In_224);
or U341 (N_341,In_644,In_1217);
nor U342 (N_342,In_606,In_87);
and U343 (N_343,In_1357,In_822);
nand U344 (N_344,In_934,In_1322);
and U345 (N_345,In_543,In_828);
nor U346 (N_346,In_1459,In_1455);
nor U347 (N_347,In_86,In_350);
or U348 (N_348,In_870,In_62);
nand U349 (N_349,In_121,In_1097);
nor U350 (N_350,In_532,In_829);
and U351 (N_351,In_259,In_390);
and U352 (N_352,In_1346,In_1385);
nand U353 (N_353,In_1259,In_453);
nor U354 (N_354,In_229,In_1048);
and U355 (N_355,In_38,In_688);
nor U356 (N_356,In_313,In_815);
nand U357 (N_357,In_257,In_192);
nand U358 (N_358,In_1450,In_16);
nor U359 (N_359,In_147,In_1050);
nand U360 (N_360,In_608,In_941);
nand U361 (N_361,In_436,In_491);
nand U362 (N_362,In_96,In_651);
and U363 (N_363,In_668,In_1119);
or U364 (N_364,In_1219,In_1304);
or U365 (N_365,In_1397,In_1180);
or U366 (N_366,In_114,In_855);
or U367 (N_367,In_1239,In_264);
nand U368 (N_368,In_465,In_1319);
or U369 (N_369,In_578,In_872);
and U370 (N_370,In_392,In_1422);
or U371 (N_371,In_82,In_1127);
or U372 (N_372,In_1432,In_580);
and U373 (N_373,In_358,In_1314);
and U374 (N_374,In_250,In_1409);
or U375 (N_375,In_1336,In_242);
nand U376 (N_376,In_412,In_1108);
and U377 (N_377,In_698,In_520);
nand U378 (N_378,In_573,In_858);
xor U379 (N_379,In_304,In_685);
and U380 (N_380,In_783,In_661);
and U381 (N_381,In_680,In_207);
nor U382 (N_382,In_586,In_1199);
or U383 (N_383,In_300,In_116);
or U384 (N_384,In_1285,In_534);
or U385 (N_385,In_776,In_802);
nand U386 (N_386,In_220,In_222);
or U387 (N_387,In_1098,In_1356);
and U388 (N_388,In_1117,In_464);
nor U389 (N_389,In_1481,In_527);
nor U390 (N_390,In_980,In_122);
nand U391 (N_391,In_716,In_602);
and U392 (N_392,In_897,In_1402);
nor U393 (N_393,In_656,In_1438);
and U394 (N_394,In_34,In_1131);
nand U395 (N_395,In_1300,In_1496);
or U396 (N_396,In_1072,In_1129);
nand U397 (N_397,In_340,In_790);
nand U398 (N_398,In_1391,In_613);
or U399 (N_399,In_244,In_153);
and U400 (N_400,In_119,In_291);
nand U401 (N_401,In_1212,In_604);
nand U402 (N_402,In_635,In_547);
and U403 (N_403,In_1284,In_276);
and U404 (N_404,In_601,In_553);
nor U405 (N_405,In_1373,In_8);
or U406 (N_406,In_476,In_1462);
and U407 (N_407,In_526,In_1155);
nor U408 (N_408,In_169,In_163);
nand U409 (N_409,In_213,In_1060);
nand U410 (N_410,In_405,In_204);
and U411 (N_411,In_552,In_1266);
nor U412 (N_412,In_810,In_1166);
nor U413 (N_413,In_761,In_303);
nor U414 (N_414,In_943,In_290);
or U415 (N_415,In_1482,In_382);
nand U416 (N_416,In_938,In_4);
nor U417 (N_417,In_1164,In_237);
or U418 (N_418,In_640,In_1454);
and U419 (N_419,In_344,In_577);
nor U420 (N_420,In_210,In_879);
nand U421 (N_421,In_130,In_323);
nand U422 (N_422,In_838,In_185);
nand U423 (N_423,In_549,In_217);
or U424 (N_424,In_72,In_429);
nand U425 (N_425,In_215,In_1170);
and U426 (N_426,In_715,In_496);
nand U427 (N_427,In_1105,In_903);
and U428 (N_428,In_1408,In_61);
and U429 (N_429,In_755,In_890);
nand U430 (N_430,In_787,In_877);
or U431 (N_431,In_1128,In_523);
nand U432 (N_432,In_189,In_1058);
or U433 (N_433,In_1406,In_519);
nor U434 (N_434,In_1485,In_255);
xnor U435 (N_435,In_327,In_624);
nand U436 (N_436,In_981,In_572);
and U437 (N_437,In_118,In_792);
nand U438 (N_438,In_699,In_769);
nand U439 (N_439,In_451,In_1330);
nor U440 (N_440,In_925,In_1256);
nand U441 (N_441,In_483,In_538);
or U442 (N_442,In_505,In_648);
nor U443 (N_443,In_1041,In_515);
nand U444 (N_444,In_1401,In_516);
or U445 (N_445,In_69,In_1445);
nand U446 (N_446,In_542,In_148);
and U447 (N_447,In_1080,In_809);
or U448 (N_448,In_772,In_336);
nor U449 (N_449,In_1191,In_80);
and U450 (N_450,In_339,In_1103);
nand U451 (N_451,In_332,In_1160);
or U452 (N_452,In_535,In_298);
and U453 (N_453,In_1074,In_1381);
nand U454 (N_454,In_383,In_177);
nand U455 (N_455,In_74,In_381);
nor U456 (N_456,In_1424,In_893);
nor U457 (N_457,In_342,In_1143);
and U458 (N_458,In_1006,In_135);
nor U459 (N_459,In_1234,In_248);
nand U460 (N_460,In_44,In_1295);
nor U461 (N_461,In_710,In_46);
or U462 (N_462,In_908,In_1360);
nand U463 (N_463,In_957,In_700);
nor U464 (N_464,In_982,In_561);
or U465 (N_465,In_431,In_287);
nand U466 (N_466,In_1001,In_1483);
nand U467 (N_467,In_1061,In_637);
and U468 (N_468,In_449,In_324);
nand U469 (N_469,In_47,In_992);
nand U470 (N_470,In_410,In_1062);
nor U471 (N_471,In_884,In_1169);
and U472 (N_472,In_201,In_1342);
nor U473 (N_473,In_466,In_843);
nor U474 (N_474,In_901,In_129);
or U475 (N_475,In_1198,In_485);
nand U476 (N_476,In_946,In_387);
or U477 (N_477,In_73,In_1310);
nand U478 (N_478,In_371,In_322);
nor U479 (N_479,In_373,In_674);
nor U480 (N_480,In_346,In_867);
nand U481 (N_481,In_1263,In_84);
nand U482 (N_482,In_544,In_949);
or U483 (N_483,In_583,In_1022);
nor U484 (N_484,In_817,In_914);
nor U485 (N_485,In_1331,In_798);
nor U486 (N_486,In_379,In_1194);
or U487 (N_487,In_403,In_110);
nand U488 (N_488,In_784,In_1126);
or U489 (N_489,In_927,In_555);
nor U490 (N_490,In_660,In_857);
nor U491 (N_491,In_619,In_803);
nor U492 (N_492,In_1478,In_876);
nand U493 (N_493,In_278,In_1243);
and U494 (N_494,In_161,In_849);
nand U495 (N_495,In_473,In_818);
nand U496 (N_496,In_1090,In_1013);
or U497 (N_497,In_1175,In_1388);
or U498 (N_498,In_211,In_751);
or U499 (N_499,In_963,In_132);
nor U500 (N_500,In_1035,In_922);
or U501 (N_501,In_1039,In_887);
and U502 (N_502,In_740,In_208);
nand U503 (N_503,In_345,In_839);
and U504 (N_504,In_987,In_78);
nand U505 (N_505,In_788,In_352);
or U506 (N_506,In_852,In_1390);
or U507 (N_507,In_693,In_1324);
and U508 (N_508,In_1085,In_1430);
nor U509 (N_509,In_1045,In_1413);
xor U510 (N_510,In_55,In_11);
nand U511 (N_511,In_1412,In_494);
nand U512 (N_512,In_1471,In_1270);
nor U513 (N_513,In_910,In_563);
nand U514 (N_514,In_1246,In_666);
or U515 (N_515,In_638,In_703);
or U516 (N_516,In_1208,In_1275);
nand U517 (N_517,In_885,In_881);
nor U518 (N_518,In_781,In_219);
and U519 (N_519,In_302,In_1383);
nand U520 (N_520,In_1435,In_1023);
or U521 (N_521,In_597,In_707);
or U522 (N_522,In_658,In_22);
nor U523 (N_523,In_627,In_576);
or U524 (N_524,In_1235,In_1070);
nand U525 (N_525,In_1261,In_1030);
or U526 (N_526,In_1203,In_271);
or U527 (N_527,In_430,In_1178);
nand U528 (N_528,In_705,In_993);
nand U529 (N_529,In_1073,In_460);
nand U530 (N_530,In_955,In_171);
and U531 (N_531,In_826,In_1029);
or U532 (N_532,In_459,In_636);
nor U533 (N_533,In_819,In_1144);
or U534 (N_534,In_1066,In_1429);
nand U535 (N_535,In_261,In_1374);
or U536 (N_536,In_56,In_191);
nand U537 (N_537,In_1444,In_1326);
nand U538 (N_538,In_1042,In_823);
nand U539 (N_539,In_1280,In_600);
or U540 (N_540,In_320,In_1124);
nor U541 (N_541,In_1245,In_894);
or U542 (N_542,In_1474,In_1433);
nor U543 (N_543,In_746,In_104);
or U544 (N_544,In_1236,In_969);
nand U545 (N_545,In_571,In_1291);
nor U546 (N_546,In_582,In_1201);
and U547 (N_547,In_330,In_448);
or U548 (N_548,In_1393,In_1416);
nand U549 (N_549,In_1018,In_612);
nand U550 (N_550,In_833,In_88);
nor U551 (N_551,In_413,In_391);
nor U552 (N_552,In_742,In_642);
nor U553 (N_553,In_1188,In_260);
and U554 (N_554,In_947,In_596);
or U555 (N_555,In_591,In_1396);
or U556 (N_556,In_501,In_615);
nor U557 (N_557,In_984,In_241);
nand U558 (N_558,In_53,In_1320);
nand U559 (N_559,In_1389,In_209);
and U560 (N_560,In_75,In_1487);
nor U561 (N_561,In_1091,In_355);
nand U562 (N_562,In_1071,In_907);
nand U563 (N_563,In_1038,In_1443);
and U564 (N_564,In_479,In_721);
nand U565 (N_565,In_1075,In_662);
nor U566 (N_566,In_1499,In_717);
nand U567 (N_567,In_1333,In_315);
and U568 (N_568,In_395,In_36);
and U569 (N_569,In_155,In_3);
nand U570 (N_570,In_677,In_198);
and U571 (N_571,In_653,In_634);
nor U572 (N_572,In_333,In_1057);
nand U573 (N_573,In_569,In_1376);
nor U574 (N_574,In_764,In_137);
or U575 (N_575,In_1466,In_279);
or U576 (N_576,In_507,In_652);
and U577 (N_577,In_386,In_1120);
nand U578 (N_578,In_414,In_1123);
or U579 (N_579,In_435,In_971);
and U580 (N_580,In_131,In_854);
or U581 (N_581,In_1028,In_745);
and U582 (N_582,In_252,In_270);
nand U583 (N_583,In_856,In_1464);
nand U584 (N_584,In_1135,In_24);
and U585 (N_585,In_1255,In_1100);
nand U586 (N_586,In_588,In_1076);
nor U587 (N_587,In_1081,In_639);
and U588 (N_588,In_444,In_1283);
and U589 (N_589,In_294,In_1332);
or U590 (N_590,In_159,In_375);
nand U591 (N_591,In_141,In_477);
or U592 (N_592,In_1021,In_1012);
or U593 (N_593,In_1040,In_1162);
nor U594 (N_594,In_1274,In_492);
or U595 (N_595,In_1186,In_808);
or U596 (N_596,In_906,In_961);
nand U597 (N_597,In_1020,In_1027);
nor U598 (N_598,In_861,In_307);
nor U599 (N_599,In_21,In_1494);
nand U600 (N_600,In_362,In_136);
or U601 (N_601,In_146,In_299);
nand U602 (N_602,In_762,In_1321);
or U603 (N_603,In_1311,In_398);
and U604 (N_604,In_187,In_1210);
or U605 (N_605,In_1003,In_1371);
nor U606 (N_606,In_1113,In_441);
nand U607 (N_607,In_1457,In_1053);
and U608 (N_608,In_50,In_1341);
nand U609 (N_609,In_1014,In_789);
and U610 (N_610,In_1358,In_314);
and U611 (N_611,In_377,In_1238);
or U612 (N_612,In_929,In_1207);
nand U613 (N_613,In_450,In_230);
or U614 (N_614,In_1379,In_288);
or U615 (N_615,In_748,In_1477);
nand U616 (N_616,In_1472,In_1299);
nor U617 (N_617,In_1446,In_1498);
or U618 (N_618,In_1287,In_2);
nand U619 (N_619,In_554,In_958);
or U620 (N_620,In_60,In_389);
or U621 (N_621,In_692,In_1005);
nand U622 (N_622,In_869,In_274);
or U623 (N_623,In_236,In_797);
nand U624 (N_624,In_574,In_736);
and U625 (N_625,In_752,In_378);
or U626 (N_626,In_418,In_221);
and U627 (N_627,In_811,In_238);
and U628 (N_628,In_81,In_1449);
and U629 (N_629,In_409,In_708);
or U630 (N_630,In_1087,In_864);
nor U631 (N_631,In_1190,In_1460);
or U632 (N_632,In_1051,In_367);
nor U633 (N_633,In_15,In_1420);
nand U634 (N_634,In_915,In_190);
nor U635 (N_635,In_1265,In_684);
or U636 (N_636,In_1136,In_1114);
nand U637 (N_637,In_1377,In_1372);
nand U638 (N_638,In_49,In_1010);
nor U639 (N_639,In_785,In_794);
xnor U640 (N_640,In_539,In_948);
and U641 (N_641,In_1140,In_913);
and U642 (N_642,In_482,In_100);
or U643 (N_643,In_1365,In_180);
or U644 (N_644,In_239,In_994);
and U645 (N_645,In_618,In_732);
and U646 (N_646,In_657,In_1230);
nor U647 (N_647,In_669,In_7);
and U648 (N_648,In_193,In_902);
and U649 (N_649,In_548,In_1142);
and U650 (N_650,In_989,In_645);
and U651 (N_651,In_107,In_445);
nor U652 (N_652,In_964,In_268);
or U653 (N_653,In_151,In_904);
nor U654 (N_654,In_396,In_1102);
and U655 (N_655,In_676,In_411);
nand U656 (N_656,In_458,In_741);
or U657 (N_657,In_286,In_495);
and U658 (N_658,In_1387,In_805);
or U659 (N_659,In_59,In_1469);
nor U660 (N_660,In_1227,In_1231);
and U661 (N_661,In_400,In_1240);
or U662 (N_662,In_434,In_374);
and U663 (N_663,In_1106,In_128);
and U664 (N_664,In_545,In_967);
nand U665 (N_665,In_616,In_1176);
nand U666 (N_666,In_895,In_1089);
and U667 (N_667,In_1197,In_1294);
nor U668 (N_668,In_1181,In_103);
nand U669 (N_669,In_991,In_1046);
or U670 (N_670,In_446,In_106);
or U671 (N_671,In_489,In_233);
nor U672 (N_672,In_1092,In_1279);
nor U673 (N_673,In_184,In_123);
and U674 (N_674,In_629,In_1195);
or U675 (N_675,In_461,In_348);
nand U676 (N_676,In_1359,In_32);
and U677 (N_677,In_366,In_93);
nand U678 (N_678,In_422,In_1196);
xor U679 (N_679,In_112,In_883);
nor U680 (N_680,In_167,In_1407);
or U681 (N_681,In_152,In_697);
and U682 (N_682,In_183,In_825);
nand U683 (N_683,In_1392,In_361);
or U684 (N_684,In_720,In_1340);
nand U685 (N_685,In_1125,In_1019);
and U686 (N_686,In_733,In_911);
nor U687 (N_687,In_246,In_814);
nor U688 (N_688,In_689,In_1168);
nand U689 (N_689,In_1047,In_228);
or U690 (N_690,In_508,In_937);
nor U691 (N_691,In_1414,In_1226);
nor U692 (N_692,In_1315,In_363);
and U693 (N_693,In_1132,In_775);
and U694 (N_694,In_457,In_1282);
and U695 (N_695,In_1189,In_1421);
or U696 (N_696,In_1480,In_33);
or U697 (N_697,In_734,In_1486);
nor U698 (N_698,In_1440,In_972);
nor U699 (N_699,In_701,In_1111);
nor U700 (N_700,In_1327,In_723);
xor U701 (N_701,In_188,In_749);
or U702 (N_702,In_1115,In_206);
and U703 (N_703,In_1083,In_1093);
nand U704 (N_704,In_284,In_419);
and U705 (N_705,In_625,In_513);
nor U706 (N_706,In_753,In_970);
or U707 (N_707,In_953,In_1493);
or U708 (N_708,In_1244,In_111);
or U709 (N_709,In_933,In_813);
nand U710 (N_710,In_170,In_263);
nor U711 (N_711,In_643,In_607);
nand U712 (N_712,In_777,In_1034);
nand U713 (N_713,In_581,In_620);
nor U714 (N_714,In_498,In_417);
and U715 (N_715,In_421,In_730);
and U716 (N_716,In_28,In_1148);
nor U717 (N_717,In_205,In_1088);
and U718 (N_718,In_889,In_214);
nor U719 (N_719,In_486,In_1161);
and U720 (N_720,In_956,In_713);
nand U721 (N_721,In_12,In_427);
and U722 (N_722,In_157,In_1069);
nand U723 (N_723,In_1174,In_1479);
nand U724 (N_724,In_1417,In_309);
nand U725 (N_725,In_1109,In_310);
and U726 (N_726,In_1153,In_1251);
or U727 (N_727,In_90,In_1099);
nand U728 (N_728,In_510,In_610);
and U729 (N_729,In_1297,In_25);
nor U730 (N_730,In_990,In_402);
nor U731 (N_731,In_42,In_504);
or U732 (N_732,In_195,In_83);
nand U733 (N_733,In_6,In_197);
and U734 (N_734,In_1167,In_1276);
or U735 (N_735,In_500,In_726);
nor U736 (N_736,In_1394,In_256);
nor U737 (N_737,In_909,In_977);
nor U738 (N_738,In_873,In_92);
and U739 (N_739,In_29,In_567);
or U740 (N_740,In_113,In_834);
nor U741 (N_741,In_5,In_1017);
nor U742 (N_742,In_678,In_614);
and U743 (N_743,In_564,In_45);
or U744 (N_744,In_1316,In_670);
nor U745 (N_745,In_1096,In_1149);
and U746 (N_746,In_108,In_1138);
or U747 (N_747,In_1154,In_919);
or U748 (N_748,In_952,In_456);
or U749 (N_749,In_1470,In_1269);
or U750 (N_750,In_429,In_189);
nor U751 (N_751,In_958,In_10);
nor U752 (N_752,In_856,In_893);
nor U753 (N_753,In_240,In_100);
or U754 (N_754,In_915,In_623);
and U755 (N_755,In_1047,In_504);
nand U756 (N_756,In_1019,In_633);
and U757 (N_757,In_264,In_760);
nand U758 (N_758,In_140,In_1211);
and U759 (N_759,In_529,In_407);
and U760 (N_760,In_364,In_978);
or U761 (N_761,In_456,In_1065);
and U762 (N_762,In_543,In_339);
nor U763 (N_763,In_89,In_1044);
nand U764 (N_764,In_157,In_222);
and U765 (N_765,In_1478,In_479);
and U766 (N_766,In_1043,In_701);
nor U767 (N_767,In_361,In_202);
or U768 (N_768,In_964,In_760);
or U769 (N_769,In_554,In_728);
or U770 (N_770,In_1229,In_279);
or U771 (N_771,In_989,In_1076);
nor U772 (N_772,In_377,In_1195);
nor U773 (N_773,In_1231,In_1475);
nor U774 (N_774,In_844,In_597);
and U775 (N_775,In_694,In_1435);
nand U776 (N_776,In_505,In_1487);
nand U777 (N_777,In_874,In_200);
and U778 (N_778,In_667,In_80);
and U779 (N_779,In_1377,In_507);
nand U780 (N_780,In_387,In_699);
or U781 (N_781,In_1088,In_0);
nor U782 (N_782,In_337,In_1334);
and U783 (N_783,In_584,In_180);
nor U784 (N_784,In_507,In_95);
nor U785 (N_785,In_1365,In_409);
nor U786 (N_786,In_1254,In_1126);
nand U787 (N_787,In_246,In_441);
nand U788 (N_788,In_922,In_1033);
and U789 (N_789,In_972,In_9);
nor U790 (N_790,In_739,In_1362);
or U791 (N_791,In_1240,In_1341);
nand U792 (N_792,In_60,In_227);
xnor U793 (N_793,In_542,In_129);
nand U794 (N_794,In_315,In_372);
nand U795 (N_795,In_540,In_425);
nand U796 (N_796,In_898,In_239);
or U797 (N_797,In_473,In_720);
or U798 (N_798,In_559,In_1101);
or U799 (N_799,In_481,In_1325);
or U800 (N_800,In_437,In_99);
nor U801 (N_801,In_682,In_1067);
and U802 (N_802,In_620,In_153);
or U803 (N_803,In_1172,In_254);
nor U804 (N_804,In_509,In_1021);
nand U805 (N_805,In_1493,In_234);
nor U806 (N_806,In_1056,In_1408);
or U807 (N_807,In_98,In_482);
or U808 (N_808,In_503,In_38);
or U809 (N_809,In_902,In_306);
nor U810 (N_810,In_11,In_1434);
nor U811 (N_811,In_999,In_1053);
or U812 (N_812,In_275,In_305);
and U813 (N_813,In_827,In_615);
or U814 (N_814,In_873,In_424);
or U815 (N_815,In_1222,In_1085);
and U816 (N_816,In_1030,In_912);
nand U817 (N_817,In_91,In_1321);
or U818 (N_818,In_30,In_1149);
and U819 (N_819,In_1172,In_1208);
nand U820 (N_820,In_287,In_1169);
and U821 (N_821,In_631,In_90);
and U822 (N_822,In_1271,In_401);
or U823 (N_823,In_384,In_894);
nor U824 (N_824,In_1156,In_679);
nor U825 (N_825,In_482,In_67);
nand U826 (N_826,In_598,In_631);
nand U827 (N_827,In_225,In_504);
nor U828 (N_828,In_824,In_528);
nand U829 (N_829,In_120,In_1390);
and U830 (N_830,In_902,In_621);
and U831 (N_831,In_9,In_545);
or U832 (N_832,In_918,In_55);
nand U833 (N_833,In_997,In_394);
or U834 (N_834,In_1355,In_710);
nand U835 (N_835,In_97,In_380);
xor U836 (N_836,In_1106,In_44);
or U837 (N_837,In_1463,In_929);
and U838 (N_838,In_829,In_878);
or U839 (N_839,In_1053,In_1397);
or U840 (N_840,In_390,In_410);
or U841 (N_841,In_1442,In_362);
and U842 (N_842,In_557,In_1233);
nor U843 (N_843,In_1402,In_1016);
or U844 (N_844,In_972,In_306);
or U845 (N_845,In_805,In_526);
or U846 (N_846,In_1029,In_803);
and U847 (N_847,In_975,In_855);
and U848 (N_848,In_495,In_1407);
nor U849 (N_849,In_1375,In_853);
nor U850 (N_850,In_595,In_826);
or U851 (N_851,In_855,In_886);
or U852 (N_852,In_249,In_1398);
nor U853 (N_853,In_1108,In_1402);
and U854 (N_854,In_498,In_1271);
or U855 (N_855,In_213,In_411);
and U856 (N_856,In_705,In_938);
nand U857 (N_857,In_702,In_1251);
and U858 (N_858,In_101,In_244);
nor U859 (N_859,In_703,In_173);
or U860 (N_860,In_1422,In_13);
nor U861 (N_861,In_610,In_690);
or U862 (N_862,In_324,In_987);
and U863 (N_863,In_88,In_277);
nand U864 (N_864,In_507,In_831);
nor U865 (N_865,In_522,In_358);
nor U866 (N_866,In_1328,In_1068);
nand U867 (N_867,In_1180,In_574);
nand U868 (N_868,In_321,In_511);
and U869 (N_869,In_924,In_347);
nor U870 (N_870,In_633,In_1306);
nor U871 (N_871,In_848,In_795);
nand U872 (N_872,In_1237,In_905);
and U873 (N_873,In_939,In_1270);
nor U874 (N_874,In_796,In_808);
nor U875 (N_875,In_480,In_610);
and U876 (N_876,In_645,In_996);
xor U877 (N_877,In_1068,In_318);
nand U878 (N_878,In_335,In_1457);
or U879 (N_879,In_1030,In_1407);
or U880 (N_880,In_562,In_1256);
nand U881 (N_881,In_1074,In_799);
and U882 (N_882,In_904,In_167);
or U883 (N_883,In_101,In_416);
and U884 (N_884,In_1040,In_553);
nor U885 (N_885,In_1016,In_445);
and U886 (N_886,In_902,In_1104);
and U887 (N_887,In_324,In_547);
nor U888 (N_888,In_976,In_35);
and U889 (N_889,In_984,In_1420);
and U890 (N_890,In_993,In_437);
nor U891 (N_891,In_1195,In_1193);
nor U892 (N_892,In_1135,In_951);
and U893 (N_893,In_710,In_299);
or U894 (N_894,In_865,In_647);
nand U895 (N_895,In_347,In_844);
nand U896 (N_896,In_809,In_43);
nor U897 (N_897,In_1037,In_312);
or U898 (N_898,In_53,In_1174);
and U899 (N_899,In_1283,In_417);
and U900 (N_900,In_672,In_886);
and U901 (N_901,In_1241,In_1024);
nand U902 (N_902,In_596,In_37);
nor U903 (N_903,In_1225,In_1014);
or U904 (N_904,In_1196,In_1197);
or U905 (N_905,In_1255,In_1185);
or U906 (N_906,In_646,In_1143);
or U907 (N_907,In_41,In_1100);
and U908 (N_908,In_782,In_759);
and U909 (N_909,In_1041,In_855);
and U910 (N_910,In_1332,In_648);
nor U911 (N_911,In_1425,In_1020);
and U912 (N_912,In_565,In_1266);
and U913 (N_913,In_1047,In_754);
nor U914 (N_914,In_783,In_1476);
nand U915 (N_915,In_404,In_945);
and U916 (N_916,In_1407,In_579);
nor U917 (N_917,In_165,In_1273);
nor U918 (N_918,In_136,In_1345);
and U919 (N_919,In_1298,In_1306);
nor U920 (N_920,In_798,In_1110);
or U921 (N_921,In_740,In_197);
and U922 (N_922,In_761,In_1127);
nand U923 (N_923,In_778,In_902);
and U924 (N_924,In_951,In_335);
nor U925 (N_925,In_893,In_206);
nand U926 (N_926,In_261,In_493);
or U927 (N_927,In_891,In_831);
nand U928 (N_928,In_536,In_1094);
nor U929 (N_929,In_218,In_1177);
and U930 (N_930,In_699,In_6);
or U931 (N_931,In_406,In_1056);
nand U932 (N_932,In_1314,In_718);
nand U933 (N_933,In_1040,In_894);
nor U934 (N_934,In_659,In_661);
and U935 (N_935,In_1133,In_171);
nand U936 (N_936,In_165,In_812);
or U937 (N_937,In_226,In_238);
nor U938 (N_938,In_89,In_996);
and U939 (N_939,In_1164,In_54);
or U940 (N_940,In_691,In_1023);
nor U941 (N_941,In_728,In_1365);
nand U942 (N_942,In_575,In_140);
nand U943 (N_943,In_1469,In_459);
nand U944 (N_944,In_1375,In_560);
xor U945 (N_945,In_964,In_1075);
nor U946 (N_946,In_0,In_118);
or U947 (N_947,In_1101,In_1358);
and U948 (N_948,In_127,In_1418);
or U949 (N_949,In_1319,In_1350);
nor U950 (N_950,In_111,In_890);
or U951 (N_951,In_1404,In_1309);
nand U952 (N_952,In_625,In_1415);
nor U953 (N_953,In_147,In_473);
nor U954 (N_954,In_1125,In_1040);
nor U955 (N_955,In_1489,In_148);
or U956 (N_956,In_653,In_302);
or U957 (N_957,In_75,In_695);
nand U958 (N_958,In_1196,In_18);
nand U959 (N_959,In_594,In_617);
nand U960 (N_960,In_28,In_1296);
nor U961 (N_961,In_768,In_124);
nor U962 (N_962,In_672,In_41);
and U963 (N_963,In_763,In_1360);
nor U964 (N_964,In_122,In_1288);
and U965 (N_965,In_973,In_1087);
nor U966 (N_966,In_1141,In_91);
and U967 (N_967,In_767,In_1181);
or U968 (N_968,In_1297,In_715);
nand U969 (N_969,In_93,In_274);
and U970 (N_970,In_169,In_561);
nand U971 (N_971,In_1220,In_666);
nor U972 (N_972,In_664,In_932);
or U973 (N_973,In_201,In_507);
nand U974 (N_974,In_135,In_1082);
nand U975 (N_975,In_1169,In_122);
nor U976 (N_976,In_735,In_364);
nor U977 (N_977,In_102,In_812);
or U978 (N_978,In_1139,In_1169);
nand U979 (N_979,In_1422,In_718);
and U980 (N_980,In_1074,In_1462);
and U981 (N_981,In_596,In_263);
and U982 (N_982,In_530,In_949);
or U983 (N_983,In_903,In_1348);
nand U984 (N_984,In_158,In_145);
nor U985 (N_985,In_1312,In_1328);
and U986 (N_986,In_1221,In_871);
nand U987 (N_987,In_464,In_848);
nor U988 (N_988,In_753,In_101);
nor U989 (N_989,In_1207,In_873);
and U990 (N_990,In_1330,In_1087);
nand U991 (N_991,In_785,In_1270);
nand U992 (N_992,In_372,In_1115);
nand U993 (N_993,In_172,In_30);
or U994 (N_994,In_28,In_1425);
nand U995 (N_995,In_685,In_914);
and U996 (N_996,In_354,In_198);
and U997 (N_997,In_876,In_988);
and U998 (N_998,In_342,In_567);
nand U999 (N_999,In_246,In_1074);
nand U1000 (N_1000,In_608,In_67);
or U1001 (N_1001,In_443,In_1471);
or U1002 (N_1002,In_33,In_272);
nor U1003 (N_1003,In_1195,In_524);
and U1004 (N_1004,In_802,In_139);
nand U1005 (N_1005,In_1202,In_1081);
nand U1006 (N_1006,In_1459,In_744);
nand U1007 (N_1007,In_759,In_960);
nor U1008 (N_1008,In_87,In_803);
nand U1009 (N_1009,In_123,In_571);
and U1010 (N_1010,In_1234,In_266);
and U1011 (N_1011,In_1068,In_924);
or U1012 (N_1012,In_1058,In_1312);
nand U1013 (N_1013,In_1315,In_1142);
or U1014 (N_1014,In_118,In_579);
and U1015 (N_1015,In_1395,In_715);
and U1016 (N_1016,In_1498,In_961);
or U1017 (N_1017,In_985,In_735);
nand U1018 (N_1018,In_613,In_134);
nor U1019 (N_1019,In_785,In_134);
nor U1020 (N_1020,In_250,In_158);
or U1021 (N_1021,In_397,In_900);
and U1022 (N_1022,In_190,In_198);
and U1023 (N_1023,In_1099,In_1019);
nor U1024 (N_1024,In_677,In_161);
nor U1025 (N_1025,In_444,In_686);
or U1026 (N_1026,In_1188,In_1118);
and U1027 (N_1027,In_125,In_775);
nand U1028 (N_1028,In_792,In_71);
nand U1029 (N_1029,In_435,In_416);
nand U1030 (N_1030,In_1273,In_1389);
nor U1031 (N_1031,In_1096,In_31);
nor U1032 (N_1032,In_687,In_54);
or U1033 (N_1033,In_165,In_1290);
or U1034 (N_1034,In_830,In_1442);
nand U1035 (N_1035,In_934,In_1365);
nand U1036 (N_1036,In_561,In_623);
and U1037 (N_1037,In_343,In_437);
or U1038 (N_1038,In_995,In_1264);
or U1039 (N_1039,In_925,In_1076);
and U1040 (N_1040,In_1222,In_265);
and U1041 (N_1041,In_849,In_721);
nand U1042 (N_1042,In_572,In_1266);
and U1043 (N_1043,In_685,In_1053);
and U1044 (N_1044,In_1166,In_779);
or U1045 (N_1045,In_323,In_1458);
and U1046 (N_1046,In_1372,In_297);
and U1047 (N_1047,In_489,In_432);
nand U1048 (N_1048,In_531,In_507);
and U1049 (N_1049,In_855,In_118);
nor U1050 (N_1050,In_1428,In_57);
and U1051 (N_1051,In_928,In_1361);
and U1052 (N_1052,In_21,In_1386);
and U1053 (N_1053,In_1140,In_518);
and U1054 (N_1054,In_1237,In_98);
nand U1055 (N_1055,In_875,In_203);
nor U1056 (N_1056,In_444,In_14);
and U1057 (N_1057,In_733,In_406);
nand U1058 (N_1058,In_197,In_393);
or U1059 (N_1059,In_501,In_82);
or U1060 (N_1060,In_527,In_680);
and U1061 (N_1061,In_239,In_659);
nor U1062 (N_1062,In_161,In_900);
nand U1063 (N_1063,In_429,In_1006);
and U1064 (N_1064,In_188,In_1366);
or U1065 (N_1065,In_216,In_144);
or U1066 (N_1066,In_415,In_87);
or U1067 (N_1067,In_33,In_546);
nand U1068 (N_1068,In_355,In_1074);
and U1069 (N_1069,In_58,In_1273);
nand U1070 (N_1070,In_1449,In_377);
nand U1071 (N_1071,In_1260,In_202);
nor U1072 (N_1072,In_482,In_544);
and U1073 (N_1073,In_0,In_2);
or U1074 (N_1074,In_788,In_1173);
and U1075 (N_1075,In_1076,In_628);
nand U1076 (N_1076,In_218,In_800);
and U1077 (N_1077,In_335,In_535);
nand U1078 (N_1078,In_17,In_1090);
nor U1079 (N_1079,In_685,In_320);
nand U1080 (N_1080,In_583,In_1439);
and U1081 (N_1081,In_423,In_535);
nand U1082 (N_1082,In_1175,In_734);
or U1083 (N_1083,In_460,In_412);
nand U1084 (N_1084,In_481,In_1136);
nor U1085 (N_1085,In_1282,In_228);
and U1086 (N_1086,In_840,In_1377);
and U1087 (N_1087,In_289,In_1075);
nor U1088 (N_1088,In_1025,In_659);
and U1089 (N_1089,In_249,In_1205);
and U1090 (N_1090,In_1225,In_1047);
nor U1091 (N_1091,In_810,In_462);
nand U1092 (N_1092,In_308,In_651);
nand U1093 (N_1093,In_1236,In_1039);
and U1094 (N_1094,In_1397,In_897);
nand U1095 (N_1095,In_1340,In_833);
or U1096 (N_1096,In_171,In_433);
or U1097 (N_1097,In_375,In_161);
and U1098 (N_1098,In_1463,In_1184);
and U1099 (N_1099,In_664,In_763);
nor U1100 (N_1100,In_1339,In_1483);
nand U1101 (N_1101,In_348,In_899);
and U1102 (N_1102,In_1040,In_1216);
or U1103 (N_1103,In_916,In_53);
nand U1104 (N_1104,In_595,In_841);
nor U1105 (N_1105,In_1043,In_289);
nand U1106 (N_1106,In_624,In_143);
nor U1107 (N_1107,In_430,In_40);
nand U1108 (N_1108,In_863,In_1317);
or U1109 (N_1109,In_358,In_1071);
and U1110 (N_1110,In_500,In_465);
and U1111 (N_1111,In_1472,In_1131);
nand U1112 (N_1112,In_1096,In_343);
or U1113 (N_1113,In_833,In_1499);
nor U1114 (N_1114,In_450,In_525);
and U1115 (N_1115,In_1080,In_744);
nor U1116 (N_1116,In_663,In_1272);
nor U1117 (N_1117,In_70,In_109);
nand U1118 (N_1118,In_808,In_1356);
nor U1119 (N_1119,In_91,In_1330);
nor U1120 (N_1120,In_640,In_13);
and U1121 (N_1121,In_770,In_1412);
nand U1122 (N_1122,In_1295,In_1423);
nand U1123 (N_1123,In_1107,In_624);
xnor U1124 (N_1124,In_1423,In_809);
nor U1125 (N_1125,In_173,In_1202);
nand U1126 (N_1126,In_102,In_1321);
nand U1127 (N_1127,In_429,In_459);
or U1128 (N_1128,In_1488,In_1);
nand U1129 (N_1129,In_111,In_193);
nand U1130 (N_1130,In_388,In_346);
nand U1131 (N_1131,In_1477,In_27);
nor U1132 (N_1132,In_138,In_730);
nor U1133 (N_1133,In_655,In_1100);
or U1134 (N_1134,In_958,In_233);
nor U1135 (N_1135,In_1362,In_318);
nand U1136 (N_1136,In_681,In_1330);
and U1137 (N_1137,In_370,In_808);
or U1138 (N_1138,In_688,In_1011);
nand U1139 (N_1139,In_819,In_1389);
xor U1140 (N_1140,In_1144,In_490);
and U1141 (N_1141,In_1260,In_220);
and U1142 (N_1142,In_676,In_884);
and U1143 (N_1143,In_1282,In_400);
nand U1144 (N_1144,In_920,In_778);
or U1145 (N_1145,In_226,In_995);
nor U1146 (N_1146,In_1046,In_666);
nor U1147 (N_1147,In_128,In_1429);
and U1148 (N_1148,In_1294,In_91);
or U1149 (N_1149,In_1132,In_1082);
nor U1150 (N_1150,In_1060,In_32);
nor U1151 (N_1151,In_813,In_528);
or U1152 (N_1152,In_978,In_178);
nor U1153 (N_1153,In_739,In_162);
and U1154 (N_1154,In_6,In_45);
and U1155 (N_1155,In_1187,In_562);
and U1156 (N_1156,In_1112,In_73);
nor U1157 (N_1157,In_1036,In_707);
and U1158 (N_1158,In_955,In_1040);
nand U1159 (N_1159,In_211,In_1151);
nand U1160 (N_1160,In_1486,In_383);
xor U1161 (N_1161,In_275,In_1154);
and U1162 (N_1162,In_546,In_74);
nor U1163 (N_1163,In_627,In_488);
and U1164 (N_1164,In_544,In_998);
nor U1165 (N_1165,In_1011,In_218);
nand U1166 (N_1166,In_1064,In_844);
nor U1167 (N_1167,In_720,In_714);
nand U1168 (N_1168,In_1118,In_562);
and U1169 (N_1169,In_716,In_764);
or U1170 (N_1170,In_631,In_1334);
nand U1171 (N_1171,In_114,In_196);
nand U1172 (N_1172,In_262,In_389);
nor U1173 (N_1173,In_183,In_526);
or U1174 (N_1174,In_1286,In_1174);
or U1175 (N_1175,In_702,In_1064);
nand U1176 (N_1176,In_95,In_6);
nor U1177 (N_1177,In_491,In_1384);
nand U1178 (N_1178,In_394,In_492);
nand U1179 (N_1179,In_377,In_1472);
or U1180 (N_1180,In_963,In_723);
or U1181 (N_1181,In_1484,In_1275);
or U1182 (N_1182,In_179,In_1407);
nand U1183 (N_1183,In_641,In_1341);
or U1184 (N_1184,In_422,In_902);
nand U1185 (N_1185,In_904,In_629);
nand U1186 (N_1186,In_472,In_1);
nor U1187 (N_1187,In_19,In_120);
nor U1188 (N_1188,In_1179,In_1414);
nor U1189 (N_1189,In_296,In_404);
nand U1190 (N_1190,In_950,In_734);
nand U1191 (N_1191,In_820,In_446);
and U1192 (N_1192,In_951,In_237);
or U1193 (N_1193,In_1493,In_1294);
or U1194 (N_1194,In_756,In_1217);
and U1195 (N_1195,In_1115,In_241);
nand U1196 (N_1196,In_945,In_1123);
and U1197 (N_1197,In_399,In_18);
and U1198 (N_1198,In_1135,In_1197);
or U1199 (N_1199,In_515,In_324);
nor U1200 (N_1200,In_1330,In_475);
or U1201 (N_1201,In_303,In_1018);
nand U1202 (N_1202,In_1427,In_1016);
nand U1203 (N_1203,In_447,In_1057);
nand U1204 (N_1204,In_985,In_974);
nand U1205 (N_1205,In_1257,In_884);
nand U1206 (N_1206,In_391,In_636);
nor U1207 (N_1207,In_789,In_1275);
or U1208 (N_1208,In_395,In_591);
nor U1209 (N_1209,In_718,In_1440);
nand U1210 (N_1210,In_121,In_995);
and U1211 (N_1211,In_1424,In_1317);
or U1212 (N_1212,In_1310,In_155);
or U1213 (N_1213,In_683,In_891);
nor U1214 (N_1214,In_304,In_1361);
and U1215 (N_1215,In_620,In_308);
nand U1216 (N_1216,In_639,In_330);
nor U1217 (N_1217,In_44,In_880);
nor U1218 (N_1218,In_1142,In_921);
nor U1219 (N_1219,In_887,In_93);
nand U1220 (N_1220,In_625,In_656);
nand U1221 (N_1221,In_360,In_741);
nor U1222 (N_1222,In_1178,In_356);
and U1223 (N_1223,In_1215,In_832);
nand U1224 (N_1224,In_680,In_588);
or U1225 (N_1225,In_1173,In_513);
nand U1226 (N_1226,In_1170,In_786);
or U1227 (N_1227,In_651,In_732);
nor U1228 (N_1228,In_1345,In_232);
nand U1229 (N_1229,In_830,In_1248);
nor U1230 (N_1230,In_1167,In_1291);
and U1231 (N_1231,In_1439,In_100);
and U1232 (N_1232,In_966,In_440);
nor U1233 (N_1233,In_286,In_210);
and U1234 (N_1234,In_331,In_1397);
nand U1235 (N_1235,In_1350,In_709);
and U1236 (N_1236,In_456,In_1128);
nor U1237 (N_1237,In_1073,In_1034);
or U1238 (N_1238,In_1030,In_105);
nor U1239 (N_1239,In_395,In_1171);
or U1240 (N_1240,In_1032,In_273);
and U1241 (N_1241,In_85,In_1017);
and U1242 (N_1242,In_901,In_109);
and U1243 (N_1243,In_1299,In_117);
nor U1244 (N_1244,In_495,In_593);
and U1245 (N_1245,In_414,In_1056);
and U1246 (N_1246,In_652,In_1187);
and U1247 (N_1247,In_180,In_1369);
nand U1248 (N_1248,In_635,In_571);
nand U1249 (N_1249,In_299,In_1394);
or U1250 (N_1250,In_181,In_1477);
nand U1251 (N_1251,In_83,In_729);
or U1252 (N_1252,In_716,In_690);
nor U1253 (N_1253,In_115,In_52);
and U1254 (N_1254,In_993,In_855);
and U1255 (N_1255,In_72,In_263);
nor U1256 (N_1256,In_347,In_1458);
and U1257 (N_1257,In_454,In_679);
or U1258 (N_1258,In_681,In_1000);
or U1259 (N_1259,In_740,In_170);
and U1260 (N_1260,In_566,In_324);
and U1261 (N_1261,In_734,In_989);
or U1262 (N_1262,In_405,In_542);
nor U1263 (N_1263,In_793,In_131);
nand U1264 (N_1264,In_973,In_1205);
or U1265 (N_1265,In_878,In_157);
nor U1266 (N_1266,In_781,In_1475);
or U1267 (N_1267,In_1453,In_1088);
nor U1268 (N_1268,In_1190,In_148);
or U1269 (N_1269,In_568,In_1273);
and U1270 (N_1270,In_844,In_633);
nor U1271 (N_1271,In_600,In_800);
or U1272 (N_1272,In_567,In_862);
nand U1273 (N_1273,In_641,In_634);
or U1274 (N_1274,In_361,In_1206);
nand U1275 (N_1275,In_488,In_331);
and U1276 (N_1276,In_585,In_571);
nor U1277 (N_1277,In_839,In_1304);
nor U1278 (N_1278,In_1353,In_514);
nor U1279 (N_1279,In_1486,In_1411);
nand U1280 (N_1280,In_286,In_334);
nor U1281 (N_1281,In_242,In_1256);
nor U1282 (N_1282,In_1329,In_991);
nand U1283 (N_1283,In_964,In_583);
and U1284 (N_1284,In_1195,In_134);
nand U1285 (N_1285,In_489,In_1282);
nand U1286 (N_1286,In_261,In_950);
and U1287 (N_1287,In_464,In_483);
and U1288 (N_1288,In_224,In_520);
nor U1289 (N_1289,In_599,In_1015);
and U1290 (N_1290,In_37,In_595);
nor U1291 (N_1291,In_501,In_1371);
or U1292 (N_1292,In_1302,In_203);
nand U1293 (N_1293,In_1356,In_437);
or U1294 (N_1294,In_1308,In_1255);
nand U1295 (N_1295,In_300,In_844);
nor U1296 (N_1296,In_1149,In_1395);
nand U1297 (N_1297,In_1288,In_1388);
and U1298 (N_1298,In_389,In_1102);
nand U1299 (N_1299,In_807,In_532);
nand U1300 (N_1300,In_129,In_1265);
and U1301 (N_1301,In_481,In_906);
or U1302 (N_1302,In_379,In_945);
nand U1303 (N_1303,In_1283,In_901);
nand U1304 (N_1304,In_876,In_1118);
nand U1305 (N_1305,In_439,In_40);
and U1306 (N_1306,In_109,In_821);
nand U1307 (N_1307,In_783,In_1207);
or U1308 (N_1308,In_1158,In_272);
or U1309 (N_1309,In_1205,In_131);
and U1310 (N_1310,In_1394,In_1451);
and U1311 (N_1311,In_63,In_1361);
or U1312 (N_1312,In_45,In_599);
and U1313 (N_1313,In_914,In_811);
and U1314 (N_1314,In_1159,In_383);
nor U1315 (N_1315,In_86,In_42);
or U1316 (N_1316,In_843,In_766);
and U1317 (N_1317,In_968,In_182);
or U1318 (N_1318,In_107,In_698);
nor U1319 (N_1319,In_342,In_936);
and U1320 (N_1320,In_146,In_1185);
and U1321 (N_1321,In_664,In_676);
nand U1322 (N_1322,In_1275,In_385);
nand U1323 (N_1323,In_1308,In_300);
nor U1324 (N_1324,In_113,In_1224);
or U1325 (N_1325,In_1054,In_1262);
and U1326 (N_1326,In_21,In_335);
and U1327 (N_1327,In_306,In_1308);
nor U1328 (N_1328,In_688,In_815);
and U1329 (N_1329,In_1497,In_617);
nor U1330 (N_1330,In_126,In_509);
and U1331 (N_1331,In_1217,In_1072);
nor U1332 (N_1332,In_1394,In_52);
and U1333 (N_1333,In_327,In_1463);
nand U1334 (N_1334,In_1194,In_1375);
nor U1335 (N_1335,In_818,In_346);
and U1336 (N_1336,In_763,In_17);
nor U1337 (N_1337,In_939,In_652);
and U1338 (N_1338,In_610,In_263);
and U1339 (N_1339,In_657,In_1441);
nand U1340 (N_1340,In_979,In_1233);
and U1341 (N_1341,In_395,In_1112);
and U1342 (N_1342,In_698,In_530);
xor U1343 (N_1343,In_1310,In_1053);
and U1344 (N_1344,In_285,In_639);
and U1345 (N_1345,In_1240,In_440);
nor U1346 (N_1346,In_109,In_1118);
or U1347 (N_1347,In_907,In_810);
nor U1348 (N_1348,In_263,In_327);
and U1349 (N_1349,In_726,In_1192);
nor U1350 (N_1350,In_178,In_1452);
nand U1351 (N_1351,In_1029,In_406);
or U1352 (N_1352,In_640,In_1208);
and U1353 (N_1353,In_354,In_449);
nor U1354 (N_1354,In_1444,In_1400);
and U1355 (N_1355,In_569,In_821);
nand U1356 (N_1356,In_842,In_1194);
or U1357 (N_1357,In_965,In_790);
nand U1358 (N_1358,In_1370,In_873);
or U1359 (N_1359,In_602,In_953);
or U1360 (N_1360,In_1320,In_1041);
nor U1361 (N_1361,In_1249,In_44);
nor U1362 (N_1362,In_460,In_808);
nand U1363 (N_1363,In_519,In_1079);
and U1364 (N_1364,In_1422,In_676);
and U1365 (N_1365,In_142,In_853);
nand U1366 (N_1366,In_266,In_828);
nor U1367 (N_1367,In_560,In_627);
nor U1368 (N_1368,In_195,In_1254);
or U1369 (N_1369,In_829,In_527);
or U1370 (N_1370,In_90,In_1301);
and U1371 (N_1371,In_515,In_623);
and U1372 (N_1372,In_164,In_1262);
and U1373 (N_1373,In_344,In_34);
and U1374 (N_1374,In_1128,In_1163);
and U1375 (N_1375,In_85,In_1192);
nor U1376 (N_1376,In_1016,In_423);
and U1377 (N_1377,In_1246,In_1261);
and U1378 (N_1378,In_110,In_140);
and U1379 (N_1379,In_501,In_1021);
and U1380 (N_1380,In_798,In_1404);
and U1381 (N_1381,In_1201,In_465);
and U1382 (N_1382,In_404,In_1040);
nand U1383 (N_1383,In_289,In_1132);
and U1384 (N_1384,In_186,In_252);
and U1385 (N_1385,In_1478,In_632);
nor U1386 (N_1386,In_213,In_32);
nor U1387 (N_1387,In_979,In_896);
nor U1388 (N_1388,In_606,In_145);
nand U1389 (N_1389,In_1297,In_793);
nand U1390 (N_1390,In_475,In_853);
or U1391 (N_1391,In_1379,In_8);
and U1392 (N_1392,In_335,In_1084);
and U1393 (N_1393,In_1337,In_540);
nor U1394 (N_1394,In_202,In_465);
or U1395 (N_1395,In_433,In_9);
nor U1396 (N_1396,In_713,In_883);
nor U1397 (N_1397,In_681,In_1105);
nor U1398 (N_1398,In_939,In_173);
or U1399 (N_1399,In_1441,In_58);
nand U1400 (N_1400,In_790,In_388);
nor U1401 (N_1401,In_466,In_1243);
nand U1402 (N_1402,In_319,In_571);
or U1403 (N_1403,In_26,In_784);
nor U1404 (N_1404,In_1434,In_720);
nand U1405 (N_1405,In_38,In_1392);
or U1406 (N_1406,In_1145,In_130);
and U1407 (N_1407,In_190,In_129);
nor U1408 (N_1408,In_1236,In_491);
or U1409 (N_1409,In_542,In_223);
nand U1410 (N_1410,In_1330,In_613);
and U1411 (N_1411,In_1255,In_1309);
nand U1412 (N_1412,In_403,In_329);
nand U1413 (N_1413,In_1110,In_1189);
nand U1414 (N_1414,In_359,In_1118);
nor U1415 (N_1415,In_684,In_1491);
nand U1416 (N_1416,In_25,In_1054);
nor U1417 (N_1417,In_1127,In_988);
nand U1418 (N_1418,In_673,In_172);
and U1419 (N_1419,In_1109,In_870);
nand U1420 (N_1420,In_1231,In_680);
nor U1421 (N_1421,In_520,In_928);
nor U1422 (N_1422,In_626,In_713);
and U1423 (N_1423,In_755,In_1344);
nand U1424 (N_1424,In_134,In_119);
or U1425 (N_1425,In_710,In_360);
nor U1426 (N_1426,In_1233,In_383);
nor U1427 (N_1427,In_1151,In_694);
and U1428 (N_1428,In_1420,In_1404);
and U1429 (N_1429,In_1187,In_1106);
or U1430 (N_1430,In_1210,In_702);
nor U1431 (N_1431,In_749,In_756);
and U1432 (N_1432,In_355,In_699);
or U1433 (N_1433,In_900,In_622);
nor U1434 (N_1434,In_1445,In_68);
and U1435 (N_1435,In_1164,In_950);
and U1436 (N_1436,In_423,In_1074);
nand U1437 (N_1437,In_455,In_1002);
or U1438 (N_1438,In_604,In_351);
nor U1439 (N_1439,In_1260,In_526);
and U1440 (N_1440,In_1490,In_628);
nor U1441 (N_1441,In_498,In_1482);
or U1442 (N_1442,In_829,In_1373);
nor U1443 (N_1443,In_974,In_857);
or U1444 (N_1444,In_908,In_658);
nand U1445 (N_1445,In_411,In_32);
or U1446 (N_1446,In_1194,In_736);
and U1447 (N_1447,In_1036,In_249);
nand U1448 (N_1448,In_1180,In_628);
nor U1449 (N_1449,In_1002,In_1495);
or U1450 (N_1450,In_1228,In_1365);
nand U1451 (N_1451,In_1483,In_203);
nor U1452 (N_1452,In_124,In_25);
and U1453 (N_1453,In_840,In_60);
and U1454 (N_1454,In_1266,In_1319);
or U1455 (N_1455,In_441,In_851);
and U1456 (N_1456,In_464,In_392);
and U1457 (N_1457,In_472,In_384);
nor U1458 (N_1458,In_515,In_874);
nor U1459 (N_1459,In_954,In_174);
nor U1460 (N_1460,In_31,In_996);
nor U1461 (N_1461,In_1399,In_443);
nand U1462 (N_1462,In_1244,In_1432);
nor U1463 (N_1463,In_1376,In_1216);
and U1464 (N_1464,In_725,In_650);
nand U1465 (N_1465,In_44,In_320);
or U1466 (N_1466,In_359,In_597);
nand U1467 (N_1467,In_1487,In_617);
and U1468 (N_1468,In_1055,In_1135);
nor U1469 (N_1469,In_191,In_637);
and U1470 (N_1470,In_1435,In_921);
nor U1471 (N_1471,In_1144,In_418);
xnor U1472 (N_1472,In_725,In_62);
or U1473 (N_1473,In_663,In_797);
nand U1474 (N_1474,In_1266,In_501);
nand U1475 (N_1475,In_747,In_1273);
nor U1476 (N_1476,In_45,In_1277);
and U1477 (N_1477,In_875,In_773);
nor U1478 (N_1478,In_420,In_1221);
nand U1479 (N_1479,In_1000,In_886);
nand U1480 (N_1480,In_480,In_1479);
or U1481 (N_1481,In_819,In_749);
nand U1482 (N_1482,In_248,In_1094);
nor U1483 (N_1483,In_179,In_641);
and U1484 (N_1484,In_423,In_757);
and U1485 (N_1485,In_350,In_830);
nor U1486 (N_1486,In_1453,In_225);
nor U1487 (N_1487,In_763,In_747);
nand U1488 (N_1488,In_228,In_1306);
nand U1489 (N_1489,In_158,In_631);
or U1490 (N_1490,In_357,In_1058);
nor U1491 (N_1491,In_1397,In_82);
nand U1492 (N_1492,In_244,In_1177);
or U1493 (N_1493,In_70,In_1479);
nor U1494 (N_1494,In_460,In_842);
nand U1495 (N_1495,In_1126,In_1012);
or U1496 (N_1496,In_1318,In_1016);
or U1497 (N_1497,In_350,In_1490);
nand U1498 (N_1498,In_1346,In_60);
nand U1499 (N_1499,In_875,In_953);
or U1500 (N_1500,In_1244,In_328);
or U1501 (N_1501,In_8,In_1006);
and U1502 (N_1502,In_215,In_1013);
and U1503 (N_1503,In_33,In_450);
nand U1504 (N_1504,In_805,In_1375);
nor U1505 (N_1505,In_1272,In_1142);
or U1506 (N_1506,In_304,In_1068);
and U1507 (N_1507,In_341,In_220);
nand U1508 (N_1508,In_930,In_788);
or U1509 (N_1509,In_831,In_1214);
nor U1510 (N_1510,In_1156,In_694);
nand U1511 (N_1511,In_1059,In_1085);
nand U1512 (N_1512,In_850,In_1247);
nand U1513 (N_1513,In_1452,In_498);
or U1514 (N_1514,In_1401,In_177);
nor U1515 (N_1515,In_1356,In_1354);
nand U1516 (N_1516,In_513,In_1284);
nand U1517 (N_1517,In_339,In_1381);
and U1518 (N_1518,In_488,In_951);
nand U1519 (N_1519,In_78,In_709);
nand U1520 (N_1520,In_458,In_1059);
and U1521 (N_1521,In_760,In_477);
nor U1522 (N_1522,In_7,In_914);
nand U1523 (N_1523,In_450,In_726);
nor U1524 (N_1524,In_773,In_1079);
and U1525 (N_1525,In_1445,In_483);
nand U1526 (N_1526,In_1489,In_731);
and U1527 (N_1527,In_1000,In_831);
or U1528 (N_1528,In_837,In_978);
nand U1529 (N_1529,In_1179,In_1448);
nand U1530 (N_1530,In_386,In_97);
nand U1531 (N_1531,In_1423,In_482);
or U1532 (N_1532,In_784,In_517);
nand U1533 (N_1533,In_821,In_1293);
nand U1534 (N_1534,In_273,In_142);
or U1535 (N_1535,In_1425,In_8);
nor U1536 (N_1536,In_800,In_1462);
or U1537 (N_1537,In_524,In_1207);
or U1538 (N_1538,In_1177,In_681);
and U1539 (N_1539,In_790,In_691);
nand U1540 (N_1540,In_372,In_502);
nor U1541 (N_1541,In_341,In_129);
or U1542 (N_1542,In_1391,In_674);
nor U1543 (N_1543,In_1270,In_817);
nand U1544 (N_1544,In_1353,In_1324);
nand U1545 (N_1545,In_1025,In_311);
and U1546 (N_1546,In_332,In_1114);
nor U1547 (N_1547,In_1035,In_1333);
nor U1548 (N_1548,In_183,In_373);
nand U1549 (N_1549,In_1038,In_1482);
and U1550 (N_1550,In_928,In_868);
and U1551 (N_1551,In_204,In_894);
nor U1552 (N_1552,In_261,In_686);
nor U1553 (N_1553,In_931,In_1298);
nand U1554 (N_1554,In_369,In_600);
nor U1555 (N_1555,In_84,In_1106);
or U1556 (N_1556,In_216,In_642);
and U1557 (N_1557,In_835,In_413);
nor U1558 (N_1558,In_785,In_255);
nand U1559 (N_1559,In_332,In_1020);
nand U1560 (N_1560,In_534,In_430);
nand U1561 (N_1561,In_1313,In_499);
or U1562 (N_1562,In_261,In_262);
nand U1563 (N_1563,In_300,In_569);
or U1564 (N_1564,In_120,In_947);
or U1565 (N_1565,In_510,In_50);
or U1566 (N_1566,In_784,In_951);
and U1567 (N_1567,In_880,In_609);
nor U1568 (N_1568,In_655,In_1073);
nor U1569 (N_1569,In_1012,In_685);
nand U1570 (N_1570,In_76,In_74);
nor U1571 (N_1571,In_148,In_1262);
or U1572 (N_1572,In_135,In_1108);
nor U1573 (N_1573,In_321,In_404);
or U1574 (N_1574,In_3,In_1468);
nor U1575 (N_1575,In_37,In_993);
or U1576 (N_1576,In_109,In_1226);
or U1577 (N_1577,In_1082,In_1310);
or U1578 (N_1578,In_275,In_1024);
and U1579 (N_1579,In_1171,In_1367);
or U1580 (N_1580,In_113,In_1086);
or U1581 (N_1581,In_1041,In_540);
nand U1582 (N_1582,In_1012,In_1225);
or U1583 (N_1583,In_203,In_1344);
nand U1584 (N_1584,In_970,In_1050);
and U1585 (N_1585,In_935,In_658);
nand U1586 (N_1586,In_728,In_299);
nand U1587 (N_1587,In_370,In_1118);
nor U1588 (N_1588,In_1321,In_1266);
and U1589 (N_1589,In_589,In_194);
nor U1590 (N_1590,In_656,In_129);
and U1591 (N_1591,In_872,In_513);
nand U1592 (N_1592,In_1009,In_920);
nor U1593 (N_1593,In_689,In_736);
nor U1594 (N_1594,In_804,In_50);
nand U1595 (N_1595,In_238,In_114);
and U1596 (N_1596,In_368,In_24);
and U1597 (N_1597,In_576,In_1457);
nor U1598 (N_1598,In_428,In_1112);
and U1599 (N_1599,In_1197,In_1048);
or U1600 (N_1600,In_956,In_551);
nand U1601 (N_1601,In_392,In_1127);
nand U1602 (N_1602,In_746,In_1015);
nand U1603 (N_1603,In_1489,In_769);
and U1604 (N_1604,In_616,In_313);
nand U1605 (N_1605,In_1241,In_1017);
and U1606 (N_1606,In_1410,In_518);
and U1607 (N_1607,In_1483,In_582);
nor U1608 (N_1608,In_721,In_1324);
and U1609 (N_1609,In_1001,In_140);
and U1610 (N_1610,In_2,In_894);
and U1611 (N_1611,In_580,In_1359);
or U1612 (N_1612,In_1497,In_354);
or U1613 (N_1613,In_946,In_103);
or U1614 (N_1614,In_811,In_147);
or U1615 (N_1615,In_859,In_963);
nand U1616 (N_1616,In_438,In_1028);
and U1617 (N_1617,In_864,In_372);
or U1618 (N_1618,In_1441,In_66);
or U1619 (N_1619,In_1034,In_1451);
nand U1620 (N_1620,In_961,In_1169);
or U1621 (N_1621,In_697,In_852);
nand U1622 (N_1622,In_829,In_96);
nor U1623 (N_1623,In_289,In_1060);
and U1624 (N_1624,In_1183,In_1060);
nor U1625 (N_1625,In_5,In_1010);
nand U1626 (N_1626,In_462,In_109);
or U1627 (N_1627,In_624,In_642);
nor U1628 (N_1628,In_1215,In_313);
nand U1629 (N_1629,In_1494,In_57);
or U1630 (N_1630,In_1498,In_1067);
nor U1631 (N_1631,In_658,In_160);
nand U1632 (N_1632,In_1414,In_752);
nand U1633 (N_1633,In_125,In_1153);
and U1634 (N_1634,In_1043,In_1291);
and U1635 (N_1635,In_988,In_738);
and U1636 (N_1636,In_654,In_813);
nor U1637 (N_1637,In_83,In_367);
nand U1638 (N_1638,In_292,In_1427);
nor U1639 (N_1639,In_1097,In_1088);
nand U1640 (N_1640,In_373,In_835);
nand U1641 (N_1641,In_777,In_1240);
nor U1642 (N_1642,In_1030,In_328);
or U1643 (N_1643,In_1319,In_640);
xor U1644 (N_1644,In_1241,In_61);
nor U1645 (N_1645,In_858,In_1098);
nand U1646 (N_1646,In_731,In_359);
and U1647 (N_1647,In_430,In_836);
or U1648 (N_1648,In_183,In_1377);
or U1649 (N_1649,In_1187,In_707);
or U1650 (N_1650,In_550,In_1391);
or U1651 (N_1651,In_980,In_803);
or U1652 (N_1652,In_1386,In_117);
or U1653 (N_1653,In_136,In_49);
and U1654 (N_1654,In_418,In_415);
or U1655 (N_1655,In_27,In_1221);
or U1656 (N_1656,In_562,In_1244);
or U1657 (N_1657,In_96,In_154);
or U1658 (N_1658,In_1127,In_1130);
or U1659 (N_1659,In_1207,In_1083);
nor U1660 (N_1660,In_1460,In_1336);
nor U1661 (N_1661,In_759,In_885);
nor U1662 (N_1662,In_1312,In_605);
nor U1663 (N_1663,In_1293,In_1037);
nand U1664 (N_1664,In_168,In_242);
and U1665 (N_1665,In_376,In_1464);
or U1666 (N_1666,In_1126,In_1369);
nor U1667 (N_1667,In_490,In_789);
and U1668 (N_1668,In_1482,In_1045);
and U1669 (N_1669,In_809,In_1305);
nand U1670 (N_1670,In_691,In_1449);
or U1671 (N_1671,In_959,In_830);
or U1672 (N_1672,In_1354,In_373);
and U1673 (N_1673,In_1361,In_978);
nor U1674 (N_1674,In_349,In_271);
or U1675 (N_1675,In_754,In_181);
nor U1676 (N_1676,In_52,In_1373);
nor U1677 (N_1677,In_191,In_536);
and U1678 (N_1678,In_26,In_519);
or U1679 (N_1679,In_1369,In_1304);
nand U1680 (N_1680,In_450,In_554);
and U1681 (N_1681,In_1475,In_499);
or U1682 (N_1682,In_734,In_617);
and U1683 (N_1683,In_616,In_1355);
xnor U1684 (N_1684,In_224,In_710);
nor U1685 (N_1685,In_1226,In_631);
and U1686 (N_1686,In_870,In_138);
nand U1687 (N_1687,In_66,In_38);
and U1688 (N_1688,In_252,In_1299);
or U1689 (N_1689,In_729,In_182);
nand U1690 (N_1690,In_572,In_1196);
nand U1691 (N_1691,In_803,In_837);
nor U1692 (N_1692,In_100,In_642);
and U1693 (N_1693,In_1411,In_1083);
nand U1694 (N_1694,In_320,In_871);
or U1695 (N_1695,In_410,In_758);
or U1696 (N_1696,In_112,In_776);
nor U1697 (N_1697,In_1249,In_1265);
xor U1698 (N_1698,In_154,In_1231);
nor U1699 (N_1699,In_1189,In_48);
nand U1700 (N_1700,In_1324,In_1405);
and U1701 (N_1701,In_16,In_1487);
or U1702 (N_1702,In_151,In_365);
or U1703 (N_1703,In_1141,In_592);
nand U1704 (N_1704,In_1394,In_540);
and U1705 (N_1705,In_1479,In_630);
and U1706 (N_1706,In_8,In_1434);
nand U1707 (N_1707,In_997,In_282);
nand U1708 (N_1708,In_498,In_35);
nor U1709 (N_1709,In_164,In_201);
or U1710 (N_1710,In_1342,In_1237);
or U1711 (N_1711,In_1031,In_439);
and U1712 (N_1712,In_1048,In_360);
or U1713 (N_1713,In_1327,In_238);
nor U1714 (N_1714,In_47,In_1440);
and U1715 (N_1715,In_226,In_828);
nand U1716 (N_1716,In_1127,In_1251);
or U1717 (N_1717,In_398,In_654);
nor U1718 (N_1718,In_1228,In_1068);
nand U1719 (N_1719,In_1208,In_563);
nand U1720 (N_1720,In_185,In_1257);
nor U1721 (N_1721,In_938,In_325);
nand U1722 (N_1722,In_23,In_692);
nand U1723 (N_1723,In_432,In_75);
nor U1724 (N_1724,In_1312,In_1268);
nor U1725 (N_1725,In_603,In_668);
nor U1726 (N_1726,In_1183,In_769);
or U1727 (N_1727,In_196,In_1064);
and U1728 (N_1728,In_939,In_749);
and U1729 (N_1729,In_1062,In_720);
and U1730 (N_1730,In_1479,In_798);
nor U1731 (N_1731,In_348,In_50);
or U1732 (N_1732,In_1248,In_666);
xnor U1733 (N_1733,In_1393,In_960);
and U1734 (N_1734,In_1029,In_79);
nand U1735 (N_1735,In_1496,In_590);
and U1736 (N_1736,In_850,In_146);
nor U1737 (N_1737,In_80,In_1344);
nand U1738 (N_1738,In_53,In_1068);
and U1739 (N_1739,In_136,In_1403);
and U1740 (N_1740,In_219,In_523);
and U1741 (N_1741,In_317,In_253);
nand U1742 (N_1742,In_838,In_360);
nor U1743 (N_1743,In_162,In_1110);
nor U1744 (N_1744,In_399,In_323);
nor U1745 (N_1745,In_1312,In_501);
nor U1746 (N_1746,In_134,In_753);
and U1747 (N_1747,In_1357,In_1159);
or U1748 (N_1748,In_1447,In_265);
nand U1749 (N_1749,In_812,In_352);
and U1750 (N_1750,In_207,In_426);
or U1751 (N_1751,In_771,In_50);
and U1752 (N_1752,In_1286,In_663);
nand U1753 (N_1753,In_1423,In_1358);
and U1754 (N_1754,In_563,In_985);
or U1755 (N_1755,In_1130,In_221);
and U1756 (N_1756,In_330,In_981);
or U1757 (N_1757,In_208,In_1255);
and U1758 (N_1758,In_1088,In_235);
and U1759 (N_1759,In_1432,In_328);
or U1760 (N_1760,In_30,In_126);
nand U1761 (N_1761,In_1037,In_816);
nand U1762 (N_1762,In_407,In_1419);
and U1763 (N_1763,In_505,In_138);
nor U1764 (N_1764,In_263,In_764);
nor U1765 (N_1765,In_504,In_1391);
and U1766 (N_1766,In_384,In_909);
nand U1767 (N_1767,In_286,In_1306);
and U1768 (N_1768,In_885,In_563);
and U1769 (N_1769,In_1195,In_549);
or U1770 (N_1770,In_351,In_1232);
nand U1771 (N_1771,In_1438,In_1);
nor U1772 (N_1772,In_1007,In_1240);
nor U1773 (N_1773,In_248,In_476);
or U1774 (N_1774,In_1179,In_409);
nand U1775 (N_1775,In_1149,In_372);
nand U1776 (N_1776,In_1230,In_1386);
nand U1777 (N_1777,In_565,In_83);
nand U1778 (N_1778,In_254,In_1316);
and U1779 (N_1779,In_361,In_660);
and U1780 (N_1780,In_667,In_1207);
nand U1781 (N_1781,In_1011,In_199);
and U1782 (N_1782,In_483,In_218);
nor U1783 (N_1783,In_224,In_1222);
nor U1784 (N_1784,In_1377,In_422);
nor U1785 (N_1785,In_34,In_156);
nor U1786 (N_1786,In_727,In_408);
nand U1787 (N_1787,In_564,In_1274);
nor U1788 (N_1788,In_1374,In_546);
and U1789 (N_1789,In_129,In_276);
nand U1790 (N_1790,In_1317,In_465);
and U1791 (N_1791,In_948,In_1226);
nor U1792 (N_1792,In_1038,In_719);
nand U1793 (N_1793,In_872,In_1234);
nand U1794 (N_1794,In_1055,In_903);
or U1795 (N_1795,In_592,In_1320);
nand U1796 (N_1796,In_1215,In_1499);
nor U1797 (N_1797,In_259,In_362);
or U1798 (N_1798,In_1073,In_1377);
xnor U1799 (N_1799,In_601,In_59);
nand U1800 (N_1800,In_1307,In_492);
nor U1801 (N_1801,In_806,In_1162);
and U1802 (N_1802,In_745,In_289);
and U1803 (N_1803,In_298,In_1457);
or U1804 (N_1804,In_648,In_1352);
nand U1805 (N_1805,In_267,In_425);
nand U1806 (N_1806,In_1083,In_186);
or U1807 (N_1807,In_79,In_1390);
and U1808 (N_1808,In_909,In_517);
or U1809 (N_1809,In_1115,In_59);
nor U1810 (N_1810,In_181,In_791);
nand U1811 (N_1811,In_758,In_838);
xnor U1812 (N_1812,In_285,In_220);
nor U1813 (N_1813,In_319,In_708);
or U1814 (N_1814,In_1307,In_131);
nand U1815 (N_1815,In_1396,In_969);
or U1816 (N_1816,In_393,In_903);
and U1817 (N_1817,In_82,In_1015);
and U1818 (N_1818,In_1449,In_850);
nand U1819 (N_1819,In_1351,In_607);
and U1820 (N_1820,In_1010,In_710);
nand U1821 (N_1821,In_784,In_1190);
nor U1822 (N_1822,In_851,In_1083);
xor U1823 (N_1823,In_312,In_757);
nor U1824 (N_1824,In_439,In_893);
or U1825 (N_1825,In_912,In_55);
or U1826 (N_1826,In_604,In_88);
nand U1827 (N_1827,In_409,In_1371);
nand U1828 (N_1828,In_1448,In_220);
xnor U1829 (N_1829,In_221,In_307);
or U1830 (N_1830,In_1225,In_1178);
or U1831 (N_1831,In_1330,In_571);
nand U1832 (N_1832,In_215,In_618);
or U1833 (N_1833,In_1319,In_1333);
nor U1834 (N_1834,In_525,In_598);
nor U1835 (N_1835,In_101,In_73);
nand U1836 (N_1836,In_527,In_263);
or U1837 (N_1837,In_987,In_120);
nor U1838 (N_1838,In_569,In_677);
nand U1839 (N_1839,In_278,In_1415);
nor U1840 (N_1840,In_191,In_1125);
nor U1841 (N_1841,In_871,In_361);
and U1842 (N_1842,In_488,In_125);
nor U1843 (N_1843,In_309,In_1367);
nand U1844 (N_1844,In_774,In_18);
and U1845 (N_1845,In_857,In_544);
nor U1846 (N_1846,In_88,In_1151);
nand U1847 (N_1847,In_1276,In_425);
or U1848 (N_1848,In_950,In_778);
or U1849 (N_1849,In_444,In_32);
nor U1850 (N_1850,In_420,In_520);
or U1851 (N_1851,In_401,In_1172);
and U1852 (N_1852,In_1330,In_913);
or U1853 (N_1853,In_1068,In_1334);
or U1854 (N_1854,In_1046,In_1113);
and U1855 (N_1855,In_1411,In_908);
nand U1856 (N_1856,In_821,In_50);
or U1857 (N_1857,In_949,In_1101);
and U1858 (N_1858,In_619,In_1317);
and U1859 (N_1859,In_1250,In_980);
nor U1860 (N_1860,In_968,In_408);
and U1861 (N_1861,In_855,In_385);
or U1862 (N_1862,In_1116,In_1134);
nor U1863 (N_1863,In_900,In_982);
or U1864 (N_1864,In_1256,In_1011);
nand U1865 (N_1865,In_543,In_73);
nand U1866 (N_1866,In_134,In_711);
nor U1867 (N_1867,In_468,In_161);
and U1868 (N_1868,In_127,In_978);
nor U1869 (N_1869,In_1165,In_118);
or U1870 (N_1870,In_1357,In_807);
and U1871 (N_1871,In_825,In_1084);
nand U1872 (N_1872,In_225,In_509);
or U1873 (N_1873,In_315,In_866);
nand U1874 (N_1874,In_1211,In_1338);
nand U1875 (N_1875,In_1284,In_1429);
xnor U1876 (N_1876,In_77,In_905);
nor U1877 (N_1877,In_199,In_728);
or U1878 (N_1878,In_310,In_1264);
or U1879 (N_1879,In_1336,In_1213);
or U1880 (N_1880,In_115,In_73);
nand U1881 (N_1881,In_447,In_1450);
nor U1882 (N_1882,In_809,In_294);
nand U1883 (N_1883,In_1238,In_27);
and U1884 (N_1884,In_1386,In_859);
nor U1885 (N_1885,In_234,In_1216);
nand U1886 (N_1886,In_1055,In_1234);
nor U1887 (N_1887,In_1065,In_837);
or U1888 (N_1888,In_1180,In_857);
and U1889 (N_1889,In_853,In_440);
nor U1890 (N_1890,In_1268,In_1103);
or U1891 (N_1891,In_583,In_825);
or U1892 (N_1892,In_850,In_203);
nand U1893 (N_1893,In_359,In_1137);
nor U1894 (N_1894,In_1068,In_1009);
nand U1895 (N_1895,In_1283,In_905);
nor U1896 (N_1896,In_259,In_1355);
or U1897 (N_1897,In_70,In_138);
nor U1898 (N_1898,In_1082,In_735);
or U1899 (N_1899,In_165,In_181);
and U1900 (N_1900,In_781,In_1479);
and U1901 (N_1901,In_852,In_1477);
and U1902 (N_1902,In_1332,In_1168);
nand U1903 (N_1903,In_1004,In_1460);
nor U1904 (N_1904,In_746,In_1473);
and U1905 (N_1905,In_459,In_851);
nor U1906 (N_1906,In_1380,In_573);
or U1907 (N_1907,In_221,In_1424);
nand U1908 (N_1908,In_46,In_231);
nor U1909 (N_1909,In_3,In_175);
and U1910 (N_1910,In_930,In_951);
nor U1911 (N_1911,In_803,In_519);
nand U1912 (N_1912,In_520,In_1152);
or U1913 (N_1913,In_286,In_791);
or U1914 (N_1914,In_1305,In_490);
nor U1915 (N_1915,In_605,In_1152);
nor U1916 (N_1916,In_794,In_923);
nand U1917 (N_1917,In_594,In_1038);
and U1918 (N_1918,In_612,In_610);
and U1919 (N_1919,In_892,In_289);
or U1920 (N_1920,In_214,In_210);
or U1921 (N_1921,In_741,In_1442);
and U1922 (N_1922,In_612,In_32);
nand U1923 (N_1923,In_1281,In_786);
nor U1924 (N_1924,In_1409,In_900);
nor U1925 (N_1925,In_1473,In_719);
or U1926 (N_1926,In_711,In_396);
or U1927 (N_1927,In_318,In_330);
nand U1928 (N_1928,In_1039,In_420);
and U1929 (N_1929,In_976,In_290);
or U1930 (N_1930,In_1392,In_995);
nand U1931 (N_1931,In_1054,In_1470);
nor U1932 (N_1932,In_614,In_651);
nand U1933 (N_1933,In_1287,In_862);
xnor U1934 (N_1934,In_1305,In_1279);
and U1935 (N_1935,In_897,In_1274);
nand U1936 (N_1936,In_235,In_587);
and U1937 (N_1937,In_16,In_687);
nor U1938 (N_1938,In_23,In_391);
or U1939 (N_1939,In_500,In_1036);
nand U1940 (N_1940,In_1033,In_155);
nor U1941 (N_1941,In_249,In_55);
or U1942 (N_1942,In_333,In_275);
nand U1943 (N_1943,In_1047,In_1120);
nand U1944 (N_1944,In_337,In_1021);
or U1945 (N_1945,In_218,In_1030);
nor U1946 (N_1946,In_274,In_859);
nor U1947 (N_1947,In_1413,In_436);
or U1948 (N_1948,In_248,In_1027);
and U1949 (N_1949,In_888,In_848);
and U1950 (N_1950,In_1130,In_184);
or U1951 (N_1951,In_1336,In_154);
nand U1952 (N_1952,In_1172,In_467);
nand U1953 (N_1953,In_15,In_1435);
and U1954 (N_1954,In_1406,In_1309);
nand U1955 (N_1955,In_597,In_266);
and U1956 (N_1956,In_963,In_879);
or U1957 (N_1957,In_1106,In_757);
nor U1958 (N_1958,In_1186,In_1408);
nor U1959 (N_1959,In_354,In_1216);
nor U1960 (N_1960,In_621,In_516);
nor U1961 (N_1961,In_209,In_52);
or U1962 (N_1962,In_1360,In_999);
or U1963 (N_1963,In_1333,In_1272);
nand U1964 (N_1964,In_903,In_467);
and U1965 (N_1965,In_133,In_165);
nand U1966 (N_1966,In_536,In_893);
nor U1967 (N_1967,In_825,In_167);
and U1968 (N_1968,In_936,In_621);
or U1969 (N_1969,In_181,In_919);
or U1970 (N_1970,In_652,In_845);
nand U1971 (N_1971,In_449,In_85);
nor U1972 (N_1972,In_136,In_1370);
nand U1973 (N_1973,In_1066,In_837);
or U1974 (N_1974,In_593,In_1163);
or U1975 (N_1975,In_452,In_1);
nand U1976 (N_1976,In_170,In_1156);
or U1977 (N_1977,In_1460,In_1108);
and U1978 (N_1978,In_250,In_1107);
nor U1979 (N_1979,In_1180,In_474);
nor U1980 (N_1980,In_1094,In_185);
and U1981 (N_1981,In_21,In_266);
nand U1982 (N_1982,In_1449,In_1107);
or U1983 (N_1983,In_858,In_386);
nor U1984 (N_1984,In_679,In_778);
nor U1985 (N_1985,In_53,In_1492);
nand U1986 (N_1986,In_1028,In_649);
or U1987 (N_1987,In_1485,In_844);
nand U1988 (N_1988,In_255,In_1066);
or U1989 (N_1989,In_572,In_1246);
or U1990 (N_1990,In_266,In_1075);
nand U1991 (N_1991,In_798,In_554);
nor U1992 (N_1992,In_1129,In_422);
and U1993 (N_1993,In_925,In_1267);
nand U1994 (N_1994,In_995,In_544);
nor U1995 (N_1995,In_45,In_540);
and U1996 (N_1996,In_827,In_512);
nor U1997 (N_1997,In_126,In_746);
and U1998 (N_1998,In_1271,In_83);
and U1999 (N_1999,In_1070,In_1178);
or U2000 (N_2000,In_601,In_886);
and U2001 (N_2001,In_1291,In_984);
or U2002 (N_2002,In_1183,In_278);
or U2003 (N_2003,In_993,In_1000);
or U2004 (N_2004,In_308,In_753);
or U2005 (N_2005,In_239,In_112);
and U2006 (N_2006,In_682,In_718);
nor U2007 (N_2007,In_1406,In_258);
nor U2008 (N_2008,In_1454,In_400);
or U2009 (N_2009,In_1241,In_1170);
or U2010 (N_2010,In_1006,In_177);
nor U2011 (N_2011,In_1205,In_188);
or U2012 (N_2012,In_966,In_54);
or U2013 (N_2013,In_307,In_1363);
or U2014 (N_2014,In_1243,In_1007);
nand U2015 (N_2015,In_1269,In_1005);
and U2016 (N_2016,In_1473,In_151);
nand U2017 (N_2017,In_44,In_1068);
nand U2018 (N_2018,In_871,In_787);
and U2019 (N_2019,In_807,In_1427);
nand U2020 (N_2020,In_85,In_893);
or U2021 (N_2021,In_1153,In_829);
nor U2022 (N_2022,In_1450,In_1149);
or U2023 (N_2023,In_873,In_1036);
or U2024 (N_2024,In_614,In_989);
nor U2025 (N_2025,In_666,In_1275);
and U2026 (N_2026,In_157,In_1286);
nand U2027 (N_2027,In_590,In_954);
nor U2028 (N_2028,In_592,In_464);
and U2029 (N_2029,In_455,In_317);
nand U2030 (N_2030,In_1071,In_353);
or U2031 (N_2031,In_383,In_734);
nor U2032 (N_2032,In_874,In_1275);
nand U2033 (N_2033,In_609,In_715);
and U2034 (N_2034,In_217,In_519);
or U2035 (N_2035,In_589,In_928);
nand U2036 (N_2036,In_732,In_1238);
nand U2037 (N_2037,In_748,In_197);
or U2038 (N_2038,In_1225,In_908);
or U2039 (N_2039,In_1099,In_94);
nor U2040 (N_2040,In_542,In_1489);
or U2041 (N_2041,In_1103,In_566);
and U2042 (N_2042,In_187,In_407);
and U2043 (N_2043,In_120,In_1293);
and U2044 (N_2044,In_980,In_244);
xor U2045 (N_2045,In_817,In_251);
and U2046 (N_2046,In_1035,In_117);
and U2047 (N_2047,In_400,In_1197);
or U2048 (N_2048,In_72,In_588);
nor U2049 (N_2049,In_313,In_67);
nand U2050 (N_2050,In_310,In_1155);
and U2051 (N_2051,In_229,In_1337);
nor U2052 (N_2052,In_187,In_557);
nor U2053 (N_2053,In_1158,In_1200);
and U2054 (N_2054,In_202,In_1320);
and U2055 (N_2055,In_1096,In_1414);
or U2056 (N_2056,In_631,In_1005);
nand U2057 (N_2057,In_1416,In_832);
or U2058 (N_2058,In_1205,In_1459);
nor U2059 (N_2059,In_449,In_802);
and U2060 (N_2060,In_870,In_263);
nor U2061 (N_2061,In_191,In_33);
xor U2062 (N_2062,In_48,In_704);
nor U2063 (N_2063,In_313,In_1408);
and U2064 (N_2064,In_1445,In_1249);
nand U2065 (N_2065,In_984,In_827);
and U2066 (N_2066,In_1384,In_143);
nand U2067 (N_2067,In_757,In_254);
or U2068 (N_2068,In_831,In_1456);
and U2069 (N_2069,In_672,In_1013);
nand U2070 (N_2070,In_214,In_371);
nor U2071 (N_2071,In_518,In_767);
and U2072 (N_2072,In_1489,In_650);
nand U2073 (N_2073,In_976,In_250);
and U2074 (N_2074,In_258,In_216);
nand U2075 (N_2075,In_839,In_512);
nor U2076 (N_2076,In_1040,In_692);
and U2077 (N_2077,In_910,In_310);
nand U2078 (N_2078,In_111,In_671);
nor U2079 (N_2079,In_197,In_626);
nand U2080 (N_2080,In_1172,In_772);
or U2081 (N_2081,In_174,In_687);
or U2082 (N_2082,In_328,In_422);
nor U2083 (N_2083,In_702,In_704);
and U2084 (N_2084,In_208,In_1286);
nand U2085 (N_2085,In_1051,In_334);
nor U2086 (N_2086,In_1015,In_1327);
nand U2087 (N_2087,In_118,In_206);
nand U2088 (N_2088,In_315,In_1085);
nor U2089 (N_2089,In_398,In_758);
and U2090 (N_2090,In_1345,In_958);
nor U2091 (N_2091,In_1320,In_875);
and U2092 (N_2092,In_1401,In_1316);
or U2093 (N_2093,In_181,In_1016);
and U2094 (N_2094,In_734,In_187);
xor U2095 (N_2095,In_514,In_330);
or U2096 (N_2096,In_687,In_451);
and U2097 (N_2097,In_766,In_1126);
nor U2098 (N_2098,In_1265,In_741);
and U2099 (N_2099,In_731,In_910);
nor U2100 (N_2100,In_1305,In_1363);
nand U2101 (N_2101,In_978,In_555);
or U2102 (N_2102,In_1336,In_1465);
nor U2103 (N_2103,In_1143,In_862);
nor U2104 (N_2104,In_711,In_706);
nor U2105 (N_2105,In_717,In_95);
nand U2106 (N_2106,In_536,In_751);
nand U2107 (N_2107,In_1088,In_844);
nor U2108 (N_2108,In_959,In_519);
or U2109 (N_2109,In_788,In_175);
and U2110 (N_2110,In_1051,In_16);
or U2111 (N_2111,In_708,In_27);
and U2112 (N_2112,In_999,In_335);
nor U2113 (N_2113,In_1215,In_346);
and U2114 (N_2114,In_1411,In_454);
and U2115 (N_2115,In_1354,In_1122);
and U2116 (N_2116,In_400,In_1219);
nand U2117 (N_2117,In_193,In_347);
nand U2118 (N_2118,In_676,In_103);
nor U2119 (N_2119,In_499,In_621);
nand U2120 (N_2120,In_496,In_943);
nor U2121 (N_2121,In_1323,In_217);
and U2122 (N_2122,In_313,In_135);
nand U2123 (N_2123,In_527,In_73);
nor U2124 (N_2124,In_1007,In_1241);
xor U2125 (N_2125,In_1329,In_1373);
or U2126 (N_2126,In_904,In_481);
and U2127 (N_2127,In_958,In_936);
and U2128 (N_2128,In_102,In_1165);
nor U2129 (N_2129,In_196,In_999);
or U2130 (N_2130,In_1383,In_376);
nand U2131 (N_2131,In_437,In_914);
nor U2132 (N_2132,In_333,In_950);
and U2133 (N_2133,In_1487,In_1158);
nand U2134 (N_2134,In_1236,In_385);
nand U2135 (N_2135,In_1105,In_639);
or U2136 (N_2136,In_1221,In_1280);
nand U2137 (N_2137,In_1139,In_744);
nor U2138 (N_2138,In_1236,In_1029);
nor U2139 (N_2139,In_1122,In_956);
nor U2140 (N_2140,In_555,In_1345);
nor U2141 (N_2141,In_682,In_354);
and U2142 (N_2142,In_843,In_133);
nor U2143 (N_2143,In_1158,In_790);
nand U2144 (N_2144,In_971,In_199);
nor U2145 (N_2145,In_1006,In_1268);
and U2146 (N_2146,In_1252,In_365);
or U2147 (N_2147,In_186,In_190);
nor U2148 (N_2148,In_1490,In_696);
and U2149 (N_2149,In_346,In_738);
and U2150 (N_2150,In_875,In_1427);
or U2151 (N_2151,In_876,In_924);
and U2152 (N_2152,In_1439,In_1290);
nand U2153 (N_2153,In_183,In_248);
nand U2154 (N_2154,In_1179,In_310);
or U2155 (N_2155,In_1386,In_846);
or U2156 (N_2156,In_704,In_210);
nand U2157 (N_2157,In_695,In_1292);
nand U2158 (N_2158,In_194,In_1348);
or U2159 (N_2159,In_364,In_1311);
or U2160 (N_2160,In_1226,In_618);
nor U2161 (N_2161,In_645,In_353);
nor U2162 (N_2162,In_1034,In_1056);
nor U2163 (N_2163,In_314,In_1310);
and U2164 (N_2164,In_323,In_140);
or U2165 (N_2165,In_1112,In_213);
nand U2166 (N_2166,In_176,In_641);
or U2167 (N_2167,In_9,In_502);
nor U2168 (N_2168,In_932,In_191);
and U2169 (N_2169,In_930,In_549);
nor U2170 (N_2170,In_1070,In_1228);
and U2171 (N_2171,In_16,In_973);
nor U2172 (N_2172,In_593,In_598);
or U2173 (N_2173,In_222,In_121);
nor U2174 (N_2174,In_40,In_107);
and U2175 (N_2175,In_1171,In_482);
nor U2176 (N_2176,In_137,In_154);
and U2177 (N_2177,In_322,In_1117);
nand U2178 (N_2178,In_443,In_786);
and U2179 (N_2179,In_262,In_813);
nor U2180 (N_2180,In_806,In_566);
nand U2181 (N_2181,In_1472,In_961);
xnor U2182 (N_2182,In_207,In_710);
nand U2183 (N_2183,In_849,In_142);
or U2184 (N_2184,In_27,In_377);
nor U2185 (N_2185,In_454,In_1046);
or U2186 (N_2186,In_1321,In_1100);
nand U2187 (N_2187,In_1102,In_848);
nand U2188 (N_2188,In_419,In_1343);
or U2189 (N_2189,In_709,In_223);
nor U2190 (N_2190,In_886,In_347);
and U2191 (N_2191,In_609,In_1415);
and U2192 (N_2192,In_1424,In_1330);
nor U2193 (N_2193,In_1439,In_1130);
nand U2194 (N_2194,In_383,In_473);
nand U2195 (N_2195,In_1183,In_1310);
or U2196 (N_2196,In_1397,In_1470);
nor U2197 (N_2197,In_212,In_1257);
or U2198 (N_2198,In_477,In_384);
nand U2199 (N_2199,In_485,In_820);
and U2200 (N_2200,In_582,In_473);
nor U2201 (N_2201,In_1115,In_20);
and U2202 (N_2202,In_180,In_774);
and U2203 (N_2203,In_1216,In_1430);
or U2204 (N_2204,In_417,In_1391);
and U2205 (N_2205,In_930,In_619);
or U2206 (N_2206,In_104,In_1175);
nor U2207 (N_2207,In_318,In_1293);
and U2208 (N_2208,In_1197,In_338);
nor U2209 (N_2209,In_1451,In_1489);
nand U2210 (N_2210,In_1353,In_350);
and U2211 (N_2211,In_231,In_422);
xor U2212 (N_2212,In_659,In_1415);
nand U2213 (N_2213,In_746,In_1070);
nand U2214 (N_2214,In_703,In_1392);
nor U2215 (N_2215,In_1093,In_252);
or U2216 (N_2216,In_433,In_21);
and U2217 (N_2217,In_244,In_1270);
and U2218 (N_2218,In_928,In_546);
nor U2219 (N_2219,In_1254,In_325);
or U2220 (N_2220,In_641,In_596);
nor U2221 (N_2221,In_1429,In_703);
or U2222 (N_2222,In_1306,In_411);
and U2223 (N_2223,In_128,In_769);
nand U2224 (N_2224,In_299,In_333);
nand U2225 (N_2225,In_475,In_1164);
nand U2226 (N_2226,In_824,In_384);
nor U2227 (N_2227,In_974,In_588);
nor U2228 (N_2228,In_495,In_553);
or U2229 (N_2229,In_181,In_916);
or U2230 (N_2230,In_1229,In_717);
and U2231 (N_2231,In_363,In_1170);
nand U2232 (N_2232,In_907,In_233);
nand U2233 (N_2233,In_960,In_381);
nand U2234 (N_2234,In_1444,In_1288);
and U2235 (N_2235,In_1068,In_1000);
nor U2236 (N_2236,In_1260,In_251);
and U2237 (N_2237,In_1180,In_712);
or U2238 (N_2238,In_777,In_1027);
or U2239 (N_2239,In_1449,In_1140);
nand U2240 (N_2240,In_130,In_49);
and U2241 (N_2241,In_1269,In_1483);
or U2242 (N_2242,In_781,In_150);
nand U2243 (N_2243,In_153,In_970);
nand U2244 (N_2244,In_793,In_144);
and U2245 (N_2245,In_1186,In_851);
and U2246 (N_2246,In_1417,In_62);
nor U2247 (N_2247,In_620,In_351);
or U2248 (N_2248,In_1003,In_379);
or U2249 (N_2249,In_1366,In_150);
nor U2250 (N_2250,In_379,In_480);
nand U2251 (N_2251,In_471,In_895);
and U2252 (N_2252,In_175,In_1269);
nand U2253 (N_2253,In_680,In_1251);
nor U2254 (N_2254,In_184,In_788);
nand U2255 (N_2255,In_912,In_1060);
xor U2256 (N_2256,In_608,In_619);
and U2257 (N_2257,In_611,In_1247);
nand U2258 (N_2258,In_1464,In_851);
or U2259 (N_2259,In_504,In_841);
or U2260 (N_2260,In_1330,In_1036);
nor U2261 (N_2261,In_29,In_826);
nand U2262 (N_2262,In_875,In_1193);
nor U2263 (N_2263,In_1375,In_994);
or U2264 (N_2264,In_250,In_279);
or U2265 (N_2265,In_653,In_75);
nor U2266 (N_2266,In_231,In_360);
and U2267 (N_2267,In_786,In_1369);
or U2268 (N_2268,In_1469,In_771);
or U2269 (N_2269,In_871,In_370);
nand U2270 (N_2270,In_532,In_375);
and U2271 (N_2271,In_5,In_79);
nor U2272 (N_2272,In_1417,In_44);
nor U2273 (N_2273,In_550,In_1022);
and U2274 (N_2274,In_1114,In_1368);
or U2275 (N_2275,In_1036,In_946);
nand U2276 (N_2276,In_1042,In_514);
or U2277 (N_2277,In_709,In_1265);
or U2278 (N_2278,In_632,In_563);
nor U2279 (N_2279,In_708,In_704);
nor U2280 (N_2280,In_68,In_614);
nor U2281 (N_2281,In_1283,In_1084);
and U2282 (N_2282,In_393,In_1251);
nor U2283 (N_2283,In_219,In_1442);
nand U2284 (N_2284,In_415,In_562);
or U2285 (N_2285,In_59,In_870);
nand U2286 (N_2286,In_757,In_1025);
or U2287 (N_2287,In_488,In_471);
or U2288 (N_2288,In_785,In_507);
nand U2289 (N_2289,In_1349,In_1234);
and U2290 (N_2290,In_275,In_611);
nand U2291 (N_2291,In_1074,In_828);
nand U2292 (N_2292,In_1298,In_990);
nand U2293 (N_2293,In_1418,In_671);
and U2294 (N_2294,In_832,In_169);
nand U2295 (N_2295,In_462,In_598);
nand U2296 (N_2296,In_1081,In_1175);
and U2297 (N_2297,In_316,In_973);
and U2298 (N_2298,In_340,In_155);
nor U2299 (N_2299,In_1188,In_859);
nor U2300 (N_2300,In_844,In_803);
or U2301 (N_2301,In_1110,In_506);
or U2302 (N_2302,In_1167,In_629);
or U2303 (N_2303,In_1021,In_971);
nand U2304 (N_2304,In_1036,In_200);
and U2305 (N_2305,In_770,In_1258);
nand U2306 (N_2306,In_1128,In_737);
and U2307 (N_2307,In_48,In_545);
and U2308 (N_2308,In_967,In_1064);
and U2309 (N_2309,In_1491,In_589);
or U2310 (N_2310,In_691,In_1044);
and U2311 (N_2311,In_85,In_1452);
nand U2312 (N_2312,In_685,In_461);
and U2313 (N_2313,In_9,In_1267);
nand U2314 (N_2314,In_1334,In_398);
nand U2315 (N_2315,In_415,In_1331);
nor U2316 (N_2316,In_380,In_226);
nor U2317 (N_2317,In_425,In_1303);
or U2318 (N_2318,In_1036,In_984);
and U2319 (N_2319,In_1369,In_772);
nand U2320 (N_2320,In_1408,In_522);
nand U2321 (N_2321,In_1356,In_1310);
nor U2322 (N_2322,In_337,In_417);
nor U2323 (N_2323,In_638,In_887);
nand U2324 (N_2324,In_177,In_168);
and U2325 (N_2325,In_1276,In_112);
nand U2326 (N_2326,In_560,In_328);
nand U2327 (N_2327,In_646,In_1086);
nor U2328 (N_2328,In_1354,In_1301);
and U2329 (N_2329,In_1074,In_1449);
or U2330 (N_2330,In_232,In_1480);
nand U2331 (N_2331,In_69,In_1002);
or U2332 (N_2332,In_676,In_793);
and U2333 (N_2333,In_40,In_1489);
nor U2334 (N_2334,In_428,In_121);
or U2335 (N_2335,In_479,In_787);
or U2336 (N_2336,In_1159,In_418);
or U2337 (N_2337,In_382,In_226);
or U2338 (N_2338,In_620,In_360);
or U2339 (N_2339,In_254,In_843);
nor U2340 (N_2340,In_1302,In_491);
nor U2341 (N_2341,In_1235,In_1461);
or U2342 (N_2342,In_641,In_797);
nor U2343 (N_2343,In_373,In_898);
nor U2344 (N_2344,In_1051,In_591);
and U2345 (N_2345,In_845,In_1186);
and U2346 (N_2346,In_1013,In_81);
and U2347 (N_2347,In_1122,In_557);
nor U2348 (N_2348,In_572,In_379);
nand U2349 (N_2349,In_27,In_531);
and U2350 (N_2350,In_929,In_754);
nand U2351 (N_2351,In_184,In_1299);
nand U2352 (N_2352,In_652,In_1482);
or U2353 (N_2353,In_374,In_217);
or U2354 (N_2354,In_166,In_1155);
or U2355 (N_2355,In_456,In_214);
nor U2356 (N_2356,In_879,In_138);
nor U2357 (N_2357,In_361,In_1086);
nand U2358 (N_2358,In_1400,In_1393);
nor U2359 (N_2359,In_1375,In_1101);
or U2360 (N_2360,In_1396,In_1106);
or U2361 (N_2361,In_791,In_450);
or U2362 (N_2362,In_609,In_1005);
nor U2363 (N_2363,In_1050,In_399);
and U2364 (N_2364,In_1467,In_273);
nor U2365 (N_2365,In_1201,In_283);
or U2366 (N_2366,In_1412,In_267);
nand U2367 (N_2367,In_1209,In_789);
nor U2368 (N_2368,In_142,In_814);
and U2369 (N_2369,In_903,In_971);
or U2370 (N_2370,In_1064,In_386);
nor U2371 (N_2371,In_89,In_584);
and U2372 (N_2372,In_1107,In_252);
nand U2373 (N_2373,In_1125,In_471);
and U2374 (N_2374,In_399,In_612);
nand U2375 (N_2375,In_1304,In_216);
or U2376 (N_2376,In_641,In_694);
nor U2377 (N_2377,In_698,In_961);
nand U2378 (N_2378,In_784,In_1087);
xnor U2379 (N_2379,In_156,In_943);
or U2380 (N_2380,In_1224,In_559);
and U2381 (N_2381,In_1020,In_977);
or U2382 (N_2382,In_1243,In_1330);
nor U2383 (N_2383,In_248,In_587);
nor U2384 (N_2384,In_446,In_616);
nor U2385 (N_2385,In_1306,In_241);
nor U2386 (N_2386,In_1021,In_57);
or U2387 (N_2387,In_223,In_1233);
nor U2388 (N_2388,In_110,In_236);
or U2389 (N_2389,In_741,In_200);
nand U2390 (N_2390,In_80,In_780);
nor U2391 (N_2391,In_748,In_534);
and U2392 (N_2392,In_832,In_713);
or U2393 (N_2393,In_1350,In_1200);
nand U2394 (N_2394,In_261,In_1007);
nand U2395 (N_2395,In_880,In_270);
nand U2396 (N_2396,In_1014,In_1311);
nand U2397 (N_2397,In_454,In_199);
or U2398 (N_2398,In_5,In_1305);
nor U2399 (N_2399,In_453,In_411);
and U2400 (N_2400,In_149,In_1028);
and U2401 (N_2401,In_1135,In_1195);
or U2402 (N_2402,In_29,In_107);
nand U2403 (N_2403,In_606,In_1140);
or U2404 (N_2404,In_272,In_1187);
nand U2405 (N_2405,In_1074,In_1300);
nand U2406 (N_2406,In_1204,In_901);
nand U2407 (N_2407,In_660,In_510);
nor U2408 (N_2408,In_1323,In_257);
or U2409 (N_2409,In_1212,In_1408);
or U2410 (N_2410,In_1104,In_89);
xor U2411 (N_2411,In_425,In_1118);
and U2412 (N_2412,In_328,In_1408);
nand U2413 (N_2413,In_220,In_377);
or U2414 (N_2414,In_638,In_781);
and U2415 (N_2415,In_702,In_160);
and U2416 (N_2416,In_238,In_171);
nand U2417 (N_2417,In_83,In_153);
or U2418 (N_2418,In_1385,In_348);
or U2419 (N_2419,In_1487,In_516);
and U2420 (N_2420,In_81,In_1299);
and U2421 (N_2421,In_982,In_130);
nand U2422 (N_2422,In_998,In_1364);
nor U2423 (N_2423,In_1393,In_494);
nand U2424 (N_2424,In_1285,In_336);
or U2425 (N_2425,In_105,In_52);
nand U2426 (N_2426,In_1352,In_1163);
nand U2427 (N_2427,In_5,In_1341);
nand U2428 (N_2428,In_480,In_1328);
or U2429 (N_2429,In_524,In_116);
and U2430 (N_2430,In_568,In_1135);
nand U2431 (N_2431,In_411,In_989);
and U2432 (N_2432,In_1166,In_1025);
nor U2433 (N_2433,In_107,In_50);
and U2434 (N_2434,In_192,In_526);
xnor U2435 (N_2435,In_448,In_565);
and U2436 (N_2436,In_563,In_900);
or U2437 (N_2437,In_1392,In_1318);
nor U2438 (N_2438,In_1483,In_682);
and U2439 (N_2439,In_23,In_1389);
or U2440 (N_2440,In_1064,In_522);
nand U2441 (N_2441,In_1377,In_239);
nor U2442 (N_2442,In_725,In_1024);
nor U2443 (N_2443,In_839,In_878);
and U2444 (N_2444,In_989,In_366);
nand U2445 (N_2445,In_1405,In_317);
or U2446 (N_2446,In_1116,In_14);
or U2447 (N_2447,In_150,In_789);
nor U2448 (N_2448,In_645,In_1178);
nand U2449 (N_2449,In_1155,In_884);
or U2450 (N_2450,In_872,In_1056);
nand U2451 (N_2451,In_358,In_953);
nor U2452 (N_2452,In_266,In_187);
nor U2453 (N_2453,In_1478,In_727);
nor U2454 (N_2454,In_913,In_458);
nand U2455 (N_2455,In_418,In_1443);
and U2456 (N_2456,In_1453,In_1153);
nand U2457 (N_2457,In_206,In_694);
and U2458 (N_2458,In_407,In_1165);
or U2459 (N_2459,In_1130,In_1112);
nor U2460 (N_2460,In_951,In_1034);
and U2461 (N_2461,In_582,In_704);
nand U2462 (N_2462,In_1040,In_427);
xnor U2463 (N_2463,In_1028,In_696);
nor U2464 (N_2464,In_91,In_397);
nand U2465 (N_2465,In_952,In_60);
and U2466 (N_2466,In_1322,In_647);
nor U2467 (N_2467,In_1328,In_1378);
nor U2468 (N_2468,In_1274,In_1129);
nand U2469 (N_2469,In_1325,In_35);
or U2470 (N_2470,In_684,In_204);
nand U2471 (N_2471,In_965,In_995);
nand U2472 (N_2472,In_47,In_161);
nor U2473 (N_2473,In_899,In_980);
xnor U2474 (N_2474,In_1350,In_596);
and U2475 (N_2475,In_123,In_288);
and U2476 (N_2476,In_268,In_1367);
nor U2477 (N_2477,In_1324,In_807);
and U2478 (N_2478,In_1447,In_50);
nand U2479 (N_2479,In_153,In_333);
nor U2480 (N_2480,In_700,In_1401);
and U2481 (N_2481,In_479,In_39);
nor U2482 (N_2482,In_471,In_44);
nand U2483 (N_2483,In_454,In_1283);
or U2484 (N_2484,In_659,In_8);
nor U2485 (N_2485,In_1475,In_318);
nand U2486 (N_2486,In_906,In_1311);
or U2487 (N_2487,In_622,In_852);
and U2488 (N_2488,In_475,In_213);
nand U2489 (N_2489,In_1214,In_1019);
nor U2490 (N_2490,In_982,In_690);
nand U2491 (N_2491,In_385,In_0);
nor U2492 (N_2492,In_689,In_1400);
nand U2493 (N_2493,In_1206,In_1373);
nor U2494 (N_2494,In_484,In_1354);
xor U2495 (N_2495,In_1348,In_439);
nand U2496 (N_2496,In_1121,In_1183);
nand U2497 (N_2497,In_1254,In_196);
and U2498 (N_2498,In_783,In_120);
nand U2499 (N_2499,In_155,In_894);
or U2500 (N_2500,In_643,In_540);
xor U2501 (N_2501,In_1191,In_1241);
nor U2502 (N_2502,In_406,In_131);
nand U2503 (N_2503,In_57,In_376);
nand U2504 (N_2504,In_1002,In_995);
nor U2505 (N_2505,In_1027,In_739);
or U2506 (N_2506,In_1213,In_539);
and U2507 (N_2507,In_593,In_1493);
nand U2508 (N_2508,In_476,In_287);
and U2509 (N_2509,In_715,In_1320);
nand U2510 (N_2510,In_437,In_1251);
nor U2511 (N_2511,In_625,In_1024);
nand U2512 (N_2512,In_574,In_1348);
nor U2513 (N_2513,In_1461,In_337);
nor U2514 (N_2514,In_1048,In_377);
or U2515 (N_2515,In_174,In_404);
or U2516 (N_2516,In_545,In_1408);
and U2517 (N_2517,In_942,In_866);
nor U2518 (N_2518,In_318,In_183);
nand U2519 (N_2519,In_638,In_1194);
or U2520 (N_2520,In_451,In_195);
or U2521 (N_2521,In_714,In_608);
and U2522 (N_2522,In_1026,In_1285);
or U2523 (N_2523,In_1121,In_459);
nand U2524 (N_2524,In_595,In_35);
nand U2525 (N_2525,In_1013,In_123);
nand U2526 (N_2526,In_1168,In_1011);
nand U2527 (N_2527,In_453,In_851);
nand U2528 (N_2528,In_394,In_875);
and U2529 (N_2529,In_590,In_332);
nor U2530 (N_2530,In_257,In_1382);
or U2531 (N_2531,In_1467,In_1303);
nor U2532 (N_2532,In_62,In_187);
nor U2533 (N_2533,In_625,In_1230);
or U2534 (N_2534,In_18,In_1123);
nand U2535 (N_2535,In_704,In_881);
and U2536 (N_2536,In_762,In_1241);
and U2537 (N_2537,In_271,In_355);
or U2538 (N_2538,In_1022,In_614);
nor U2539 (N_2539,In_807,In_528);
nand U2540 (N_2540,In_1009,In_663);
or U2541 (N_2541,In_877,In_822);
and U2542 (N_2542,In_1251,In_341);
nand U2543 (N_2543,In_1296,In_406);
and U2544 (N_2544,In_1070,In_1308);
and U2545 (N_2545,In_173,In_516);
and U2546 (N_2546,In_223,In_309);
and U2547 (N_2547,In_123,In_487);
nand U2548 (N_2548,In_1134,In_749);
and U2549 (N_2549,In_1101,In_939);
nor U2550 (N_2550,In_273,In_794);
or U2551 (N_2551,In_90,In_1392);
or U2552 (N_2552,In_433,In_1287);
and U2553 (N_2553,In_1103,In_13);
or U2554 (N_2554,In_1204,In_54);
and U2555 (N_2555,In_854,In_491);
nand U2556 (N_2556,In_1217,In_961);
nand U2557 (N_2557,In_1051,In_25);
nand U2558 (N_2558,In_861,In_412);
and U2559 (N_2559,In_637,In_1209);
or U2560 (N_2560,In_690,In_1081);
or U2561 (N_2561,In_1241,In_141);
nor U2562 (N_2562,In_729,In_682);
nor U2563 (N_2563,In_42,In_987);
nor U2564 (N_2564,In_1274,In_530);
and U2565 (N_2565,In_86,In_795);
nor U2566 (N_2566,In_615,In_1498);
or U2567 (N_2567,In_1328,In_727);
nor U2568 (N_2568,In_1480,In_1211);
and U2569 (N_2569,In_1352,In_1345);
and U2570 (N_2570,In_53,In_750);
nor U2571 (N_2571,In_577,In_1496);
or U2572 (N_2572,In_989,In_730);
or U2573 (N_2573,In_1272,In_1440);
nand U2574 (N_2574,In_1300,In_631);
or U2575 (N_2575,In_951,In_233);
nor U2576 (N_2576,In_1084,In_1338);
nor U2577 (N_2577,In_214,In_1089);
or U2578 (N_2578,In_923,In_477);
or U2579 (N_2579,In_760,In_306);
or U2580 (N_2580,In_271,In_964);
nor U2581 (N_2581,In_1371,In_587);
nand U2582 (N_2582,In_817,In_1);
nand U2583 (N_2583,In_630,In_1005);
nor U2584 (N_2584,In_1379,In_413);
and U2585 (N_2585,In_78,In_1452);
and U2586 (N_2586,In_926,In_1008);
or U2587 (N_2587,In_714,In_848);
and U2588 (N_2588,In_973,In_499);
nor U2589 (N_2589,In_298,In_16);
nor U2590 (N_2590,In_1311,In_104);
nor U2591 (N_2591,In_757,In_352);
or U2592 (N_2592,In_763,In_46);
or U2593 (N_2593,In_681,In_984);
nor U2594 (N_2594,In_144,In_713);
nand U2595 (N_2595,In_877,In_888);
or U2596 (N_2596,In_1211,In_355);
or U2597 (N_2597,In_854,In_552);
nand U2598 (N_2598,In_81,In_205);
and U2599 (N_2599,In_707,In_117);
nor U2600 (N_2600,In_649,In_1263);
and U2601 (N_2601,In_369,In_445);
nand U2602 (N_2602,In_150,In_760);
and U2603 (N_2603,In_499,In_1222);
nand U2604 (N_2604,In_41,In_920);
and U2605 (N_2605,In_484,In_532);
or U2606 (N_2606,In_877,In_589);
nor U2607 (N_2607,In_1253,In_765);
or U2608 (N_2608,In_755,In_95);
and U2609 (N_2609,In_1460,In_898);
or U2610 (N_2610,In_714,In_325);
nand U2611 (N_2611,In_84,In_1069);
and U2612 (N_2612,In_476,In_892);
nand U2613 (N_2613,In_382,In_66);
nor U2614 (N_2614,In_1278,In_1);
and U2615 (N_2615,In_562,In_1373);
or U2616 (N_2616,In_738,In_901);
nor U2617 (N_2617,In_1460,In_672);
or U2618 (N_2618,In_859,In_475);
nor U2619 (N_2619,In_365,In_537);
or U2620 (N_2620,In_1381,In_1446);
nor U2621 (N_2621,In_1199,In_385);
nor U2622 (N_2622,In_1471,In_77);
nand U2623 (N_2623,In_340,In_928);
nand U2624 (N_2624,In_399,In_1288);
or U2625 (N_2625,In_584,In_714);
or U2626 (N_2626,In_99,In_1391);
nand U2627 (N_2627,In_1496,In_254);
nand U2628 (N_2628,In_497,In_1431);
or U2629 (N_2629,In_913,In_795);
nor U2630 (N_2630,In_193,In_820);
nand U2631 (N_2631,In_1263,In_1364);
and U2632 (N_2632,In_445,In_855);
and U2633 (N_2633,In_1238,In_29);
nor U2634 (N_2634,In_330,In_853);
or U2635 (N_2635,In_679,In_1375);
nor U2636 (N_2636,In_762,In_1259);
nor U2637 (N_2637,In_1416,In_1129);
nand U2638 (N_2638,In_1499,In_218);
or U2639 (N_2639,In_806,In_757);
or U2640 (N_2640,In_480,In_420);
and U2641 (N_2641,In_818,In_1288);
and U2642 (N_2642,In_276,In_376);
nor U2643 (N_2643,In_563,In_1003);
nor U2644 (N_2644,In_848,In_978);
and U2645 (N_2645,In_59,In_1095);
nor U2646 (N_2646,In_1445,In_174);
nand U2647 (N_2647,In_81,In_1233);
and U2648 (N_2648,In_892,In_1295);
and U2649 (N_2649,In_1085,In_120);
nor U2650 (N_2650,In_144,In_351);
nor U2651 (N_2651,In_1050,In_250);
and U2652 (N_2652,In_535,In_136);
or U2653 (N_2653,In_562,In_224);
or U2654 (N_2654,In_614,In_100);
and U2655 (N_2655,In_1211,In_1262);
nor U2656 (N_2656,In_982,In_43);
or U2657 (N_2657,In_1063,In_707);
nand U2658 (N_2658,In_27,In_1294);
nand U2659 (N_2659,In_1493,In_545);
and U2660 (N_2660,In_1153,In_171);
and U2661 (N_2661,In_29,In_863);
nand U2662 (N_2662,In_817,In_1078);
nor U2663 (N_2663,In_1116,In_224);
or U2664 (N_2664,In_1075,In_1330);
or U2665 (N_2665,In_294,In_1162);
nand U2666 (N_2666,In_1005,In_1437);
and U2667 (N_2667,In_702,In_1180);
nor U2668 (N_2668,In_1342,In_1443);
nor U2669 (N_2669,In_980,In_310);
nand U2670 (N_2670,In_306,In_921);
nor U2671 (N_2671,In_1479,In_88);
nand U2672 (N_2672,In_716,In_1289);
or U2673 (N_2673,In_951,In_618);
nand U2674 (N_2674,In_647,In_451);
or U2675 (N_2675,In_1373,In_606);
nand U2676 (N_2676,In_629,In_485);
or U2677 (N_2677,In_965,In_99);
or U2678 (N_2678,In_250,In_409);
nor U2679 (N_2679,In_688,In_423);
and U2680 (N_2680,In_872,In_385);
and U2681 (N_2681,In_860,In_62);
and U2682 (N_2682,In_934,In_338);
nand U2683 (N_2683,In_272,In_416);
xor U2684 (N_2684,In_1031,In_436);
nor U2685 (N_2685,In_800,In_756);
nand U2686 (N_2686,In_68,In_99);
nand U2687 (N_2687,In_1161,In_1016);
nor U2688 (N_2688,In_659,In_519);
nand U2689 (N_2689,In_559,In_202);
nor U2690 (N_2690,In_1451,In_912);
nand U2691 (N_2691,In_1235,In_704);
and U2692 (N_2692,In_182,In_590);
xor U2693 (N_2693,In_989,In_1095);
or U2694 (N_2694,In_1359,In_323);
and U2695 (N_2695,In_1084,In_153);
nand U2696 (N_2696,In_107,In_358);
nand U2697 (N_2697,In_309,In_1232);
nand U2698 (N_2698,In_1057,In_639);
or U2699 (N_2699,In_1467,In_1438);
nand U2700 (N_2700,In_41,In_54);
or U2701 (N_2701,In_1301,In_774);
and U2702 (N_2702,In_132,In_1265);
nand U2703 (N_2703,In_619,In_252);
nand U2704 (N_2704,In_1066,In_1028);
nor U2705 (N_2705,In_687,In_930);
and U2706 (N_2706,In_911,In_543);
and U2707 (N_2707,In_1275,In_276);
nand U2708 (N_2708,In_1305,In_633);
and U2709 (N_2709,In_37,In_469);
nand U2710 (N_2710,In_39,In_752);
nand U2711 (N_2711,In_1482,In_1463);
or U2712 (N_2712,In_1218,In_339);
or U2713 (N_2713,In_259,In_1436);
nand U2714 (N_2714,In_1212,In_73);
xnor U2715 (N_2715,In_1343,In_710);
nor U2716 (N_2716,In_1169,In_422);
nand U2717 (N_2717,In_1353,In_624);
nor U2718 (N_2718,In_548,In_84);
and U2719 (N_2719,In_1260,In_1348);
or U2720 (N_2720,In_1426,In_647);
nand U2721 (N_2721,In_1386,In_101);
or U2722 (N_2722,In_1191,In_1316);
nor U2723 (N_2723,In_1365,In_144);
nand U2724 (N_2724,In_225,In_981);
nor U2725 (N_2725,In_1089,In_335);
and U2726 (N_2726,In_1239,In_592);
nor U2727 (N_2727,In_816,In_633);
and U2728 (N_2728,In_1366,In_693);
or U2729 (N_2729,In_726,In_1094);
and U2730 (N_2730,In_1461,In_1146);
and U2731 (N_2731,In_761,In_615);
and U2732 (N_2732,In_976,In_20);
or U2733 (N_2733,In_1098,In_223);
and U2734 (N_2734,In_1368,In_150);
nor U2735 (N_2735,In_405,In_965);
nand U2736 (N_2736,In_539,In_1441);
or U2737 (N_2737,In_159,In_801);
nand U2738 (N_2738,In_1354,In_43);
nor U2739 (N_2739,In_15,In_887);
nand U2740 (N_2740,In_116,In_158);
nor U2741 (N_2741,In_206,In_193);
nand U2742 (N_2742,In_659,In_976);
or U2743 (N_2743,In_405,In_1173);
and U2744 (N_2744,In_1253,In_722);
nor U2745 (N_2745,In_590,In_665);
nor U2746 (N_2746,In_583,In_407);
or U2747 (N_2747,In_1235,In_1125);
or U2748 (N_2748,In_1230,In_1202);
xor U2749 (N_2749,In_1174,In_577);
and U2750 (N_2750,In_615,In_1125);
nand U2751 (N_2751,In_323,In_934);
nand U2752 (N_2752,In_1320,In_1185);
nand U2753 (N_2753,In_1460,In_240);
nand U2754 (N_2754,In_1290,In_1127);
and U2755 (N_2755,In_855,In_295);
or U2756 (N_2756,In_944,In_1312);
nor U2757 (N_2757,In_1094,In_504);
nand U2758 (N_2758,In_22,In_274);
nor U2759 (N_2759,In_186,In_173);
nor U2760 (N_2760,In_775,In_140);
or U2761 (N_2761,In_428,In_1151);
nor U2762 (N_2762,In_663,In_71);
or U2763 (N_2763,In_529,In_600);
or U2764 (N_2764,In_994,In_267);
and U2765 (N_2765,In_191,In_1434);
nor U2766 (N_2766,In_984,In_1143);
or U2767 (N_2767,In_1064,In_719);
or U2768 (N_2768,In_573,In_33);
or U2769 (N_2769,In_824,In_1118);
nor U2770 (N_2770,In_53,In_292);
nor U2771 (N_2771,In_1474,In_391);
nor U2772 (N_2772,In_65,In_837);
nor U2773 (N_2773,In_372,In_379);
or U2774 (N_2774,In_464,In_1202);
nor U2775 (N_2775,In_935,In_1232);
nand U2776 (N_2776,In_170,In_382);
nand U2777 (N_2777,In_473,In_805);
and U2778 (N_2778,In_999,In_932);
and U2779 (N_2779,In_187,In_149);
nor U2780 (N_2780,In_939,In_571);
or U2781 (N_2781,In_1495,In_849);
and U2782 (N_2782,In_684,In_1485);
nand U2783 (N_2783,In_834,In_784);
and U2784 (N_2784,In_709,In_1323);
nor U2785 (N_2785,In_1378,In_697);
nand U2786 (N_2786,In_1377,In_1472);
nor U2787 (N_2787,In_277,In_1335);
nand U2788 (N_2788,In_718,In_492);
nor U2789 (N_2789,In_376,In_993);
nand U2790 (N_2790,In_980,In_1097);
nor U2791 (N_2791,In_960,In_1047);
nand U2792 (N_2792,In_884,In_273);
or U2793 (N_2793,In_334,In_875);
nand U2794 (N_2794,In_778,In_554);
nand U2795 (N_2795,In_970,In_294);
nor U2796 (N_2796,In_1374,In_931);
nand U2797 (N_2797,In_9,In_1159);
nand U2798 (N_2798,In_837,In_1429);
nor U2799 (N_2799,In_738,In_438);
or U2800 (N_2800,In_588,In_501);
nor U2801 (N_2801,In_1442,In_1383);
nand U2802 (N_2802,In_1398,In_1089);
and U2803 (N_2803,In_377,In_1224);
nand U2804 (N_2804,In_1296,In_50);
nor U2805 (N_2805,In_73,In_1463);
and U2806 (N_2806,In_152,In_1156);
nor U2807 (N_2807,In_113,In_1348);
and U2808 (N_2808,In_753,In_1070);
nand U2809 (N_2809,In_891,In_586);
nor U2810 (N_2810,In_655,In_1396);
or U2811 (N_2811,In_570,In_1493);
or U2812 (N_2812,In_93,In_1237);
nand U2813 (N_2813,In_45,In_1377);
nand U2814 (N_2814,In_1272,In_1308);
nand U2815 (N_2815,In_1350,In_433);
nor U2816 (N_2816,In_374,In_250);
nand U2817 (N_2817,In_564,In_1492);
nor U2818 (N_2818,In_1421,In_1038);
and U2819 (N_2819,In_637,In_1263);
nor U2820 (N_2820,In_108,In_632);
nor U2821 (N_2821,In_61,In_779);
nand U2822 (N_2822,In_324,In_971);
and U2823 (N_2823,In_310,In_922);
nor U2824 (N_2824,In_580,In_1466);
nand U2825 (N_2825,In_333,In_524);
nor U2826 (N_2826,In_41,In_1405);
and U2827 (N_2827,In_459,In_871);
or U2828 (N_2828,In_396,In_108);
nand U2829 (N_2829,In_1301,In_1427);
and U2830 (N_2830,In_1346,In_164);
and U2831 (N_2831,In_1230,In_199);
or U2832 (N_2832,In_747,In_1268);
and U2833 (N_2833,In_534,In_844);
and U2834 (N_2834,In_1021,In_533);
nor U2835 (N_2835,In_790,In_1030);
or U2836 (N_2836,In_583,In_862);
and U2837 (N_2837,In_745,In_343);
or U2838 (N_2838,In_1182,In_369);
or U2839 (N_2839,In_1068,In_468);
nand U2840 (N_2840,In_290,In_1302);
nand U2841 (N_2841,In_893,In_491);
nor U2842 (N_2842,In_1071,In_108);
and U2843 (N_2843,In_345,In_338);
and U2844 (N_2844,In_653,In_1418);
or U2845 (N_2845,In_545,In_110);
nand U2846 (N_2846,In_819,In_1205);
or U2847 (N_2847,In_944,In_258);
nand U2848 (N_2848,In_900,In_1138);
or U2849 (N_2849,In_293,In_339);
and U2850 (N_2850,In_2,In_23);
nor U2851 (N_2851,In_1098,In_899);
nor U2852 (N_2852,In_1443,In_519);
nor U2853 (N_2853,In_393,In_730);
nand U2854 (N_2854,In_1124,In_664);
nor U2855 (N_2855,In_1336,In_798);
or U2856 (N_2856,In_534,In_257);
and U2857 (N_2857,In_1279,In_544);
and U2858 (N_2858,In_1434,In_713);
nand U2859 (N_2859,In_481,In_80);
nand U2860 (N_2860,In_698,In_537);
nand U2861 (N_2861,In_1153,In_1244);
and U2862 (N_2862,In_136,In_1163);
and U2863 (N_2863,In_387,In_512);
or U2864 (N_2864,In_577,In_923);
nor U2865 (N_2865,In_1101,In_1034);
or U2866 (N_2866,In_1019,In_1120);
and U2867 (N_2867,In_1052,In_771);
nor U2868 (N_2868,In_505,In_601);
or U2869 (N_2869,In_896,In_201);
or U2870 (N_2870,In_973,In_888);
and U2871 (N_2871,In_1183,In_312);
and U2872 (N_2872,In_236,In_455);
or U2873 (N_2873,In_1178,In_1012);
nor U2874 (N_2874,In_125,In_510);
and U2875 (N_2875,In_289,In_32);
nand U2876 (N_2876,In_1056,In_790);
and U2877 (N_2877,In_258,In_767);
nand U2878 (N_2878,In_563,In_503);
nand U2879 (N_2879,In_528,In_1313);
nand U2880 (N_2880,In_34,In_161);
nand U2881 (N_2881,In_789,In_985);
nor U2882 (N_2882,In_1171,In_1064);
nand U2883 (N_2883,In_90,In_421);
and U2884 (N_2884,In_1279,In_824);
nand U2885 (N_2885,In_1465,In_797);
nor U2886 (N_2886,In_155,In_1201);
and U2887 (N_2887,In_1221,In_838);
nand U2888 (N_2888,In_1406,In_482);
and U2889 (N_2889,In_271,In_1027);
nand U2890 (N_2890,In_1296,In_932);
nor U2891 (N_2891,In_1014,In_740);
nand U2892 (N_2892,In_897,In_575);
nor U2893 (N_2893,In_1245,In_808);
and U2894 (N_2894,In_1157,In_826);
and U2895 (N_2895,In_1,In_700);
nor U2896 (N_2896,In_552,In_554);
nor U2897 (N_2897,In_988,In_449);
or U2898 (N_2898,In_878,In_637);
and U2899 (N_2899,In_1194,In_44);
nand U2900 (N_2900,In_119,In_259);
nor U2901 (N_2901,In_220,In_1385);
nor U2902 (N_2902,In_948,In_242);
and U2903 (N_2903,In_1366,In_142);
nand U2904 (N_2904,In_519,In_809);
nor U2905 (N_2905,In_146,In_448);
and U2906 (N_2906,In_1118,In_505);
or U2907 (N_2907,In_331,In_1368);
or U2908 (N_2908,In_366,In_643);
or U2909 (N_2909,In_1379,In_1030);
and U2910 (N_2910,In_260,In_522);
and U2911 (N_2911,In_841,In_189);
nor U2912 (N_2912,In_537,In_642);
nor U2913 (N_2913,In_1161,In_79);
or U2914 (N_2914,In_1029,In_404);
nand U2915 (N_2915,In_348,In_343);
or U2916 (N_2916,In_273,In_1411);
or U2917 (N_2917,In_602,In_1363);
nand U2918 (N_2918,In_1414,In_1157);
nor U2919 (N_2919,In_1097,In_1168);
nor U2920 (N_2920,In_1087,In_179);
or U2921 (N_2921,In_1200,In_827);
or U2922 (N_2922,In_198,In_652);
nor U2923 (N_2923,In_887,In_1375);
nor U2924 (N_2924,In_1450,In_576);
nor U2925 (N_2925,In_169,In_1332);
and U2926 (N_2926,In_704,In_1475);
nand U2927 (N_2927,In_80,In_1070);
and U2928 (N_2928,In_1388,In_767);
and U2929 (N_2929,In_421,In_1056);
nand U2930 (N_2930,In_344,In_1323);
and U2931 (N_2931,In_1235,In_0);
and U2932 (N_2932,In_937,In_1449);
or U2933 (N_2933,In_636,In_881);
nor U2934 (N_2934,In_769,In_420);
and U2935 (N_2935,In_547,In_463);
nor U2936 (N_2936,In_1214,In_1491);
nand U2937 (N_2937,In_511,In_887);
or U2938 (N_2938,In_318,In_533);
nor U2939 (N_2939,In_1086,In_1374);
nor U2940 (N_2940,In_1411,In_169);
nand U2941 (N_2941,In_1359,In_1125);
or U2942 (N_2942,In_813,In_1212);
or U2943 (N_2943,In_893,In_1328);
nor U2944 (N_2944,In_799,In_784);
and U2945 (N_2945,In_1304,In_1172);
nand U2946 (N_2946,In_234,In_628);
and U2947 (N_2947,In_930,In_81);
or U2948 (N_2948,In_404,In_888);
and U2949 (N_2949,In_661,In_675);
nor U2950 (N_2950,In_29,In_314);
nand U2951 (N_2951,In_814,In_1036);
nor U2952 (N_2952,In_271,In_942);
and U2953 (N_2953,In_291,In_490);
nor U2954 (N_2954,In_322,In_373);
and U2955 (N_2955,In_681,In_1204);
or U2956 (N_2956,In_753,In_330);
nand U2957 (N_2957,In_870,In_1341);
or U2958 (N_2958,In_1324,In_763);
nor U2959 (N_2959,In_885,In_262);
or U2960 (N_2960,In_331,In_1484);
or U2961 (N_2961,In_873,In_323);
nand U2962 (N_2962,In_633,In_209);
and U2963 (N_2963,In_368,In_45);
and U2964 (N_2964,In_414,In_948);
nand U2965 (N_2965,In_39,In_612);
and U2966 (N_2966,In_1184,In_1128);
and U2967 (N_2967,In_216,In_950);
nand U2968 (N_2968,In_1058,In_1436);
and U2969 (N_2969,In_1381,In_959);
or U2970 (N_2970,In_1135,In_442);
nor U2971 (N_2971,In_705,In_713);
or U2972 (N_2972,In_730,In_300);
nor U2973 (N_2973,In_46,In_251);
nand U2974 (N_2974,In_505,In_1347);
nand U2975 (N_2975,In_673,In_1354);
nand U2976 (N_2976,In_44,In_380);
and U2977 (N_2977,In_313,In_971);
nor U2978 (N_2978,In_574,In_1267);
nor U2979 (N_2979,In_723,In_99);
and U2980 (N_2980,In_1077,In_1388);
or U2981 (N_2981,In_1370,In_741);
or U2982 (N_2982,In_1146,In_596);
nor U2983 (N_2983,In_522,In_490);
or U2984 (N_2984,In_962,In_1477);
or U2985 (N_2985,In_1155,In_1098);
nor U2986 (N_2986,In_314,In_244);
nand U2987 (N_2987,In_999,In_529);
or U2988 (N_2988,In_25,In_338);
or U2989 (N_2989,In_1391,In_186);
or U2990 (N_2990,In_211,In_800);
nand U2991 (N_2991,In_1486,In_81);
nor U2992 (N_2992,In_1363,In_647);
or U2993 (N_2993,In_1054,In_1342);
and U2994 (N_2994,In_483,In_1416);
nand U2995 (N_2995,In_551,In_924);
nand U2996 (N_2996,In_117,In_750);
or U2997 (N_2997,In_1319,In_1393);
nand U2998 (N_2998,In_243,In_837);
nor U2999 (N_2999,In_454,In_1013);
and U3000 (N_3000,N_460,N_1415);
nand U3001 (N_3001,N_2392,N_1118);
and U3002 (N_3002,N_2778,N_1401);
and U3003 (N_3003,N_961,N_2021);
and U3004 (N_3004,N_639,N_2361);
or U3005 (N_3005,N_2044,N_516);
nand U3006 (N_3006,N_1352,N_1110);
nand U3007 (N_3007,N_329,N_503);
nor U3008 (N_3008,N_2360,N_395);
or U3009 (N_3009,N_2086,N_724);
nand U3010 (N_3010,N_349,N_2090);
nor U3011 (N_3011,N_167,N_1731);
and U3012 (N_3012,N_1987,N_12);
or U3013 (N_3013,N_2550,N_2559);
or U3014 (N_3014,N_376,N_975);
nand U3015 (N_3015,N_856,N_46);
and U3016 (N_3016,N_2137,N_1019);
nor U3017 (N_3017,N_345,N_1932);
nand U3018 (N_3018,N_325,N_1866);
nor U3019 (N_3019,N_2910,N_2930);
or U3020 (N_3020,N_2454,N_2878);
nor U3021 (N_3021,N_1641,N_176);
and U3022 (N_3022,N_1599,N_314);
and U3023 (N_3023,N_2192,N_923);
and U3024 (N_3024,N_1432,N_2885);
or U3025 (N_3025,N_1361,N_2453);
nand U3026 (N_3026,N_2526,N_508);
and U3027 (N_3027,N_1742,N_2490);
nor U3028 (N_3028,N_1616,N_2950);
or U3029 (N_3029,N_571,N_2436);
and U3030 (N_3030,N_773,N_1840);
or U3031 (N_3031,N_1714,N_201);
nand U3032 (N_3032,N_2790,N_792);
or U3033 (N_3033,N_755,N_788);
or U3034 (N_3034,N_2714,N_2398);
and U3035 (N_3035,N_1382,N_2025);
and U3036 (N_3036,N_860,N_0);
and U3037 (N_3037,N_1071,N_207);
and U3038 (N_3038,N_271,N_2040);
nand U3039 (N_3039,N_2418,N_1765);
nand U3040 (N_3040,N_2853,N_2792);
and U3041 (N_3041,N_946,N_1752);
or U3042 (N_3042,N_1972,N_631);
and U3043 (N_3043,N_132,N_1052);
nor U3044 (N_3044,N_2250,N_1409);
or U3045 (N_3045,N_763,N_184);
or U3046 (N_3046,N_1706,N_1702);
nand U3047 (N_3047,N_2095,N_2277);
or U3048 (N_3048,N_972,N_1903);
and U3049 (N_3049,N_509,N_1751);
nor U3050 (N_3050,N_124,N_2652);
or U3051 (N_3051,N_283,N_699);
nand U3052 (N_3052,N_796,N_1721);
nor U3053 (N_3053,N_1555,N_2340);
nor U3054 (N_3054,N_1615,N_2585);
nor U3055 (N_3055,N_781,N_636);
nand U3056 (N_3056,N_1654,N_483);
and U3057 (N_3057,N_664,N_1506);
or U3058 (N_3058,N_1399,N_214);
or U3059 (N_3059,N_1929,N_1077);
and U3060 (N_3060,N_1716,N_2178);
or U3061 (N_3061,N_2576,N_739);
nor U3062 (N_3062,N_307,N_1210);
or U3063 (N_3063,N_2305,N_2688);
or U3064 (N_3064,N_497,N_2111);
and U3065 (N_3065,N_530,N_2868);
or U3066 (N_3066,N_710,N_2510);
and U3067 (N_3067,N_162,N_2329);
or U3068 (N_3068,N_1509,N_2933);
nor U3069 (N_3069,N_1355,N_1519);
nor U3070 (N_3070,N_2261,N_354);
or U3071 (N_3071,N_2531,N_2975);
and U3072 (N_3072,N_1180,N_1434);
and U3073 (N_3073,N_1737,N_364);
and U3074 (N_3074,N_1523,N_2046);
or U3075 (N_3075,N_2404,N_709);
nand U3076 (N_3076,N_1013,N_125);
and U3077 (N_3077,N_1146,N_900);
or U3078 (N_3078,N_1833,N_926);
or U3079 (N_3079,N_2027,N_154);
nor U3080 (N_3080,N_2851,N_2801);
or U3081 (N_3081,N_2982,N_2496);
nor U3082 (N_3082,N_1113,N_1472);
nor U3083 (N_3083,N_2249,N_750);
or U3084 (N_3084,N_308,N_1111);
and U3085 (N_3085,N_2057,N_2405);
nand U3086 (N_3086,N_1839,N_1418);
or U3087 (N_3087,N_2946,N_2687);
and U3088 (N_3088,N_2254,N_1307);
nand U3089 (N_3089,N_2581,N_2050);
nor U3090 (N_3090,N_1535,N_960);
nor U3091 (N_3091,N_1952,N_1186);
and U3092 (N_3092,N_617,N_358);
or U3093 (N_3093,N_1796,N_1167);
nand U3094 (N_3094,N_1539,N_2798);
nor U3095 (N_3095,N_396,N_2140);
or U3096 (N_3096,N_295,N_1480);
nor U3097 (N_3097,N_1996,N_2932);
nand U3098 (N_3098,N_2587,N_776);
and U3099 (N_3099,N_1898,N_1375);
or U3100 (N_3100,N_1760,N_920);
nor U3101 (N_3101,N_1958,N_2474);
nand U3102 (N_3102,N_821,N_2690);
and U3103 (N_3103,N_2502,N_2596);
and U3104 (N_3104,N_217,N_1142);
or U3105 (N_3105,N_1131,N_870);
nor U3106 (N_3106,N_2219,N_1703);
nor U3107 (N_3107,N_749,N_2547);
or U3108 (N_3108,N_1129,N_1379);
and U3109 (N_3109,N_2700,N_1465);
nor U3110 (N_3110,N_524,N_1384);
or U3111 (N_3111,N_2552,N_1886);
or U3112 (N_3112,N_2609,N_2574);
and U3113 (N_3113,N_2895,N_580);
nor U3114 (N_3114,N_2958,N_743);
and U3115 (N_3115,N_536,N_526);
or U3116 (N_3116,N_2266,N_1607);
and U3117 (N_3117,N_1450,N_789);
and U3118 (N_3118,N_474,N_1713);
and U3119 (N_3119,N_986,N_1152);
nor U3120 (N_3120,N_1137,N_621);
nor U3121 (N_3121,N_2936,N_2091);
nand U3122 (N_3122,N_312,N_79);
nand U3123 (N_3123,N_2055,N_2566);
nor U3124 (N_3124,N_1466,N_1340);
nor U3125 (N_3125,N_212,N_787);
and U3126 (N_3126,N_414,N_772);
nand U3127 (N_3127,N_93,N_447);
nand U3128 (N_3128,N_2684,N_1857);
and U3129 (N_3129,N_2287,N_456);
nor U3130 (N_3130,N_604,N_2886);
nand U3131 (N_3131,N_386,N_630);
or U3132 (N_3132,N_2108,N_1205);
nor U3133 (N_3133,N_1968,N_2839);
nand U3134 (N_3134,N_2168,N_2522);
or U3135 (N_3135,N_725,N_1481);
and U3136 (N_3136,N_1718,N_2296);
nor U3137 (N_3137,N_704,N_1049);
or U3138 (N_3138,N_1638,N_1622);
nand U3139 (N_3139,N_531,N_1688);
nor U3140 (N_3140,N_2015,N_1172);
nand U3141 (N_3141,N_2291,N_23);
nor U3142 (N_3142,N_653,N_2204);
and U3143 (N_3143,N_2170,N_284);
nand U3144 (N_3144,N_1921,N_1732);
or U3145 (N_3145,N_566,N_1918);
nor U3146 (N_3146,N_2176,N_2473);
and U3147 (N_3147,N_593,N_27);
nor U3148 (N_3148,N_2664,N_1588);
nand U3149 (N_3149,N_1561,N_352);
nor U3150 (N_3150,N_2008,N_2925);
or U3151 (N_3151,N_1610,N_611);
and U3152 (N_3152,N_826,N_1670);
nor U3153 (N_3153,N_2110,N_2626);
nor U3154 (N_3154,N_2974,N_2921);
nand U3155 (N_3155,N_2191,N_385);
and U3156 (N_3156,N_1281,N_1133);
nand U3157 (N_3157,N_2029,N_1032);
xor U3158 (N_3158,N_600,N_1749);
and U3159 (N_3159,N_2653,N_478);
or U3160 (N_3160,N_771,N_2363);
nand U3161 (N_3161,N_2075,N_472);
nand U3162 (N_3162,N_1837,N_2376);
nand U3163 (N_3163,N_2832,N_1912);
nor U3164 (N_3164,N_16,N_1206);
nor U3165 (N_3165,N_717,N_113);
and U3166 (N_3166,N_2309,N_964);
nand U3167 (N_3167,N_2460,N_371);
nor U3168 (N_3168,N_1030,N_2583);
nand U3169 (N_3169,N_1427,N_2628);
nor U3170 (N_3170,N_2618,N_1603);
xor U3171 (N_3171,N_150,N_2466);
and U3172 (N_3172,N_1977,N_457);
nor U3173 (N_3173,N_1067,N_1302);
nand U3174 (N_3174,N_2301,N_2282);
or U3175 (N_3175,N_1404,N_2794);
nor U3176 (N_3176,N_1242,N_2634);
nor U3177 (N_3177,N_2318,N_1999);
and U3178 (N_3178,N_1288,N_1832);
nor U3179 (N_3179,N_2004,N_2594);
or U3180 (N_3180,N_1087,N_1849);
nand U3181 (N_3181,N_2088,N_1687);
nor U3182 (N_3182,N_1123,N_1882);
nor U3183 (N_3183,N_2399,N_1863);
nand U3184 (N_3184,N_436,N_1347);
nand U3185 (N_3185,N_823,N_1493);
and U3186 (N_3186,N_2469,N_519);
nand U3187 (N_3187,N_1130,N_2968);
or U3188 (N_3188,N_2880,N_1967);
nor U3189 (N_3189,N_673,N_2630);
or U3190 (N_3190,N_1754,N_1011);
nor U3191 (N_3191,N_2380,N_911);
nor U3192 (N_3192,N_1161,N_2633);
and U3193 (N_3193,N_2299,N_1150);
nor U3194 (N_3194,N_225,N_1997);
or U3195 (N_3195,N_323,N_2573);
nor U3196 (N_3196,N_85,N_387);
and U3197 (N_3197,N_1693,N_161);
nand U3198 (N_3198,N_609,N_126);
or U3199 (N_3199,N_904,N_2455);
nand U3200 (N_3200,N_2118,N_1144);
or U3201 (N_3201,N_2214,N_2553);
nand U3202 (N_3202,N_432,N_2079);
and U3203 (N_3203,N_953,N_2283);
or U3204 (N_3204,N_1510,N_390);
or U3205 (N_3205,N_1109,N_2348);
or U3206 (N_3206,N_2124,N_1847);
or U3207 (N_3207,N_1257,N_2441);
xor U3208 (N_3208,N_695,N_2195);
nor U3209 (N_3209,N_2406,N_263);
nand U3210 (N_3210,N_989,N_1444);
or U3211 (N_3211,N_2963,N_1983);
or U3212 (N_3212,N_2740,N_2847);
and U3213 (N_3213,N_2674,N_1566);
nand U3214 (N_3214,N_671,N_66);
nand U3215 (N_3215,N_342,N_452);
and U3216 (N_3216,N_619,N_869);
xor U3217 (N_3217,N_799,N_2290);
or U3218 (N_3218,N_2023,N_2916);
nand U3219 (N_3219,N_769,N_2658);
or U3220 (N_3220,N_562,N_1774);
nor U3221 (N_3221,N_2678,N_1892);
nor U3222 (N_3222,N_927,N_2820);
and U3223 (N_3223,N_293,N_242);
or U3224 (N_3224,N_1888,N_2943);
nor U3225 (N_3225,N_505,N_2720);
and U3226 (N_3226,N_982,N_1571);
nor U3227 (N_3227,N_2164,N_1679);
nand U3228 (N_3228,N_2842,N_2386);
nor U3229 (N_3229,N_1894,N_373);
and U3230 (N_3230,N_2659,N_1790);
and U3231 (N_3231,N_1101,N_2661);
or U3232 (N_3232,N_2312,N_644);
nor U3233 (N_3233,N_1798,N_175);
nor U3234 (N_3234,N_163,N_2985);
nor U3235 (N_3235,N_2369,N_1018);
and U3236 (N_3236,N_1239,N_2796);
nor U3237 (N_3237,N_2210,N_267);
nor U3238 (N_3238,N_2148,N_2648);
nand U3239 (N_3239,N_2888,N_1826);
or U3240 (N_3240,N_2288,N_1148);
nand U3241 (N_3241,N_2774,N_2285);
or U3242 (N_3242,N_1364,N_2962);
and U3243 (N_3243,N_196,N_909);
nand U3244 (N_3244,N_430,N_885);
nand U3245 (N_3245,N_694,N_1717);
nand U3246 (N_3246,N_864,N_1422);
nand U3247 (N_3247,N_2988,N_542);
nand U3248 (N_3248,N_102,N_1669);
or U3249 (N_3249,N_337,N_1272);
or U3250 (N_3250,N_1395,N_997);
and U3251 (N_3251,N_1026,N_59);
nand U3252 (N_3252,N_1407,N_663);
and U3253 (N_3253,N_1378,N_2912);
and U3254 (N_3254,N_2651,N_2158);
and U3255 (N_3255,N_440,N_2415);
nor U3256 (N_3256,N_2072,N_2252);
nor U3257 (N_3257,N_1175,N_412);
nand U3258 (N_3258,N_667,N_1700);
and U3259 (N_3259,N_902,N_177);
nor U3260 (N_3260,N_827,N_2059);
and U3261 (N_3261,N_1672,N_1515);
nand U3262 (N_3262,N_896,N_2253);
and U3263 (N_3263,N_221,N_2591);
and U3264 (N_3264,N_1315,N_544);
or U3265 (N_3265,N_363,N_2414);
and U3266 (N_3266,N_328,N_2101);
and U3267 (N_3267,N_1746,N_9);
nand U3268 (N_3268,N_25,N_518);
nor U3269 (N_3269,N_626,N_1969);
or U3270 (N_3270,N_2139,N_983);
or U3271 (N_3271,N_2759,N_924);
nand U3272 (N_3272,N_1514,N_319);
and U3273 (N_3273,N_1033,N_991);
nor U3274 (N_3274,N_2434,N_91);
nand U3275 (N_3275,N_2131,N_1621);
and U3276 (N_3276,N_2697,N_1995);
and U3277 (N_3277,N_2843,N_1102);
or U3278 (N_3278,N_2903,N_2133);
or U3279 (N_3279,N_867,N_1015);
and U3280 (N_3280,N_1601,N_2443);
nand U3281 (N_3281,N_1244,N_1369);
or U3282 (N_3282,N_874,N_1310);
and U3283 (N_3283,N_728,N_2727);
and U3284 (N_3284,N_1188,N_662);
or U3285 (N_3285,N_2544,N_259);
and U3286 (N_3286,N_2677,N_2138);
nor U3287 (N_3287,N_1517,N_228);
nand U3288 (N_3288,N_2813,N_2855);
or U3289 (N_3289,N_592,N_1660);
nor U3290 (N_3290,N_2987,N_2292);
nand U3291 (N_3291,N_2150,N_830);
nor U3292 (N_3292,N_73,N_500);
nor U3293 (N_3293,N_1631,N_1443);
and U3294 (N_3294,N_2507,N_852);
and U3295 (N_3295,N_384,N_875);
and U3296 (N_3296,N_1014,N_2222);
nand U3297 (N_3297,N_58,N_1248);
or U3298 (N_3298,N_669,N_2734);
nand U3299 (N_3299,N_1750,N_2572);
nand U3300 (N_3300,N_1372,N_1096);
or U3301 (N_3301,N_485,N_1483);
and U3302 (N_3302,N_1667,N_1416);
and U3303 (N_3303,N_2848,N_1125);
or U3304 (N_3304,N_1695,N_1990);
and U3305 (N_3305,N_2738,N_206);
or U3306 (N_3306,N_2773,N_2497);
nor U3307 (N_3307,N_1545,N_173);
or U3308 (N_3308,N_2387,N_324);
nand U3309 (N_3309,N_601,N_2647);
nand U3310 (N_3310,N_2731,N_2324);
or U3311 (N_3311,N_2772,N_2718);
and U3312 (N_3312,N_1006,N_584);
nor U3313 (N_3313,N_2006,N_149);
nand U3314 (N_3314,N_2042,N_2297);
nor U3315 (N_3315,N_970,N_321);
and U3316 (N_3316,N_894,N_1512);
or U3317 (N_3317,N_468,N_1270);
or U3318 (N_3318,N_2821,N_800);
nor U3319 (N_3319,N_1157,N_2877);
or U3320 (N_3320,N_916,N_866);
nor U3321 (N_3321,N_2498,N_2230);
nand U3322 (N_3322,N_759,N_1277);
nand U3323 (N_3323,N_2263,N_41);
nor U3324 (N_3324,N_565,N_15);
or U3325 (N_3325,N_1652,N_2109);
and U3326 (N_3326,N_1226,N_2120);
nor U3327 (N_3327,N_1504,N_1808);
or U3328 (N_3328,N_1452,N_49);
nand U3329 (N_3329,N_1901,N_1273);
nand U3330 (N_3330,N_2597,N_1214);
nor U3331 (N_3331,N_2940,N_344);
and U3332 (N_3332,N_825,N_2979);
and U3333 (N_3333,N_2881,N_726);
or U3334 (N_3334,N_2425,N_1484);
or U3335 (N_3335,N_540,N_2556);
or U3336 (N_3336,N_2532,N_1072);
and U3337 (N_3337,N_637,N_1985);
nand U3338 (N_3338,N_968,N_816);
nand U3339 (N_3339,N_370,N_1389);
or U3340 (N_3340,N_218,N_736);
and U3341 (N_3341,N_133,N_2711);
nor U3342 (N_3342,N_401,N_2273);
or U3343 (N_3343,N_2493,N_697);
and U3344 (N_3344,N_2756,N_1000);
or U3345 (N_3345,N_1394,N_2602);
and U3346 (N_3346,N_420,N_2331);
or U3347 (N_3347,N_383,N_164);
nand U3348 (N_3348,N_480,N_2314);
and U3349 (N_3349,N_67,N_2799);
and U3350 (N_3350,N_2657,N_606);
nand U3351 (N_3351,N_494,N_1485);
and U3352 (N_3352,N_1457,N_1341);
and U3353 (N_3353,N_1575,N_2592);
nand U3354 (N_3354,N_1329,N_2354);
or U3355 (N_3355,N_2478,N_17);
or U3356 (N_3356,N_1656,N_490);
or U3357 (N_3357,N_131,N_2529);
nand U3358 (N_3358,N_368,N_1028);
nand U3359 (N_3359,N_1779,N_993);
nand U3360 (N_3360,N_2588,N_252);
or U3361 (N_3361,N_1936,N_757);
nor U3362 (N_3362,N_2216,N_2571);
or U3363 (N_3363,N_466,N_2394);
nor U3364 (N_3364,N_2112,N_2514);
and U3365 (N_3365,N_340,N_719);
nor U3366 (N_3366,N_931,N_2048);
nor U3367 (N_3367,N_1313,N_1091);
and U3368 (N_3368,N_2680,N_1838);
and U3369 (N_3369,N_411,N_2402);
nand U3370 (N_3370,N_1973,N_303);
and U3371 (N_3371,N_461,N_1678);
nand U3372 (N_3372,N_2969,N_2945);
or U3373 (N_3373,N_2879,N_2508);
or U3374 (N_3374,N_1040,N_1354);
and U3375 (N_3375,N_521,N_1078);
xnor U3376 (N_3376,N_2181,N_31);
nand U3377 (N_3377,N_2791,N_279);
or U3378 (N_3378,N_1020,N_2561);
nor U3379 (N_3379,N_1441,N_685);
nor U3380 (N_3380,N_810,N_1256);
nand U3381 (N_3381,N_1628,N_2052);
nand U3382 (N_3382,N_678,N_680);
nor U3383 (N_3383,N_226,N_2769);
nand U3384 (N_3384,N_1035,N_602);
nand U3385 (N_3385,N_425,N_2347);
nand U3386 (N_3386,N_1637,N_2906);
or U3387 (N_3387,N_1223,N_120);
and U3388 (N_3388,N_199,N_2683);
nor U3389 (N_3389,N_1100,N_389);
nand U3390 (N_3390,N_2450,N_2952);
nor U3391 (N_3391,N_747,N_1964);
or U3392 (N_3392,N_2377,N_2670);
or U3393 (N_3393,N_266,N_555);
nand U3394 (N_3394,N_1112,N_2442);
nor U3395 (N_3395,N_610,N_11);
or U3396 (N_3396,N_2231,N_1715);
or U3397 (N_3397,N_2857,N_2279);
and U3398 (N_3398,N_2825,N_2736);
nor U3399 (N_3399,N_36,N_462);
nor U3400 (N_3400,N_97,N_243);
and U3401 (N_3401,N_1423,N_424);
nor U3402 (N_3402,N_1358,N_1899);
or U3403 (N_3403,N_1170,N_236);
nand U3404 (N_3404,N_907,N_1994);
nor U3405 (N_3405,N_1199,N_2874);
nor U3406 (N_3406,N_1353,N_260);
and U3407 (N_3407,N_1828,N_2548);
nor U3408 (N_3408,N_512,N_282);
or U3409 (N_3409,N_969,N_2146);
or U3410 (N_3410,N_2622,N_2056);
and U3411 (N_3411,N_375,N_34);
or U3412 (N_3412,N_634,N_1594);
and U3413 (N_3413,N_2365,N_1464);
nor U3414 (N_3414,N_878,N_1897);
and U3415 (N_3415,N_2890,N_1103);
or U3416 (N_3416,N_1547,N_121);
nor U3417 (N_3417,N_1806,N_984);
or U3418 (N_3418,N_1500,N_733);
nor U3419 (N_3419,N_1408,N_1513);
nor U3420 (N_3420,N_1876,N_30);
or U3421 (N_3421,N_1862,N_1497);
or U3422 (N_3422,N_152,N_1386);
nand U3423 (N_3423,N_2893,N_2335);
nand U3424 (N_3424,N_2580,N_1986);
or U3425 (N_3425,N_2149,N_1377);
xnor U3426 (N_3426,N_372,N_82);
nand U3427 (N_3427,N_831,N_679);
nor U3428 (N_3428,N_253,N_889);
nand U3429 (N_3429,N_2777,N_2949);
nor U3430 (N_3430,N_1117,N_1088);
nor U3431 (N_3431,N_1580,N_2616);
and U3432 (N_3432,N_2197,N_1044);
or U3433 (N_3433,N_2440,N_1546);
or U3434 (N_3434,N_1324,N_1570);
and U3435 (N_3435,N_1646,N_893);
xnor U3436 (N_3436,N_940,N_2388);
or U3437 (N_3437,N_598,N_613);
or U3438 (N_3438,N_2613,N_838);
nand U3439 (N_3439,N_2698,N_2465);
nor U3440 (N_3440,N_409,N_361);
nor U3441 (N_3441,N_966,N_1351);
nand U3442 (N_3442,N_2787,N_1680);
and U3443 (N_3443,N_1825,N_476);
nand U3444 (N_3444,N_742,N_2489);
or U3445 (N_3445,N_2991,N_220);
or U3446 (N_3446,N_1048,N_2937);
nor U3447 (N_3447,N_2517,N_1733);
or U3448 (N_3448,N_209,N_1783);
and U3449 (N_3449,N_2492,N_317);
nor U3450 (N_3450,N_1081,N_2681);
nand U3451 (N_3451,N_905,N_577);
and U3452 (N_3452,N_819,N_1151);
nor U3453 (N_3453,N_453,N_37);
and U3454 (N_3454,N_2518,N_1595);
and U3455 (N_3455,N_2030,N_1748);
nand U3456 (N_3456,N_1182,N_24);
or U3457 (N_3457,N_1951,N_2830);
or U3458 (N_3458,N_189,N_1822);
or U3459 (N_3459,N_2795,N_2433);
nor U3460 (N_3460,N_720,N_1259);
and U3461 (N_3461,N_247,N_2693);
nand U3462 (N_3462,N_675,N_1767);
nor U3463 (N_3463,N_1282,N_1286);
nor U3464 (N_3464,N_1446,N_2141);
or U3465 (N_3465,N_2852,N_441);
or U3466 (N_3466,N_2833,N_1727);
nor U3467 (N_3467,N_366,N_676);
nand U3468 (N_3468,N_915,N_1400);
nor U3469 (N_3469,N_2073,N_2332);
nand U3470 (N_3470,N_2488,N_1577);
nand U3471 (N_3471,N_2353,N_2128);
and U3472 (N_3472,N_129,N_336);
nand U3473 (N_3473,N_570,N_886);
nor U3474 (N_3474,N_98,N_2132);
or U3475 (N_3475,N_795,N_513);
nand U3476 (N_3476,N_638,N_222);
nand U3477 (N_3477,N_1203,N_1173);
or U3478 (N_3478,N_1469,N_433);
nand U3479 (N_3479,N_90,N_2523);
and U3480 (N_3480,N_1902,N_1690);
or U3481 (N_3481,N_2814,N_1770);
nand U3482 (N_3482,N_2336,N_1850);
nor U3483 (N_3483,N_1883,N_589);
nor U3484 (N_3484,N_1271,N_791);
or U3485 (N_3485,N_1114,N_934);
nor U3486 (N_3486,N_702,N_273);
nand U3487 (N_3487,N_1177,N_1880);
nand U3488 (N_3488,N_2311,N_691);
nor U3489 (N_3489,N_2470,N_2998);
or U3490 (N_3490,N_84,N_2822);
or U3491 (N_3491,N_2728,N_2077);
or U3492 (N_3492,N_1005,N_2351);
nand U3493 (N_3493,N_1881,N_2366);
nand U3494 (N_3494,N_1705,N_471);
nand U3495 (N_3495,N_2130,N_1209);
nor U3496 (N_3496,N_2505,N_326);
nor U3497 (N_3497,N_654,N_879);
and U3498 (N_3498,N_155,N_465);
nand U3499 (N_3499,N_2157,N_2907);
nor U3500 (N_3500,N_1107,N_2174);
nand U3501 (N_3501,N_665,N_2604);
or U3502 (N_3502,N_1193,N_2154);
or U3503 (N_3503,N_1604,N_919);
nand U3504 (N_3504,N_2001,N_369);
nand U3505 (N_3505,N_95,N_2121);
or U3506 (N_3506,N_347,N_1771);
nor U3507 (N_3507,N_2205,N_391);
nor U3508 (N_3508,N_1245,N_705);
nand U3509 (N_3509,N_1805,N_2016);
nor U3510 (N_3510,N_1022,N_1009);
or U3511 (N_3511,N_2815,N_620);
or U3512 (N_3512,N_2169,N_1879);
and U3513 (N_3513,N_402,N_1079);
or U3514 (N_3514,N_559,N_958);
or U3515 (N_3515,N_2114,N_1537);
nand U3516 (N_3516,N_1950,N_2913);
nand U3517 (N_3517,N_2463,N_1316);
and U3518 (N_3518,N_1492,N_2918);
nor U3519 (N_3519,N_2603,N_2229);
nor U3520 (N_3520,N_2612,N_1417);
or U3521 (N_3521,N_535,N_1224);
nor U3522 (N_3522,N_2758,N_1978);
nor U3523 (N_3523,N_1873,N_1907);
nand U3524 (N_3524,N_2126,N_29);
nor U3525 (N_3525,N_52,N_681);
and U3526 (N_3526,N_94,N_2793);
and U3527 (N_3527,N_1053,N_1845);
nand U3528 (N_3528,N_1608,N_2649);
and U3529 (N_3529,N_1891,N_2135);
nor U3530 (N_3530,N_1947,N_240);
or U3531 (N_3531,N_1734,N_2185);
nand U3532 (N_3532,N_2558,N_877);
nor U3533 (N_3533,N_2540,N_1699);
nand U3534 (N_3534,N_1183,N_2246);
nand U3535 (N_3535,N_115,N_2341);
nor U3536 (N_3536,N_281,N_398);
and U3537 (N_3537,N_2512,N_288);
or U3538 (N_3538,N_567,N_1955);
or U3539 (N_3539,N_895,N_2504);
nor U3540 (N_3540,N_2076,N_297);
nand U3541 (N_3541,N_2565,N_2391);
nand U3542 (N_3542,N_1885,N_1916);
xor U3543 (N_3543,N_2064,N_545);
or U3544 (N_3544,N_2213,N_1772);
and U3545 (N_3545,N_2644,N_1335);
or U3546 (N_3546,N_1121,N_917);
or U3547 (N_3547,N_2837,N_2965);
nor U3548 (N_3548,N_841,N_119);
nor U3549 (N_3549,N_1128,N_2509);
nor U3550 (N_3550,N_1991,N_1581);
and U3551 (N_3551,N_2092,N_1083);
nand U3552 (N_3552,N_2276,N_2448);
or U3553 (N_3553,N_1719,N_1777);
and U3554 (N_3554,N_2663,N_1478);
nor U3555 (N_3555,N_534,N_2407);
or U3556 (N_3556,N_624,N_734);
nor U3557 (N_3557,N_2543,N_2901);
nand U3558 (N_3558,N_2600,N_285);
nand U3559 (N_3559,N_1196,N_1312);
nand U3560 (N_3560,N_2383,N_1507);
nand U3561 (N_3561,N_2033,N_1208);
xnor U3562 (N_3562,N_1917,N_2546);
or U3563 (N_3563,N_2269,N_507);
and U3564 (N_3564,N_1764,N_2632);
nand U3565 (N_3565,N_2476,N_1305);
nor U3566 (N_3566,N_523,N_110);
nand U3567 (N_3567,N_127,N_2082);
or U3568 (N_3568,N_2104,N_2749);
or U3569 (N_3569,N_157,N_2430);
nand U3570 (N_3570,N_1155,N_1747);
nor U3571 (N_3571,N_2608,N_2062);
and U3572 (N_3572,N_1642,N_511);
and U3573 (N_3573,N_2039,N_1782);
xnor U3574 (N_3574,N_2705,N_208);
nor U3575 (N_3575,N_692,N_2447);
or U3576 (N_3576,N_1532,N_1585);
nor U3577 (N_3577,N_55,N_756);
and U3578 (N_3578,N_21,N_857);
and U3579 (N_3579,N_2374,N_2941);
nor U3580 (N_3580,N_205,N_959);
nor U3581 (N_3581,N_1762,N_2143);
nand U3582 (N_3582,N_77,N_2875);
nor U3583 (N_3583,N_2849,N_2646);
or U3584 (N_3584,N_1290,N_197);
or U3585 (N_3585,N_1410,N_2970);
or U3586 (N_3586,N_627,N_1623);
or U3587 (N_3587,N_2527,N_1047);
or U3588 (N_3588,N_1893,N_1859);
nor U3589 (N_3589,N_2530,N_2317);
or U3590 (N_3590,N_701,N_2202);
or U3591 (N_3591,N_1120,N_186);
nor U3592 (N_3592,N_117,N_467);
or U3593 (N_3593,N_1412,N_1390);
and U3594 (N_3594,N_1090,N_1237);
nand U3595 (N_3595,N_1970,N_988);
or U3596 (N_3596,N_1851,N_2007);
nand U3597 (N_3597,N_1494,N_1197);
nand U3598 (N_3598,N_845,N_707);
nand U3599 (N_3599,N_582,N_2173);
and U3600 (N_3600,N_393,N_381);
nor U3601 (N_3601,N_1473,N_463);
and U3602 (N_3602,N_2810,N_2475);
or U3603 (N_3603,N_556,N_753);
or U3604 (N_3604,N_1613,N_1370);
or U3605 (N_3605,N_945,N_2058);
or U3606 (N_3606,N_123,N_195);
and U3607 (N_3607,N_1802,N_2741);
and U3608 (N_3608,N_802,N_1166);
nand U3609 (N_3609,N_1984,N_995);
and U3610 (N_3610,N_213,N_2395);
and U3611 (N_3611,N_1381,N_2797);
nand U3612 (N_3612,N_153,N_901);
or U3613 (N_3613,N_2992,N_537);
and U3614 (N_3614,N_320,N_1348);
and U3615 (N_3615,N_899,N_2719);
nor U3616 (N_3616,N_2535,N_2268);
and U3617 (N_3617,N_258,N_1651);
nor U3618 (N_3618,N_238,N_26);
and U3619 (N_3619,N_1874,N_625);
or U3620 (N_3620,N_276,N_2765);
nor U3621 (N_3621,N_1686,N_1174);
or U3622 (N_3622,N_357,N_1818);
or U3623 (N_3623,N_172,N_1253);
or U3624 (N_3624,N_812,N_1439);
or U3625 (N_3625,N_2919,N_751);
and U3626 (N_3626,N_2066,N_146);
nor U3627 (N_3627,N_2043,N_99);
or U3628 (N_3628,N_847,N_1592);
nor U3629 (N_3629,N_2624,N_1403);
xor U3630 (N_3630,N_2145,N_1948);
and U3631 (N_3631,N_1322,N_1711);
or U3632 (N_3632,N_1051,N_811);
nor U3633 (N_3633,N_2645,N_2827);
nor U3634 (N_3634,N_2818,N_1331);
or U3635 (N_3635,N_105,N_1159);
nor U3636 (N_3636,N_374,N_2545);
and U3637 (N_3637,N_543,N_2980);
nor U3638 (N_3638,N_1761,N_950);
nand U3639 (N_3639,N_1065,N_1816);
nand U3640 (N_3640,N_2241,N_2270);
nand U3641 (N_3641,N_1299,N_1896);
or U3642 (N_3642,N_2917,N_491);
and U3643 (N_3643,N_829,N_1753);
nor U3644 (N_3644,N_2831,N_778);
nor U3645 (N_3645,N_2631,N_2259);
and U3646 (N_3646,N_2242,N_2152);
nor U3647 (N_3647,N_2844,N_180);
or U3648 (N_3648,N_1528,N_2541);
and U3649 (N_3649,N_2401,N_981);
or U3650 (N_3650,N_1975,N_2069);
nor U3651 (N_3651,N_1620,N_1491);
and U3652 (N_3652,N_10,N_640);
or U3653 (N_3653,N_248,N_1046);
or U3654 (N_3654,N_2716,N_2549);
nor U3655 (N_3655,N_2867,N_147);
or U3656 (N_3656,N_1204,N_820);
and U3657 (N_3657,N_2134,N_2171);
and U3658 (N_3658,N_2417,N_890);
or U3659 (N_3659,N_2676,N_1756);
nor U3660 (N_3660,N_1425,N_2358);
nand U3661 (N_3661,N_1658,N_1831);
and U3662 (N_3662,N_313,N_1864);
nor U3663 (N_3663,N_2826,N_938);
and U3664 (N_3664,N_871,N_318);
nand U3665 (N_3665,N_403,N_45);
nand U3666 (N_3666,N_1007,N_1192);
nor U3667 (N_3667,N_1787,N_1105);
nor U3668 (N_3668,N_1373,N_2051);
or U3669 (N_3669,N_2996,N_2557);
nand U3670 (N_3670,N_745,N_1550);
nor U3671 (N_3671,N_1935,N_930);
xnor U3672 (N_3672,N_2188,N_1066);
and U3673 (N_3673,N_2233,N_290);
or U3674 (N_3674,N_274,N_484);
nand U3675 (N_3675,N_2577,N_92);
and U3676 (N_3676,N_1911,N_2590);
nand U3677 (N_3677,N_760,N_1156);
and U3678 (N_3678,N_13,N_1908);
and U3679 (N_3679,N_74,N_2060);
or U3680 (N_3680,N_2375,N_850);
nor U3681 (N_3681,N_2359,N_2026);
or U3682 (N_3682,N_1360,N_2902);
nor U3683 (N_3683,N_1168,N_2944);
or U3684 (N_3684,N_2239,N_1291);
nor U3685 (N_3685,N_2163,N_233);
nand U3686 (N_3686,N_2009,N_338);
or U3687 (N_3687,N_839,N_1836);
xnor U3688 (N_3688,N_784,N_2554);
nand U3689 (N_3689,N_1942,N_2500);
or U3690 (N_3690,N_1073,N_2303);
nor U3691 (N_3691,N_351,N_1396);
or U3692 (N_3692,N_1383,N_1824);
or U3693 (N_3693,N_1689,N_56);
nand U3694 (N_3694,N_330,N_1600);
nor U3695 (N_3695,N_2638,N_1933);
and U3696 (N_3696,N_862,N_730);
and U3697 (N_3697,N_19,N_1225);
nor U3698 (N_3698,N_136,N_2662);
and U3699 (N_3699,N_775,N_1356);
or U3700 (N_3700,N_1050,N_2726);
nor U3701 (N_3701,N_2144,N_2656);
xnor U3702 (N_3702,N_428,N_32);
or U3703 (N_3703,N_1008,N_2882);
or U3704 (N_3704,N_2579,N_479);
nand U3705 (N_3705,N_1323,N_170);
and U3706 (N_3706,N_1829,N_554);
nor U3707 (N_3707,N_2629,N_1596);
and U3708 (N_3708,N_2177,N_1122);
nor U3709 (N_3709,N_1819,N_1140);
nor U3710 (N_3710,N_698,N_2668);
and U3711 (N_3711,N_608,N_686);
or U3712 (N_3712,N_723,N_2054);
nand U3713 (N_3713,N_2472,N_81);
and U3714 (N_3714,N_1855,N_586);
nand U3715 (N_3715,N_1459,N_994);
or U3716 (N_3716,N_2161,N_855);
nand U3717 (N_3717,N_1701,N_2200);
or U3718 (N_3718,N_2870,N_2215);
and U3719 (N_3719,N_688,N_632);
nand U3720 (N_3720,N_2973,N_956);
or U3721 (N_3721,N_1433,N_649);
or U3722 (N_3722,N_1293,N_1222);
and U3723 (N_3723,N_670,N_1380);
or U3724 (N_3724,N_1939,N_1966);
nor U3725 (N_3725,N_2993,N_1426);
nor U3726 (N_3726,N_1579,N_1846);
or U3727 (N_3727,N_612,N_532);
nand U3728 (N_3728,N_2125,N_144);
nand U3729 (N_3729,N_941,N_933);
nor U3730 (N_3730,N_2486,N_1560);
nor U3731 (N_3731,N_353,N_2325);
nor U3732 (N_3732,N_168,N_289);
nor U3733 (N_3733,N_2483,N_100);
nor U3734 (N_3734,N_1184,N_1227);
or U3735 (N_3735,N_744,N_735);
nand U3736 (N_3736,N_135,N_1673);
nand U3737 (N_3737,N_499,N_1190);
nor U3738 (N_3738,N_2182,N_2458);
or U3739 (N_3739,N_1564,N_729);
nand U3740 (N_3740,N_450,N_2094);
or U3741 (N_3741,N_2589,N_1582);
and U3742 (N_3742,N_2682,N_2999);
and U3743 (N_3743,N_764,N_1058);
and U3744 (N_3744,N_2685,N_1858);
and U3745 (N_3745,N_2003,N_1421);
or U3746 (N_3746,N_1076,N_1165);
and U3747 (N_3747,N_1854,N_2551);
or U3748 (N_3748,N_2788,N_1392);
or U3749 (N_3749,N_2623,N_2513);
and U3750 (N_3750,N_2538,N_2753);
and U3751 (N_3751,N_310,N_2819);
or U3752 (N_3752,N_2696,N_2097);
nor U3753 (N_3753,N_1763,N_1247);
or U3754 (N_3754,N_2706,N_2083);
nand U3755 (N_3755,N_269,N_797);
nor U3756 (N_3756,N_2775,N_897);
or U3757 (N_3757,N_1944,N_2704);
or U3758 (N_3758,N_2098,N_2274);
nand U3759 (N_3759,N_156,N_2203);
nor U3760 (N_3760,N_844,N_1021);
or U3761 (N_3761,N_2984,N_2762);
and U3762 (N_3762,N_2569,N_1776);
or U3763 (N_3763,N_2829,N_2802);
nand U3764 (N_3764,N_1811,N_590);
nand U3765 (N_3765,N_50,N_2295);
nand U3766 (N_3766,N_400,N_2155);
nor U3767 (N_3767,N_1219,N_1803);
nor U3768 (N_3768,N_2479,N_487);
and U3769 (N_3769,N_853,N_1261);
and U3770 (N_3770,N_2534,N_2713);
or U3771 (N_3771,N_1249,N_108);
nor U3772 (N_3772,N_2976,N_1463);
or U3773 (N_3773,N_2920,N_191);
nand U3774 (N_3774,N_859,N_1720);
and U3775 (N_3775,N_300,N_996);
or U3776 (N_3776,N_2914,N_422);
nand U3777 (N_3777,N_2953,N_498);
or U3778 (N_3778,N_415,N_1871);
or U3779 (N_3779,N_642,N_2370);
or U3780 (N_3780,N_1298,N_903);
or U3781 (N_3781,N_2342,N_801);
nand U3782 (N_3782,N_454,N_696);
and U3783 (N_3783,N_1189,N_1960);
or U3784 (N_3784,N_672,N_2672);
nand U3785 (N_3785,N_2735,N_38);
and U3786 (N_3786,N_1029,N_331);
or U3787 (N_3787,N_2212,N_421);
nor U3788 (N_3788,N_1910,N_517);
and U3789 (N_3789,N_1475,N_1438);
and U3790 (N_3790,N_2304,N_211);
and U3791 (N_3791,N_2960,N_2896);
or U3792 (N_3792,N_2087,N_1094);
or U3793 (N_3793,N_684,N_1914);
nand U3794 (N_3794,N_87,N_1758);
nor U3795 (N_3795,N_643,N_1630);
nor U3796 (N_3796,N_2757,N_1865);
or U3797 (N_3797,N_394,N_1357);
nand U3798 (N_3798,N_1640,N_198);
xor U3799 (N_3799,N_1612,N_2032);
or U3800 (N_3800,N_417,N_2223);
nor U3801 (N_3801,N_1963,N_2828);
nand U3802 (N_3802,N_2665,N_1844);
and U3803 (N_3803,N_1735,N_1424);
nor U3804 (N_3804,N_762,N_1179);
nor U3805 (N_3805,N_367,N_2255);
or U3806 (N_3806,N_1726,N_786);
or U3807 (N_3807,N_215,N_2116);
nand U3808 (N_3808,N_2807,N_2840);
nand U3809 (N_3809,N_2014,N_1268);
nor U3810 (N_3810,N_1576,N_522);
or U3811 (N_3811,N_2935,N_1141);
nand U3812 (N_3812,N_182,N_1723);
nand U3813 (N_3813,N_846,N_2211);
or U3814 (N_3814,N_2671,N_2593);
nor U3815 (N_3815,N_2897,N_2400);
or U3816 (N_3816,N_722,N_2686);
and U3817 (N_3817,N_2760,N_2586);
nor U3818 (N_3818,N_914,N_2811);
nor U3819 (N_3819,N_1287,N_83);
nand U3820 (N_3820,N_2724,N_2403);
nor U3821 (N_3821,N_75,N_2699);
and U3822 (N_3822,N_305,N_1201);
or U3823 (N_3823,N_1233,N_2694);
nor U3824 (N_3824,N_551,N_714);
nor U3825 (N_3825,N_731,N_1974);
and U3826 (N_3826,N_936,N_219);
and U3827 (N_3827,N_1792,N_1365);
nand U3828 (N_3828,N_1980,N_2494);
nand U3829 (N_3829,N_1784,N_1559);
nor U3830 (N_3830,N_2385,N_2344);
nor U3831 (N_3831,N_1949,N_2117);
nand U3832 (N_3832,N_2183,N_89);
nand U3833 (N_3833,N_22,N_1682);
or U3834 (N_3834,N_547,N_2511);
nand U3835 (N_3835,N_327,N_2859);
or U3836 (N_3836,N_2107,N_1778);
and U3837 (N_3837,N_1086,N_268);
or U3838 (N_3838,N_587,N_1406);
or U3839 (N_3839,N_2099,N_560);
nor U3840 (N_3840,N_1773,N_502);
or U3841 (N_3841,N_1254,N_2865);
nand U3842 (N_3842,N_2892,N_1971);
or U3843 (N_3843,N_1301,N_1842);
xor U3844 (N_3844,N_1627,N_1362);
and U3845 (N_3845,N_746,N_2234);
or U3846 (N_3846,N_1572,N_449);
and U3847 (N_3847,N_1332,N_1488);
nor U3848 (N_3848,N_2338,N_482);
or U3849 (N_3849,N_111,N_2217);
or U3850 (N_3850,N_1267,N_647);
or U3851 (N_3851,N_1336,N_2449);
nand U3852 (N_3852,N_2378,N_1289);
or U3853 (N_3853,N_882,N_1662);
nand U3854 (N_3854,N_379,N_1419);
nand U3855 (N_3855,N_1531,N_1031);
and U3856 (N_3856,N_635,N_2605);
or U3857 (N_3857,N_142,N_2034);
nand U3858 (N_3858,N_455,N_2971);
and U3859 (N_3859,N_2339,N_2272);
nand U3860 (N_3860,N_2424,N_2275);
and U3861 (N_3861,N_2218,N_2715);
nor U3862 (N_3862,N_2428,N_2345);
or U3863 (N_3863,N_1325,N_2221);
nor U3864 (N_3864,N_1558,N_525);
nand U3865 (N_3865,N_1448,N_1470);
xnor U3866 (N_3866,N_122,N_1023);
or U3867 (N_3867,N_1835,N_1685);
or U3868 (N_3868,N_140,N_1584);
and U3869 (N_3869,N_346,N_134);
nand U3870 (N_3870,N_718,N_47);
and U3871 (N_3871,N_1106,N_2931);
and U3872 (N_3872,N_1527,N_668);
or U3873 (N_3873,N_785,N_1229);
nor U3874 (N_3874,N_716,N_979);
nand U3875 (N_3875,N_64,N_572);
or U3876 (N_3876,N_1578,N_2459);
or U3877 (N_3877,N_359,N_1661);
nor U3878 (N_3878,N_343,N_1522);
nor U3879 (N_3879,N_2899,N_597);
nor U3880 (N_3880,N_277,N_1471);
and U3881 (N_3881,N_204,N_2499);
or U3882 (N_3882,N_2781,N_700);
nand U3883 (N_3883,N_287,N_1038);
nand U3884 (N_3884,N_2501,N_2575);
or U3885 (N_3885,N_533,N_1216);
nor U3886 (N_3886,N_2081,N_3);
nand U3887 (N_3887,N_1126,N_2994);
nand U3888 (N_3888,N_721,N_2190);
nand U3889 (N_3889,N_2480,N_2883);
nand U3890 (N_3890,N_1074,N_579);
nor U3891 (N_3891,N_1860,N_2435);
and U3892 (N_3892,N_929,N_2621);
and U3893 (N_3893,N_264,N_458);
nor U3894 (N_3894,N_834,N_1024);
or U3895 (N_3895,N_957,N_2528);
nand U3896 (N_3896,N_1691,N_103);
and U3897 (N_3897,N_661,N_2627);
and U3898 (N_3898,N_2412,N_779);
nor U3899 (N_3899,N_2900,N_448);
or U3900 (N_3900,N_1549,N_2655);
or U3901 (N_3901,N_2611,N_515);
nor U3902 (N_3902,N_2089,N_558);
nand U3903 (N_3903,N_2783,N_1568);
or U3904 (N_3904,N_967,N_362);
or U3905 (N_3905,N_1202,N_1795);
or U3906 (N_3906,N_356,N_1320);
and U3907 (N_3907,N_1162,N_407);
nand U3908 (N_3908,N_1520,N_1655);
nor U3909 (N_3909,N_1132,N_183);
and U3910 (N_3910,N_564,N_1875);
nand U3911 (N_3911,N_552,N_241);
nand U3912 (N_3912,N_2873,N_2113);
nor U3913 (N_3913,N_943,N_2967);
nand U3914 (N_3914,N_1736,N_404);
nand U3915 (N_3915,N_1793,N_1965);
xnor U3916 (N_3916,N_291,N_677);
nor U3917 (N_3917,N_2800,N_1556);
nor U3918 (N_3918,N_1292,N_962);
and U3919 (N_3919,N_2068,N_1294);
nand U3920 (N_3920,N_223,N_2036);
and U3921 (N_3921,N_2166,N_193);
or U3922 (N_3922,N_306,N_1725);
or U3923 (N_3923,N_1136,N_2321);
and U3924 (N_3924,N_2349,N_2429);
nor U3925 (N_3925,N_2568,N_2834);
nor U3926 (N_3926,N_2328,N_1187);
and U3927 (N_3927,N_1704,N_840);
and U3928 (N_3928,N_2063,N_40);
nand U3929 (N_3929,N_2989,N_1877);
or U3930 (N_3930,N_246,N_1775);
nand U3931 (N_3931,N_652,N_1398);
and U3932 (N_3932,N_591,N_2491);
and U3933 (N_3933,N_2172,N_1124);
or U3934 (N_3934,N_1041,N_2495);
nand U3935 (N_3935,N_1342,N_1853);
and U3936 (N_3936,N_1436,N_851);
or U3937 (N_3937,N_2238,N_1252);
or U3938 (N_3938,N_2256,N_2159);
nand U3939 (N_3939,N_1388,N_475);
and U3940 (N_3940,N_1653,N_774);
nor U3941 (N_3941,N_539,N_2516);
or U3942 (N_3942,N_2084,N_496);
or U3943 (N_3943,N_116,N_399);
nand U3944 (N_3944,N_2983,N_72);
nor U3945 (N_3945,N_767,N_629);
nand U3946 (N_3946,N_2226,N_1447);
and U3947 (N_3947,N_1241,N_1565);
or U3948 (N_3948,N_1260,N_2964);
nor U3949 (N_3949,N_2948,N_2995);
and U3950 (N_3950,N_169,N_2393);
or U3951 (N_3951,N_495,N_835);
or U3952 (N_3952,N_166,N_244);
or U3953 (N_3953,N_1573,N_262);
nand U3954 (N_3954,N_63,N_1012);
and U3955 (N_3955,N_2308,N_477);
or U3956 (N_3956,N_332,N_1437);
nand U3957 (N_3957,N_898,N_1092);
and U3958 (N_3958,N_1218,N_814);
or U3959 (N_3959,N_2926,N_1143);
and U3960 (N_3960,N_486,N_1815);
nor U3961 (N_3961,N_1843,N_2789);
and U3962 (N_3962,N_1799,N_489);
nor U3963 (N_3963,N_1827,N_658);
nor U3964 (N_3964,N_1171,N_2410);
or U3965 (N_3965,N_1195,N_2220);
or U3966 (N_3966,N_1017,N_578);
nand U3967 (N_3967,N_683,N_538);
and U3968 (N_3968,N_1198,N_1145);
and U3969 (N_3969,N_1215,N_14);
and U3970 (N_3970,N_1037,N_657);
or U3971 (N_3971,N_1263,N_1574);
nand U3972 (N_3972,N_2481,N_2520);
or U3973 (N_3973,N_1922,N_2928);
nand U3974 (N_3974,N_392,N_143);
nand U3975 (N_3975,N_2240,N_824);
nor U3976 (N_3976,N_1533,N_408);
and U3977 (N_3977,N_1789,N_1296);
nor U3978 (N_3978,N_1895,N_1743);
nor U3979 (N_3979,N_2709,N_2564);
and U3980 (N_3980,N_1283,N_1285);
nor U3981 (N_3981,N_2737,N_2614);
and U3982 (N_3982,N_2850,N_2041);
nor U3983 (N_3983,N_2180,N_2426);
nor U3984 (N_3984,N_2271,N_299);
and U3985 (N_3985,N_1780,N_2236);
nand U3986 (N_3986,N_837,N_2281);
and U3987 (N_3987,N_596,N_1269);
or U3988 (N_3988,N_963,N_2539);
nor U3989 (N_3989,N_1841,N_2193);
or U3990 (N_3990,N_158,N_80);
nor U3991 (N_3991,N_2142,N_2280);
or U3992 (N_3992,N_1158,N_1303);
nor U3993 (N_3993,N_1057,N_1084);
nor U3994 (N_3994,N_2729,N_174);
xor U3995 (N_3995,N_2355,N_1583);
and U3996 (N_3996,N_1255,N_2869);
or U3997 (N_3997,N_2227,N_178);
or U3998 (N_3998,N_2457,N_883);
nand U3999 (N_3999,N_2357,N_2986);
or U4000 (N_4000,N_1309,N_1486);
nand U4001 (N_4001,N_2924,N_442);
nor U4002 (N_4002,N_1391,N_60);
nor U4003 (N_4003,N_382,N_2805);
and U4004 (N_4004,N_2445,N_954);
and U4005 (N_4005,N_1943,N_2432);
nand U4006 (N_4006,N_2625,N_1657);
and U4007 (N_4007,N_280,N_803);
and U4008 (N_4008,N_2477,N_2934);
or U4009 (N_4009,N_833,N_2766);
and U4010 (N_4010,N_2637,N_1598);
or U4011 (N_4011,N_2232,N_2364);
or U4012 (N_4012,N_1643,N_2005);
nand U4013 (N_4013,N_1609,N_2750);
xor U4014 (N_4014,N_2666,N_2327);
or U4015 (N_4015,N_687,N_1440);
nand U4016 (N_4016,N_2761,N_2396);
nor U4017 (N_4017,N_1280,N_1684);
xor U4018 (N_4018,N_2536,N_1626);
and U4019 (N_4019,N_1739,N_2444);
nand U4020 (N_4020,N_2884,N_1449);
nand U4021 (N_4021,N_69,N_1722);
nor U4022 (N_4022,N_1814,N_1923);
nor U4023 (N_4023,N_224,N_1905);
nand U4024 (N_4024,N_2235,N_1926);
nand U4025 (N_4025,N_1200,N_1430);
and U4026 (N_4026,N_470,N_1232);
nand U4027 (N_4027,N_2100,N_1346);
or U4028 (N_4028,N_2468,N_2990);
nand U4029 (N_4029,N_439,N_2225);
and U4030 (N_4030,N_1569,N_2835);
and U4031 (N_4031,N_1632,N_2782);
and U4032 (N_4032,N_942,N_2382);
nor U4033 (N_4033,N_1445,N_561);
or U4034 (N_4034,N_2446,N_216);
nor U4035 (N_4035,N_1063,N_378);
nand U4036 (N_4036,N_2080,N_1317);
and U4037 (N_4037,N_1479,N_2584);
nand U4038 (N_4038,N_1376,N_1337);
nor U4039 (N_4039,N_645,N_2320);
nor U4040 (N_4040,N_858,N_1692);
nand U4041 (N_4041,N_54,N_1169);
and U4042 (N_4042,N_2024,N_510);
nand U4043 (N_4043,N_1235,N_2767);
nand U4044 (N_4044,N_2343,N_2102);
nor U4045 (N_4045,N_880,N_881);
or U4046 (N_4046,N_1097,N_1645);
nand U4047 (N_4047,N_2286,N_1413);
and U4048 (N_4048,N_1089,N_2115);
and U4049 (N_4049,N_2031,N_118);
and U4050 (N_4050,N_2854,N_2175);
and U4051 (N_4051,N_1668,N_1297);
nor U4052 (N_4052,N_1878,N_1181);
nand U4053 (N_4053,N_808,N_2228);
nor U4054 (N_4054,N_2598,N_1813);
nand U4055 (N_4055,N_107,N_2515);
nand U4056 (N_4056,N_1070,N_413);
and U4057 (N_4057,N_187,N_1516);
nor U4058 (N_4058,N_2423,N_906);
and U4059 (N_4059,N_646,N_527);
and U4060 (N_4060,N_553,N_2601);
nand U4061 (N_4061,N_2871,N_1741);
and U4062 (N_4062,N_1405,N_1314);
nor U4063 (N_4063,N_1548,N_2804);
and U4064 (N_4064,N_2533,N_768);
nor U4065 (N_4065,N_39,N_529);
or U4066 (N_4066,N_727,N_1634);
and U4067 (N_4067,N_2771,N_1306);
or U4068 (N_4068,N_2722,N_2754);
nor U4069 (N_4069,N_2306,N_2184);
nor U4070 (N_4070,N_1525,N_2752);
nand U4071 (N_4071,N_1414,N_815);
nor U4072 (N_4072,N_2784,N_1246);
and U4073 (N_4073,N_514,N_192);
nor U4074 (N_4074,N_239,N_1698);
nand U4075 (N_4075,N_1659,N_805);
nor U4076 (N_4076,N_2939,N_1797);
nand U4077 (N_4077,N_2356,N_2923);
nor U4078 (N_4078,N_377,N_112);
nor U4079 (N_4079,N_418,N_1639);
or U4080 (N_4080,N_1085,N_2570);
nand U4081 (N_4081,N_2431,N_1108);
or U4082 (N_4082,N_573,N_1387);
nand U4083 (N_4083,N_2635,N_1498);
xnor U4084 (N_4084,N_2409,N_1834);
and U4085 (N_4085,N_234,N_656);
and U4086 (N_4086,N_1884,N_2846);
nor U4087 (N_4087,N_42,N_2817);
nand U4088 (N_4088,N_818,N_2105);
or U4089 (N_4089,N_2260,N_2067);
and U4090 (N_4090,N_2725,N_2521);
and U4091 (N_4091,N_434,N_2905);
nor U4092 (N_4092,N_1104,N_1553);
nor U4093 (N_4093,N_2894,N_585);
nand U4094 (N_4094,N_588,N_1534);
or U4095 (N_4095,N_944,N_2751);
and U4096 (N_4096,N_2482,N_2779);
nor U4097 (N_4097,N_2002,N_1318);
or U4098 (N_4098,N_1663,N_548);
nand U4099 (N_4099,N_1467,N_1442);
nor U4100 (N_4100,N_1119,N_437);
nand U4101 (N_4101,N_2978,N_350);
or U4102 (N_4102,N_1618,N_1508);
or U4103 (N_4103,N_255,N_2411);
nor U4104 (N_4104,N_2413,N_595);
nor U4105 (N_4105,N_190,N_2641);
nand U4106 (N_4106,N_1039,N_2153);
or U4107 (N_4107,N_171,N_2313);
and U4108 (N_4108,N_2419,N_1149);
and U4109 (N_4109,N_568,N_139);
nor U4110 (N_4110,N_1295,N_1276);
or U4111 (N_4111,N_1338,N_1788);
nor U4112 (N_4112,N_1350,N_1420);
nand U4113 (N_4113,N_2689,N_1586);
and U4114 (N_4114,N_1931,N_732);
or U4115 (N_4115,N_1766,N_1544);
xor U4116 (N_4116,N_335,N_581);
nor U4117 (N_4117,N_1957,N_1524);
nor U4118 (N_4118,N_53,N_2519);
nor U4119 (N_4119,N_939,N_2642);
or U4120 (N_4120,N_633,N_1940);
or U4121 (N_4121,N_1153,N_2070);
or U4122 (N_4122,N_2786,N_1551);
or U4123 (N_4123,N_227,N_2702);
nor U4124 (N_4124,N_1934,N_2165);
nand U4125 (N_4125,N_922,N_2416);
nor U4126 (N_4126,N_2972,N_2768);
nor U4127 (N_4127,N_1633,N_690);
nor U4128 (N_4128,N_1363,N_1989);
nand U4129 (N_4129,N_48,N_141);
or U4130 (N_4130,N_1738,N_2451);
and U4131 (N_4131,N_1082,N_1794);
nand U4132 (N_4132,N_1724,N_2294);
xor U4133 (N_4133,N_766,N_2542);
and U4134 (N_4134,N_4,N_2922);
and U4135 (N_4135,N_848,N_2701);
nand U4136 (N_4136,N_2456,N_1240);
or U4137 (N_4137,N_6,N_1069);
or U4138 (N_4138,N_57,N_2379);
or U4139 (N_4139,N_2889,N_473);
nor U4140 (N_4140,N_1557,N_309);
nand U4141 (N_4141,N_1453,N_1062);
nor U4142 (N_4142,N_316,N_1330);
nor U4143 (N_4143,N_651,N_2462);
nor U4144 (N_4144,N_1431,N_1683);
nand U4145 (N_4145,N_51,N_419);
nand U4146 (N_4146,N_2013,N_1160);
or U4147 (N_4147,N_1636,N_35);
or U4148 (N_4148,N_1988,N_2997);
or U4149 (N_4149,N_1915,N_660);
nor U4150 (N_4150,N_1059,N_949);
or U4151 (N_4151,N_2438,N_1677);
nand U4152 (N_4152,N_230,N_2326);
nor U4153 (N_4153,N_798,N_2695);
or U4154 (N_4154,N_1538,N_1061);
and U4155 (N_4155,N_1495,N_1904);
or U4156 (N_4156,N_1998,N_842);
nor U4157 (N_4157,N_1868,N_2372);
nand U4158 (N_4158,N_563,N_445);
or U4159 (N_4159,N_2464,N_2262);
nand U4160 (N_4160,N_2582,N_1311);
or U4161 (N_4161,N_2675,N_689);
nor U4162 (N_4162,N_1138,N_2106);
nor U4163 (N_4163,N_145,N_918);
nor U4164 (N_4164,N_2723,N_1666);
and U4165 (N_4165,N_1251,N_1800);
or U4166 (N_4166,N_738,N_1769);
nand U4167 (N_4167,N_2362,N_971);
nor U4168 (N_4168,N_2764,N_1333);
or U4169 (N_4169,N_1696,N_2555);
and U4170 (N_4170,N_2,N_380);
or U4171 (N_4171,N_1258,N_1648);
nor U4172 (N_4172,N_1135,N_2739);
and U4173 (N_4173,N_2776,N_1243);
nand U4174 (N_4174,N_2129,N_2606);
and U4175 (N_4175,N_607,N_333);
or U4176 (N_4176,N_1274,N_2248);
or U4177 (N_4177,N_1591,N_1962);
or U4178 (N_4178,N_151,N_1068);
nand U4179 (N_4179,N_2620,N_2243);
and U4180 (N_4180,N_2371,N_1919);
or U4181 (N_4181,N_1055,N_2337);
and U4182 (N_4182,N_1002,N_659);
nor U4183 (N_4183,N_71,N_952);
nor U4184 (N_4184,N_999,N_1593);
nand U4185 (N_4185,N_2300,N_1953);
or U4186 (N_4186,N_2710,N_807);
or U4187 (N_4187,N_1697,N_315);
nand U4188 (N_4188,N_355,N_1712);
nor U4189 (N_4189,N_210,N_1625);
and U4190 (N_4190,N_254,N_481);
nor U4191 (N_4191,N_1397,N_1502);
nor U4192 (N_4192,N_2323,N_492);
nor U4193 (N_4193,N_2189,N_1675);
and U4194 (N_4194,N_2487,N_1676);
and U4195 (N_4195,N_397,N_2836);
and U4196 (N_4196,N_2408,N_188);
and U4197 (N_4197,N_615,N_2224);
nor U4198 (N_4198,N_2467,N_873);
and U4199 (N_4199,N_294,N_1530);
nor U4200 (N_4200,N_2278,N_594);
nor U4201 (N_4201,N_1900,N_1755);
and U4202 (N_4202,N_2876,N_298);
nand U4203 (N_4203,N_832,N_2824);
nand U4204 (N_4204,N_286,N_910);
and U4205 (N_4205,N_2421,N_261);
nand U4206 (N_4206,N_2595,N_334);
or U4207 (N_4207,N_711,N_2703);
or U4208 (N_4208,N_2506,N_1567);
nor U4209 (N_4209,N_2927,N_1455);
and U4210 (N_4210,N_674,N_955);
nor U4211 (N_4211,N_464,N_1262);
or U4212 (N_4212,N_1402,N_2712);
and U4213 (N_4213,N_2812,N_708);
and U4214 (N_4214,N_1460,N_980);
or U4215 (N_4215,N_872,N_1821);
and U4216 (N_4216,N_1671,N_2862);
nor U4217 (N_4217,N_549,N_2732);
or U4218 (N_4218,N_2119,N_603);
nand U4219 (N_4219,N_504,N_1890);
or U4220 (N_4220,N_782,N_622);
and U4221 (N_4221,N_794,N_20);
nand U4222 (N_4222,N_623,N_1909);
nand U4223 (N_4223,N_2691,N_2333);
nor U4224 (N_4224,N_2898,N_2667);
nand U4225 (N_4225,N_501,N_1319);
nor U4226 (N_4226,N_2809,N_2258);
nor U4227 (N_4227,N_1278,N_2045);
nor U4228 (N_4228,N_2770,N_5);
and U4229 (N_4229,N_137,N_2942);
nor U4230 (N_4230,N_2265,N_2000);
and U4231 (N_4231,N_2389,N_2640);
and U4232 (N_4232,N_2748,N_748);
and U4233 (N_4233,N_836,N_546);
or U4234 (N_4234,N_44,N_304);
and U4235 (N_4235,N_2607,N_2864);
and U4236 (N_4236,N_2160,N_2156);
or U4237 (N_4237,N_1477,N_2298);
nor U4238 (N_4238,N_1300,N_783);
and U4239 (N_4239,N_666,N_148);
nand U4240 (N_4240,N_249,N_752);
nand U4241 (N_4241,N_1694,N_2267);
xor U4242 (N_4242,N_7,N_1543);
nor U4243 (N_4243,N_1264,N_2284);
or U4244 (N_4244,N_2047,N_2151);
nand U4245 (N_4245,N_528,N_410);
nor U4246 (N_4246,N_1034,N_1981);
or U4247 (N_4247,N_1617,N_2206);
or U4248 (N_4248,N_2319,N_2959);
nand U4249 (N_4249,N_231,N_2194);
and U4250 (N_4250,N_2721,N_109);
nand U4251 (N_4251,N_921,N_2011);
and U4252 (N_4252,N_1328,N_2316);
nand U4253 (N_4253,N_1221,N_1946);
or U4254 (N_4254,N_106,N_2264);
nor U4255 (N_4255,N_165,N_1856);
nor U4256 (N_4256,N_2615,N_1228);
and U4257 (N_4257,N_1054,N_1385);
nor U4258 (N_4258,N_977,N_2167);
nand U4259 (N_4259,N_1979,N_1820);
nand U4260 (N_4260,N_1759,N_2247);
nor U4261 (N_4261,N_1359,N_1781);
nand U4262 (N_4262,N_557,N_1729);
nor U4263 (N_4263,N_520,N_493);
nand U4264 (N_4264,N_947,N_2966);
or U4265 (N_4265,N_2763,N_1650);
nor U4266 (N_4266,N_908,N_1937);
and U4267 (N_4267,N_2310,N_1154);
and U4268 (N_4268,N_2207,N_985);
or U4269 (N_4269,N_438,N_641);
nor U4270 (N_4270,N_459,N_1606);
and U4271 (N_4271,N_429,N_793);
nor U4272 (N_4272,N_2856,N_1250);
or U4273 (N_4273,N_2293,N_1511);
nand U4274 (N_4274,N_777,N_1945);
and U4275 (N_4275,N_235,N_1930);
nand U4276 (N_4276,N_1127,N_2244);
nand U4277 (N_4277,N_426,N_76);
and U4278 (N_4278,N_1518,N_2485);
or U4279 (N_4279,N_1468,N_451);
or U4280 (N_4280,N_2619,N_265);
nand U4281 (N_4281,N_250,N_1541);
nand U4282 (N_4282,N_8,N_2390);
nand U4283 (N_4283,N_1867,N_2186);
nor U4284 (N_4284,N_2179,N_569);
nand U4285 (N_4285,N_2707,N_2017);
or U4286 (N_4286,N_1010,N_2384);
nand U4287 (N_4287,N_2484,N_2471);
and U4288 (N_4288,N_1924,N_203);
or U4289 (N_4289,N_828,N_1817);
nand U4290 (N_4290,N_928,N_61);
or U4291 (N_4291,N_1490,N_2037);
and U4292 (N_4292,N_1326,N_416);
and U4293 (N_4293,N_1454,N_311);
and U4294 (N_4294,N_2915,N_599);
or U4295 (N_4295,N_1956,N_935);
nand U4296 (N_4296,N_2891,N_1619);
nor U4297 (N_4297,N_2257,N_1462);
or U4298 (N_4298,N_854,N_2599);
or U4299 (N_4299,N_2954,N_2322);
nor U4300 (N_4300,N_443,N_138);
and U4301 (N_4301,N_1927,N_973);
nand U4302 (N_4302,N_1064,N_2199);
nand U4303 (N_4303,N_159,N_1339);
or U4304 (N_4304,N_1745,N_104);
or U4305 (N_4305,N_130,N_1629);
and U4306 (N_4306,N_1279,N_1207);
and U4307 (N_4307,N_2887,N_1238);
or U4308 (N_4308,N_435,N_2816);
nor U4309 (N_4309,N_229,N_1501);
and U4310 (N_4310,N_2537,N_202);
and U4311 (N_4311,N_1321,N_469);
or U4312 (N_4312,N_754,N_2636);
and U4313 (N_4313,N_405,N_18);
nor U4314 (N_4314,N_822,N_1);
nand U4315 (N_4315,N_2909,N_2673);
nand U4316 (N_4316,N_1234,N_2610);
or U4317 (N_4317,N_1080,N_1499);
nor U4318 (N_4318,N_2198,N_1791);
or U4319 (N_4319,N_2122,N_1042);
and U4320 (N_4320,N_2196,N_804);
nand U4321 (N_4321,N_1872,N_761);
and U4322 (N_4322,N_2861,N_181);
and U4323 (N_4323,N_2743,N_2352);
nand U4324 (N_4324,N_1757,N_278);
nand U4325 (N_4325,N_912,N_574);
nor U4326 (N_4326,N_2977,N_2955);
nor U4327 (N_4327,N_1147,N_1552);
nor U4328 (N_4328,N_70,N_1213);
or U4329 (N_4329,N_861,N_2904);
nor U4330 (N_4330,N_1194,N_2123);
nand U4331 (N_4331,N_2845,N_88);
nor U4332 (N_4332,N_1740,N_1982);
nand U4333 (N_4333,N_2368,N_1807);
or U4334 (N_4334,N_1211,N_1664);
or U4335 (N_4335,N_33,N_2237);
and U4336 (N_4336,N_1976,N_650);
and U4337 (N_4337,N_406,N_976);
or U4338 (N_4338,N_712,N_78);
nand U4339 (N_4339,N_583,N_2746);
nor U4340 (N_4340,N_2078,N_2841);
nand U4341 (N_4341,N_2669,N_2136);
nand U4342 (N_4342,N_2639,N_1098);
nor U4343 (N_4343,N_2654,N_1093);
nor U4344 (N_4344,N_1563,N_1496);
or U4345 (N_4345,N_1304,N_1830);
or U4346 (N_4346,N_2208,N_2452);
and U4347 (N_4347,N_2018,N_2860);
and U4348 (N_4348,N_1134,N_2187);
nor U4349 (N_4349,N_817,N_1367);
and U4350 (N_4350,N_884,N_2563);
nor U4351 (N_4351,N_576,N_2035);
nor U4352 (N_4352,N_1810,N_1099);
nor U4353 (N_4353,N_1889,N_2617);
nand U4354 (N_4354,N_1605,N_1429);
nand U4355 (N_4355,N_388,N_1540);
xor U4356 (N_4356,N_2022,N_1597);
nand U4357 (N_4357,N_1536,N_1435);
nor U4358 (N_4358,N_1681,N_1635);
nand U4359 (N_4359,N_1027,N_813);
or U4360 (N_4360,N_1941,N_2147);
and U4361 (N_4361,N_865,N_1045);
nor U4362 (N_4362,N_2330,N_965);
nand U4363 (N_4363,N_998,N_1614);
or U4364 (N_4364,N_275,N_1230);
and U4365 (N_4365,N_1489,N_2562);
nand U4366 (N_4366,N_2717,N_1728);
xor U4367 (N_4367,N_1928,N_1178);
nand U4368 (N_4368,N_1056,N_2747);
nand U4369 (N_4369,N_992,N_1164);
and U4370 (N_4370,N_655,N_892);
and U4371 (N_4371,N_2334,N_1163);
or U4372 (N_4372,N_1371,N_1611);
or U4373 (N_4373,N_1461,N_713);
nor U4374 (N_4374,N_2744,N_2525);
nor U4375 (N_4375,N_2302,N_1993);
nand U4376 (N_4376,N_974,N_2803);
and U4377 (N_4377,N_1521,N_2162);
or U4378 (N_4378,N_1587,N_741);
nand U4379 (N_4379,N_2823,N_427);
or U4380 (N_4380,N_1920,N_1823);
or U4381 (N_4381,N_1474,N_1554);
nand U4382 (N_4382,N_2209,N_1393);
nand U4383 (N_4383,N_891,N_1003);
and U4384 (N_4384,N_925,N_1913);
nand U4385 (N_4385,N_780,N_2439);
and U4386 (N_4386,N_1036,N_65);
nor U4387 (N_4387,N_978,N_2381);
or U4388 (N_4388,N_1115,N_1217);
and U4389 (N_4389,N_2938,N_2785);
nand U4390 (N_4390,N_506,N_68);
nand U4391 (N_4391,N_1275,N_1709);
or U4392 (N_4392,N_1647,N_2019);
or U4393 (N_4393,N_876,N_1768);
nand U4394 (N_4394,N_1327,N_2245);
and U4395 (N_4395,N_2806,N_1060);
and U4396 (N_4396,N_1308,N_1025);
nor U4397 (N_4397,N_2692,N_2650);
nor U4398 (N_4398,N_1334,N_715);
nand U4399 (N_4399,N_444,N_62);
and U4400 (N_4400,N_740,N_1368);
nand U4401 (N_4401,N_616,N_2708);
and U4402 (N_4402,N_2437,N_1482);
nand U4403 (N_4403,N_292,N_2578);
nand U4404 (N_4404,N_2049,N_990);
nand U4405 (N_4405,N_1176,N_2567);
nor U4406 (N_4406,N_1708,N_2201);
and U4407 (N_4407,N_2346,N_1191);
nand U4408 (N_4408,N_2780,N_937);
or U4409 (N_4409,N_693,N_1458);
or U4410 (N_4410,N_1804,N_1786);
or U4411 (N_4411,N_1870,N_758);
and U4412 (N_4412,N_1644,N_1503);
xnor U4413 (N_4413,N_194,N_1220);
nor U4414 (N_4414,N_256,N_1284);
or U4415 (N_4415,N_2427,N_809);
and U4416 (N_4416,N_179,N_2061);
or U4417 (N_4417,N_1411,N_2679);
nand U4418 (N_4418,N_2289,N_888);
nand U4419 (N_4419,N_185,N_1801);
nand U4420 (N_4420,N_237,N_128);
or U4421 (N_4421,N_360,N_1542);
nor U4422 (N_4422,N_849,N_1016);
and U4423 (N_4423,N_2012,N_1526);
nand U4424 (N_4424,N_1665,N_1812);
nor U4425 (N_4425,N_101,N_575);
or U4426 (N_4426,N_160,N_948);
nor U4427 (N_4427,N_2957,N_913);
nor U4428 (N_4428,N_1906,N_1231);
or U4429 (N_4429,N_1649,N_1848);
xnor U4430 (N_4430,N_1451,N_1001);
or U4431 (N_4431,N_272,N_541);
nor U4432 (N_4432,N_706,N_1710);
nor U4433 (N_4433,N_423,N_1212);
or U4434 (N_4434,N_301,N_614);
nand U4435 (N_4435,N_1236,N_2981);
nor U4436 (N_4436,N_2461,N_2315);
or U4437 (N_4437,N_1374,N_1004);
or U4438 (N_4438,N_2858,N_43);
nor U4439 (N_4439,N_765,N_2956);
nor U4440 (N_4440,N_1343,N_251);
nand U4441 (N_4441,N_2071,N_446);
nor U4442 (N_4442,N_28,N_2503);
nand U4443 (N_4443,N_302,N_1887);
and U4444 (N_4444,N_1505,N_2733);
nand U4445 (N_4445,N_2028,N_245);
nand U4446 (N_4446,N_1869,N_2745);
nand U4447 (N_4447,N_2660,N_2420);
and U4448 (N_4448,N_341,N_790);
or U4449 (N_4449,N_2074,N_2560);
and U4450 (N_4450,N_2808,N_770);
or U4451 (N_4451,N_322,N_1590);
nor U4452 (N_4452,N_2127,N_2093);
or U4453 (N_4453,N_737,N_1095);
nand U4454 (N_4454,N_1602,N_2951);
or U4455 (N_4455,N_1674,N_1344);
or U4456 (N_4456,N_431,N_2103);
nor U4457 (N_4457,N_2367,N_2053);
nand U4458 (N_4458,N_932,N_1116);
or U4459 (N_4459,N_2947,N_951);
and U4460 (N_4460,N_1562,N_200);
nand U4461 (N_4461,N_648,N_1938);
or U4462 (N_4462,N_2422,N_605);
nor U4463 (N_4463,N_987,N_682);
or U4464 (N_4464,N_1961,N_1959);
or U4465 (N_4465,N_1861,N_296);
or U4466 (N_4466,N_2643,N_1925);
and U4467 (N_4467,N_2251,N_96);
xor U4468 (N_4468,N_2524,N_1345);
nand U4469 (N_4469,N_1529,N_2872);
nand U4470 (N_4470,N_2730,N_2929);
and U4471 (N_4471,N_1707,N_1785);
and U4472 (N_4472,N_1852,N_232);
and U4473 (N_4473,N_1043,N_270);
nand U4474 (N_4474,N_488,N_1185);
nand U4475 (N_4475,N_887,N_1428);
and U4476 (N_4476,N_2038,N_2065);
and U4477 (N_4477,N_618,N_2908);
or U4478 (N_4478,N_1809,N_550);
or U4479 (N_4479,N_1589,N_806);
nand U4480 (N_4480,N_1992,N_1139);
and U4481 (N_4481,N_1476,N_2961);
nor U4482 (N_4482,N_2020,N_339);
nand U4483 (N_4483,N_1456,N_1954);
or U4484 (N_4484,N_863,N_2863);
and U4485 (N_4485,N_348,N_2911);
nand U4486 (N_4486,N_86,N_2755);
and U4487 (N_4487,N_868,N_1744);
and U4488 (N_4488,N_114,N_1366);
nor U4489 (N_4489,N_2096,N_257);
nand U4490 (N_4490,N_2838,N_1075);
and U4491 (N_4491,N_703,N_1349);
and U4492 (N_4492,N_2866,N_2350);
or U4493 (N_4493,N_2742,N_1265);
and U4494 (N_4494,N_1624,N_2085);
or U4495 (N_4495,N_2397,N_365);
nand U4496 (N_4496,N_2307,N_2373);
and U4497 (N_4497,N_2010,N_628);
nand U4498 (N_4498,N_1730,N_1266);
nand U4499 (N_4499,N_1487,N_843);
nand U4500 (N_4500,N_2569,N_1249);
nand U4501 (N_4501,N_1641,N_2867);
or U4502 (N_4502,N_723,N_2037);
nor U4503 (N_4503,N_2806,N_598);
and U4504 (N_4504,N_208,N_371);
nor U4505 (N_4505,N_7,N_1606);
or U4506 (N_4506,N_1929,N_2341);
or U4507 (N_4507,N_2997,N_2948);
and U4508 (N_4508,N_1399,N_1414);
nand U4509 (N_4509,N_1173,N_2869);
and U4510 (N_4510,N_363,N_1170);
or U4511 (N_4511,N_1833,N_2717);
nand U4512 (N_4512,N_1041,N_262);
nor U4513 (N_4513,N_1739,N_1738);
nand U4514 (N_4514,N_1697,N_831);
or U4515 (N_4515,N_563,N_244);
and U4516 (N_4516,N_394,N_43);
and U4517 (N_4517,N_432,N_184);
nand U4518 (N_4518,N_952,N_2686);
nand U4519 (N_4519,N_1349,N_2722);
or U4520 (N_4520,N_1902,N_998);
or U4521 (N_4521,N_1935,N_1975);
nor U4522 (N_4522,N_1286,N_84);
or U4523 (N_4523,N_845,N_2816);
nand U4524 (N_4524,N_1543,N_2128);
and U4525 (N_4525,N_1099,N_1434);
or U4526 (N_4526,N_768,N_2743);
or U4527 (N_4527,N_2527,N_2416);
or U4528 (N_4528,N_1912,N_1688);
and U4529 (N_4529,N_929,N_918);
nor U4530 (N_4530,N_2990,N_1961);
nor U4531 (N_4531,N_2023,N_2755);
or U4532 (N_4532,N_655,N_2940);
and U4533 (N_4533,N_1128,N_1488);
and U4534 (N_4534,N_685,N_647);
and U4535 (N_4535,N_323,N_1373);
nand U4536 (N_4536,N_1705,N_1453);
nand U4537 (N_4537,N_1009,N_2292);
or U4538 (N_4538,N_550,N_1201);
or U4539 (N_4539,N_441,N_828);
or U4540 (N_4540,N_2351,N_2902);
or U4541 (N_4541,N_1049,N_2181);
nor U4542 (N_4542,N_974,N_2390);
nand U4543 (N_4543,N_1033,N_536);
nand U4544 (N_4544,N_1608,N_995);
or U4545 (N_4545,N_2797,N_2811);
nand U4546 (N_4546,N_2014,N_1783);
nor U4547 (N_4547,N_149,N_281);
and U4548 (N_4548,N_1170,N_1655);
nand U4549 (N_4549,N_979,N_2497);
and U4550 (N_4550,N_1887,N_890);
nor U4551 (N_4551,N_2224,N_2317);
nor U4552 (N_4552,N_119,N_2228);
or U4553 (N_4553,N_324,N_2878);
or U4554 (N_4554,N_2082,N_381);
and U4555 (N_4555,N_702,N_2604);
or U4556 (N_4556,N_1887,N_526);
and U4557 (N_4557,N_29,N_1347);
or U4558 (N_4558,N_2668,N_1864);
or U4559 (N_4559,N_1332,N_1018);
or U4560 (N_4560,N_1535,N_2361);
nand U4561 (N_4561,N_995,N_194);
nor U4562 (N_4562,N_46,N_1776);
and U4563 (N_4563,N_2466,N_962);
and U4564 (N_4564,N_2528,N_1077);
nand U4565 (N_4565,N_2706,N_2044);
nor U4566 (N_4566,N_82,N_1050);
or U4567 (N_4567,N_2061,N_478);
or U4568 (N_4568,N_783,N_1231);
or U4569 (N_4569,N_2211,N_1831);
nor U4570 (N_4570,N_544,N_1312);
xnor U4571 (N_4571,N_1349,N_55);
and U4572 (N_4572,N_1566,N_1578);
nand U4573 (N_4573,N_1454,N_1266);
nand U4574 (N_4574,N_411,N_124);
nor U4575 (N_4575,N_2653,N_1645);
and U4576 (N_4576,N_2043,N_1175);
nor U4577 (N_4577,N_2777,N_359);
nor U4578 (N_4578,N_1685,N_2530);
nor U4579 (N_4579,N_1594,N_1080);
nor U4580 (N_4580,N_2318,N_372);
and U4581 (N_4581,N_587,N_604);
and U4582 (N_4582,N_970,N_595);
and U4583 (N_4583,N_2323,N_1631);
or U4584 (N_4584,N_2657,N_2764);
and U4585 (N_4585,N_1429,N_305);
nor U4586 (N_4586,N_234,N_550);
nor U4587 (N_4587,N_1391,N_486);
nand U4588 (N_4588,N_1384,N_807);
nor U4589 (N_4589,N_901,N_628);
or U4590 (N_4590,N_2623,N_366);
or U4591 (N_4591,N_690,N_2951);
or U4592 (N_4592,N_526,N_2038);
or U4593 (N_4593,N_40,N_594);
nand U4594 (N_4594,N_120,N_2632);
nand U4595 (N_4595,N_801,N_591);
nor U4596 (N_4596,N_256,N_977);
nor U4597 (N_4597,N_1624,N_402);
nand U4598 (N_4598,N_1490,N_644);
and U4599 (N_4599,N_974,N_1040);
and U4600 (N_4600,N_1516,N_2985);
or U4601 (N_4601,N_2793,N_814);
or U4602 (N_4602,N_1118,N_1686);
nand U4603 (N_4603,N_689,N_2046);
nor U4604 (N_4604,N_283,N_600);
or U4605 (N_4605,N_25,N_2645);
and U4606 (N_4606,N_1728,N_979);
or U4607 (N_4607,N_1748,N_2315);
or U4608 (N_4608,N_374,N_826);
and U4609 (N_4609,N_2984,N_2851);
or U4610 (N_4610,N_597,N_312);
and U4611 (N_4611,N_96,N_2187);
or U4612 (N_4612,N_1938,N_2097);
or U4613 (N_4613,N_139,N_2008);
nor U4614 (N_4614,N_98,N_446);
nand U4615 (N_4615,N_1544,N_2295);
and U4616 (N_4616,N_1499,N_1898);
and U4617 (N_4617,N_2967,N_621);
and U4618 (N_4618,N_528,N_906);
nand U4619 (N_4619,N_2532,N_2775);
nand U4620 (N_4620,N_1200,N_1578);
nor U4621 (N_4621,N_2479,N_1175);
or U4622 (N_4622,N_1142,N_2411);
nand U4623 (N_4623,N_1893,N_2645);
nor U4624 (N_4624,N_1190,N_1061);
or U4625 (N_4625,N_2224,N_476);
and U4626 (N_4626,N_49,N_2318);
nor U4627 (N_4627,N_1607,N_2685);
and U4628 (N_4628,N_1271,N_302);
and U4629 (N_4629,N_1544,N_719);
and U4630 (N_4630,N_1187,N_2764);
nand U4631 (N_4631,N_356,N_2186);
and U4632 (N_4632,N_1183,N_2345);
and U4633 (N_4633,N_1380,N_402);
and U4634 (N_4634,N_1302,N_2374);
and U4635 (N_4635,N_624,N_2822);
and U4636 (N_4636,N_1264,N_2957);
nor U4637 (N_4637,N_1591,N_1669);
or U4638 (N_4638,N_107,N_614);
or U4639 (N_4639,N_1932,N_617);
nor U4640 (N_4640,N_1643,N_1937);
xor U4641 (N_4641,N_2175,N_2465);
nor U4642 (N_4642,N_901,N_753);
nand U4643 (N_4643,N_478,N_1502);
and U4644 (N_4644,N_353,N_1492);
nor U4645 (N_4645,N_577,N_1685);
and U4646 (N_4646,N_369,N_1238);
or U4647 (N_4647,N_2785,N_799);
and U4648 (N_4648,N_2666,N_1095);
and U4649 (N_4649,N_262,N_789);
nor U4650 (N_4650,N_433,N_175);
nand U4651 (N_4651,N_897,N_2547);
and U4652 (N_4652,N_1356,N_748);
nand U4653 (N_4653,N_627,N_2523);
or U4654 (N_4654,N_372,N_529);
and U4655 (N_4655,N_2248,N_2423);
nand U4656 (N_4656,N_1473,N_2024);
nor U4657 (N_4657,N_2377,N_1562);
and U4658 (N_4658,N_2057,N_1621);
or U4659 (N_4659,N_1201,N_713);
and U4660 (N_4660,N_1016,N_2352);
or U4661 (N_4661,N_2110,N_1071);
nand U4662 (N_4662,N_2925,N_2002);
nor U4663 (N_4663,N_966,N_2033);
nand U4664 (N_4664,N_1059,N_1959);
or U4665 (N_4665,N_1059,N_1262);
nor U4666 (N_4666,N_852,N_1309);
nand U4667 (N_4667,N_2586,N_1212);
and U4668 (N_4668,N_1528,N_2613);
nand U4669 (N_4669,N_128,N_160);
nor U4670 (N_4670,N_2636,N_677);
and U4671 (N_4671,N_1235,N_1345);
nand U4672 (N_4672,N_2767,N_223);
nor U4673 (N_4673,N_771,N_163);
nor U4674 (N_4674,N_1395,N_244);
nand U4675 (N_4675,N_2225,N_1593);
and U4676 (N_4676,N_1828,N_746);
and U4677 (N_4677,N_599,N_1036);
and U4678 (N_4678,N_435,N_1039);
nand U4679 (N_4679,N_2291,N_884);
nand U4680 (N_4680,N_454,N_2118);
nor U4681 (N_4681,N_1036,N_1796);
nand U4682 (N_4682,N_278,N_1079);
nand U4683 (N_4683,N_1730,N_1666);
nor U4684 (N_4684,N_446,N_2561);
or U4685 (N_4685,N_213,N_2400);
and U4686 (N_4686,N_78,N_1974);
or U4687 (N_4687,N_2388,N_2862);
and U4688 (N_4688,N_1826,N_2222);
and U4689 (N_4689,N_1271,N_1925);
and U4690 (N_4690,N_2526,N_1722);
and U4691 (N_4691,N_2414,N_1239);
nor U4692 (N_4692,N_2395,N_756);
and U4693 (N_4693,N_1766,N_119);
and U4694 (N_4694,N_1456,N_2387);
nor U4695 (N_4695,N_1241,N_1228);
nor U4696 (N_4696,N_687,N_994);
or U4697 (N_4697,N_1308,N_1839);
and U4698 (N_4698,N_1742,N_1168);
nand U4699 (N_4699,N_1441,N_2049);
nor U4700 (N_4700,N_1495,N_1308);
nor U4701 (N_4701,N_2373,N_700);
or U4702 (N_4702,N_1487,N_726);
or U4703 (N_4703,N_748,N_1069);
or U4704 (N_4704,N_1105,N_1885);
and U4705 (N_4705,N_1475,N_94);
nor U4706 (N_4706,N_974,N_313);
and U4707 (N_4707,N_1082,N_419);
or U4708 (N_4708,N_1334,N_473);
and U4709 (N_4709,N_1832,N_1556);
nor U4710 (N_4710,N_411,N_2457);
nor U4711 (N_4711,N_2848,N_1503);
nor U4712 (N_4712,N_499,N_2025);
or U4713 (N_4713,N_2674,N_499);
nand U4714 (N_4714,N_865,N_788);
nor U4715 (N_4715,N_381,N_435);
or U4716 (N_4716,N_2365,N_662);
nand U4717 (N_4717,N_2714,N_735);
nor U4718 (N_4718,N_2001,N_2897);
nand U4719 (N_4719,N_856,N_2855);
nand U4720 (N_4720,N_1356,N_1980);
nor U4721 (N_4721,N_1653,N_670);
nand U4722 (N_4722,N_513,N_1462);
nand U4723 (N_4723,N_2873,N_2175);
and U4724 (N_4724,N_744,N_2250);
or U4725 (N_4725,N_2440,N_2576);
nor U4726 (N_4726,N_1730,N_579);
or U4727 (N_4727,N_2400,N_1121);
nor U4728 (N_4728,N_576,N_1262);
nor U4729 (N_4729,N_2102,N_1291);
nor U4730 (N_4730,N_2046,N_1215);
nor U4731 (N_4731,N_1923,N_802);
and U4732 (N_4732,N_2861,N_1590);
or U4733 (N_4733,N_906,N_1787);
nand U4734 (N_4734,N_1836,N_2945);
nor U4735 (N_4735,N_150,N_200);
and U4736 (N_4736,N_2928,N_1895);
or U4737 (N_4737,N_2580,N_405);
nand U4738 (N_4738,N_1054,N_41);
nor U4739 (N_4739,N_2234,N_1334);
nand U4740 (N_4740,N_2932,N_939);
and U4741 (N_4741,N_647,N_631);
nand U4742 (N_4742,N_937,N_691);
nand U4743 (N_4743,N_2723,N_2267);
nor U4744 (N_4744,N_1438,N_66);
or U4745 (N_4745,N_113,N_1572);
nand U4746 (N_4746,N_162,N_2216);
and U4747 (N_4747,N_413,N_804);
nand U4748 (N_4748,N_1322,N_946);
and U4749 (N_4749,N_1613,N_10);
nor U4750 (N_4750,N_993,N_2474);
nor U4751 (N_4751,N_1633,N_2050);
xnor U4752 (N_4752,N_2853,N_1654);
nand U4753 (N_4753,N_2605,N_332);
nand U4754 (N_4754,N_1519,N_1786);
nor U4755 (N_4755,N_612,N_900);
nand U4756 (N_4756,N_533,N_2685);
or U4757 (N_4757,N_867,N_2690);
or U4758 (N_4758,N_2195,N_1919);
and U4759 (N_4759,N_2489,N_2404);
nand U4760 (N_4760,N_2798,N_393);
and U4761 (N_4761,N_2022,N_1100);
or U4762 (N_4762,N_1252,N_2061);
and U4763 (N_4763,N_142,N_1664);
and U4764 (N_4764,N_2050,N_2122);
or U4765 (N_4765,N_597,N_2942);
and U4766 (N_4766,N_2626,N_2928);
or U4767 (N_4767,N_1468,N_1134);
nor U4768 (N_4768,N_2453,N_2571);
and U4769 (N_4769,N_2897,N_1701);
nand U4770 (N_4770,N_53,N_270);
or U4771 (N_4771,N_1015,N_409);
nand U4772 (N_4772,N_1364,N_1004);
and U4773 (N_4773,N_1654,N_1385);
nand U4774 (N_4774,N_2554,N_2468);
nor U4775 (N_4775,N_1453,N_1878);
or U4776 (N_4776,N_2860,N_2272);
nor U4777 (N_4777,N_2040,N_1866);
nand U4778 (N_4778,N_1488,N_2261);
or U4779 (N_4779,N_958,N_1266);
and U4780 (N_4780,N_1921,N_970);
nor U4781 (N_4781,N_52,N_970);
nand U4782 (N_4782,N_2886,N_2524);
nand U4783 (N_4783,N_112,N_223);
nand U4784 (N_4784,N_1052,N_861);
nand U4785 (N_4785,N_1773,N_1650);
xnor U4786 (N_4786,N_2756,N_1561);
and U4787 (N_4787,N_1002,N_2636);
nor U4788 (N_4788,N_79,N_1988);
xor U4789 (N_4789,N_1870,N_45);
nand U4790 (N_4790,N_1543,N_2278);
and U4791 (N_4791,N_1406,N_1908);
nand U4792 (N_4792,N_1048,N_316);
or U4793 (N_4793,N_567,N_1078);
and U4794 (N_4794,N_266,N_2969);
and U4795 (N_4795,N_605,N_1616);
nor U4796 (N_4796,N_2259,N_1453);
nor U4797 (N_4797,N_428,N_2280);
nand U4798 (N_4798,N_238,N_1079);
nor U4799 (N_4799,N_2887,N_1218);
or U4800 (N_4800,N_1021,N_2816);
nor U4801 (N_4801,N_425,N_1862);
nor U4802 (N_4802,N_2146,N_2537);
nand U4803 (N_4803,N_1761,N_448);
nand U4804 (N_4804,N_1149,N_877);
nor U4805 (N_4805,N_697,N_805);
nor U4806 (N_4806,N_1022,N_481);
nand U4807 (N_4807,N_2871,N_2616);
nand U4808 (N_4808,N_1568,N_557);
nand U4809 (N_4809,N_469,N_2998);
and U4810 (N_4810,N_368,N_2235);
nand U4811 (N_4811,N_2297,N_2251);
nor U4812 (N_4812,N_2294,N_2736);
and U4813 (N_4813,N_860,N_1377);
nand U4814 (N_4814,N_884,N_2172);
or U4815 (N_4815,N_2896,N_2081);
or U4816 (N_4816,N_608,N_2775);
nand U4817 (N_4817,N_2044,N_745);
or U4818 (N_4818,N_534,N_464);
or U4819 (N_4819,N_215,N_1977);
and U4820 (N_4820,N_2211,N_1394);
nand U4821 (N_4821,N_2779,N_2669);
nor U4822 (N_4822,N_725,N_1423);
nor U4823 (N_4823,N_967,N_995);
or U4824 (N_4824,N_465,N_711);
nor U4825 (N_4825,N_954,N_2167);
or U4826 (N_4826,N_313,N_2902);
nand U4827 (N_4827,N_2291,N_1213);
and U4828 (N_4828,N_948,N_2311);
nand U4829 (N_4829,N_60,N_768);
nor U4830 (N_4830,N_1916,N_422);
or U4831 (N_4831,N_2546,N_1979);
or U4832 (N_4832,N_1233,N_2545);
and U4833 (N_4833,N_641,N_2507);
nor U4834 (N_4834,N_69,N_605);
nor U4835 (N_4835,N_1684,N_1035);
nor U4836 (N_4836,N_2931,N_1473);
nor U4837 (N_4837,N_61,N_809);
and U4838 (N_4838,N_599,N_1934);
and U4839 (N_4839,N_760,N_301);
nand U4840 (N_4840,N_1940,N_2635);
nor U4841 (N_4841,N_2850,N_1068);
and U4842 (N_4842,N_2623,N_539);
and U4843 (N_4843,N_2099,N_173);
nand U4844 (N_4844,N_2711,N_2565);
nor U4845 (N_4845,N_2163,N_610);
nor U4846 (N_4846,N_2261,N_1610);
nor U4847 (N_4847,N_2659,N_681);
or U4848 (N_4848,N_2575,N_2110);
and U4849 (N_4849,N_2828,N_795);
or U4850 (N_4850,N_1825,N_2747);
nand U4851 (N_4851,N_2052,N_950);
or U4852 (N_4852,N_1139,N_1185);
and U4853 (N_4853,N_1280,N_797);
nand U4854 (N_4854,N_1819,N_2786);
nor U4855 (N_4855,N_941,N_1873);
or U4856 (N_4856,N_1921,N_2260);
nor U4857 (N_4857,N_2818,N_724);
and U4858 (N_4858,N_71,N_1290);
or U4859 (N_4859,N_2849,N_977);
nand U4860 (N_4860,N_2339,N_1918);
nand U4861 (N_4861,N_1867,N_1403);
nor U4862 (N_4862,N_528,N_848);
nand U4863 (N_4863,N_1920,N_1527);
nand U4864 (N_4864,N_384,N_543);
nand U4865 (N_4865,N_2952,N_825);
nor U4866 (N_4866,N_2283,N_700);
and U4867 (N_4867,N_1605,N_2466);
or U4868 (N_4868,N_1899,N_1513);
nor U4869 (N_4869,N_1325,N_1266);
nor U4870 (N_4870,N_1171,N_1857);
nor U4871 (N_4871,N_1761,N_2221);
nor U4872 (N_4872,N_370,N_939);
nor U4873 (N_4873,N_33,N_2214);
nor U4874 (N_4874,N_328,N_1705);
or U4875 (N_4875,N_1969,N_2225);
nand U4876 (N_4876,N_1900,N_238);
nand U4877 (N_4877,N_528,N_1838);
nand U4878 (N_4878,N_2010,N_116);
nand U4879 (N_4879,N_2354,N_1580);
nand U4880 (N_4880,N_752,N_1206);
and U4881 (N_4881,N_2547,N_1287);
and U4882 (N_4882,N_1408,N_124);
and U4883 (N_4883,N_19,N_857);
or U4884 (N_4884,N_2373,N_1401);
or U4885 (N_4885,N_175,N_375);
nor U4886 (N_4886,N_1930,N_238);
or U4887 (N_4887,N_2033,N_1624);
nor U4888 (N_4888,N_1877,N_2580);
and U4889 (N_4889,N_415,N_2232);
or U4890 (N_4890,N_2747,N_2314);
and U4891 (N_4891,N_86,N_1102);
or U4892 (N_4892,N_727,N_733);
xnor U4893 (N_4893,N_1202,N_29);
nor U4894 (N_4894,N_106,N_1451);
nand U4895 (N_4895,N_1803,N_1437);
nor U4896 (N_4896,N_1596,N_2225);
or U4897 (N_4897,N_2360,N_1698);
nor U4898 (N_4898,N_1285,N_1610);
nand U4899 (N_4899,N_1705,N_1645);
or U4900 (N_4900,N_281,N_590);
and U4901 (N_4901,N_1715,N_1764);
and U4902 (N_4902,N_2790,N_286);
nand U4903 (N_4903,N_2457,N_600);
or U4904 (N_4904,N_1069,N_261);
nand U4905 (N_4905,N_2456,N_2056);
and U4906 (N_4906,N_1882,N_506);
or U4907 (N_4907,N_1156,N_312);
nor U4908 (N_4908,N_548,N_875);
and U4909 (N_4909,N_1818,N_2961);
nor U4910 (N_4910,N_724,N_1851);
and U4911 (N_4911,N_184,N_874);
nand U4912 (N_4912,N_2287,N_1385);
and U4913 (N_4913,N_104,N_140);
nor U4914 (N_4914,N_1157,N_206);
and U4915 (N_4915,N_1688,N_1183);
or U4916 (N_4916,N_1164,N_2484);
nor U4917 (N_4917,N_2348,N_2682);
and U4918 (N_4918,N_2456,N_238);
or U4919 (N_4919,N_837,N_1617);
nor U4920 (N_4920,N_2179,N_782);
and U4921 (N_4921,N_1012,N_1201);
or U4922 (N_4922,N_2650,N_2856);
or U4923 (N_4923,N_2660,N_2591);
and U4924 (N_4924,N_224,N_1424);
or U4925 (N_4925,N_1797,N_886);
nor U4926 (N_4926,N_884,N_419);
and U4927 (N_4927,N_2682,N_2234);
nand U4928 (N_4928,N_2566,N_1418);
and U4929 (N_4929,N_874,N_2572);
and U4930 (N_4930,N_102,N_241);
and U4931 (N_4931,N_2911,N_488);
nor U4932 (N_4932,N_1779,N_427);
and U4933 (N_4933,N_2042,N_2764);
nand U4934 (N_4934,N_1525,N_2478);
or U4935 (N_4935,N_301,N_157);
nand U4936 (N_4936,N_705,N_1138);
xnor U4937 (N_4937,N_541,N_2088);
and U4938 (N_4938,N_1033,N_479);
and U4939 (N_4939,N_876,N_501);
and U4940 (N_4940,N_1019,N_2683);
or U4941 (N_4941,N_2691,N_1474);
nand U4942 (N_4942,N_1315,N_1771);
and U4943 (N_4943,N_2104,N_4);
nor U4944 (N_4944,N_1757,N_1029);
nor U4945 (N_4945,N_2022,N_1320);
nor U4946 (N_4946,N_2188,N_1029);
nor U4947 (N_4947,N_1619,N_1252);
and U4948 (N_4948,N_2117,N_1197);
nand U4949 (N_4949,N_2470,N_33);
and U4950 (N_4950,N_2988,N_2804);
or U4951 (N_4951,N_2479,N_1597);
nand U4952 (N_4952,N_2071,N_2365);
nor U4953 (N_4953,N_587,N_2401);
and U4954 (N_4954,N_2988,N_2827);
nand U4955 (N_4955,N_2047,N_1671);
and U4956 (N_4956,N_2861,N_519);
and U4957 (N_4957,N_454,N_691);
or U4958 (N_4958,N_613,N_976);
or U4959 (N_4959,N_1435,N_2299);
or U4960 (N_4960,N_2371,N_1336);
and U4961 (N_4961,N_1959,N_867);
nand U4962 (N_4962,N_589,N_2652);
or U4963 (N_4963,N_1967,N_209);
nand U4964 (N_4964,N_158,N_2269);
or U4965 (N_4965,N_2734,N_1046);
or U4966 (N_4966,N_1078,N_1702);
nor U4967 (N_4967,N_1225,N_1420);
nor U4968 (N_4968,N_948,N_971);
nor U4969 (N_4969,N_1361,N_1400);
or U4970 (N_4970,N_1938,N_1451);
and U4971 (N_4971,N_737,N_891);
nor U4972 (N_4972,N_114,N_787);
or U4973 (N_4973,N_1304,N_2559);
or U4974 (N_4974,N_2647,N_1227);
or U4975 (N_4975,N_1837,N_1845);
nor U4976 (N_4976,N_291,N_567);
nor U4977 (N_4977,N_1351,N_814);
and U4978 (N_4978,N_1009,N_2006);
and U4979 (N_4979,N_357,N_121);
or U4980 (N_4980,N_2713,N_1454);
or U4981 (N_4981,N_424,N_1473);
nor U4982 (N_4982,N_2169,N_2881);
or U4983 (N_4983,N_2048,N_228);
or U4984 (N_4984,N_2195,N_1181);
or U4985 (N_4985,N_2144,N_2476);
nor U4986 (N_4986,N_2068,N_1970);
nand U4987 (N_4987,N_2189,N_1398);
or U4988 (N_4988,N_1600,N_359);
or U4989 (N_4989,N_2088,N_300);
nand U4990 (N_4990,N_1068,N_2011);
nor U4991 (N_4991,N_675,N_2897);
or U4992 (N_4992,N_880,N_2237);
nor U4993 (N_4993,N_2495,N_295);
xnor U4994 (N_4994,N_1309,N_355);
or U4995 (N_4995,N_1770,N_1911);
nor U4996 (N_4996,N_2103,N_2749);
or U4997 (N_4997,N_24,N_2881);
and U4998 (N_4998,N_614,N_2975);
nor U4999 (N_4999,N_2402,N_2885);
xnor U5000 (N_5000,N_686,N_1541);
or U5001 (N_5001,N_2918,N_2834);
and U5002 (N_5002,N_2905,N_1025);
or U5003 (N_5003,N_2432,N_780);
or U5004 (N_5004,N_2126,N_548);
and U5005 (N_5005,N_2341,N_532);
and U5006 (N_5006,N_2995,N_2554);
and U5007 (N_5007,N_2823,N_376);
nor U5008 (N_5008,N_1112,N_2114);
nand U5009 (N_5009,N_1840,N_1497);
and U5010 (N_5010,N_1480,N_714);
and U5011 (N_5011,N_2059,N_2801);
and U5012 (N_5012,N_2343,N_1321);
nor U5013 (N_5013,N_2192,N_2535);
nor U5014 (N_5014,N_498,N_1128);
nand U5015 (N_5015,N_2834,N_2596);
nor U5016 (N_5016,N_2264,N_223);
nand U5017 (N_5017,N_2186,N_1181);
xnor U5018 (N_5018,N_2854,N_367);
and U5019 (N_5019,N_1049,N_2161);
nand U5020 (N_5020,N_1671,N_701);
nor U5021 (N_5021,N_2410,N_1538);
or U5022 (N_5022,N_2335,N_1564);
or U5023 (N_5023,N_1069,N_452);
nor U5024 (N_5024,N_1205,N_62);
nand U5025 (N_5025,N_1656,N_1375);
and U5026 (N_5026,N_328,N_2127);
or U5027 (N_5027,N_231,N_2393);
nor U5028 (N_5028,N_2222,N_1946);
or U5029 (N_5029,N_666,N_1283);
nor U5030 (N_5030,N_2954,N_665);
or U5031 (N_5031,N_1881,N_1545);
and U5032 (N_5032,N_109,N_10);
or U5033 (N_5033,N_1052,N_66);
or U5034 (N_5034,N_660,N_2127);
xnor U5035 (N_5035,N_709,N_2550);
and U5036 (N_5036,N_856,N_1724);
nand U5037 (N_5037,N_31,N_820);
and U5038 (N_5038,N_1589,N_398);
nor U5039 (N_5039,N_1322,N_1162);
nor U5040 (N_5040,N_1505,N_2079);
nand U5041 (N_5041,N_141,N_678);
and U5042 (N_5042,N_1825,N_2071);
or U5043 (N_5043,N_2094,N_2675);
and U5044 (N_5044,N_2387,N_2059);
nand U5045 (N_5045,N_1530,N_2677);
nor U5046 (N_5046,N_2866,N_1333);
nor U5047 (N_5047,N_2660,N_346);
and U5048 (N_5048,N_811,N_1065);
nor U5049 (N_5049,N_2638,N_325);
and U5050 (N_5050,N_467,N_1483);
or U5051 (N_5051,N_1420,N_1466);
and U5052 (N_5052,N_722,N_2327);
nand U5053 (N_5053,N_187,N_2170);
and U5054 (N_5054,N_1548,N_847);
nor U5055 (N_5055,N_1897,N_2127);
nor U5056 (N_5056,N_2621,N_1178);
and U5057 (N_5057,N_2273,N_914);
nor U5058 (N_5058,N_1410,N_61);
nor U5059 (N_5059,N_1713,N_1779);
nor U5060 (N_5060,N_2159,N_1169);
nand U5061 (N_5061,N_1197,N_532);
nand U5062 (N_5062,N_2865,N_651);
and U5063 (N_5063,N_1948,N_450);
and U5064 (N_5064,N_1742,N_750);
or U5065 (N_5065,N_151,N_284);
nand U5066 (N_5066,N_1591,N_2491);
or U5067 (N_5067,N_21,N_615);
or U5068 (N_5068,N_1066,N_68);
or U5069 (N_5069,N_2045,N_2358);
nand U5070 (N_5070,N_2998,N_786);
and U5071 (N_5071,N_1429,N_1338);
or U5072 (N_5072,N_2214,N_864);
nor U5073 (N_5073,N_703,N_1548);
and U5074 (N_5074,N_596,N_1567);
and U5075 (N_5075,N_981,N_2800);
nand U5076 (N_5076,N_2714,N_1652);
nand U5077 (N_5077,N_1017,N_1683);
or U5078 (N_5078,N_2660,N_224);
nand U5079 (N_5079,N_1474,N_2151);
and U5080 (N_5080,N_1065,N_666);
nand U5081 (N_5081,N_2093,N_972);
nor U5082 (N_5082,N_4,N_1150);
or U5083 (N_5083,N_1112,N_491);
nor U5084 (N_5084,N_1305,N_1129);
or U5085 (N_5085,N_797,N_200);
nand U5086 (N_5086,N_898,N_661);
nand U5087 (N_5087,N_886,N_125);
or U5088 (N_5088,N_2812,N_2259);
or U5089 (N_5089,N_2010,N_787);
nor U5090 (N_5090,N_2498,N_884);
nor U5091 (N_5091,N_2156,N_202);
nor U5092 (N_5092,N_1073,N_168);
nand U5093 (N_5093,N_937,N_2341);
nor U5094 (N_5094,N_1307,N_890);
nor U5095 (N_5095,N_10,N_1713);
nor U5096 (N_5096,N_2261,N_1406);
nand U5097 (N_5097,N_138,N_2462);
nor U5098 (N_5098,N_2594,N_2788);
and U5099 (N_5099,N_2852,N_112);
and U5100 (N_5100,N_1396,N_2508);
nand U5101 (N_5101,N_1249,N_519);
and U5102 (N_5102,N_191,N_1138);
nor U5103 (N_5103,N_1916,N_2989);
nand U5104 (N_5104,N_808,N_234);
nand U5105 (N_5105,N_2902,N_1070);
or U5106 (N_5106,N_2299,N_2910);
and U5107 (N_5107,N_915,N_2941);
and U5108 (N_5108,N_555,N_1435);
nand U5109 (N_5109,N_784,N_1633);
and U5110 (N_5110,N_90,N_460);
or U5111 (N_5111,N_1328,N_712);
nor U5112 (N_5112,N_1723,N_581);
nand U5113 (N_5113,N_2270,N_1911);
nor U5114 (N_5114,N_2119,N_1405);
or U5115 (N_5115,N_2002,N_648);
and U5116 (N_5116,N_2178,N_2120);
nand U5117 (N_5117,N_2739,N_1699);
and U5118 (N_5118,N_2650,N_131);
nor U5119 (N_5119,N_1910,N_2583);
nor U5120 (N_5120,N_1484,N_1998);
nor U5121 (N_5121,N_750,N_2887);
nand U5122 (N_5122,N_2389,N_1164);
nor U5123 (N_5123,N_1018,N_118);
nand U5124 (N_5124,N_2181,N_923);
or U5125 (N_5125,N_1097,N_2228);
nor U5126 (N_5126,N_270,N_251);
or U5127 (N_5127,N_1278,N_569);
and U5128 (N_5128,N_2746,N_2010);
nor U5129 (N_5129,N_168,N_862);
nand U5130 (N_5130,N_612,N_1069);
or U5131 (N_5131,N_1110,N_2824);
nand U5132 (N_5132,N_619,N_1532);
or U5133 (N_5133,N_73,N_2033);
nand U5134 (N_5134,N_2165,N_2589);
and U5135 (N_5135,N_299,N_1286);
nor U5136 (N_5136,N_1048,N_1761);
or U5137 (N_5137,N_189,N_1692);
or U5138 (N_5138,N_93,N_657);
nor U5139 (N_5139,N_1438,N_2566);
nand U5140 (N_5140,N_2068,N_776);
or U5141 (N_5141,N_749,N_1955);
and U5142 (N_5142,N_75,N_141);
nor U5143 (N_5143,N_2490,N_1003);
or U5144 (N_5144,N_2467,N_1826);
and U5145 (N_5145,N_2599,N_2998);
nor U5146 (N_5146,N_313,N_1655);
nor U5147 (N_5147,N_2996,N_1466);
nor U5148 (N_5148,N_330,N_291);
or U5149 (N_5149,N_1708,N_2991);
nor U5150 (N_5150,N_452,N_430);
and U5151 (N_5151,N_1118,N_2008);
and U5152 (N_5152,N_2881,N_1006);
and U5153 (N_5153,N_1223,N_1581);
nand U5154 (N_5154,N_2235,N_2719);
or U5155 (N_5155,N_493,N_1452);
nor U5156 (N_5156,N_2368,N_373);
nor U5157 (N_5157,N_1207,N_1985);
nand U5158 (N_5158,N_1056,N_1389);
and U5159 (N_5159,N_2519,N_1703);
or U5160 (N_5160,N_2506,N_327);
nor U5161 (N_5161,N_2555,N_59);
nor U5162 (N_5162,N_752,N_179);
nor U5163 (N_5163,N_2382,N_1091);
or U5164 (N_5164,N_1184,N_148);
or U5165 (N_5165,N_746,N_2021);
or U5166 (N_5166,N_2952,N_686);
nand U5167 (N_5167,N_426,N_1859);
nor U5168 (N_5168,N_2345,N_1520);
or U5169 (N_5169,N_1358,N_1444);
nand U5170 (N_5170,N_849,N_2686);
and U5171 (N_5171,N_1415,N_76);
or U5172 (N_5172,N_2664,N_1943);
or U5173 (N_5173,N_342,N_1469);
and U5174 (N_5174,N_1882,N_2911);
and U5175 (N_5175,N_911,N_166);
nor U5176 (N_5176,N_2987,N_2259);
or U5177 (N_5177,N_206,N_365);
or U5178 (N_5178,N_1755,N_2892);
nand U5179 (N_5179,N_411,N_859);
nand U5180 (N_5180,N_103,N_212);
nand U5181 (N_5181,N_1756,N_432);
or U5182 (N_5182,N_619,N_2594);
or U5183 (N_5183,N_989,N_365);
nand U5184 (N_5184,N_1764,N_1140);
or U5185 (N_5185,N_1307,N_1346);
nand U5186 (N_5186,N_2958,N_2722);
or U5187 (N_5187,N_2614,N_2091);
or U5188 (N_5188,N_2561,N_2383);
and U5189 (N_5189,N_1150,N_1204);
nor U5190 (N_5190,N_2158,N_2620);
xor U5191 (N_5191,N_227,N_2843);
or U5192 (N_5192,N_189,N_1511);
nor U5193 (N_5193,N_1724,N_1614);
nor U5194 (N_5194,N_1750,N_697);
or U5195 (N_5195,N_1118,N_1220);
nand U5196 (N_5196,N_2399,N_1076);
and U5197 (N_5197,N_2843,N_655);
or U5198 (N_5198,N_2236,N_1088);
nor U5199 (N_5199,N_2566,N_1855);
nor U5200 (N_5200,N_2743,N_2181);
nand U5201 (N_5201,N_1106,N_819);
nand U5202 (N_5202,N_2966,N_868);
and U5203 (N_5203,N_919,N_1579);
and U5204 (N_5204,N_1492,N_1673);
nand U5205 (N_5205,N_893,N_1119);
or U5206 (N_5206,N_2374,N_661);
and U5207 (N_5207,N_2260,N_62);
and U5208 (N_5208,N_8,N_2388);
nand U5209 (N_5209,N_866,N_2092);
or U5210 (N_5210,N_2604,N_699);
nand U5211 (N_5211,N_2126,N_2989);
nor U5212 (N_5212,N_451,N_1845);
or U5213 (N_5213,N_1975,N_2203);
or U5214 (N_5214,N_2896,N_447);
nor U5215 (N_5215,N_2398,N_2695);
or U5216 (N_5216,N_2342,N_2525);
or U5217 (N_5217,N_900,N_244);
nor U5218 (N_5218,N_2932,N_190);
and U5219 (N_5219,N_2470,N_2010);
nor U5220 (N_5220,N_2983,N_2231);
and U5221 (N_5221,N_1049,N_1212);
nor U5222 (N_5222,N_1156,N_677);
nand U5223 (N_5223,N_93,N_144);
nand U5224 (N_5224,N_2039,N_1211);
and U5225 (N_5225,N_1420,N_2360);
nand U5226 (N_5226,N_484,N_65);
nand U5227 (N_5227,N_968,N_1625);
nor U5228 (N_5228,N_61,N_2237);
and U5229 (N_5229,N_432,N_832);
nand U5230 (N_5230,N_2564,N_2212);
nor U5231 (N_5231,N_632,N_1848);
nor U5232 (N_5232,N_1241,N_1809);
nor U5233 (N_5233,N_2883,N_2780);
or U5234 (N_5234,N_1402,N_693);
nand U5235 (N_5235,N_2323,N_1700);
and U5236 (N_5236,N_2924,N_1522);
nand U5237 (N_5237,N_1221,N_1672);
or U5238 (N_5238,N_2572,N_1354);
nand U5239 (N_5239,N_2900,N_2288);
or U5240 (N_5240,N_2909,N_2221);
or U5241 (N_5241,N_2555,N_286);
and U5242 (N_5242,N_2690,N_1009);
nor U5243 (N_5243,N_1018,N_866);
nand U5244 (N_5244,N_787,N_2812);
nor U5245 (N_5245,N_2728,N_942);
or U5246 (N_5246,N_2651,N_647);
nor U5247 (N_5247,N_2160,N_2380);
and U5248 (N_5248,N_2336,N_2418);
or U5249 (N_5249,N_1173,N_714);
or U5250 (N_5250,N_2792,N_2105);
or U5251 (N_5251,N_1648,N_519);
nor U5252 (N_5252,N_162,N_947);
or U5253 (N_5253,N_1215,N_2148);
or U5254 (N_5254,N_212,N_888);
xnor U5255 (N_5255,N_1349,N_1235);
nand U5256 (N_5256,N_1882,N_858);
or U5257 (N_5257,N_2001,N_1369);
nor U5258 (N_5258,N_820,N_300);
nor U5259 (N_5259,N_715,N_353);
nand U5260 (N_5260,N_2531,N_1150);
or U5261 (N_5261,N_2499,N_1385);
nor U5262 (N_5262,N_818,N_1371);
nand U5263 (N_5263,N_595,N_2242);
nand U5264 (N_5264,N_1229,N_459);
or U5265 (N_5265,N_29,N_1547);
or U5266 (N_5266,N_18,N_2791);
nor U5267 (N_5267,N_1446,N_2511);
and U5268 (N_5268,N_1246,N_484);
nor U5269 (N_5269,N_2257,N_1919);
or U5270 (N_5270,N_1265,N_1569);
or U5271 (N_5271,N_2473,N_2149);
nor U5272 (N_5272,N_1199,N_1099);
or U5273 (N_5273,N_1742,N_2852);
and U5274 (N_5274,N_1665,N_1578);
nand U5275 (N_5275,N_2008,N_1080);
nor U5276 (N_5276,N_1869,N_1521);
nand U5277 (N_5277,N_1660,N_1602);
nor U5278 (N_5278,N_606,N_2447);
and U5279 (N_5279,N_131,N_911);
nor U5280 (N_5280,N_2818,N_1835);
nor U5281 (N_5281,N_1305,N_336);
nor U5282 (N_5282,N_498,N_755);
nand U5283 (N_5283,N_1926,N_163);
or U5284 (N_5284,N_215,N_411);
and U5285 (N_5285,N_525,N_1125);
or U5286 (N_5286,N_2590,N_1798);
or U5287 (N_5287,N_1998,N_2862);
and U5288 (N_5288,N_533,N_2150);
nand U5289 (N_5289,N_68,N_1984);
nor U5290 (N_5290,N_2514,N_1028);
nor U5291 (N_5291,N_2512,N_2622);
nor U5292 (N_5292,N_2239,N_803);
and U5293 (N_5293,N_951,N_2407);
nand U5294 (N_5294,N_1052,N_2904);
or U5295 (N_5295,N_1184,N_930);
nor U5296 (N_5296,N_2981,N_328);
nor U5297 (N_5297,N_1584,N_1854);
nand U5298 (N_5298,N_1365,N_196);
nand U5299 (N_5299,N_130,N_2348);
nand U5300 (N_5300,N_571,N_2207);
or U5301 (N_5301,N_110,N_2655);
or U5302 (N_5302,N_1378,N_778);
nand U5303 (N_5303,N_730,N_2705);
or U5304 (N_5304,N_1085,N_963);
and U5305 (N_5305,N_41,N_2717);
or U5306 (N_5306,N_2805,N_716);
nand U5307 (N_5307,N_1816,N_1327);
nor U5308 (N_5308,N_2384,N_785);
and U5309 (N_5309,N_1489,N_1011);
and U5310 (N_5310,N_83,N_2092);
nand U5311 (N_5311,N_670,N_2153);
nor U5312 (N_5312,N_1113,N_1125);
nor U5313 (N_5313,N_656,N_1106);
nand U5314 (N_5314,N_222,N_2851);
or U5315 (N_5315,N_184,N_1688);
and U5316 (N_5316,N_2173,N_434);
or U5317 (N_5317,N_1661,N_2262);
nand U5318 (N_5318,N_1867,N_553);
and U5319 (N_5319,N_1841,N_2005);
and U5320 (N_5320,N_447,N_1611);
nand U5321 (N_5321,N_2463,N_2223);
and U5322 (N_5322,N_1283,N_2906);
nand U5323 (N_5323,N_917,N_660);
xnor U5324 (N_5324,N_591,N_2176);
nor U5325 (N_5325,N_2299,N_2218);
nand U5326 (N_5326,N_2404,N_1246);
and U5327 (N_5327,N_2876,N_2368);
or U5328 (N_5328,N_350,N_988);
and U5329 (N_5329,N_2612,N_2504);
nand U5330 (N_5330,N_2883,N_1401);
and U5331 (N_5331,N_970,N_2031);
or U5332 (N_5332,N_2959,N_1423);
nand U5333 (N_5333,N_1575,N_2044);
nor U5334 (N_5334,N_2787,N_1676);
xor U5335 (N_5335,N_2961,N_1270);
or U5336 (N_5336,N_2354,N_2048);
or U5337 (N_5337,N_2595,N_126);
and U5338 (N_5338,N_1755,N_493);
nand U5339 (N_5339,N_1804,N_1471);
xor U5340 (N_5340,N_2527,N_2849);
nand U5341 (N_5341,N_1891,N_2378);
and U5342 (N_5342,N_1338,N_1033);
nor U5343 (N_5343,N_100,N_2788);
nand U5344 (N_5344,N_1766,N_860);
nor U5345 (N_5345,N_2111,N_1317);
and U5346 (N_5346,N_2446,N_2905);
nor U5347 (N_5347,N_1652,N_1862);
nor U5348 (N_5348,N_2495,N_1861);
and U5349 (N_5349,N_0,N_2962);
nand U5350 (N_5350,N_629,N_2393);
nand U5351 (N_5351,N_1161,N_1939);
nor U5352 (N_5352,N_597,N_1353);
nor U5353 (N_5353,N_2068,N_114);
nand U5354 (N_5354,N_1187,N_917);
or U5355 (N_5355,N_1492,N_2809);
nor U5356 (N_5356,N_564,N_90);
nand U5357 (N_5357,N_2272,N_1525);
or U5358 (N_5358,N_24,N_738);
and U5359 (N_5359,N_451,N_129);
nand U5360 (N_5360,N_1753,N_1632);
and U5361 (N_5361,N_2220,N_533);
nor U5362 (N_5362,N_2477,N_540);
and U5363 (N_5363,N_1171,N_99);
and U5364 (N_5364,N_349,N_2695);
and U5365 (N_5365,N_1700,N_1160);
or U5366 (N_5366,N_2781,N_1764);
or U5367 (N_5367,N_121,N_474);
and U5368 (N_5368,N_1182,N_1815);
xor U5369 (N_5369,N_1778,N_2056);
and U5370 (N_5370,N_2151,N_2737);
or U5371 (N_5371,N_928,N_2550);
and U5372 (N_5372,N_682,N_2189);
nand U5373 (N_5373,N_2876,N_813);
or U5374 (N_5374,N_1697,N_1963);
or U5375 (N_5375,N_316,N_815);
nor U5376 (N_5376,N_679,N_880);
xnor U5377 (N_5377,N_2175,N_374);
and U5378 (N_5378,N_385,N_2994);
or U5379 (N_5379,N_1627,N_891);
nand U5380 (N_5380,N_579,N_2498);
or U5381 (N_5381,N_572,N_2930);
or U5382 (N_5382,N_1848,N_1351);
nand U5383 (N_5383,N_901,N_161);
or U5384 (N_5384,N_2111,N_430);
nand U5385 (N_5385,N_1445,N_1355);
nor U5386 (N_5386,N_82,N_2668);
nor U5387 (N_5387,N_0,N_2302);
or U5388 (N_5388,N_1898,N_1761);
and U5389 (N_5389,N_445,N_1454);
nand U5390 (N_5390,N_1635,N_2132);
and U5391 (N_5391,N_1695,N_1268);
nor U5392 (N_5392,N_307,N_287);
nand U5393 (N_5393,N_2875,N_2119);
and U5394 (N_5394,N_1199,N_825);
and U5395 (N_5395,N_4,N_634);
or U5396 (N_5396,N_562,N_1752);
and U5397 (N_5397,N_2342,N_284);
or U5398 (N_5398,N_1746,N_1968);
and U5399 (N_5399,N_2198,N_2688);
and U5400 (N_5400,N_1295,N_1383);
nor U5401 (N_5401,N_2841,N_377);
or U5402 (N_5402,N_2425,N_2140);
nand U5403 (N_5403,N_1688,N_365);
or U5404 (N_5404,N_1378,N_178);
nand U5405 (N_5405,N_539,N_643);
nand U5406 (N_5406,N_1870,N_1991);
or U5407 (N_5407,N_2757,N_2434);
or U5408 (N_5408,N_309,N_1260);
or U5409 (N_5409,N_2766,N_382);
nor U5410 (N_5410,N_1456,N_705);
nand U5411 (N_5411,N_9,N_2180);
and U5412 (N_5412,N_2790,N_939);
nor U5413 (N_5413,N_1675,N_1446);
nand U5414 (N_5414,N_1747,N_108);
nor U5415 (N_5415,N_451,N_1569);
or U5416 (N_5416,N_2363,N_1473);
nor U5417 (N_5417,N_1360,N_2835);
nor U5418 (N_5418,N_879,N_2264);
and U5419 (N_5419,N_2951,N_1747);
nand U5420 (N_5420,N_1976,N_558);
or U5421 (N_5421,N_461,N_546);
or U5422 (N_5422,N_92,N_140);
nor U5423 (N_5423,N_12,N_1998);
or U5424 (N_5424,N_2727,N_1155);
or U5425 (N_5425,N_2285,N_952);
or U5426 (N_5426,N_938,N_1468);
nor U5427 (N_5427,N_2404,N_2607);
and U5428 (N_5428,N_2727,N_1891);
and U5429 (N_5429,N_1456,N_22);
nand U5430 (N_5430,N_807,N_1558);
or U5431 (N_5431,N_865,N_2361);
nand U5432 (N_5432,N_2760,N_2456);
nand U5433 (N_5433,N_964,N_112);
or U5434 (N_5434,N_111,N_1779);
nand U5435 (N_5435,N_660,N_820);
xor U5436 (N_5436,N_1510,N_2033);
and U5437 (N_5437,N_1361,N_1990);
and U5438 (N_5438,N_337,N_684);
and U5439 (N_5439,N_240,N_821);
or U5440 (N_5440,N_80,N_331);
or U5441 (N_5441,N_670,N_818);
and U5442 (N_5442,N_929,N_2851);
nor U5443 (N_5443,N_464,N_37);
nor U5444 (N_5444,N_2688,N_876);
and U5445 (N_5445,N_1413,N_774);
and U5446 (N_5446,N_161,N_707);
nand U5447 (N_5447,N_193,N_1861);
nor U5448 (N_5448,N_2679,N_1505);
or U5449 (N_5449,N_1166,N_2496);
nand U5450 (N_5450,N_845,N_2731);
nor U5451 (N_5451,N_2912,N_1732);
nand U5452 (N_5452,N_956,N_2709);
or U5453 (N_5453,N_2082,N_475);
nor U5454 (N_5454,N_2644,N_559);
nand U5455 (N_5455,N_551,N_1774);
nor U5456 (N_5456,N_2632,N_2394);
and U5457 (N_5457,N_1034,N_387);
nand U5458 (N_5458,N_586,N_1208);
nand U5459 (N_5459,N_2550,N_1774);
and U5460 (N_5460,N_2001,N_664);
or U5461 (N_5461,N_1298,N_1103);
nand U5462 (N_5462,N_850,N_1259);
and U5463 (N_5463,N_2387,N_2348);
nor U5464 (N_5464,N_951,N_2464);
nand U5465 (N_5465,N_205,N_2283);
and U5466 (N_5466,N_2335,N_1036);
and U5467 (N_5467,N_1456,N_514);
nor U5468 (N_5468,N_2809,N_1953);
and U5469 (N_5469,N_1157,N_2714);
and U5470 (N_5470,N_1590,N_2274);
and U5471 (N_5471,N_1433,N_2247);
nand U5472 (N_5472,N_2238,N_1225);
nor U5473 (N_5473,N_1905,N_1820);
nor U5474 (N_5474,N_1165,N_30);
nor U5475 (N_5475,N_2755,N_803);
nand U5476 (N_5476,N_1472,N_2808);
nand U5477 (N_5477,N_2933,N_1530);
nor U5478 (N_5478,N_2693,N_970);
nor U5479 (N_5479,N_1505,N_1966);
xor U5480 (N_5480,N_331,N_679);
or U5481 (N_5481,N_2460,N_2127);
and U5482 (N_5482,N_2977,N_1845);
nor U5483 (N_5483,N_1444,N_1156);
or U5484 (N_5484,N_2986,N_2375);
nor U5485 (N_5485,N_1389,N_2880);
nor U5486 (N_5486,N_1851,N_1705);
and U5487 (N_5487,N_2742,N_569);
nand U5488 (N_5488,N_54,N_834);
nand U5489 (N_5489,N_920,N_2455);
nand U5490 (N_5490,N_2964,N_355);
nor U5491 (N_5491,N_821,N_977);
and U5492 (N_5492,N_2671,N_603);
and U5493 (N_5493,N_2132,N_2426);
nand U5494 (N_5494,N_359,N_2791);
nor U5495 (N_5495,N_2009,N_567);
and U5496 (N_5496,N_1185,N_1575);
nor U5497 (N_5497,N_1981,N_2395);
or U5498 (N_5498,N_1834,N_1037);
and U5499 (N_5499,N_274,N_794);
and U5500 (N_5500,N_1270,N_1195);
nand U5501 (N_5501,N_114,N_539);
nand U5502 (N_5502,N_1895,N_1681);
nand U5503 (N_5503,N_1501,N_731);
nor U5504 (N_5504,N_261,N_526);
and U5505 (N_5505,N_2973,N_1555);
nand U5506 (N_5506,N_2603,N_1765);
nor U5507 (N_5507,N_914,N_1093);
nor U5508 (N_5508,N_2616,N_1910);
nand U5509 (N_5509,N_2363,N_2696);
nor U5510 (N_5510,N_884,N_596);
or U5511 (N_5511,N_1204,N_95);
nand U5512 (N_5512,N_1940,N_1194);
and U5513 (N_5513,N_909,N_2918);
and U5514 (N_5514,N_1685,N_953);
nor U5515 (N_5515,N_2974,N_2090);
nor U5516 (N_5516,N_1738,N_1461);
and U5517 (N_5517,N_1479,N_1202);
nor U5518 (N_5518,N_2170,N_2595);
nor U5519 (N_5519,N_587,N_2007);
nor U5520 (N_5520,N_273,N_724);
and U5521 (N_5521,N_1159,N_2572);
and U5522 (N_5522,N_2887,N_1543);
nand U5523 (N_5523,N_1369,N_473);
or U5524 (N_5524,N_1507,N_2196);
and U5525 (N_5525,N_36,N_1156);
and U5526 (N_5526,N_1683,N_1894);
and U5527 (N_5527,N_1342,N_1900);
nor U5528 (N_5528,N_2666,N_158);
nand U5529 (N_5529,N_1547,N_2049);
and U5530 (N_5530,N_1489,N_2052);
nand U5531 (N_5531,N_1461,N_1834);
nor U5532 (N_5532,N_2753,N_2145);
nor U5533 (N_5533,N_906,N_836);
nor U5534 (N_5534,N_1531,N_1247);
nand U5535 (N_5535,N_2123,N_1853);
nor U5536 (N_5536,N_2719,N_897);
and U5537 (N_5537,N_75,N_2673);
nor U5538 (N_5538,N_22,N_90);
nand U5539 (N_5539,N_476,N_1802);
nand U5540 (N_5540,N_1130,N_183);
nor U5541 (N_5541,N_1267,N_1949);
and U5542 (N_5542,N_1748,N_2429);
nor U5543 (N_5543,N_283,N_705);
nor U5544 (N_5544,N_334,N_1266);
and U5545 (N_5545,N_1725,N_2535);
nand U5546 (N_5546,N_2528,N_2406);
nor U5547 (N_5547,N_2204,N_419);
nor U5548 (N_5548,N_1662,N_40);
nand U5549 (N_5549,N_242,N_1817);
nor U5550 (N_5550,N_2066,N_2675);
and U5551 (N_5551,N_813,N_2607);
nor U5552 (N_5552,N_1128,N_1045);
or U5553 (N_5553,N_2531,N_752);
nand U5554 (N_5554,N_157,N_1436);
or U5555 (N_5555,N_262,N_2823);
and U5556 (N_5556,N_2243,N_1426);
or U5557 (N_5557,N_459,N_1896);
or U5558 (N_5558,N_2415,N_753);
nand U5559 (N_5559,N_2665,N_928);
nand U5560 (N_5560,N_384,N_681);
nor U5561 (N_5561,N_270,N_1017);
nand U5562 (N_5562,N_610,N_2870);
and U5563 (N_5563,N_1848,N_224);
nor U5564 (N_5564,N_2834,N_2736);
or U5565 (N_5565,N_559,N_794);
or U5566 (N_5566,N_2367,N_1536);
and U5567 (N_5567,N_968,N_142);
and U5568 (N_5568,N_2604,N_2338);
or U5569 (N_5569,N_2967,N_1522);
nor U5570 (N_5570,N_472,N_1843);
nor U5571 (N_5571,N_960,N_1480);
or U5572 (N_5572,N_1137,N_2925);
or U5573 (N_5573,N_2096,N_804);
nand U5574 (N_5574,N_1618,N_147);
and U5575 (N_5575,N_2464,N_1513);
nand U5576 (N_5576,N_2636,N_1505);
nor U5577 (N_5577,N_1546,N_1312);
nor U5578 (N_5578,N_635,N_445);
and U5579 (N_5579,N_1030,N_263);
nand U5580 (N_5580,N_2383,N_2135);
and U5581 (N_5581,N_1278,N_2681);
nor U5582 (N_5582,N_674,N_1999);
nor U5583 (N_5583,N_614,N_1395);
and U5584 (N_5584,N_2346,N_1981);
or U5585 (N_5585,N_1812,N_370);
or U5586 (N_5586,N_1717,N_1210);
nand U5587 (N_5587,N_1819,N_1415);
nand U5588 (N_5588,N_505,N_1329);
nor U5589 (N_5589,N_2615,N_1433);
nor U5590 (N_5590,N_85,N_1349);
nor U5591 (N_5591,N_2674,N_2952);
nor U5592 (N_5592,N_1572,N_1570);
nand U5593 (N_5593,N_1663,N_2028);
nand U5594 (N_5594,N_1637,N_2681);
and U5595 (N_5595,N_544,N_1858);
and U5596 (N_5596,N_1363,N_1288);
or U5597 (N_5597,N_245,N_324);
or U5598 (N_5598,N_1763,N_2870);
nor U5599 (N_5599,N_442,N_79);
nor U5600 (N_5600,N_998,N_1810);
nand U5601 (N_5601,N_339,N_799);
or U5602 (N_5602,N_260,N_2938);
and U5603 (N_5603,N_2230,N_991);
nor U5604 (N_5604,N_1728,N_597);
nor U5605 (N_5605,N_1191,N_455);
nand U5606 (N_5606,N_2410,N_729);
or U5607 (N_5607,N_259,N_1519);
and U5608 (N_5608,N_2517,N_2271);
and U5609 (N_5609,N_2738,N_346);
nand U5610 (N_5610,N_2932,N_1762);
nor U5611 (N_5611,N_2229,N_1396);
nand U5612 (N_5612,N_1334,N_2312);
nor U5613 (N_5613,N_2983,N_2801);
nor U5614 (N_5614,N_1492,N_2617);
or U5615 (N_5615,N_57,N_1358);
nand U5616 (N_5616,N_2968,N_718);
and U5617 (N_5617,N_1008,N_2936);
or U5618 (N_5618,N_772,N_163);
or U5619 (N_5619,N_371,N_2684);
or U5620 (N_5620,N_102,N_2098);
nand U5621 (N_5621,N_906,N_340);
nand U5622 (N_5622,N_859,N_330);
nor U5623 (N_5623,N_497,N_2794);
nor U5624 (N_5624,N_598,N_2630);
nor U5625 (N_5625,N_905,N_1643);
and U5626 (N_5626,N_1347,N_2858);
and U5627 (N_5627,N_2733,N_1662);
nor U5628 (N_5628,N_2892,N_675);
nor U5629 (N_5629,N_2271,N_2326);
and U5630 (N_5630,N_2815,N_690);
nor U5631 (N_5631,N_2329,N_2345);
nor U5632 (N_5632,N_20,N_406);
nand U5633 (N_5633,N_2749,N_1997);
nor U5634 (N_5634,N_280,N_2379);
nand U5635 (N_5635,N_401,N_1725);
nand U5636 (N_5636,N_1507,N_2966);
and U5637 (N_5637,N_2736,N_525);
or U5638 (N_5638,N_2350,N_2025);
nand U5639 (N_5639,N_2825,N_1199);
or U5640 (N_5640,N_126,N_2709);
or U5641 (N_5641,N_1675,N_1089);
or U5642 (N_5642,N_1262,N_2064);
nor U5643 (N_5643,N_392,N_38);
and U5644 (N_5644,N_2454,N_2350);
nand U5645 (N_5645,N_705,N_2160);
nand U5646 (N_5646,N_357,N_1002);
or U5647 (N_5647,N_283,N_2260);
nand U5648 (N_5648,N_355,N_1863);
and U5649 (N_5649,N_439,N_1287);
or U5650 (N_5650,N_999,N_2928);
or U5651 (N_5651,N_1692,N_762);
and U5652 (N_5652,N_2856,N_1573);
nand U5653 (N_5653,N_663,N_2676);
nor U5654 (N_5654,N_771,N_1940);
nand U5655 (N_5655,N_1407,N_680);
nand U5656 (N_5656,N_407,N_2693);
nand U5657 (N_5657,N_1230,N_1625);
nor U5658 (N_5658,N_38,N_1567);
and U5659 (N_5659,N_805,N_2473);
and U5660 (N_5660,N_1760,N_2874);
nand U5661 (N_5661,N_417,N_2426);
and U5662 (N_5662,N_2538,N_1800);
nand U5663 (N_5663,N_694,N_2954);
or U5664 (N_5664,N_2734,N_887);
nand U5665 (N_5665,N_249,N_1374);
nor U5666 (N_5666,N_1800,N_73);
and U5667 (N_5667,N_1228,N_2160);
nand U5668 (N_5668,N_1903,N_232);
nand U5669 (N_5669,N_1313,N_2364);
or U5670 (N_5670,N_2332,N_2824);
and U5671 (N_5671,N_604,N_2785);
nor U5672 (N_5672,N_1062,N_2897);
or U5673 (N_5673,N_1464,N_1767);
and U5674 (N_5674,N_572,N_2330);
nor U5675 (N_5675,N_1478,N_2330);
nand U5676 (N_5676,N_2472,N_564);
and U5677 (N_5677,N_2041,N_2303);
and U5678 (N_5678,N_382,N_1299);
nand U5679 (N_5679,N_992,N_718);
nand U5680 (N_5680,N_1363,N_1094);
nand U5681 (N_5681,N_2479,N_2329);
nor U5682 (N_5682,N_222,N_767);
nand U5683 (N_5683,N_962,N_1182);
nor U5684 (N_5684,N_2906,N_1195);
and U5685 (N_5685,N_743,N_366);
nand U5686 (N_5686,N_2631,N_2744);
nand U5687 (N_5687,N_2028,N_1524);
nor U5688 (N_5688,N_351,N_788);
or U5689 (N_5689,N_987,N_308);
and U5690 (N_5690,N_1238,N_231);
nor U5691 (N_5691,N_1707,N_2657);
nor U5692 (N_5692,N_1406,N_669);
or U5693 (N_5693,N_1694,N_2661);
or U5694 (N_5694,N_567,N_444);
nor U5695 (N_5695,N_2169,N_943);
nand U5696 (N_5696,N_1264,N_553);
or U5697 (N_5697,N_525,N_749);
nand U5698 (N_5698,N_1519,N_2014);
nor U5699 (N_5699,N_1609,N_1467);
nand U5700 (N_5700,N_1811,N_2738);
or U5701 (N_5701,N_1230,N_2445);
nor U5702 (N_5702,N_211,N_1960);
or U5703 (N_5703,N_1135,N_1711);
and U5704 (N_5704,N_1802,N_2170);
or U5705 (N_5705,N_2366,N_295);
or U5706 (N_5706,N_1432,N_196);
or U5707 (N_5707,N_1546,N_1652);
nor U5708 (N_5708,N_1546,N_2699);
and U5709 (N_5709,N_1823,N_2604);
and U5710 (N_5710,N_1399,N_1369);
and U5711 (N_5711,N_1458,N_2991);
and U5712 (N_5712,N_700,N_2298);
nor U5713 (N_5713,N_850,N_1478);
or U5714 (N_5714,N_100,N_1102);
nor U5715 (N_5715,N_2019,N_2502);
or U5716 (N_5716,N_436,N_2992);
nor U5717 (N_5717,N_1493,N_2329);
nand U5718 (N_5718,N_1198,N_1096);
nand U5719 (N_5719,N_1482,N_1262);
or U5720 (N_5720,N_500,N_1576);
nor U5721 (N_5721,N_1084,N_1749);
and U5722 (N_5722,N_258,N_1885);
or U5723 (N_5723,N_930,N_2579);
and U5724 (N_5724,N_201,N_2979);
nor U5725 (N_5725,N_1612,N_1653);
and U5726 (N_5726,N_2806,N_1970);
nand U5727 (N_5727,N_230,N_2969);
and U5728 (N_5728,N_2931,N_267);
xor U5729 (N_5729,N_2521,N_151);
nand U5730 (N_5730,N_2957,N_765);
and U5731 (N_5731,N_1740,N_1386);
or U5732 (N_5732,N_2561,N_2517);
nor U5733 (N_5733,N_1606,N_531);
and U5734 (N_5734,N_1537,N_171);
and U5735 (N_5735,N_403,N_572);
and U5736 (N_5736,N_1320,N_1256);
nand U5737 (N_5737,N_1427,N_1984);
or U5738 (N_5738,N_669,N_539);
and U5739 (N_5739,N_1512,N_1186);
nand U5740 (N_5740,N_29,N_1359);
or U5741 (N_5741,N_1023,N_2806);
and U5742 (N_5742,N_2055,N_1565);
or U5743 (N_5743,N_1766,N_2089);
nand U5744 (N_5744,N_515,N_917);
and U5745 (N_5745,N_2941,N_1949);
nor U5746 (N_5746,N_1378,N_2301);
and U5747 (N_5747,N_1891,N_2681);
nand U5748 (N_5748,N_1,N_2817);
and U5749 (N_5749,N_751,N_2712);
nand U5750 (N_5750,N_1379,N_498);
nand U5751 (N_5751,N_1516,N_430);
nor U5752 (N_5752,N_2850,N_1555);
nor U5753 (N_5753,N_2677,N_802);
or U5754 (N_5754,N_1244,N_2589);
xor U5755 (N_5755,N_2203,N_2404);
nor U5756 (N_5756,N_216,N_2974);
or U5757 (N_5757,N_1527,N_772);
or U5758 (N_5758,N_2968,N_2223);
nand U5759 (N_5759,N_738,N_1156);
nand U5760 (N_5760,N_1260,N_396);
nor U5761 (N_5761,N_888,N_2361);
and U5762 (N_5762,N_1308,N_2541);
nand U5763 (N_5763,N_1543,N_595);
and U5764 (N_5764,N_2452,N_351);
nor U5765 (N_5765,N_1583,N_1040);
nand U5766 (N_5766,N_968,N_1516);
and U5767 (N_5767,N_1163,N_1290);
and U5768 (N_5768,N_35,N_234);
nand U5769 (N_5769,N_2601,N_124);
nand U5770 (N_5770,N_2386,N_1279);
and U5771 (N_5771,N_2001,N_1577);
and U5772 (N_5772,N_2181,N_299);
nor U5773 (N_5773,N_1288,N_2157);
and U5774 (N_5774,N_1769,N_315);
nor U5775 (N_5775,N_997,N_2226);
and U5776 (N_5776,N_1886,N_2024);
or U5777 (N_5777,N_976,N_1734);
nand U5778 (N_5778,N_1438,N_2422);
nor U5779 (N_5779,N_63,N_2187);
or U5780 (N_5780,N_1760,N_1060);
or U5781 (N_5781,N_1635,N_2197);
nand U5782 (N_5782,N_2257,N_1569);
nand U5783 (N_5783,N_180,N_1304);
or U5784 (N_5784,N_2098,N_1163);
or U5785 (N_5785,N_2992,N_653);
nand U5786 (N_5786,N_1939,N_322);
and U5787 (N_5787,N_2180,N_2413);
or U5788 (N_5788,N_2460,N_1357);
and U5789 (N_5789,N_1713,N_2945);
or U5790 (N_5790,N_1806,N_1919);
or U5791 (N_5791,N_1305,N_1553);
or U5792 (N_5792,N_718,N_729);
nand U5793 (N_5793,N_1279,N_2269);
and U5794 (N_5794,N_1446,N_1381);
nand U5795 (N_5795,N_2978,N_1162);
and U5796 (N_5796,N_242,N_133);
nand U5797 (N_5797,N_1741,N_641);
nor U5798 (N_5798,N_307,N_2886);
nor U5799 (N_5799,N_2735,N_2298);
nor U5800 (N_5800,N_2972,N_2141);
nand U5801 (N_5801,N_90,N_1122);
and U5802 (N_5802,N_33,N_1899);
and U5803 (N_5803,N_1283,N_2397);
nand U5804 (N_5804,N_1922,N_1285);
or U5805 (N_5805,N_1292,N_2867);
or U5806 (N_5806,N_2873,N_1022);
and U5807 (N_5807,N_1810,N_744);
or U5808 (N_5808,N_2165,N_994);
xnor U5809 (N_5809,N_521,N_1279);
or U5810 (N_5810,N_2876,N_303);
or U5811 (N_5811,N_1502,N_2966);
and U5812 (N_5812,N_962,N_2244);
nand U5813 (N_5813,N_1417,N_808);
and U5814 (N_5814,N_189,N_1724);
and U5815 (N_5815,N_2178,N_1763);
nor U5816 (N_5816,N_1374,N_1237);
nor U5817 (N_5817,N_979,N_1029);
nand U5818 (N_5818,N_2038,N_1819);
or U5819 (N_5819,N_1512,N_1082);
nand U5820 (N_5820,N_1081,N_2880);
or U5821 (N_5821,N_1992,N_1221);
nor U5822 (N_5822,N_1804,N_2865);
nand U5823 (N_5823,N_2846,N_2);
nor U5824 (N_5824,N_155,N_246);
or U5825 (N_5825,N_444,N_1126);
nand U5826 (N_5826,N_1111,N_2314);
or U5827 (N_5827,N_878,N_1809);
and U5828 (N_5828,N_967,N_1162);
or U5829 (N_5829,N_2687,N_34);
or U5830 (N_5830,N_2033,N_1963);
nand U5831 (N_5831,N_2234,N_410);
nand U5832 (N_5832,N_1094,N_1603);
nand U5833 (N_5833,N_794,N_1917);
and U5834 (N_5834,N_2302,N_1981);
nand U5835 (N_5835,N_1748,N_2137);
nor U5836 (N_5836,N_2435,N_1545);
xor U5837 (N_5837,N_2400,N_2552);
and U5838 (N_5838,N_2912,N_980);
and U5839 (N_5839,N_230,N_1771);
and U5840 (N_5840,N_2203,N_2716);
nand U5841 (N_5841,N_1498,N_520);
and U5842 (N_5842,N_691,N_1483);
and U5843 (N_5843,N_1839,N_2250);
nor U5844 (N_5844,N_2557,N_2169);
or U5845 (N_5845,N_2603,N_2574);
and U5846 (N_5846,N_2620,N_954);
nor U5847 (N_5847,N_351,N_712);
nand U5848 (N_5848,N_1288,N_143);
nor U5849 (N_5849,N_2384,N_639);
and U5850 (N_5850,N_279,N_1154);
or U5851 (N_5851,N_2737,N_156);
or U5852 (N_5852,N_1363,N_1938);
nor U5853 (N_5853,N_1878,N_818);
or U5854 (N_5854,N_1246,N_1182);
nor U5855 (N_5855,N_585,N_2921);
nor U5856 (N_5856,N_2767,N_670);
or U5857 (N_5857,N_896,N_290);
nand U5858 (N_5858,N_345,N_172);
and U5859 (N_5859,N_1713,N_2074);
nor U5860 (N_5860,N_2993,N_1325);
or U5861 (N_5861,N_1327,N_445);
nor U5862 (N_5862,N_811,N_2251);
nand U5863 (N_5863,N_1349,N_25);
or U5864 (N_5864,N_184,N_2554);
nor U5865 (N_5865,N_928,N_1166);
and U5866 (N_5866,N_1882,N_2520);
and U5867 (N_5867,N_2057,N_909);
nor U5868 (N_5868,N_1681,N_199);
or U5869 (N_5869,N_435,N_254);
nand U5870 (N_5870,N_974,N_2799);
nor U5871 (N_5871,N_1988,N_1018);
or U5872 (N_5872,N_950,N_290);
or U5873 (N_5873,N_2818,N_1014);
nor U5874 (N_5874,N_2691,N_2612);
nor U5875 (N_5875,N_2887,N_2798);
and U5876 (N_5876,N_1631,N_1544);
nand U5877 (N_5877,N_388,N_664);
nor U5878 (N_5878,N_1004,N_2099);
nor U5879 (N_5879,N_1586,N_160);
or U5880 (N_5880,N_769,N_2339);
nand U5881 (N_5881,N_444,N_2029);
nand U5882 (N_5882,N_463,N_1221);
or U5883 (N_5883,N_1951,N_2334);
and U5884 (N_5884,N_2444,N_701);
or U5885 (N_5885,N_1255,N_2222);
nor U5886 (N_5886,N_1087,N_2392);
and U5887 (N_5887,N_673,N_1166);
nand U5888 (N_5888,N_1201,N_2080);
xnor U5889 (N_5889,N_394,N_1932);
and U5890 (N_5890,N_2443,N_2223);
or U5891 (N_5891,N_1255,N_12);
and U5892 (N_5892,N_721,N_2487);
or U5893 (N_5893,N_1749,N_1070);
or U5894 (N_5894,N_2730,N_1509);
nand U5895 (N_5895,N_1489,N_1776);
and U5896 (N_5896,N_2099,N_1944);
nand U5897 (N_5897,N_143,N_1870);
nand U5898 (N_5898,N_2408,N_2867);
nand U5899 (N_5899,N_997,N_459);
nor U5900 (N_5900,N_374,N_2646);
and U5901 (N_5901,N_2778,N_2790);
or U5902 (N_5902,N_144,N_2065);
or U5903 (N_5903,N_124,N_770);
nand U5904 (N_5904,N_2593,N_906);
nor U5905 (N_5905,N_1039,N_1872);
nand U5906 (N_5906,N_2003,N_645);
and U5907 (N_5907,N_543,N_1457);
nor U5908 (N_5908,N_190,N_663);
or U5909 (N_5909,N_32,N_502);
and U5910 (N_5910,N_682,N_547);
and U5911 (N_5911,N_861,N_1694);
nor U5912 (N_5912,N_757,N_923);
or U5913 (N_5913,N_2245,N_318);
nor U5914 (N_5914,N_1048,N_2670);
or U5915 (N_5915,N_2354,N_1321);
and U5916 (N_5916,N_747,N_1741);
or U5917 (N_5917,N_2934,N_2336);
and U5918 (N_5918,N_1843,N_52);
nand U5919 (N_5919,N_2101,N_1385);
nand U5920 (N_5920,N_980,N_1744);
or U5921 (N_5921,N_1331,N_1800);
or U5922 (N_5922,N_2046,N_1471);
nand U5923 (N_5923,N_401,N_1091);
nor U5924 (N_5924,N_46,N_1883);
nand U5925 (N_5925,N_973,N_433);
nand U5926 (N_5926,N_717,N_460);
and U5927 (N_5927,N_181,N_1832);
and U5928 (N_5928,N_62,N_1682);
nor U5929 (N_5929,N_2640,N_526);
and U5930 (N_5930,N_2989,N_1018);
nand U5931 (N_5931,N_196,N_2276);
or U5932 (N_5932,N_2726,N_1996);
nor U5933 (N_5933,N_2429,N_428);
or U5934 (N_5934,N_2387,N_1944);
or U5935 (N_5935,N_1388,N_760);
and U5936 (N_5936,N_49,N_2590);
or U5937 (N_5937,N_2572,N_2092);
or U5938 (N_5938,N_590,N_188);
and U5939 (N_5939,N_2756,N_1082);
or U5940 (N_5940,N_470,N_2966);
and U5941 (N_5941,N_2157,N_375);
nor U5942 (N_5942,N_820,N_587);
xor U5943 (N_5943,N_962,N_872);
nor U5944 (N_5944,N_1375,N_653);
nand U5945 (N_5945,N_1206,N_1532);
nor U5946 (N_5946,N_2281,N_767);
or U5947 (N_5947,N_298,N_1993);
nor U5948 (N_5948,N_548,N_2626);
nand U5949 (N_5949,N_2497,N_2991);
and U5950 (N_5950,N_2088,N_2352);
nor U5951 (N_5951,N_2628,N_1309);
nor U5952 (N_5952,N_2440,N_1284);
nor U5953 (N_5953,N_745,N_1444);
nor U5954 (N_5954,N_2222,N_191);
nor U5955 (N_5955,N_410,N_195);
and U5956 (N_5956,N_2874,N_304);
nor U5957 (N_5957,N_991,N_2500);
nand U5958 (N_5958,N_1386,N_2969);
nand U5959 (N_5959,N_324,N_1463);
and U5960 (N_5960,N_281,N_2918);
and U5961 (N_5961,N_1585,N_2127);
nor U5962 (N_5962,N_2670,N_1571);
or U5963 (N_5963,N_2828,N_1530);
and U5964 (N_5964,N_2810,N_869);
or U5965 (N_5965,N_2865,N_2023);
nand U5966 (N_5966,N_2873,N_2046);
and U5967 (N_5967,N_720,N_2258);
nor U5968 (N_5968,N_301,N_1973);
or U5969 (N_5969,N_1017,N_352);
nand U5970 (N_5970,N_1635,N_1415);
nor U5971 (N_5971,N_1469,N_2970);
or U5972 (N_5972,N_1779,N_2770);
nand U5973 (N_5973,N_548,N_826);
nand U5974 (N_5974,N_1510,N_154);
or U5975 (N_5975,N_2846,N_2882);
and U5976 (N_5976,N_432,N_1516);
xor U5977 (N_5977,N_1433,N_257);
nand U5978 (N_5978,N_553,N_2010);
nor U5979 (N_5979,N_565,N_2981);
nor U5980 (N_5980,N_251,N_2449);
nor U5981 (N_5981,N_2439,N_2661);
and U5982 (N_5982,N_2218,N_2210);
and U5983 (N_5983,N_1532,N_269);
nor U5984 (N_5984,N_947,N_2406);
and U5985 (N_5985,N_800,N_2946);
nand U5986 (N_5986,N_103,N_1322);
nor U5987 (N_5987,N_1526,N_1843);
or U5988 (N_5988,N_958,N_1261);
nor U5989 (N_5989,N_1582,N_2417);
and U5990 (N_5990,N_2015,N_2462);
and U5991 (N_5991,N_1468,N_2475);
and U5992 (N_5992,N_2180,N_2187);
nand U5993 (N_5993,N_1314,N_2858);
and U5994 (N_5994,N_2702,N_1724);
and U5995 (N_5995,N_2989,N_2478);
and U5996 (N_5996,N_507,N_1487);
and U5997 (N_5997,N_1365,N_512);
or U5998 (N_5998,N_2517,N_19);
nand U5999 (N_5999,N_1620,N_130);
or U6000 (N_6000,N_3956,N_5950);
or U6001 (N_6001,N_5301,N_4079);
nor U6002 (N_6002,N_3149,N_3836);
nor U6003 (N_6003,N_5134,N_4440);
nor U6004 (N_6004,N_5784,N_4738);
xnor U6005 (N_6005,N_5399,N_5251);
nand U6006 (N_6006,N_5548,N_4802);
and U6007 (N_6007,N_4182,N_4644);
nor U6008 (N_6008,N_4107,N_5882);
nand U6009 (N_6009,N_3804,N_4080);
or U6010 (N_6010,N_4768,N_3318);
nor U6011 (N_6011,N_3617,N_4563);
and U6012 (N_6012,N_4942,N_4286);
nor U6013 (N_6013,N_4600,N_3779);
nor U6014 (N_6014,N_3583,N_4064);
nand U6015 (N_6015,N_3600,N_5462);
or U6016 (N_6016,N_5569,N_3047);
or U6017 (N_6017,N_4884,N_5035);
or U6018 (N_6018,N_4908,N_3287);
nor U6019 (N_6019,N_4835,N_3139);
or U6020 (N_6020,N_3850,N_3688);
or U6021 (N_6021,N_5335,N_4566);
nor U6022 (N_6022,N_3672,N_3557);
and U6023 (N_6023,N_3699,N_3213);
or U6024 (N_6024,N_5832,N_5000);
nor U6025 (N_6025,N_5895,N_4420);
xor U6026 (N_6026,N_5991,N_4159);
and U6027 (N_6027,N_5065,N_4972);
nand U6028 (N_6028,N_4329,N_5810);
and U6029 (N_6029,N_3878,N_3016);
nand U6030 (N_6030,N_3169,N_4293);
nand U6031 (N_6031,N_3800,N_5336);
and U6032 (N_6032,N_4921,N_3320);
or U6033 (N_6033,N_4669,N_5532);
and U6034 (N_6034,N_3368,N_4624);
nand U6035 (N_6035,N_5677,N_5738);
or U6036 (N_6036,N_5406,N_4788);
nor U6037 (N_6037,N_5373,N_5706);
or U6038 (N_6038,N_3685,N_3412);
or U6039 (N_6039,N_4887,N_5740);
nor U6040 (N_6040,N_4785,N_5854);
nor U6041 (N_6041,N_4983,N_3994);
or U6042 (N_6042,N_5542,N_5675);
nor U6043 (N_6043,N_3783,N_3290);
nor U6044 (N_6044,N_5288,N_4550);
nand U6045 (N_6045,N_5010,N_5951);
or U6046 (N_6046,N_3604,N_3306);
nor U6047 (N_6047,N_4599,N_3934);
nor U6048 (N_6048,N_5001,N_4089);
and U6049 (N_6049,N_5683,N_3853);
or U6050 (N_6050,N_3032,N_3955);
nor U6051 (N_6051,N_3868,N_4055);
xnor U6052 (N_6052,N_3326,N_4341);
nor U6053 (N_6053,N_3455,N_4358);
and U6054 (N_6054,N_4122,N_3974);
nand U6055 (N_6055,N_4243,N_3612);
and U6056 (N_6056,N_3282,N_3474);
and U6057 (N_6057,N_3402,N_3593);
xnor U6058 (N_6058,N_3852,N_3664);
nand U6059 (N_6059,N_5702,N_3095);
nor U6060 (N_6060,N_4502,N_5521);
and U6061 (N_6061,N_3351,N_3297);
nor U6062 (N_6062,N_4086,N_4779);
nor U6063 (N_6063,N_3827,N_4536);
nor U6064 (N_6064,N_4244,N_4132);
nand U6065 (N_6065,N_4213,N_4965);
nor U6066 (N_6066,N_3772,N_4652);
nor U6067 (N_6067,N_5489,N_4354);
or U6068 (N_6068,N_4288,N_3810);
and U6069 (N_6069,N_4104,N_3922);
nand U6070 (N_6070,N_5312,N_5761);
and U6071 (N_6071,N_4390,N_3870);
nor U6072 (N_6072,N_3892,N_3837);
and U6073 (N_6073,N_5719,N_3425);
or U6074 (N_6074,N_5831,N_3982);
and U6075 (N_6075,N_5528,N_3533);
nor U6076 (N_6076,N_3219,N_5783);
nor U6077 (N_6077,N_4742,N_3648);
or U6078 (N_6078,N_4202,N_5496);
and U6079 (N_6079,N_5613,N_5184);
nor U6080 (N_6080,N_4548,N_4479);
and U6081 (N_6081,N_5989,N_3038);
nand U6082 (N_6082,N_3556,N_4228);
and U6083 (N_6083,N_4749,N_5865);
nor U6084 (N_6084,N_3854,N_4095);
nand U6085 (N_6085,N_4350,N_4953);
and U6086 (N_6086,N_5013,N_5529);
or U6087 (N_6087,N_4602,N_3792);
and U6088 (N_6088,N_3833,N_3541);
and U6089 (N_6089,N_3714,N_4445);
xor U6090 (N_6090,N_4611,N_3773);
or U6091 (N_6091,N_5705,N_4667);
and U6092 (N_6092,N_4625,N_3034);
or U6093 (N_6093,N_4336,N_5632);
and U6094 (N_6094,N_4844,N_5033);
and U6095 (N_6095,N_5370,N_5094);
nor U6096 (N_6096,N_4920,N_3592);
nand U6097 (N_6097,N_4333,N_5123);
nor U6098 (N_6098,N_5670,N_5599);
and U6099 (N_6099,N_3945,N_3177);
nand U6100 (N_6100,N_5735,N_4853);
nand U6101 (N_6101,N_4156,N_3285);
nor U6102 (N_6102,N_4585,N_4808);
or U6103 (N_6103,N_4342,N_4403);
nand U6104 (N_6104,N_5631,N_5728);
and U6105 (N_6105,N_3909,N_4000);
or U6106 (N_6106,N_5612,N_3023);
and U6107 (N_6107,N_3029,N_3226);
nor U6108 (N_6108,N_4805,N_5485);
and U6109 (N_6109,N_3159,N_4995);
nor U6110 (N_6110,N_5760,N_4395);
nand U6111 (N_6111,N_5525,N_3188);
or U6112 (N_6112,N_4813,N_5781);
and U6113 (N_6113,N_4928,N_3782);
or U6114 (N_6114,N_3230,N_3729);
and U6115 (N_6115,N_3420,N_5699);
and U6116 (N_6116,N_3633,N_4396);
nor U6117 (N_6117,N_3401,N_4949);
nand U6118 (N_6118,N_4485,N_5499);
nand U6119 (N_6119,N_4367,N_5465);
nand U6120 (N_6120,N_3698,N_3597);
or U6121 (N_6121,N_3722,N_3786);
or U6122 (N_6122,N_3618,N_5736);
nor U6123 (N_6123,N_5642,N_4145);
or U6124 (N_6124,N_4637,N_3116);
nand U6125 (N_6125,N_3927,N_5311);
and U6126 (N_6126,N_4128,N_4021);
nand U6127 (N_6127,N_3136,N_3280);
nand U6128 (N_6128,N_5063,N_4411);
and U6129 (N_6129,N_4981,N_5125);
and U6130 (N_6130,N_5050,N_4684);
and U6131 (N_6131,N_5064,N_4814);
and U6132 (N_6132,N_3579,N_4385);
and U6133 (N_6133,N_3052,N_4454);
nor U6134 (N_6134,N_4061,N_5137);
nand U6135 (N_6135,N_3665,N_3971);
or U6136 (N_6136,N_3405,N_5237);
and U6137 (N_6137,N_3216,N_4909);
nand U6138 (N_6138,N_3614,N_4362);
or U6139 (N_6139,N_3299,N_4489);
nand U6140 (N_6140,N_3577,N_5358);
nand U6141 (N_6141,N_4185,N_5165);
or U6142 (N_6142,N_4277,N_4007);
nor U6143 (N_6143,N_5585,N_4508);
nor U6144 (N_6144,N_4733,N_3527);
nor U6145 (N_6145,N_5955,N_5083);
and U6146 (N_6146,N_3210,N_4425);
and U6147 (N_6147,N_5303,N_3908);
or U6148 (N_6148,N_3910,N_3466);
or U6149 (N_6149,N_3179,N_5342);
nor U6150 (N_6150,N_4514,N_3742);
or U6151 (N_6151,N_4778,N_4859);
nand U6152 (N_6152,N_3814,N_3995);
nand U6153 (N_6153,N_4631,N_4278);
nand U6154 (N_6154,N_4346,N_4923);
nand U6155 (N_6155,N_4456,N_3375);
nand U6156 (N_6156,N_4063,N_4424);
and U6157 (N_6157,N_3166,N_3671);
nand U6158 (N_6158,N_3129,N_3142);
nor U6159 (N_6159,N_5162,N_3099);
or U6160 (N_6160,N_4961,N_4894);
and U6161 (N_6161,N_3239,N_5754);
and U6162 (N_6162,N_5648,N_5930);
nor U6163 (N_6163,N_3113,N_3434);
nand U6164 (N_6164,N_5669,N_5988);
or U6165 (N_6165,N_3015,N_4711);
or U6166 (N_6166,N_5115,N_3350);
and U6167 (N_6167,N_4708,N_4427);
nor U6168 (N_6168,N_4460,N_4946);
nor U6169 (N_6169,N_3638,N_4639);
and U6170 (N_6170,N_4221,N_4301);
nand U6171 (N_6171,N_5794,N_5449);
or U6172 (N_6172,N_4381,N_4579);
nand U6173 (N_6173,N_3738,N_4470);
and U6174 (N_6174,N_5331,N_3992);
nor U6175 (N_6175,N_3242,N_4555);
and U6176 (N_6176,N_4592,N_4591);
and U6177 (N_6177,N_3358,N_5554);
nand U6178 (N_6178,N_3330,N_4025);
nor U6179 (N_6179,N_5104,N_5444);
nor U6180 (N_6180,N_5961,N_5626);
nand U6181 (N_6181,N_5688,N_4292);
nand U6182 (N_6182,N_4051,N_3866);
and U6183 (N_6183,N_4604,N_5505);
and U6184 (N_6184,N_5809,N_4557);
nor U6185 (N_6185,N_4222,N_3082);
nand U6186 (N_6186,N_5332,N_4726);
and U6187 (N_6187,N_3925,N_3252);
nor U6188 (N_6188,N_5493,N_5179);
nor U6189 (N_6189,N_5696,N_3205);
or U6190 (N_6190,N_3173,N_4932);
or U6191 (N_6191,N_3568,N_4009);
nor U6192 (N_6192,N_5200,N_3947);
nand U6193 (N_6193,N_4931,N_4473);
nor U6194 (N_6194,N_3090,N_3885);
nor U6195 (N_6195,N_5112,N_5919);
or U6196 (N_6196,N_4183,N_3413);
or U6197 (N_6197,N_3333,N_4906);
or U6198 (N_6198,N_5518,N_5963);
or U6199 (N_6199,N_4694,N_5058);
nor U6200 (N_6200,N_4318,N_3826);
nor U6201 (N_6201,N_4515,N_3138);
or U6202 (N_6202,N_3549,N_4098);
and U6203 (N_6203,N_4247,N_3865);
and U6204 (N_6204,N_5440,N_5595);
nand U6205 (N_6205,N_3567,N_3377);
nand U6206 (N_6206,N_3632,N_4534);
nor U6207 (N_6207,N_5531,N_5119);
nand U6208 (N_6208,N_3378,N_3697);
and U6209 (N_6209,N_5384,N_5533);
nor U6210 (N_6210,N_3585,N_4116);
or U6211 (N_6211,N_5899,N_5016);
nand U6212 (N_6212,N_3392,N_4576);
nand U6213 (N_6213,N_5752,N_5435);
or U6214 (N_6214,N_3325,N_3973);
or U6215 (N_6215,N_4302,N_5775);
or U6216 (N_6216,N_4646,N_5026);
nor U6217 (N_6217,N_3211,N_4806);
nor U6218 (N_6218,N_4927,N_4203);
and U6219 (N_6219,N_3171,N_4809);
nand U6220 (N_6220,N_3332,N_3979);
nor U6221 (N_6221,N_4874,N_3884);
and U6222 (N_6222,N_5059,N_5944);
nor U6223 (N_6223,N_3978,N_5223);
and U6224 (N_6224,N_3367,N_5196);
and U6225 (N_6225,N_5733,N_5806);
nor U6226 (N_6226,N_3468,N_4135);
nand U6227 (N_6227,N_3707,N_3206);
nand U6228 (N_6228,N_3143,N_4355);
and U6229 (N_6229,N_4106,N_5984);
nand U6230 (N_6230,N_3644,N_3506);
nand U6231 (N_6231,N_4728,N_3106);
and U6232 (N_6232,N_5821,N_5971);
and U6233 (N_6233,N_3728,N_5615);
nor U6234 (N_6234,N_5429,N_4616);
nor U6235 (N_6235,N_3667,N_4560);
or U6236 (N_6236,N_5928,N_3319);
and U6237 (N_6237,N_4028,N_4648);
nor U6238 (N_6238,N_3340,N_4880);
nor U6239 (N_6239,N_5602,N_5351);
nand U6240 (N_6240,N_5708,N_5557);
nor U6241 (N_6241,N_4149,N_3675);
or U6242 (N_6242,N_5153,N_4745);
nand U6243 (N_6243,N_5594,N_3511);
and U6244 (N_6244,N_3003,N_5828);
nor U6245 (N_6245,N_4412,N_3057);
nand U6246 (N_6246,N_4864,N_3238);
nand U6247 (N_6247,N_5262,N_4663);
and U6248 (N_6248,N_3382,N_3235);
or U6249 (N_6249,N_3555,N_4488);
and U6250 (N_6250,N_3469,N_3510);
xnor U6251 (N_6251,N_5394,N_3119);
and U6252 (N_6252,N_3240,N_4042);
or U6253 (N_6253,N_3220,N_5036);
nand U6254 (N_6254,N_4672,N_3341);
nor U6255 (N_6255,N_5504,N_3643);
nor U6256 (N_6256,N_5427,N_5870);
or U6257 (N_6257,N_4752,N_5645);
nand U6258 (N_6258,N_5187,N_4328);
and U6259 (N_6259,N_4230,N_4282);
or U6260 (N_6260,N_5106,N_5866);
nand U6261 (N_6261,N_3861,N_5244);
and U6262 (N_6262,N_3396,N_3492);
nand U6263 (N_6263,N_5779,N_3938);
and U6264 (N_6264,N_5634,N_4034);
xnor U6265 (N_6265,N_4590,N_5417);
and U6266 (N_6266,N_3819,N_4759);
or U6267 (N_6267,N_4922,N_5097);
and U6268 (N_6268,N_3088,N_5679);
or U6269 (N_6269,N_4510,N_3383);
nor U6270 (N_6270,N_4316,N_4374);
and U6271 (N_6271,N_4498,N_5913);
nand U6272 (N_6272,N_5791,N_3441);
or U6273 (N_6273,N_4723,N_3011);
nor U6274 (N_6274,N_3508,N_5433);
xnor U6275 (N_6275,N_4163,N_4526);
nand U6276 (N_6276,N_5715,N_5932);
or U6277 (N_6277,N_3867,N_3463);
nor U6278 (N_6278,N_3362,N_5346);
nand U6279 (N_6279,N_3303,N_5713);
and U6280 (N_6280,N_5676,N_4559);
and U6281 (N_6281,N_3208,N_5609);
nor U6282 (N_6282,N_4349,N_5726);
nand U6283 (N_6283,N_3569,N_4210);
nor U6284 (N_6284,N_4685,N_3739);
and U6285 (N_6285,N_5297,N_5091);
nor U6286 (N_6286,N_4584,N_3020);
and U6287 (N_6287,N_5302,N_4661);
nand U6288 (N_6288,N_4391,N_5183);
nor U6289 (N_6289,N_5490,N_3127);
and U6290 (N_6290,N_4945,N_3635);
nor U6291 (N_6291,N_5694,N_4597);
xnor U6292 (N_6292,N_5575,N_4455);
nand U6293 (N_6293,N_4180,N_3077);
nand U6294 (N_6294,N_3869,N_4012);
nor U6295 (N_6295,N_3515,N_4044);
or U6296 (N_6296,N_3754,N_3493);
nor U6297 (N_6297,N_3831,N_3897);
nand U6298 (N_6298,N_4799,N_3223);
nor U6299 (N_6299,N_5966,N_3312);
or U6300 (N_6300,N_5170,N_5933);
nand U6301 (N_6301,N_3603,N_3845);
and U6302 (N_6302,N_3611,N_3460);
or U6303 (N_6303,N_3946,N_5566);
nor U6304 (N_6304,N_4308,N_5603);
nand U6305 (N_6305,N_5028,N_5689);
nor U6306 (N_6306,N_4429,N_3112);
and U6307 (N_6307,N_4982,N_4251);
or U6308 (N_6308,N_5375,N_3091);
or U6309 (N_6309,N_3051,N_3905);
or U6310 (N_6310,N_3962,N_3181);
and U6311 (N_6311,N_4573,N_5473);
nor U6312 (N_6312,N_3912,N_4992);
or U6313 (N_6313,N_5942,N_3929);
xor U6314 (N_6314,N_5885,N_3153);
nand U6315 (N_6315,N_5144,N_3305);
nand U6316 (N_6316,N_4193,N_4314);
and U6317 (N_6317,N_3704,N_5099);
and U6318 (N_6318,N_3735,N_3941);
nand U6319 (N_6319,N_3162,N_3572);
and U6320 (N_6320,N_3674,N_5999);
or U6321 (N_6321,N_4140,N_3763);
or U6322 (N_6322,N_5629,N_5041);
and U6323 (N_6323,N_5608,N_3989);
nor U6324 (N_6324,N_4139,N_3203);
nor U6325 (N_6325,N_5328,N_3295);
nand U6326 (N_6326,N_4925,N_5729);
nand U6327 (N_6327,N_3943,N_3651);
or U6328 (N_6328,N_3744,N_4101);
and U6329 (N_6329,N_4129,N_4975);
nor U6330 (N_6330,N_3496,N_3229);
nand U6331 (N_6331,N_4587,N_4376);
nand U6332 (N_6332,N_5839,N_4197);
nand U6333 (N_6333,N_3394,N_4580);
or U6334 (N_6334,N_3265,N_4120);
or U6335 (N_6335,N_4141,N_4311);
nand U6336 (N_6336,N_4653,N_5032);
nor U6337 (N_6337,N_5363,N_5453);
nor U6338 (N_6338,N_3209,N_5527);
and U6339 (N_6339,N_3264,N_3544);
nand U6340 (N_6340,N_3446,N_3634);
nor U6341 (N_6341,N_5168,N_3900);
or U6342 (N_6342,N_5926,N_5310);
or U6343 (N_6343,N_5567,N_5261);
or U6344 (N_6344,N_5847,N_5546);
or U6345 (N_6345,N_5901,N_5247);
xor U6346 (N_6346,N_5222,N_5717);
nor U6347 (N_6347,N_3288,N_3871);
nand U6348 (N_6348,N_3385,N_3680);
and U6349 (N_6349,N_4735,N_3178);
and U6350 (N_6350,N_4369,N_3694);
or U6351 (N_6351,N_3953,N_3231);
nor U6352 (N_6352,N_5344,N_5309);
nand U6353 (N_6353,N_5239,N_5927);
or U6354 (N_6354,N_5484,N_5763);
or U6355 (N_6355,N_3050,N_5579);
or U6356 (N_6356,N_3349,N_5042);
and U6357 (N_6357,N_5408,N_3566);
or U6358 (N_6358,N_4124,N_5886);
and U6359 (N_6359,N_4053,N_3993);
nand U6360 (N_6360,N_3610,N_4237);
and U6361 (N_6361,N_3608,N_3967);
or U6362 (N_6362,N_5737,N_4561);
or U6363 (N_6363,N_4645,N_3484);
or U6364 (N_6364,N_5205,N_3135);
nand U6365 (N_6365,N_5007,N_5843);
or U6366 (N_6366,N_3789,N_3207);
and U6367 (N_6367,N_5896,N_4383);
nor U6368 (N_6368,N_5568,N_3311);
nor U6369 (N_6369,N_5638,N_5418);
or U6370 (N_6370,N_3073,N_5559);
and U6371 (N_6371,N_3234,N_4966);
nand U6372 (N_6372,N_4207,N_3085);
nand U6373 (N_6373,N_3898,N_3684);
nand U6374 (N_6374,N_4245,N_4365);
nand U6375 (N_6375,N_3344,N_4954);
nor U6376 (N_6376,N_3840,N_4939);
nand U6377 (N_6377,N_4831,N_3501);
and U6378 (N_6378,N_5338,N_3903);
and U6379 (N_6379,N_5392,N_4650);
nand U6380 (N_6380,N_4709,N_5700);
nand U6381 (N_6381,N_4327,N_5122);
xnor U6382 (N_6382,N_4447,N_4643);
nand U6383 (N_6383,N_4937,N_5234);
nor U6384 (N_6384,N_5053,N_4360);
nor U6385 (N_6385,N_5691,N_3727);
nand U6386 (N_6386,N_5714,N_4505);
nor U6387 (N_6387,N_4168,N_3645);
or U6388 (N_6388,N_4705,N_3761);
or U6389 (N_6389,N_5003,N_3649);
and U6390 (N_6390,N_4236,N_3580);
or U6391 (N_6391,N_4770,N_4732);
nor U6392 (N_6392,N_4895,N_4165);
and U6393 (N_6393,N_3829,N_5098);
and U6394 (N_6394,N_4774,N_4513);
nor U6395 (N_6395,N_4442,N_5758);
or U6396 (N_6396,N_4626,N_4309);
nand U6397 (N_6397,N_3278,N_3111);
and U6398 (N_6398,N_5169,N_5259);
nor U6399 (N_6399,N_4013,N_5684);
and U6400 (N_6400,N_5159,N_4551);
and U6401 (N_6401,N_5152,N_3182);
nor U6402 (N_6402,N_5537,N_5080);
nand U6403 (N_6403,N_4876,N_5350);
nor U6404 (N_6404,N_4431,N_5863);
and U6405 (N_6405,N_3808,N_4541);
and U6406 (N_6406,N_4615,N_3110);
and U6407 (N_6407,N_4636,N_4969);
nor U6408 (N_6408,N_3855,N_5596);
nand U6409 (N_6409,N_3801,N_5658);
nor U6410 (N_6410,N_3048,N_4421);
and U6411 (N_6411,N_4003,N_4727);
and U6412 (N_6412,N_5628,N_5040);
and U6413 (N_6413,N_5678,N_5268);
nand U6414 (N_6414,N_3626,N_5514);
nand U6415 (N_6415,N_3118,N_5512);
and U6416 (N_6416,N_3530,N_4899);
or U6417 (N_6417,N_3309,N_4389);
and U6418 (N_6418,N_3594,N_5477);
nand U6419 (N_6419,N_4674,N_5280);
or U6420 (N_6420,N_4205,N_5687);
nand U6421 (N_6421,N_3408,N_4570);
nor U6422 (N_6422,N_3454,N_3335);
nand U6423 (N_6423,N_3010,N_5037);
or U6424 (N_6424,N_5869,N_4756);
nor U6425 (N_6425,N_3355,N_5903);
or U6426 (N_6426,N_3079,N_5052);
nand U6427 (N_6427,N_4257,N_3163);
and U6428 (N_6428,N_3915,N_3361);
and U6429 (N_6429,N_5747,N_4138);
nor U6430 (N_6430,N_5166,N_4529);
nor U6431 (N_6431,N_3721,N_4158);
nor U6432 (N_6432,N_5413,N_4109);
or U6433 (N_6433,N_3894,N_5255);
and U6434 (N_6434,N_4148,N_3954);
or U6435 (N_6435,N_5103,N_3609);
nor U6436 (N_6436,N_3637,N_4402);
nor U6437 (N_6437,N_4268,N_5133);
and U6438 (N_6438,N_5952,N_4273);
xnor U6439 (N_6439,N_3433,N_3862);
or U6440 (N_6440,N_3526,N_4860);
or U6441 (N_6441,N_4338,N_5421);
nand U6442 (N_6442,N_5136,N_4875);
nor U6443 (N_6443,N_4495,N_5466);
nand U6444 (N_6444,N_4234,N_5401);
nand U6445 (N_6445,N_3777,N_5293);
or U6446 (N_6446,N_3768,N_5150);
and U6447 (N_6447,N_3940,N_4803);
nor U6448 (N_6448,N_4994,N_4100);
nand U6449 (N_6449,N_5539,N_3719);
nand U6450 (N_6450,N_5432,N_4056);
and U6451 (N_6451,N_3660,N_5285);
nand U6452 (N_6452,N_4067,N_5154);
nand U6453 (N_6453,N_4815,N_3123);
or U6454 (N_6454,N_5057,N_5235);
nor U6455 (N_6455,N_5348,N_5386);
nor U6456 (N_6456,N_5858,N_3370);
or U6457 (N_6457,N_3830,N_4285);
nor U6458 (N_6458,N_5793,N_4816);
nor U6459 (N_6459,N_4487,N_5667);
nor U6460 (N_6460,N_4010,N_5476);
or U6461 (N_6461,N_3384,N_4522);
nand U6462 (N_6462,N_3710,N_3558);
or U6463 (N_6463,N_4941,N_3294);
or U6464 (N_6464,N_5853,N_5107);
or U6465 (N_6465,N_4692,N_3167);
and U6466 (N_6466,N_3559,N_5622);
or U6467 (N_6467,N_4558,N_5522);
and U6468 (N_6468,N_3314,N_4608);
and U6469 (N_6469,N_5398,N_4673);
nor U6470 (N_6470,N_5047,N_5197);
nand U6471 (N_6471,N_3199,N_3150);
nor U6472 (N_6472,N_4690,N_3409);
and U6473 (N_6473,N_4220,N_4085);
xnor U6474 (N_6474,N_3832,N_4571);
nor U6475 (N_6475,N_3793,N_5495);
nand U6476 (N_6476,N_3961,N_4229);
or U6477 (N_6477,N_4492,N_4112);
xnor U6478 (N_6478,N_4170,N_3730);
or U6479 (N_6479,N_4885,N_5232);
nor U6480 (N_6480,N_5448,N_4322);
nor U6481 (N_6481,N_4361,N_5402);
or U6482 (N_6482,N_5323,N_3658);
nor U6483 (N_6483,N_4613,N_3273);
nand U6484 (N_6484,N_4696,N_3522);
nor U6485 (N_6485,N_5390,N_5551);
nor U6486 (N_6486,N_3596,N_4532);
nor U6487 (N_6487,N_4710,N_3485);
and U6488 (N_6488,N_5250,N_4486);
nor U6489 (N_6489,N_5871,N_5175);
or U6490 (N_6490,N_3045,N_5282);
and U6491 (N_6491,N_4832,N_4054);
and U6492 (N_6492,N_5653,N_4845);
nand U6493 (N_6493,N_4271,N_3125);
nor U6494 (N_6494,N_3743,N_4430);
nor U6495 (N_6495,N_3751,N_3061);
nor U6496 (N_6496,N_5308,N_4688);
nor U6497 (N_6497,N_4800,N_3712);
xnor U6498 (N_6498,N_3121,N_5487);
nor U6499 (N_6499,N_4962,N_4320);
or U6500 (N_6500,N_4950,N_3194);
nor U6501 (N_6501,N_3165,N_3507);
or U6502 (N_6502,N_4680,N_5674);
and U6503 (N_6503,N_4699,N_3711);
or U6504 (N_6504,N_4114,N_5884);
nor U6505 (N_6505,N_4415,N_4693);
nand U6506 (N_6506,N_4232,N_4484);
or U6507 (N_6507,N_4675,N_3505);
or U6508 (N_6508,N_4629,N_3520);
nand U6509 (N_6509,N_3232,N_5666);
nor U6510 (N_6510,N_3578,N_4724);
and U6511 (N_6511,N_3966,N_5787);
nand U6512 (N_6512,N_4393,N_5266);
nand U6513 (N_6513,N_5359,N_5580);
nor U6514 (N_6514,N_5269,N_5074);
nor U6515 (N_6515,N_4744,N_4047);
and U6516 (N_6516,N_3775,N_4521);
and U6517 (N_6517,N_3310,N_3835);
or U6518 (N_6518,N_5424,N_3005);
or U6519 (N_6519,N_4839,N_4188);
and U6520 (N_6520,N_3689,N_3004);
nand U6521 (N_6521,N_4397,N_5108);
and U6522 (N_6522,N_5274,N_3075);
nand U6523 (N_6523,N_3184,N_4782);
and U6524 (N_6524,N_4166,N_4910);
nand U6525 (N_6525,N_4016,N_4960);
or U6526 (N_6526,N_3902,N_5723);
and U6527 (N_6527,N_4538,N_3322);
nand U6528 (N_6528,N_4714,N_4248);
nor U6529 (N_6529,N_3481,N_3981);
and U6530 (N_6530,N_5639,N_4968);
nor U6531 (N_6531,N_3987,N_5840);
nor U6532 (N_6532,N_3054,N_3859);
xnor U6533 (N_6533,N_5770,N_5786);
and U6534 (N_6534,N_3937,N_5617);
or U6535 (N_6535,N_3233,N_3126);
nand U6536 (N_6536,N_4984,N_4605);
nor U6537 (N_6537,N_5409,N_4052);
or U6538 (N_6538,N_4997,N_5535);
or U6539 (N_6539,N_4072,N_4583);
or U6540 (N_6540,N_4419,N_4443);
nor U6541 (N_6541,N_5464,N_4235);
or U6542 (N_6542,N_4111,N_4824);
or U6543 (N_6543,N_5983,N_4208);
nor U6544 (N_6544,N_5271,N_4147);
nand U6545 (N_6545,N_4270,N_3251);
and U6546 (N_6546,N_5056,N_3292);
or U6547 (N_6547,N_3620,N_4088);
nor U6548 (N_6548,N_4134,N_3906);
and U6549 (N_6549,N_4882,N_5668);
nand U6550 (N_6550,N_3274,N_4015);
or U6551 (N_6551,N_3822,N_5388);
nor U6552 (N_6552,N_5654,N_5078);
nor U6553 (N_6553,N_5004,N_3070);
nand U6554 (N_6554,N_3646,N_4062);
and U6555 (N_6555,N_3942,N_4433);
or U6556 (N_6556,N_4986,N_5656);
and U6557 (N_6557,N_4018,N_3078);
or U6558 (N_6558,N_3964,N_3042);
or U6559 (N_6559,N_5383,N_3803);
or U6560 (N_6560,N_5181,N_5367);
or U6561 (N_6561,N_3191,N_4356);
nand U6562 (N_6562,N_5724,N_4703);
or U6563 (N_6563,N_3570,N_4115);
nor U6564 (N_6564,N_5278,N_4936);
or U6565 (N_6565,N_4843,N_4797);
and U6566 (N_6566,N_5534,N_5426);
nand U6567 (N_6567,N_5826,N_5965);
nand U6568 (N_6568,N_5650,N_3124);
or U6569 (N_6569,N_3214,N_5226);
nand U6570 (N_6570,N_5956,N_4905);
nand U6571 (N_6571,N_5949,N_5252);
nor U6572 (N_6572,N_3186,N_5396);
nand U6573 (N_6573,N_3502,N_5637);
nand U6574 (N_6574,N_5818,N_3849);
and U6575 (N_6575,N_3053,N_4697);
or U6576 (N_6576,N_3702,N_5290);
or U6577 (N_6577,N_5354,N_3930);
and U6578 (N_6578,N_4276,N_3838);
nor U6579 (N_6579,N_5541,N_4174);
or U6580 (N_6580,N_3025,N_3115);
or U6581 (N_6581,N_4252,N_5996);
nand U6582 (N_6582,N_3130,N_4090);
nor U6583 (N_6583,N_3598,N_5193);
nor U6584 (N_6584,N_3676,N_4640);
and U6585 (N_6585,N_4623,N_5459);
and U6586 (N_6586,N_3324,N_5973);
nor U6587 (N_6587,N_3696,N_3062);
or U6588 (N_6588,N_4204,N_5501);
nand U6589 (N_6589,N_5046,N_3323);
or U6590 (N_6590,N_3261,N_5701);
nand U6591 (N_6591,N_3448,N_3331);
nand U6592 (N_6592,N_3753,N_4030);
nand U6593 (N_6593,N_3403,N_5540);
and U6594 (N_6594,N_4416,N_3740);
or U6595 (N_6595,N_3788,N_3356);
or U6596 (N_6596,N_4312,N_5439);
or U6597 (N_6597,N_5883,N_3197);
and U6598 (N_6598,N_3543,N_3345);
xnor U6599 (N_6599,N_5757,N_4105);
nand U6600 (N_6600,N_4610,N_3872);
nor U6601 (N_6601,N_4533,N_5238);
nor U6602 (N_6602,N_3464,N_3300);
nor U6603 (N_6603,N_5876,N_4630);
or U6604 (N_6604,N_5646,N_3107);
and U6605 (N_6605,N_5993,N_3263);
and U6606 (N_6606,N_4904,N_3796);
nand U6607 (N_6607,N_4857,N_5571);
or U6608 (N_6608,N_4041,N_3026);
nor U6609 (N_6609,N_5703,N_3039);
nand U6610 (N_6610,N_5389,N_4450);
nand U6611 (N_6611,N_5836,N_5267);
nand U6612 (N_6612,N_5012,N_4729);
or U6613 (N_6613,N_4544,N_3784);
nor U6614 (N_6614,N_5697,N_5024);
nor U6615 (N_6615,N_3161,N_3540);
and U6616 (N_6616,N_5834,N_3440);
or U6617 (N_6617,N_4295,N_5921);
and U6618 (N_6618,N_5355,N_5563);
and U6619 (N_6619,N_3926,N_3874);
nor U6620 (N_6620,N_5085,N_3427);
nand U6621 (N_6621,N_4066,N_5570);
and U6622 (N_6622,N_3007,N_3516);
nor U6623 (N_6623,N_3030,N_3647);
and U6624 (N_6624,N_5782,N_3266);
xor U6625 (N_6625,N_3602,N_4266);
or U6626 (N_6626,N_4957,N_5910);
xor U6627 (N_6627,N_5385,N_4664);
nor U6628 (N_6628,N_5422,N_3542);
nor U6629 (N_6629,N_5908,N_4441);
and U6630 (N_6630,N_3058,N_4594);
nor U6631 (N_6631,N_3489,N_3066);
nand U6632 (N_6632,N_3997,N_3825);
or U6633 (N_6633,N_4930,N_4747);
or U6634 (N_6634,N_5589,N_4238);
or U6635 (N_6635,N_5864,N_4279);
or U6636 (N_6636,N_5372,N_3247);
and U6637 (N_6637,N_5220,N_5326);
or U6638 (N_6638,N_3301,N_5822);
or U6639 (N_6639,N_3895,N_3488);
or U6640 (N_6640,N_3764,N_4934);
and U6641 (N_6641,N_5415,N_4294);
nor U6642 (N_6642,N_5002,N_5281);
nand U6643 (N_6643,N_3277,N_4092);
and U6644 (N_6644,N_5588,N_4171);
nand U6645 (N_6645,N_4913,N_5147);
nand U6646 (N_6646,N_3093,N_3436);
and U6647 (N_6647,N_4741,N_3695);
nand U6648 (N_6648,N_5544,N_4049);
nor U6649 (N_6649,N_4043,N_3131);
and U6650 (N_6650,N_3636,N_5460);
nand U6651 (N_6651,N_4209,N_5048);
nor U6652 (N_6652,N_4005,N_4951);
or U6653 (N_6653,N_4856,N_3512);
nand U6654 (N_6654,N_3094,N_3587);
and U6655 (N_6655,N_5815,N_5657);
and U6656 (N_6656,N_4979,N_3584);
or U6657 (N_6657,N_5777,N_3518);
or U6658 (N_6658,N_5077,N_5089);
or U6659 (N_6659,N_4914,N_5210);
nor U6660 (N_6660,N_4475,N_3858);
nand U6661 (N_6661,N_5550,N_3400);
or U6662 (N_6662,N_5746,N_5019);
and U6663 (N_6663,N_5241,N_3426);
nand U6664 (N_6664,N_5076,N_5124);
nand U6665 (N_6665,N_3769,N_4911);
nor U6666 (N_6666,N_5900,N_5368);
or U6667 (N_6667,N_4372,N_5874);
nor U6668 (N_6668,N_4796,N_4472);
nand U6669 (N_6669,N_5206,N_4506);
or U6670 (N_6670,N_4263,N_4363);
nand U6671 (N_6671,N_3140,N_4087);
nand U6672 (N_6672,N_5405,N_5143);
or U6673 (N_6673,N_3490,N_5482);
nor U6674 (N_6674,N_5954,N_3074);
nor U6675 (N_6675,N_3883,N_5817);
nor U6676 (N_6676,N_5498,N_5188);
and U6677 (N_6677,N_3687,N_3619);
or U6678 (N_6678,N_4357,N_4289);
or U6679 (N_6679,N_5739,N_3360);
and U6680 (N_6680,N_3456,N_3438);
nor U6681 (N_6681,N_5769,N_5022);
or U6682 (N_6682,N_4463,N_3771);
nor U6683 (N_6683,N_4461,N_5618);
nor U6684 (N_6684,N_3797,N_4084);
nor U6685 (N_6685,N_3650,N_5315);
and U6686 (N_6686,N_4601,N_4280);
nand U6687 (N_6687,N_3313,N_5938);
and U6688 (N_6688,N_4339,N_4126);
nor U6689 (N_6689,N_4706,N_4507);
and U6690 (N_6690,N_3758,N_4315);
or U6691 (N_6691,N_5463,N_4058);
nand U6692 (N_6692,N_5395,N_5176);
or U6693 (N_6693,N_3098,N_5621);
and U6694 (N_6694,N_4110,N_4448);
nand U6695 (N_6695,N_4720,N_4689);
nor U6696 (N_6696,N_5102,N_4303);
and U6697 (N_6697,N_4117,N_5998);
and U6698 (N_6698,N_4539,N_4503);
and U6699 (N_6699,N_4748,N_4352);
and U6700 (N_6700,N_3795,N_3044);
nand U6701 (N_6701,N_4400,N_4348);
nor U6702 (N_6702,N_3439,N_5664);
nand U6703 (N_6703,N_5256,N_5920);
nand U6704 (N_6704,N_3726,N_3725);
and U6705 (N_6705,N_3731,N_5471);
and U6706 (N_6706,N_3141,N_4133);
nor U6707 (N_6707,N_4099,N_5140);
xor U6708 (N_6708,N_3380,N_4162);
nand U6709 (N_6709,N_5199,N_5709);
nor U6710 (N_6710,N_5564,N_5291);
xnor U6711 (N_6711,N_3591,N_5092);
or U6712 (N_6712,N_5730,N_4572);
nor U6713 (N_6713,N_5149,N_4666);
nand U6714 (N_6714,N_5827,N_4467);
and U6715 (N_6715,N_5587,N_5227);
nor U6716 (N_6716,N_3221,N_3663);
or U6717 (N_6717,N_5470,N_4501);
nor U6718 (N_6718,N_3709,N_5819);
nor U6719 (N_6719,N_5880,N_5911);
or U6720 (N_6720,N_5488,N_3969);
nand U6721 (N_6721,N_3755,N_3374);
and U6722 (N_6722,N_4256,N_4578);
xnor U6723 (N_6723,N_3774,N_5081);
or U6724 (N_6724,N_4033,N_4491);
or U6725 (N_6725,N_4811,N_4031);
and U6726 (N_6726,N_5069,N_5204);
or U6727 (N_6727,N_4436,N_4635);
and U6728 (N_6728,N_3972,N_4048);
nor U6729 (N_6729,N_4649,N_4094);
or U6730 (N_6730,N_3573,N_4214);
nor U6731 (N_6731,N_4588,N_5841);
or U6732 (N_6732,N_4980,N_5055);
nor U6733 (N_6733,N_3500,N_5855);
nand U6734 (N_6734,N_4973,N_3901);
or U6735 (N_6735,N_4985,N_5096);
nor U6736 (N_6736,N_3415,N_3933);
nand U6737 (N_6737,N_4497,N_5034);
or U6738 (N_6738,N_3478,N_5095);
nor U6739 (N_6739,N_4304,N_3886);
and U6740 (N_6740,N_3873,N_4186);
and U6741 (N_6741,N_3407,N_5443);
nor U6742 (N_6742,N_4524,N_3037);
nand U6743 (N_6743,N_4763,N_3834);
nor U6744 (N_6744,N_4651,N_3002);
nor U6745 (N_6745,N_3613,N_5231);
and U6746 (N_6746,N_3423,N_3628);
or U6747 (N_6747,N_4617,N_3601);
nand U6748 (N_6748,N_3068,N_3387);
and U6749 (N_6749,N_4375,N_4240);
and U6750 (N_6750,N_3701,N_3089);
nor U6751 (N_6751,N_5295,N_5148);
nand U6752 (N_6752,N_5378,N_4704);
nor U6753 (N_6753,N_3035,N_5614);
or U6754 (N_6754,N_3575,N_3913);
or U6755 (N_6755,N_5593,N_4671);
nand U6756 (N_6756,N_5929,N_5180);
or U6757 (N_6757,N_3398,N_3262);
nor U6758 (N_6758,N_5643,N_3395);
and U6759 (N_6759,N_4725,N_5414);
xor U6760 (N_6760,N_4736,N_5314);
nor U6761 (N_6761,N_4812,N_4823);
nand U6762 (N_6762,N_5404,N_3256);
nor U6763 (N_6763,N_5649,N_5474);
and U6764 (N_6764,N_4272,N_4596);
and U6765 (N_6765,N_3847,N_4537);
nand U6766 (N_6766,N_4078,N_4216);
and U6767 (N_6767,N_4881,N_4035);
or U6768 (N_6768,N_3662,N_3655);
and U6769 (N_6769,N_4801,N_3154);
and U6770 (N_6770,N_4001,N_5986);
or U6771 (N_6771,N_3321,N_5073);
or U6772 (N_6772,N_5497,N_3562);
and U6773 (N_6773,N_3806,N_3548);
and U6774 (N_6774,N_3641,N_4172);
nor U6775 (N_6775,N_3482,N_4408);
nand U6776 (N_6776,N_3736,N_5105);
or U6777 (N_6777,N_4940,N_4900);
or U6778 (N_6778,N_3734,N_3843);
or U6779 (N_6779,N_5712,N_5194);
and U6780 (N_6780,N_3316,N_3022);
nor U6781 (N_6781,N_4196,N_5857);
and U6782 (N_6782,N_4353,N_3778);
nand U6783 (N_6783,N_5325,N_5859);
xor U6784 (N_6784,N_5682,N_5451);
or U6785 (N_6785,N_5129,N_4218);
nor U6786 (N_6786,N_3281,N_4718);
and U6787 (N_6787,N_4449,N_3960);
nor U6788 (N_6788,N_4854,N_4173);
or U6789 (N_6789,N_4493,N_4231);
or U6790 (N_6790,N_4634,N_3465);
or U6791 (N_6791,N_5079,N_5319);
or U6792 (N_6792,N_5289,N_4879);
or U6793 (N_6793,N_3588,N_4260);
nor U6794 (N_6794,N_3794,N_5214);
nor U6795 (N_6795,N_5330,N_4780);
nor U6796 (N_6796,N_4317,N_3134);
nand U6797 (N_6797,N_3390,N_4828);
nand U6798 (N_6798,N_3391,N_3365);
nor U6799 (N_6799,N_4190,N_4761);
nand U6800 (N_6800,N_5767,N_5054);
nor U6801 (N_6801,N_4130,N_3673);
or U6802 (N_6802,N_4877,N_4458);
and U6803 (N_6803,N_4096,N_5038);
nor U6804 (N_6804,N_3419,N_4437);
nand U6805 (N_6805,N_5647,N_5975);
nor U6806 (N_6806,N_4091,N_4713);
nand U6807 (N_6807,N_5573,N_4211);
nand U6808 (N_6808,N_4682,N_4019);
nand U6809 (N_6809,N_4478,N_3275);
or U6810 (N_6810,N_3693,N_5862);
or U6811 (N_6811,N_3339,N_3092);
or U6812 (N_6812,N_5155,N_3120);
nand U6813 (N_6813,N_3957,N_3479);
nand U6814 (N_6814,N_4660,N_3733);
nor U6815 (N_6815,N_4791,N_4841);
or U6816 (N_6816,N_4568,N_4261);
nor U6817 (N_6817,N_5100,N_4902);
nand U6818 (N_6818,N_3245,N_3017);
and U6819 (N_6819,N_3158,N_4123);
or U6820 (N_6820,N_5468,N_5327);
nand U6821 (N_6821,N_4603,N_5520);
or U6822 (N_6822,N_5627,N_3371);
nand U6823 (N_6823,N_3629,N_5720);
nand U6824 (N_6824,N_4556,N_3805);
nor U6825 (N_6825,N_4781,N_4848);
or U6826 (N_6826,N_5364,N_4306);
nand U6827 (N_6827,N_5800,N_3257);
nor U6828 (N_6828,N_4434,N_3080);
and U6829 (N_6829,N_5380,N_5867);
and U6830 (N_6830,N_5114,N_3244);
nand U6831 (N_6831,N_3315,N_5510);
nand U6832 (N_6832,N_4771,N_4577);
nand U6833 (N_6833,N_4952,N_3681);
and U6834 (N_6834,N_4574,N_5254);
or U6835 (N_6835,N_5695,N_3013);
or U6836 (N_6836,N_5860,N_3864);
nor U6837 (N_6837,N_5582,N_3893);
and U6838 (N_6838,N_3748,N_3406);
or U6839 (N_6839,N_5031,N_5765);
or U6840 (N_6840,N_4017,N_3828);
nand U6841 (N_6841,N_5229,N_3352);
and U6842 (N_6842,N_4167,N_3364);
nor U6843 (N_6843,N_5116,N_5716);
or U6844 (N_6844,N_3813,N_4773);
nor U6845 (N_6845,N_5890,N_4175);
nor U6846 (N_6846,N_4826,N_3535);
or U6847 (N_6847,N_5978,N_5916);
or U6848 (N_6848,N_5341,N_5692);
nand U6849 (N_6849,N_3453,N_3217);
nor U6850 (N_6850,N_3999,N_4784);
nand U6851 (N_6851,N_5797,N_3065);
and U6852 (N_6852,N_3574,N_4686);
or U6853 (N_6853,N_3616,N_4766);
nand U6854 (N_6854,N_3713,N_4737);
nor U6855 (N_6855,N_3877,N_3504);
and U6856 (N_6856,N_3204,N_5833);
nor U6857 (N_6857,N_3586,N_4681);
nor U6858 (N_6858,N_5011,N_5263);
nor U6859 (N_6859,N_3146,N_3152);
nor U6860 (N_6860,N_4281,N_3424);
nor U6861 (N_6861,N_3248,N_4212);
or U6862 (N_6862,N_4977,N_4739);
nand U6863 (N_6863,N_5049,N_4407);
nand U6864 (N_6864,N_4332,N_5798);
nand U6865 (N_6865,N_4545,N_3590);
nor U6866 (N_6866,N_3951,N_5307);
or U6867 (N_6867,N_5759,N_3006);
or U6868 (N_6868,N_4399,N_5294);
and U6869 (N_6869,N_5936,N_5279);
nor U6870 (N_6870,N_3986,N_3625);
or U6871 (N_6871,N_5808,N_5875);
nor U6872 (N_6872,N_5878,N_3475);
nand U6873 (N_6873,N_4284,N_3338);
or U6874 (N_6874,N_3703,N_4511);
nor U6875 (N_6875,N_5640,N_3984);
and U6876 (N_6876,N_5872,N_5379);
or U6877 (N_6877,N_4873,N_5352);
and U6878 (N_6878,N_4633,N_4948);
nand U6879 (N_6879,N_5578,N_5663);
or U6880 (N_6880,N_4901,N_4386);
or U6881 (N_6881,N_4380,N_5624);
and U6882 (N_6882,N_5958,N_5120);
or U6883 (N_6883,N_3899,N_3963);
nor U6884 (N_6884,N_5959,N_3914);
nor U6885 (N_6885,N_3747,N_4020);
and U6886 (N_6886,N_4988,N_3534);
nor U6887 (N_6887,N_4519,N_3414);
nor U6888 (N_6888,N_5732,N_5178);
nor U6889 (N_6889,N_4422,N_5655);
nor U6890 (N_6890,N_5992,N_3737);
nor U6891 (N_6891,N_4772,N_3958);
nand U6892 (N_6892,N_5948,N_3581);
or U6893 (N_6893,N_5776,N_3514);
or U6894 (N_6894,N_3347,N_4036);
and U6895 (N_6895,N_5635,N_4423);
nand U6896 (N_6896,N_3008,N_3532);
nor U6897 (N_6897,N_3480,N_4068);
or U6898 (N_6898,N_5680,N_4990);
nand U6899 (N_6899,N_3807,N_4083);
nor U6900 (N_6900,N_4153,N_4413);
or U6901 (N_6901,N_4071,N_5852);
and U6902 (N_6902,N_4792,N_5407);
nor U6903 (N_6903,N_5045,N_4074);
nand U6904 (N_6904,N_5286,N_5127);
nand U6905 (N_6905,N_3105,N_3393);
or U6906 (N_6906,N_3189,N_5611);
or U6907 (N_6907,N_5607,N_4565);
or U6908 (N_6908,N_5524,N_3881);
nand U6909 (N_6909,N_3627,N_5762);
nor U6910 (N_6910,N_5318,N_4225);
nand U6911 (N_6911,N_3196,N_5813);
nand U6912 (N_6912,N_5851,N_4337);
and U6913 (N_6913,N_5905,N_5316);
nor U6914 (N_6914,N_5185,N_3790);
nor U6915 (N_6915,N_3890,N_4943);
nand U6916 (N_6916,N_5718,N_4482);
nor U6917 (N_6917,N_5939,N_4959);
or U6918 (N_6918,N_4269,N_4804);
and U6919 (N_6919,N_5146,N_5017);
nand U6920 (N_6920,N_5067,N_4589);
nor U6921 (N_6921,N_5277,N_3304);
or U6922 (N_6922,N_3056,N_5075);
nand U6923 (N_6923,N_4750,N_4569);
xnor U6924 (N_6924,N_4552,N_5925);
or U6925 (N_6925,N_3677,N_3546);
nor U6926 (N_6926,N_4564,N_3151);
nand U6927 (N_6927,N_4275,N_5774);
nor U6928 (N_6928,N_4516,N_4575);
or U6929 (N_6929,N_4394,N_5411);
nor U6930 (N_6930,N_5132,N_3630);
nand U6931 (N_6931,N_3547,N_5478);
and U6932 (N_6932,N_3968,N_3097);
nand U6933 (N_6933,N_4897,N_4287);
nor U6934 (N_6934,N_5592,N_4893);
or U6935 (N_6935,N_5523,N_4863);
and U6936 (N_6936,N_4187,N_3752);
or U6937 (N_6937,N_3428,N_5242);
nor U6938 (N_6938,N_5230,N_3991);
nor U6939 (N_6939,N_4226,N_4609);
nor U6940 (N_6940,N_4032,N_3296);
nor U6941 (N_6941,N_4978,N_4483);
nand U6942 (N_6942,N_5381,N_5764);
or U6943 (N_6943,N_4468,N_5753);
or U6944 (N_6944,N_5940,N_4598);
or U6945 (N_6945,N_5829,N_5850);
nor U6946 (N_6946,N_4702,N_5519);
nor U6947 (N_6947,N_3175,N_5698);
and U6948 (N_6948,N_5844,N_5560);
or U6949 (N_6949,N_5051,N_3228);
nor U6950 (N_6950,N_3983,N_5467);
nor U6951 (N_6951,N_5249,N_3715);
and U6952 (N_6952,N_4654,N_3018);
nor U6953 (N_6953,N_5693,N_3486);
nand U6954 (N_6954,N_5445,N_5785);
or U6955 (N_6955,N_4889,N_5749);
nand U6956 (N_6956,N_4073,N_4976);
nor U6957 (N_6957,N_3176,N_3308);
nand U6958 (N_6958,N_5090,N_4958);
nand U6959 (N_6959,N_4146,N_4490);
nand U6960 (N_6960,N_4258,N_4787);
nor U6961 (N_6961,N_3137,N_3444);
or U6962 (N_6962,N_4632,N_5935);
or U6963 (N_6963,N_5486,N_5213);
or U6964 (N_6964,N_4045,N_5792);
nor U6965 (N_6965,N_5877,N_4371);
and U6966 (N_6966,N_3397,N_4734);
and U6967 (N_6967,N_5377,N_3459);
nand U6968 (N_6968,N_5015,N_5438);
and U6969 (N_6969,N_5283,N_3471);
nor U6970 (N_6970,N_3642,N_5209);
nand U6971 (N_6971,N_4754,N_3064);
nor U6972 (N_6972,N_5907,N_4776);
nor U6973 (N_6973,N_4821,N_3072);
or U6974 (N_6974,N_3172,N_3621);
nand U6975 (N_6975,N_4239,N_5061);
nand U6976 (N_6976,N_4647,N_5135);
nand U6977 (N_6977,N_3531,N_4359);
nor U6978 (N_6978,N_3525,N_4793);
nor U6979 (N_6979,N_5914,N_3334);
or U6980 (N_6980,N_5898,N_5397);
nor U6981 (N_6981,N_3148,N_4050);
and U6982 (N_6982,N_5766,N_4612);
nand U6983 (N_6983,N_3336,N_5967);
nor U6984 (N_6984,N_5425,N_4525);
and U6985 (N_6985,N_4918,N_3720);
nor U6986 (N_6986,N_5419,N_5562);
nor U6987 (N_6987,N_3949,N_4466);
nand U6988 (N_6988,N_4662,N_4722);
nor U6989 (N_6989,N_4872,N_5620);
nand U6990 (N_6990,N_3222,N_5366);
xor U6991 (N_6991,N_3271,N_4102);
or U6992 (N_6992,N_5163,N_3576);
and U6993 (N_6993,N_4944,N_3122);
nand U6994 (N_6994,N_5805,N_3200);
and U6995 (N_6995,N_4103,N_5731);
nor U6996 (N_6996,N_5299,N_3357);
and U6997 (N_6997,N_4757,N_4967);
or U6998 (N_6998,N_4496,N_4683);
nand U6999 (N_6999,N_3639,N_5500);
nand U7000 (N_7000,N_4075,N_3509);
or U7001 (N_7001,N_4432,N_4323);
and U7002 (N_7002,N_4378,N_4767);
or U7003 (N_7003,N_5553,N_5018);
nor U7004 (N_7004,N_5324,N_4655);
nor U7005 (N_7005,N_3911,N_5450);
nand U7006 (N_7006,N_5734,N_3431);
nor U7007 (N_7007,N_5814,N_5934);
nor U7008 (N_7008,N_5660,N_3785);
nand U7009 (N_7009,N_4476,N_3668);
or U7010 (N_7010,N_5189,N_3939);
nand U7011 (N_7011,N_3605,N_4866);
nor U7012 (N_7012,N_4819,N_4670);
xnor U7013 (N_7013,N_3536,N_5236);
or U7014 (N_7014,N_5586,N_4868);
or U7015 (N_7015,N_3343,N_5437);
nand U7016 (N_7016,N_4157,N_5888);
xor U7017 (N_7017,N_3190,N_3366);
or U7018 (N_7018,N_4504,N_3959);
nor U7019 (N_7019,N_3888,N_3652);
xor U7020 (N_7020,N_5861,N_4029);
or U7021 (N_7021,N_5636,N_3669);
or U7022 (N_7022,N_5109,N_4715);
and U7023 (N_7023,N_4321,N_3521);
nand U7024 (N_7024,N_5043,N_3327);
or U7025 (N_7025,N_3283,N_3218);
nor U7026 (N_7026,N_4842,N_5969);
and U7027 (N_7027,N_5796,N_3657);
and U7028 (N_7028,N_4999,N_5192);
or U7029 (N_7029,N_5245,N_5804);
and U7030 (N_7030,N_4405,N_3749);
or U7031 (N_7031,N_4870,N_4926);
nor U7032 (N_7032,N_5987,N_5909);
nand U7033 (N_7033,N_3117,N_4298);
and U7034 (N_7034,N_3924,N_3690);
and U7035 (N_7035,N_4192,N_4540);
and U7036 (N_7036,N_5849,N_3388);
nand U7037 (N_7037,N_3691,N_3437);
or U7038 (N_7038,N_5816,N_4274);
nand U7039 (N_7039,N_5306,N_3988);
or U7040 (N_7040,N_5789,N_5253);
or U7041 (N_7041,N_4343,N_3430);
nor U7042 (N_7042,N_4523,N_5369);
nor U7043 (N_7043,N_3561,N_3529);
nand U7044 (N_7044,N_3147,N_4169);
nor U7045 (N_7045,N_5101,N_4777);
or U7046 (N_7046,N_3024,N_5773);
nand U7047 (N_7047,N_5685,N_5516);
or U7048 (N_7048,N_4924,N_3084);
nand U7049 (N_7049,N_5494,N_3249);
or U7050 (N_7050,N_4730,N_3083);
or U7051 (N_7051,N_5807,N_5376);
nor U7052 (N_7052,N_4886,N_4989);
nor U7053 (N_7053,N_5802,N_3724);
and U7054 (N_7054,N_5918,N_4142);
and U7055 (N_7055,N_4347,N_4500);
and U7056 (N_7056,N_3399,N_4345);
and U7057 (N_7057,N_5456,N_5820);
nand U7058 (N_7058,N_5768,N_4335);
nor U7059 (N_7059,N_5062,N_3410);
or U7060 (N_7060,N_5881,N_4871);
or U7061 (N_7061,N_4567,N_5964);
nor U7062 (N_7062,N_4038,N_3928);
nand U7063 (N_7063,N_3760,N_5472);
or U7064 (N_7064,N_3102,N_5558);
nor U7065 (N_7065,N_4404,N_4195);
nand U7066 (N_7066,N_3517,N_4081);
or U7067 (N_7067,N_5665,N_4076);
and U7068 (N_7068,N_5347,N_4668);
and U7069 (N_7069,N_3155,N_4283);
and U7070 (N_7070,N_5812,N_5304);
nor U7071 (N_7071,N_4794,N_3732);
nand U7072 (N_7072,N_5260,N_3009);
nor U7073 (N_7073,N_5985,N_3875);
nand U7074 (N_7074,N_3823,N_4721);
or U7075 (N_7075,N_4520,N_4008);
nor U7076 (N_7076,N_5771,N_5172);
or U7077 (N_7077,N_5228,N_5458);
nand U7078 (N_7078,N_5317,N_4716);
nor U7079 (N_7079,N_3809,N_4700);
nand U7080 (N_7080,N_5212,N_3686);
and U7081 (N_7081,N_4253,N_5431);
and U7082 (N_7082,N_5174,N_3595);
and U7083 (N_7083,N_5284,N_3503);
and U7084 (N_7084,N_5117,N_3811);
and U7085 (N_7085,N_3846,N_4528);
nand U7086 (N_7086,N_5513,N_4549);
nor U7087 (N_7087,N_3552,N_5572);
or U7088 (N_7088,N_5221,N_3498);
nand U7089 (N_7089,N_4368,N_5707);
nand U7090 (N_7090,N_5502,N_3537);
nand U7091 (N_7091,N_5530,N_3457);
nor U7092 (N_7092,N_5182,N_3920);
or U7093 (N_7093,N_5158,N_5276);
nor U7094 (N_7094,N_5481,N_4642);
nor U7095 (N_7095,N_4465,N_4758);
nor U7096 (N_7096,N_3379,N_4191);
nor U7097 (N_7097,N_4659,N_3286);
or U7098 (N_7098,N_4719,N_5217);
nor U7099 (N_7099,N_3081,N_3907);
nor U7100 (N_7100,N_5246,N_4535);
nor U7101 (N_7101,N_5605,N_4446);
or U7102 (N_7102,N_3100,N_5131);
and U7103 (N_7103,N_5025,N_4242);
and U7104 (N_7104,N_4364,N_4858);
nor U7105 (N_7105,N_5887,N_5547);
or U7106 (N_7106,N_5681,N_5320);
nand U7107 (N_7107,N_5842,N_5976);
or U7108 (N_7108,N_3027,N_3241);
and U7109 (N_7109,N_3476,N_3882);
nand U7110 (N_7110,N_4740,N_3272);
nor U7111 (N_7111,N_5795,N_4970);
nand U7112 (N_7112,N_4113,N_5906);
nand U7113 (N_7113,N_3133,N_5606);
or U7114 (N_7114,N_4452,N_4387);
nand U7115 (N_7115,N_5780,N_3128);
and U7116 (N_7116,N_5161,N_4290);
nand U7117 (N_7117,N_5430,N_5970);
nand U7118 (N_7118,N_4267,N_4888);
nand U7119 (N_7119,N_5475,N_5968);
or U7120 (N_7120,N_5060,N_5727);
or U7121 (N_7121,N_5846,N_3700);
nand U7122 (N_7122,N_5322,N_5941);
and U7123 (N_7123,N_5087,N_3746);
nand U7124 (N_7124,N_4119,N_3236);
nand U7125 (N_7125,N_4790,N_3404);
and U7126 (N_7126,N_5340,N_3844);
or U7127 (N_7127,N_3539,N_5538);
nand U7128 (N_7128,N_3923,N_3921);
nand U7129 (N_7129,N_4818,N_3891);
nor U7130 (N_7130,N_5894,N_3063);
and U7131 (N_7131,N_5009,N_5897);
and U7132 (N_7132,N_4582,N_3373);
or U7133 (N_7133,N_5219,N_3049);
or U7134 (N_7134,N_5068,N_5492);
nor U7135 (N_7135,N_4150,N_5721);
and U7136 (N_7136,N_3977,N_5503);
and U7137 (N_7137,N_5511,N_4919);
nor U7138 (N_7138,N_3654,N_4751);
or U7139 (N_7139,N_3513,N_5337);
or U7140 (N_7140,N_5565,N_4765);
nand U7141 (N_7141,N_4677,N_5756);
nor U7142 (N_7142,N_3164,N_4907);
or U7143 (N_7143,N_3193,N_4464);
and U7144 (N_7144,N_5591,N_4161);
nand U7145 (N_7145,N_3495,N_3192);
nor U7146 (N_7146,N_3225,N_5145);
and U7147 (N_7147,N_5339,N_3417);
nor U7148 (N_7148,N_3565,N_3114);
nand U7149 (N_7149,N_4606,N_3770);
and U7150 (N_7150,N_5434,N_5265);
nand U7151 (N_7151,N_4929,N_3267);
and U7152 (N_7152,N_4125,N_5243);
and U7153 (N_7153,N_5960,N_5946);
nor U7154 (N_7154,N_3451,N_5224);
and U7155 (N_7155,N_3551,N_3180);
and U7156 (N_7156,N_4691,N_3215);
and U7157 (N_7157,N_4851,N_5130);
and U7158 (N_7158,N_3187,N_3670);
or U7159 (N_7159,N_3692,N_5391);
and U7160 (N_7160,N_4011,N_3253);
or U7161 (N_7161,N_3104,N_4798);
or U7162 (N_7162,N_4127,N_5912);
nand U7163 (N_7163,N_4082,N_3461);
nand U7164 (N_7164,N_4215,N_5509);
and U7165 (N_7165,N_4998,N_4935);
nor U7166 (N_7166,N_5778,N_3227);
or U7167 (N_7167,N_4869,N_5423);
or U7168 (N_7168,N_3346,N_3990);
or U7169 (N_7169,N_4517,N_3422);
nand U7170 (N_7170,N_3996,N_4836);
or U7171 (N_7171,N_4417,N_4753);
nor U7172 (N_7172,N_3756,N_4344);
nand U7173 (N_7173,N_5027,N_3000);
or U7174 (N_7174,N_3059,N_3087);
and U7175 (N_7175,N_3452,N_4830);
or U7176 (N_7176,N_3798,N_4418);
nand U7177 (N_7177,N_4201,N_3363);
nand U7178 (N_7178,N_4698,N_5507);
or U7179 (N_7179,N_5371,N_5483);
nor U7180 (N_7180,N_4553,N_4996);
nor U7181 (N_7181,N_4701,N_3269);
or U7182 (N_7182,N_4291,N_3683);
nor U7183 (N_7183,N_5982,N_4607);
or U7184 (N_7184,N_5305,N_5480);
nor U7185 (N_7185,N_3919,N_3041);
nand U7186 (N_7186,N_3851,N_4152);
or U7187 (N_7187,N_4194,N_3717);
or U7188 (N_7188,N_5070,N_4947);
or U7189 (N_7189,N_3328,N_4593);
or U7190 (N_7190,N_5296,N_4223);
and U7191 (N_7191,N_4176,N_4862);
nand U7192 (N_7192,N_5110,N_5454);
or U7193 (N_7193,N_3975,N_3372);
nand U7194 (N_7194,N_5604,N_5902);
nand U7195 (N_7195,N_3848,N_4070);
and U7196 (N_7196,N_3857,N_5006);
and U7197 (N_7197,N_3258,N_4224);
or U7198 (N_7198,N_4250,N_5225);
nand U7199 (N_7199,N_4453,N_5275);
or U7200 (N_7200,N_3254,N_5157);
nand U7201 (N_7201,N_4093,N_4938);
nand U7202 (N_7202,N_4746,N_4377);
nor U7203 (N_7203,N_5208,N_4898);
and U7204 (N_7204,N_4543,N_5917);
nand U7205 (N_7205,N_5616,N_5248);
nand U7206 (N_7206,N_5126,N_4002);
and U7207 (N_7207,N_3170,N_3985);
nand U7208 (N_7208,N_4695,N_5066);
and U7209 (N_7209,N_3564,N_5173);
and U7210 (N_7210,N_5215,N_4760);
or U7211 (N_7211,N_3879,N_3524);
or U7212 (N_7212,N_3821,N_4319);
nor U7213 (N_7213,N_5138,N_3185);
nor U7214 (N_7214,N_3156,N_3432);
and U7215 (N_7215,N_5171,N_5270);
nor U7216 (N_7216,N_5823,N_4004);
and U7217 (N_7217,N_4890,N_5113);
and U7218 (N_7218,N_4439,N_4023);
nand U7219 (N_7219,N_5552,N_5362);
nor U7220 (N_7220,N_5139,N_4820);
nor U7221 (N_7221,N_5577,N_4144);
nand U7222 (N_7222,N_5020,N_3623);
or U7223 (N_7223,N_5452,N_4562);
nand U7224 (N_7224,N_5008,N_5357);
nand U7225 (N_7225,N_5313,N_5979);
nand U7226 (N_7226,N_3931,N_4077);
nand U7227 (N_7227,N_5164,N_3816);
and U7228 (N_7228,N_3487,N_4143);
and U7229 (N_7229,N_5788,N_3376);
xnor U7230 (N_7230,N_4131,N_3103);
or U7231 (N_7231,N_5561,N_3776);
and U7232 (N_7232,N_5597,N_3012);
or U7233 (N_7233,N_5211,N_3168);
or U7234 (N_7234,N_5021,N_3359);
and U7235 (N_7235,N_5623,N_4406);
nand U7236 (N_7236,N_5990,N_5755);
and U7237 (N_7237,N_5711,N_3435);
or U7238 (N_7238,N_4641,N_4326);
nand U7239 (N_7239,N_4060,N_3418);
and U7240 (N_7240,N_4494,N_5142);
or U7241 (N_7241,N_4838,N_3445);
nor U7242 (N_7242,N_5039,N_5630);
nor U7243 (N_7243,N_4262,N_3563);
nor U7244 (N_7244,N_4679,N_3824);
or U7245 (N_7245,N_4676,N_3708);
nor U7246 (N_7246,N_5584,N_5349);
nor U7247 (N_7247,N_5581,N_3615);
and U7248 (N_7248,N_4160,N_5641);
or U7249 (N_7249,N_4118,N_4227);
nor U7250 (N_7250,N_5690,N_4477);
and U7251 (N_7251,N_3656,N_5743);
or U7252 (N_7252,N_3904,N_5345);
and U7253 (N_7253,N_5873,N_3291);
or U7254 (N_7254,N_4764,N_5334);
and U7255 (N_7255,N_5491,N_4481);
nor U7256 (N_7256,N_3381,N_4254);
nor U7257 (N_7257,N_3948,N_4542);
nand U7258 (N_7258,N_5725,N_5555);
nand U7259 (N_7259,N_5374,N_3818);
nand U7260 (N_7260,N_4903,N_5811);
nor U7261 (N_7261,N_4620,N_4370);
and U7262 (N_7262,N_4409,N_3607);
nand U7263 (N_7263,N_3860,N_3935);
or U7264 (N_7264,N_4531,N_5360);
nand U7265 (N_7265,N_5361,N_4039);
and U7266 (N_7266,N_5014,N_5343);
and U7267 (N_7267,N_5526,N_5257);
nor U7268 (N_7268,N_3160,N_4334);
and U7269 (N_7269,N_4206,N_5772);
nor U7270 (N_7270,N_4883,N_5298);
and U7271 (N_7271,N_4330,N_3183);
and U7272 (N_7272,N_4628,N_3757);
and U7273 (N_7273,N_4987,N_3787);
and U7274 (N_7274,N_3980,N_3101);
nand U7275 (N_7275,N_5923,N_5742);
nand U7276 (N_7276,N_4480,N_4847);
or U7277 (N_7277,N_3289,N_3348);
and U7278 (N_7278,N_3270,N_4249);
and U7279 (N_7279,N_3246,N_5264);
and U7280 (N_7280,N_4233,N_4459);
or U7281 (N_7281,N_5044,N_5837);
and U7282 (N_7282,N_3841,N_5574);
or U7283 (N_7283,N_4678,N_3071);
and U7284 (N_7284,N_4428,N_4325);
or U7285 (N_7285,N_3631,N_5151);
nor U7286 (N_7286,N_4554,N_4121);
nor U7287 (N_7287,N_5835,N_4955);
nor U7288 (N_7288,N_3880,N_3896);
nor U7289 (N_7289,N_5671,N_4426);
nand U7290 (N_7290,N_4731,N_4296);
or U7291 (N_7291,N_3820,N_5868);
nand U7292 (N_7292,N_5673,N_5387);
or U7293 (N_7293,N_3458,N_4849);
and U7294 (N_7294,N_5879,N_3033);
nand U7295 (N_7295,N_3523,N_5801);
or U7296 (N_7296,N_4184,N_5751);
nor U7297 (N_7297,N_3554,N_3750);
nor U7298 (N_7298,N_3965,N_5272);
nor U7299 (N_7299,N_5508,N_4712);
nor U7300 (N_7300,N_3876,N_5748);
nor U7301 (N_7301,N_4707,N_3863);
and U7302 (N_7302,N_5601,N_5218);
nor U7303 (N_7303,N_3293,N_3317);
nand U7304 (N_7304,N_4509,N_4933);
nor U7305 (N_7305,N_3661,N_3040);
nand U7306 (N_7306,N_5191,N_5977);
nand U7307 (N_7307,N_4462,N_5686);
and U7308 (N_7308,N_3132,N_3528);
nor U7309 (N_7309,N_4810,N_5177);
nor U7310 (N_7310,N_5904,N_3519);
nand U7311 (N_7311,N_3202,N_5838);
nand U7312 (N_7312,N_4069,N_5924);
or U7313 (N_7313,N_5160,N_3307);
nand U7314 (N_7314,N_3916,N_3976);
or U7315 (N_7315,N_4027,N_5029);
or U7316 (N_7316,N_5167,N_5598);
and U7317 (N_7317,N_5845,N_4916);
nand U7318 (N_7318,N_5198,N_3705);
nor U7319 (N_7319,N_5088,N_4833);
nor U7320 (N_7320,N_5442,N_3622);
nor U7321 (N_7321,N_4865,N_4324);
or U7322 (N_7322,N_4026,N_3624);
or U7323 (N_7323,N_5662,N_4305);
nand U7324 (N_7324,N_5121,N_5889);
nand U7325 (N_7325,N_4373,N_4846);
nor U7326 (N_7326,N_5365,N_3212);
or U7327 (N_7327,N_3198,N_5292);
or U7328 (N_7328,N_5201,N_4154);
and U7329 (N_7329,N_4181,N_4219);
and U7330 (N_7330,N_5994,N_3918);
nand U7331 (N_7331,N_4299,N_5084);
nor U7332 (N_7332,N_5943,N_4825);
nand U7333 (N_7333,N_4057,N_3762);
nand U7334 (N_7334,N_4622,N_4657);
nand U7335 (N_7335,N_3195,N_3014);
and U7336 (N_7336,N_3571,N_5972);
nor U7337 (N_7337,N_4217,N_3678);
and U7338 (N_7338,N_3550,N_4264);
or U7339 (N_7339,N_5922,N_5652);
nor U7340 (N_7340,N_3337,N_5428);
and U7341 (N_7341,N_5830,N_3069);
or U7342 (N_7342,N_4991,N_4586);
nor U7343 (N_7343,N_3545,N_4822);
nor U7344 (N_7344,N_4241,N_3369);
nor U7345 (N_7345,N_5651,N_3470);
and U7346 (N_7346,N_5446,N_4300);
and U7347 (N_7347,N_3284,N_3499);
or U7348 (N_7348,N_5353,N_3780);
or U7349 (N_7349,N_4065,N_4547);
xor U7350 (N_7350,N_4246,N_5416);
nand U7351 (N_7351,N_3950,N_3599);
nand U7352 (N_7352,N_4638,N_4530);
or U7353 (N_7353,N_3450,N_5957);
nor U7354 (N_7354,N_4840,N_4164);
or U7355 (N_7355,N_5892,N_5329);
nor U7356 (N_7356,N_3443,N_3353);
nand U7357 (N_7357,N_4861,N_5403);
or U7358 (N_7358,N_4059,N_4658);
nand U7359 (N_7359,N_5382,N_4834);
nand U7360 (N_7360,N_5447,N_4807);
and U7361 (N_7361,N_5744,N_4014);
nand U7362 (N_7362,N_4817,N_4786);
and U7363 (N_7363,N_5856,N_3682);
or U7364 (N_7364,N_3802,N_5945);
nor U7365 (N_7365,N_3666,N_5659);
nor U7366 (N_7366,N_4307,N_5543);
nand U7367 (N_7367,N_4384,N_3449);
or U7368 (N_7368,N_4891,N_5093);
or U7369 (N_7369,N_4265,N_5745);
or U7370 (N_7370,N_4471,N_3329);
nor U7371 (N_7371,N_4401,N_3145);
nand U7372 (N_7372,N_3174,N_5590);
and U7373 (N_7373,N_5005,N_5704);
or U7374 (N_7374,N_4595,N_3706);
nand U7375 (N_7375,N_5195,N_5072);
and U7376 (N_7376,N_4618,N_4136);
nand U7377 (N_7377,N_3494,N_4619);
nand U7378 (N_7378,N_4392,N_4340);
nand U7379 (N_7379,N_5216,N_3856);
or U7380 (N_7380,N_3342,N_5915);
or U7381 (N_7381,N_5436,N_4896);
nand U7382 (N_7382,N_4912,N_5420);
nand U7383 (N_7383,N_3201,N_4388);
and U7384 (N_7384,N_5156,N_4351);
or U7385 (N_7385,N_5995,N_3060);
and U7386 (N_7386,N_4974,N_3259);
nand U7387 (N_7387,N_3302,N_5461);
nand U7388 (N_7388,N_4474,N_3718);
or U7389 (N_7389,N_3582,N_4993);
nor U7390 (N_7390,N_5556,N_5071);
nor U7391 (N_7391,N_3491,N_3389);
nor U7392 (N_7392,N_5333,N_4457);
and U7393 (N_7393,N_3766,N_4137);
or U7394 (N_7394,N_4451,N_4518);
or U7395 (N_7395,N_5517,N_4037);
nand U7396 (N_7396,N_3817,N_5393);
or U7397 (N_7397,N_3553,N_3723);
xnor U7398 (N_7398,N_4687,N_4199);
and U7399 (N_7399,N_3799,N_4915);
nor U7400 (N_7400,N_3606,N_5186);
nor U7401 (N_7401,N_4151,N_5722);
nor U7402 (N_7402,N_5469,N_5625);
and U7403 (N_7403,N_3442,N_5947);
nor U7404 (N_7404,N_5202,N_5410);
or U7405 (N_7405,N_4717,N_5803);
nor U7406 (N_7406,N_5848,N_3483);
or U7407 (N_7407,N_5141,N_5506);
nor U7408 (N_7408,N_4527,N_4963);
or U7409 (N_7409,N_4155,N_5891);
and U7410 (N_7410,N_5619,N_5203);
xnor U7411 (N_7411,N_3086,N_3055);
nor U7412 (N_7412,N_4414,N_5207);
or U7413 (N_7413,N_3386,N_5799);
or U7414 (N_7414,N_3998,N_3889);
and U7415 (N_7415,N_4614,N_4964);
or U7416 (N_7416,N_5479,N_5962);
xnor U7417 (N_7417,N_4837,N_5128);
or U7418 (N_7418,N_5515,N_3812);
or U7419 (N_7419,N_3046,N_3411);
and U7420 (N_7420,N_4499,N_4469);
nor U7421 (N_7421,N_3462,N_4892);
nor U7422 (N_7422,N_5023,N_4656);
or U7423 (N_7423,N_3043,N_4795);
nand U7424 (N_7424,N_5273,N_3887);
nand U7425 (N_7425,N_3109,N_3716);
or U7426 (N_7426,N_4046,N_4850);
nor U7427 (N_7427,N_4621,N_4775);
and U7428 (N_7428,N_4178,N_4762);
or U7429 (N_7429,N_3477,N_4546);
nand U7430 (N_7430,N_5997,N_4665);
or U7431 (N_7431,N_3076,N_4297);
nand U7432 (N_7432,N_5710,N_3538);
or U7433 (N_7433,N_4867,N_4827);
nor U7434 (N_7434,N_3472,N_3279);
and U7435 (N_7435,N_4006,N_4410);
nor U7436 (N_7436,N_4852,N_3745);
and U7437 (N_7437,N_5661,N_3421);
nor U7438 (N_7438,N_4331,N_5086);
or U7439 (N_7439,N_4108,N_4743);
and U7440 (N_7440,N_5455,N_3021);
and U7441 (N_7441,N_4255,N_3679);
nand U7442 (N_7442,N_3936,N_5931);
or U7443 (N_7443,N_3952,N_3255);
and U7444 (N_7444,N_4769,N_3917);
or U7445 (N_7445,N_5545,N_3276);
or U7446 (N_7446,N_3781,N_4438);
nor U7447 (N_7447,N_3243,N_3759);
nand U7448 (N_7448,N_3224,N_4179);
xor U7449 (N_7449,N_3640,N_3467);
or U7450 (N_7450,N_4200,N_3429);
nor U7451 (N_7451,N_4398,N_4581);
nor U7452 (N_7452,N_5111,N_3096);
and U7453 (N_7453,N_5576,N_3447);
nand U7454 (N_7454,N_5549,N_4627);
nand U7455 (N_7455,N_3473,N_3144);
and U7456 (N_7456,N_4789,N_5356);
or U7457 (N_7457,N_3839,N_3815);
and U7458 (N_7458,N_5672,N_4444);
or U7459 (N_7459,N_5457,N_4971);
nand U7460 (N_7460,N_5790,N_5741);
nand U7461 (N_7461,N_3842,N_4024);
nand U7462 (N_7462,N_3970,N_3497);
nand U7463 (N_7463,N_5400,N_5287);
nand U7464 (N_7464,N_4956,N_4379);
nand U7465 (N_7465,N_5750,N_5412);
nor U7466 (N_7466,N_3653,N_4435);
or U7467 (N_7467,N_5633,N_5321);
nor U7468 (N_7468,N_4177,N_4829);
nor U7469 (N_7469,N_3019,N_5441);
and U7470 (N_7470,N_3765,N_3791);
and U7471 (N_7471,N_3028,N_4189);
nor U7472 (N_7472,N_5937,N_5953);
or U7473 (N_7473,N_4198,N_3659);
and U7474 (N_7474,N_3298,N_5300);
nand U7475 (N_7475,N_3268,N_5600);
or U7476 (N_7476,N_5240,N_3036);
or U7477 (N_7477,N_3067,N_3237);
nor U7478 (N_7478,N_5974,N_4878);
or U7479 (N_7479,N_4783,N_3767);
or U7480 (N_7480,N_3250,N_3157);
and U7481 (N_7481,N_5233,N_3354);
nand U7482 (N_7482,N_4512,N_5825);
and U7483 (N_7483,N_3260,N_3560);
and U7484 (N_7484,N_5258,N_3589);
nor U7485 (N_7485,N_5824,N_5030);
or U7486 (N_7486,N_5644,N_3031);
nor U7487 (N_7487,N_4755,N_3108);
and U7488 (N_7488,N_4917,N_3416);
and U7489 (N_7489,N_4259,N_5118);
or U7490 (N_7490,N_4382,N_4855);
and U7491 (N_7491,N_4310,N_5082);
and U7492 (N_7492,N_5980,N_4097);
and U7493 (N_7493,N_5190,N_5610);
nor U7494 (N_7494,N_4022,N_3944);
or U7495 (N_7495,N_4313,N_3001);
nand U7496 (N_7496,N_3741,N_3932);
xor U7497 (N_7497,N_4040,N_5583);
nand U7498 (N_7498,N_4366,N_5893);
or U7499 (N_7499,N_5536,N_5981);
and U7500 (N_7500,N_4156,N_5064);
and U7501 (N_7501,N_5983,N_4332);
xor U7502 (N_7502,N_4416,N_3852);
xor U7503 (N_7503,N_3229,N_4571);
nor U7504 (N_7504,N_5130,N_4955);
nor U7505 (N_7505,N_3890,N_5389);
and U7506 (N_7506,N_4053,N_4583);
nor U7507 (N_7507,N_5719,N_3443);
nor U7508 (N_7508,N_3913,N_4349);
and U7509 (N_7509,N_3318,N_4364);
nand U7510 (N_7510,N_5091,N_5988);
and U7511 (N_7511,N_5634,N_5108);
and U7512 (N_7512,N_5206,N_4431);
and U7513 (N_7513,N_5743,N_3783);
and U7514 (N_7514,N_3156,N_4643);
and U7515 (N_7515,N_5138,N_5211);
and U7516 (N_7516,N_4659,N_5988);
nand U7517 (N_7517,N_3571,N_3159);
and U7518 (N_7518,N_4994,N_5280);
nor U7519 (N_7519,N_5373,N_5181);
nor U7520 (N_7520,N_5360,N_4393);
and U7521 (N_7521,N_5149,N_5658);
and U7522 (N_7522,N_5214,N_4551);
nand U7523 (N_7523,N_3378,N_4163);
and U7524 (N_7524,N_5635,N_4198);
nor U7525 (N_7525,N_5664,N_5899);
or U7526 (N_7526,N_3506,N_5556);
and U7527 (N_7527,N_3758,N_4299);
and U7528 (N_7528,N_5374,N_5011);
nand U7529 (N_7529,N_3925,N_3757);
nor U7530 (N_7530,N_4999,N_5884);
and U7531 (N_7531,N_4606,N_5120);
or U7532 (N_7532,N_5964,N_5241);
or U7533 (N_7533,N_5685,N_4652);
nor U7534 (N_7534,N_4924,N_4700);
nor U7535 (N_7535,N_4156,N_4762);
or U7536 (N_7536,N_3224,N_5035);
nand U7537 (N_7537,N_5792,N_4888);
or U7538 (N_7538,N_4431,N_3287);
and U7539 (N_7539,N_5778,N_3061);
and U7540 (N_7540,N_4094,N_4001);
nor U7541 (N_7541,N_5121,N_3266);
or U7542 (N_7542,N_3244,N_3889);
nor U7543 (N_7543,N_4992,N_3319);
or U7544 (N_7544,N_3061,N_4074);
and U7545 (N_7545,N_5251,N_3446);
nand U7546 (N_7546,N_3770,N_5077);
nand U7547 (N_7547,N_3727,N_3962);
or U7548 (N_7548,N_4523,N_5985);
nor U7549 (N_7549,N_4828,N_3929);
and U7550 (N_7550,N_3101,N_4034);
nor U7551 (N_7551,N_3381,N_4119);
or U7552 (N_7552,N_3056,N_4985);
nor U7553 (N_7553,N_3592,N_5171);
nor U7554 (N_7554,N_3639,N_3331);
nand U7555 (N_7555,N_3074,N_3219);
and U7556 (N_7556,N_5285,N_5715);
nand U7557 (N_7557,N_5495,N_4481);
nand U7558 (N_7558,N_3498,N_4328);
nor U7559 (N_7559,N_4917,N_5914);
nand U7560 (N_7560,N_3134,N_5215);
xor U7561 (N_7561,N_4915,N_4749);
and U7562 (N_7562,N_4611,N_3725);
nor U7563 (N_7563,N_5561,N_3445);
and U7564 (N_7564,N_5926,N_4880);
nand U7565 (N_7565,N_4816,N_4622);
nand U7566 (N_7566,N_3946,N_3960);
nand U7567 (N_7567,N_3889,N_4295);
and U7568 (N_7568,N_3984,N_5460);
or U7569 (N_7569,N_5417,N_3691);
or U7570 (N_7570,N_3610,N_3786);
nor U7571 (N_7571,N_4680,N_5315);
nand U7572 (N_7572,N_5068,N_3278);
nor U7573 (N_7573,N_4845,N_5496);
nand U7574 (N_7574,N_3733,N_4810);
and U7575 (N_7575,N_5441,N_5311);
nor U7576 (N_7576,N_5157,N_5382);
nand U7577 (N_7577,N_4613,N_5098);
nor U7578 (N_7578,N_4902,N_5616);
nor U7579 (N_7579,N_4657,N_4940);
or U7580 (N_7580,N_4098,N_3469);
and U7581 (N_7581,N_5848,N_4368);
nor U7582 (N_7582,N_5016,N_3292);
nor U7583 (N_7583,N_3631,N_4672);
or U7584 (N_7584,N_5187,N_3885);
nand U7585 (N_7585,N_4404,N_5924);
and U7586 (N_7586,N_4285,N_4168);
xor U7587 (N_7587,N_5966,N_5126);
nor U7588 (N_7588,N_3855,N_3521);
xnor U7589 (N_7589,N_4165,N_5649);
nand U7590 (N_7590,N_3435,N_4285);
nand U7591 (N_7591,N_3557,N_4622);
nor U7592 (N_7592,N_4890,N_4846);
nand U7593 (N_7593,N_4293,N_4970);
nor U7594 (N_7594,N_5746,N_3912);
or U7595 (N_7595,N_5186,N_4890);
nand U7596 (N_7596,N_4772,N_5288);
nor U7597 (N_7597,N_3765,N_4580);
nor U7598 (N_7598,N_5844,N_3612);
and U7599 (N_7599,N_4029,N_5178);
nor U7600 (N_7600,N_4655,N_4265);
nand U7601 (N_7601,N_4945,N_3489);
nand U7602 (N_7602,N_4008,N_3906);
nor U7603 (N_7603,N_3113,N_4643);
nand U7604 (N_7604,N_5834,N_3580);
nand U7605 (N_7605,N_5325,N_5473);
and U7606 (N_7606,N_5184,N_5519);
and U7607 (N_7607,N_3014,N_5397);
and U7608 (N_7608,N_4062,N_4076);
and U7609 (N_7609,N_5075,N_4021);
and U7610 (N_7610,N_4845,N_5008);
nor U7611 (N_7611,N_3016,N_3216);
and U7612 (N_7612,N_4349,N_4195);
or U7613 (N_7613,N_3296,N_4130);
and U7614 (N_7614,N_5687,N_5391);
or U7615 (N_7615,N_4761,N_4517);
or U7616 (N_7616,N_4684,N_4112);
nor U7617 (N_7617,N_5275,N_3079);
and U7618 (N_7618,N_5885,N_3926);
and U7619 (N_7619,N_4601,N_4390);
nor U7620 (N_7620,N_5896,N_5902);
and U7621 (N_7621,N_5119,N_5569);
or U7622 (N_7622,N_5610,N_4022);
or U7623 (N_7623,N_4256,N_4371);
nor U7624 (N_7624,N_4714,N_3081);
or U7625 (N_7625,N_5441,N_3814);
and U7626 (N_7626,N_4967,N_3396);
nand U7627 (N_7627,N_3338,N_5478);
nor U7628 (N_7628,N_5704,N_4615);
and U7629 (N_7629,N_3941,N_4023);
nor U7630 (N_7630,N_3187,N_3308);
or U7631 (N_7631,N_5202,N_5023);
or U7632 (N_7632,N_3214,N_3636);
nand U7633 (N_7633,N_3239,N_4699);
and U7634 (N_7634,N_5648,N_3448);
nor U7635 (N_7635,N_3761,N_4555);
or U7636 (N_7636,N_3857,N_4368);
or U7637 (N_7637,N_4334,N_5088);
nand U7638 (N_7638,N_5015,N_3661);
or U7639 (N_7639,N_5620,N_3060);
and U7640 (N_7640,N_3562,N_5227);
nor U7641 (N_7641,N_5430,N_3995);
nor U7642 (N_7642,N_3263,N_4522);
nor U7643 (N_7643,N_4650,N_3377);
nor U7644 (N_7644,N_3799,N_5857);
and U7645 (N_7645,N_4291,N_4899);
and U7646 (N_7646,N_4907,N_3640);
or U7647 (N_7647,N_3224,N_5465);
nand U7648 (N_7648,N_5459,N_4841);
or U7649 (N_7649,N_5908,N_4077);
and U7650 (N_7650,N_4488,N_3057);
or U7651 (N_7651,N_3565,N_4303);
nand U7652 (N_7652,N_5516,N_4675);
nor U7653 (N_7653,N_3277,N_5203);
and U7654 (N_7654,N_5568,N_4626);
and U7655 (N_7655,N_4134,N_4155);
or U7656 (N_7656,N_3035,N_3619);
nor U7657 (N_7657,N_3854,N_4545);
nand U7658 (N_7658,N_5863,N_5159);
and U7659 (N_7659,N_5858,N_4567);
nor U7660 (N_7660,N_3920,N_3674);
or U7661 (N_7661,N_3988,N_3848);
or U7662 (N_7662,N_4837,N_3842);
and U7663 (N_7663,N_3625,N_5102);
and U7664 (N_7664,N_5857,N_3791);
nand U7665 (N_7665,N_3045,N_3700);
or U7666 (N_7666,N_4185,N_5415);
nor U7667 (N_7667,N_5896,N_5729);
nor U7668 (N_7668,N_4101,N_4264);
and U7669 (N_7669,N_5422,N_3751);
and U7670 (N_7670,N_4374,N_3577);
nand U7671 (N_7671,N_4839,N_4354);
and U7672 (N_7672,N_4980,N_3695);
and U7673 (N_7673,N_3028,N_5158);
and U7674 (N_7674,N_4754,N_4110);
nand U7675 (N_7675,N_4498,N_3731);
nand U7676 (N_7676,N_3776,N_3447);
or U7677 (N_7677,N_4971,N_5000);
nor U7678 (N_7678,N_5798,N_3917);
nor U7679 (N_7679,N_5754,N_3323);
or U7680 (N_7680,N_5836,N_3755);
and U7681 (N_7681,N_3305,N_3810);
and U7682 (N_7682,N_4326,N_4983);
nand U7683 (N_7683,N_5507,N_5491);
nor U7684 (N_7684,N_3358,N_4749);
nor U7685 (N_7685,N_3154,N_3284);
and U7686 (N_7686,N_4817,N_3195);
nor U7687 (N_7687,N_5199,N_5473);
xor U7688 (N_7688,N_4659,N_4807);
nand U7689 (N_7689,N_5518,N_4224);
nor U7690 (N_7690,N_5829,N_3604);
nor U7691 (N_7691,N_4271,N_3851);
nand U7692 (N_7692,N_4894,N_4774);
nand U7693 (N_7693,N_5566,N_5596);
nor U7694 (N_7694,N_3591,N_5081);
xnor U7695 (N_7695,N_5085,N_4817);
or U7696 (N_7696,N_3188,N_3693);
nor U7697 (N_7697,N_4776,N_3770);
or U7698 (N_7698,N_4572,N_5912);
nand U7699 (N_7699,N_4000,N_5733);
or U7700 (N_7700,N_5992,N_5817);
nand U7701 (N_7701,N_4565,N_5679);
nand U7702 (N_7702,N_3569,N_3239);
nor U7703 (N_7703,N_4652,N_4636);
nor U7704 (N_7704,N_5757,N_4556);
and U7705 (N_7705,N_3219,N_4922);
nand U7706 (N_7706,N_5015,N_5743);
nor U7707 (N_7707,N_4027,N_3711);
nand U7708 (N_7708,N_3671,N_5284);
and U7709 (N_7709,N_4245,N_4231);
or U7710 (N_7710,N_3704,N_4422);
nor U7711 (N_7711,N_3518,N_5108);
and U7712 (N_7712,N_3225,N_4271);
or U7713 (N_7713,N_4040,N_5257);
or U7714 (N_7714,N_5308,N_3084);
nand U7715 (N_7715,N_5490,N_4668);
or U7716 (N_7716,N_3617,N_4892);
nor U7717 (N_7717,N_3725,N_4792);
nor U7718 (N_7718,N_5972,N_4103);
nand U7719 (N_7719,N_5497,N_3200);
nor U7720 (N_7720,N_3036,N_3999);
nand U7721 (N_7721,N_4084,N_5541);
nor U7722 (N_7722,N_5785,N_3339);
nand U7723 (N_7723,N_4317,N_4899);
nor U7724 (N_7724,N_3740,N_4873);
nor U7725 (N_7725,N_3401,N_3120);
nand U7726 (N_7726,N_4808,N_3239);
or U7727 (N_7727,N_4997,N_4701);
or U7728 (N_7728,N_4139,N_4181);
or U7729 (N_7729,N_5269,N_4420);
nand U7730 (N_7730,N_4728,N_4927);
or U7731 (N_7731,N_3894,N_5266);
nor U7732 (N_7732,N_4916,N_3885);
or U7733 (N_7733,N_5527,N_4570);
nor U7734 (N_7734,N_5252,N_3210);
or U7735 (N_7735,N_3998,N_3969);
xnor U7736 (N_7736,N_5821,N_5000);
and U7737 (N_7737,N_4651,N_5945);
nor U7738 (N_7738,N_3410,N_5689);
or U7739 (N_7739,N_5812,N_3694);
or U7740 (N_7740,N_4763,N_5331);
or U7741 (N_7741,N_5003,N_5991);
nand U7742 (N_7742,N_3208,N_5295);
nand U7743 (N_7743,N_4287,N_3717);
and U7744 (N_7744,N_4456,N_4478);
and U7745 (N_7745,N_3264,N_3051);
or U7746 (N_7746,N_4845,N_4638);
nand U7747 (N_7747,N_3347,N_4065);
nor U7748 (N_7748,N_4167,N_5080);
nor U7749 (N_7749,N_4343,N_3071);
nand U7750 (N_7750,N_4568,N_5646);
and U7751 (N_7751,N_4154,N_3381);
or U7752 (N_7752,N_5335,N_3973);
nand U7753 (N_7753,N_5413,N_5080);
or U7754 (N_7754,N_5086,N_4486);
nor U7755 (N_7755,N_5243,N_3553);
nor U7756 (N_7756,N_4211,N_4677);
nand U7757 (N_7757,N_3095,N_3930);
and U7758 (N_7758,N_3526,N_4753);
or U7759 (N_7759,N_3718,N_3279);
nand U7760 (N_7760,N_3247,N_4819);
nor U7761 (N_7761,N_3172,N_4812);
and U7762 (N_7762,N_4983,N_4274);
and U7763 (N_7763,N_5904,N_5010);
nor U7764 (N_7764,N_3826,N_5405);
nand U7765 (N_7765,N_4908,N_3590);
nand U7766 (N_7766,N_4590,N_3084);
nand U7767 (N_7767,N_5229,N_4216);
or U7768 (N_7768,N_4433,N_3561);
nor U7769 (N_7769,N_5544,N_3937);
or U7770 (N_7770,N_4204,N_4972);
nand U7771 (N_7771,N_5419,N_3491);
or U7772 (N_7772,N_4188,N_4390);
nand U7773 (N_7773,N_4693,N_4629);
nand U7774 (N_7774,N_4070,N_3852);
nand U7775 (N_7775,N_3611,N_5780);
nand U7776 (N_7776,N_4845,N_4087);
and U7777 (N_7777,N_4427,N_3107);
and U7778 (N_7778,N_3599,N_5186);
or U7779 (N_7779,N_5951,N_4009);
nor U7780 (N_7780,N_5991,N_4509);
and U7781 (N_7781,N_3082,N_3457);
or U7782 (N_7782,N_4373,N_4321);
nor U7783 (N_7783,N_4700,N_5444);
and U7784 (N_7784,N_3882,N_3682);
nand U7785 (N_7785,N_3115,N_3884);
nand U7786 (N_7786,N_3441,N_4933);
nand U7787 (N_7787,N_5784,N_4733);
nand U7788 (N_7788,N_3293,N_4184);
and U7789 (N_7789,N_5974,N_4152);
or U7790 (N_7790,N_3429,N_5975);
nand U7791 (N_7791,N_5539,N_4958);
or U7792 (N_7792,N_5876,N_3724);
or U7793 (N_7793,N_3853,N_5027);
nor U7794 (N_7794,N_3633,N_4417);
nand U7795 (N_7795,N_4267,N_5814);
or U7796 (N_7796,N_5437,N_4327);
nand U7797 (N_7797,N_3698,N_4921);
nand U7798 (N_7798,N_3070,N_3605);
and U7799 (N_7799,N_3937,N_5832);
and U7800 (N_7800,N_3500,N_5919);
nand U7801 (N_7801,N_5320,N_4301);
or U7802 (N_7802,N_3671,N_5083);
and U7803 (N_7803,N_4855,N_3513);
nor U7804 (N_7804,N_3241,N_4552);
nor U7805 (N_7805,N_3932,N_4328);
or U7806 (N_7806,N_4366,N_4476);
and U7807 (N_7807,N_3876,N_3101);
nor U7808 (N_7808,N_3681,N_4017);
nor U7809 (N_7809,N_5237,N_3393);
or U7810 (N_7810,N_3116,N_3460);
nand U7811 (N_7811,N_5412,N_4846);
nor U7812 (N_7812,N_3603,N_4910);
or U7813 (N_7813,N_3082,N_3228);
nand U7814 (N_7814,N_3277,N_5606);
nor U7815 (N_7815,N_3098,N_5914);
nor U7816 (N_7816,N_4422,N_3337);
or U7817 (N_7817,N_5880,N_5272);
nor U7818 (N_7818,N_3278,N_5475);
nand U7819 (N_7819,N_5119,N_4176);
or U7820 (N_7820,N_4967,N_3714);
and U7821 (N_7821,N_4284,N_4501);
nor U7822 (N_7822,N_4367,N_3670);
and U7823 (N_7823,N_4539,N_3034);
nor U7824 (N_7824,N_3275,N_5353);
nand U7825 (N_7825,N_5051,N_5887);
nor U7826 (N_7826,N_4872,N_5910);
nor U7827 (N_7827,N_5095,N_3155);
and U7828 (N_7828,N_5587,N_5232);
and U7829 (N_7829,N_5449,N_5248);
nor U7830 (N_7830,N_5372,N_4233);
nor U7831 (N_7831,N_4574,N_4800);
nand U7832 (N_7832,N_3277,N_5867);
and U7833 (N_7833,N_5911,N_3887);
or U7834 (N_7834,N_3497,N_4277);
or U7835 (N_7835,N_5592,N_3271);
or U7836 (N_7836,N_5678,N_5373);
xnor U7837 (N_7837,N_3112,N_3237);
or U7838 (N_7838,N_4338,N_4689);
nor U7839 (N_7839,N_4736,N_4433);
or U7840 (N_7840,N_4109,N_3106);
nand U7841 (N_7841,N_4940,N_4630);
nand U7842 (N_7842,N_4779,N_5817);
nand U7843 (N_7843,N_4394,N_3717);
nor U7844 (N_7844,N_4537,N_4726);
and U7845 (N_7845,N_3906,N_4426);
or U7846 (N_7846,N_5527,N_5652);
or U7847 (N_7847,N_4652,N_4954);
nand U7848 (N_7848,N_5641,N_4543);
nor U7849 (N_7849,N_3428,N_5223);
nor U7850 (N_7850,N_3754,N_5558);
and U7851 (N_7851,N_5737,N_3907);
nand U7852 (N_7852,N_3475,N_5638);
or U7853 (N_7853,N_4151,N_3071);
nor U7854 (N_7854,N_3135,N_3164);
nand U7855 (N_7855,N_3875,N_5974);
or U7856 (N_7856,N_3645,N_5995);
or U7857 (N_7857,N_4161,N_3882);
nand U7858 (N_7858,N_5666,N_4900);
or U7859 (N_7859,N_3369,N_5699);
nand U7860 (N_7860,N_3723,N_3558);
nand U7861 (N_7861,N_3447,N_5116);
nand U7862 (N_7862,N_5255,N_3840);
nor U7863 (N_7863,N_3160,N_4227);
and U7864 (N_7864,N_4761,N_5979);
nor U7865 (N_7865,N_5786,N_3737);
nor U7866 (N_7866,N_4818,N_4886);
or U7867 (N_7867,N_5995,N_5173);
nor U7868 (N_7868,N_4790,N_3051);
and U7869 (N_7869,N_4647,N_3177);
nor U7870 (N_7870,N_5460,N_3136);
or U7871 (N_7871,N_4217,N_4256);
and U7872 (N_7872,N_5941,N_5832);
nor U7873 (N_7873,N_4888,N_4352);
or U7874 (N_7874,N_4898,N_3495);
and U7875 (N_7875,N_3725,N_3046);
nand U7876 (N_7876,N_5474,N_4344);
nand U7877 (N_7877,N_5557,N_5664);
nand U7878 (N_7878,N_4395,N_5776);
and U7879 (N_7879,N_4319,N_5303);
nand U7880 (N_7880,N_4438,N_4075);
nor U7881 (N_7881,N_4848,N_4452);
nand U7882 (N_7882,N_4180,N_4850);
and U7883 (N_7883,N_3496,N_5706);
nand U7884 (N_7884,N_5581,N_4814);
nand U7885 (N_7885,N_3657,N_5291);
or U7886 (N_7886,N_3019,N_3533);
nand U7887 (N_7887,N_5746,N_3566);
or U7888 (N_7888,N_3440,N_5176);
or U7889 (N_7889,N_4970,N_3465);
nand U7890 (N_7890,N_3420,N_3204);
nor U7891 (N_7891,N_5958,N_5842);
and U7892 (N_7892,N_4175,N_4109);
and U7893 (N_7893,N_3027,N_4159);
or U7894 (N_7894,N_5569,N_5447);
and U7895 (N_7895,N_3574,N_4863);
nor U7896 (N_7896,N_4238,N_3349);
nand U7897 (N_7897,N_5969,N_5088);
and U7898 (N_7898,N_3528,N_5902);
nor U7899 (N_7899,N_3404,N_4975);
nand U7900 (N_7900,N_4436,N_4592);
nor U7901 (N_7901,N_4761,N_5027);
and U7902 (N_7902,N_4280,N_3606);
and U7903 (N_7903,N_5459,N_4361);
nor U7904 (N_7904,N_5378,N_3086);
nor U7905 (N_7905,N_4708,N_5073);
and U7906 (N_7906,N_4383,N_4608);
or U7907 (N_7907,N_4693,N_3506);
nand U7908 (N_7908,N_4517,N_5871);
nand U7909 (N_7909,N_3214,N_4280);
nand U7910 (N_7910,N_4145,N_5928);
nand U7911 (N_7911,N_5269,N_3101);
nand U7912 (N_7912,N_4229,N_3501);
and U7913 (N_7913,N_3872,N_5844);
nor U7914 (N_7914,N_5485,N_3738);
and U7915 (N_7915,N_4842,N_3187);
nor U7916 (N_7916,N_5882,N_3649);
and U7917 (N_7917,N_5454,N_5625);
nor U7918 (N_7918,N_5291,N_4257);
or U7919 (N_7919,N_4624,N_5360);
nor U7920 (N_7920,N_4208,N_3077);
or U7921 (N_7921,N_3051,N_3505);
and U7922 (N_7922,N_4776,N_3156);
nor U7923 (N_7923,N_5804,N_3819);
and U7924 (N_7924,N_4394,N_5477);
or U7925 (N_7925,N_5419,N_4240);
and U7926 (N_7926,N_4990,N_5542);
nand U7927 (N_7927,N_5938,N_3985);
nor U7928 (N_7928,N_5338,N_5870);
nand U7929 (N_7929,N_3663,N_3713);
or U7930 (N_7930,N_5131,N_5534);
and U7931 (N_7931,N_3173,N_4322);
and U7932 (N_7932,N_4006,N_3182);
and U7933 (N_7933,N_4817,N_4383);
nor U7934 (N_7934,N_3854,N_3011);
nand U7935 (N_7935,N_3673,N_3974);
or U7936 (N_7936,N_3800,N_4031);
nand U7937 (N_7937,N_3575,N_4191);
and U7938 (N_7938,N_5943,N_4010);
nor U7939 (N_7939,N_5134,N_3637);
nor U7940 (N_7940,N_5587,N_5929);
nor U7941 (N_7941,N_4783,N_5166);
nand U7942 (N_7942,N_4107,N_4510);
or U7943 (N_7943,N_3716,N_5998);
or U7944 (N_7944,N_4321,N_5715);
nand U7945 (N_7945,N_3840,N_3193);
or U7946 (N_7946,N_3972,N_4471);
and U7947 (N_7947,N_4627,N_3794);
and U7948 (N_7948,N_3089,N_4854);
or U7949 (N_7949,N_3963,N_4429);
nand U7950 (N_7950,N_4941,N_5101);
nor U7951 (N_7951,N_4413,N_3538);
nor U7952 (N_7952,N_3109,N_5446);
nor U7953 (N_7953,N_5992,N_5127);
and U7954 (N_7954,N_4120,N_4881);
nor U7955 (N_7955,N_5216,N_4311);
and U7956 (N_7956,N_5934,N_5460);
or U7957 (N_7957,N_5870,N_4049);
and U7958 (N_7958,N_4292,N_3518);
nand U7959 (N_7959,N_3767,N_4859);
or U7960 (N_7960,N_5520,N_4241);
and U7961 (N_7961,N_5017,N_3301);
nor U7962 (N_7962,N_4290,N_4672);
or U7963 (N_7963,N_5812,N_4801);
and U7964 (N_7964,N_4469,N_3325);
or U7965 (N_7965,N_4344,N_4767);
nor U7966 (N_7966,N_5897,N_4449);
nor U7967 (N_7967,N_4220,N_3961);
nand U7968 (N_7968,N_5064,N_3474);
nor U7969 (N_7969,N_5207,N_5282);
nand U7970 (N_7970,N_4178,N_3780);
nand U7971 (N_7971,N_4139,N_3352);
nor U7972 (N_7972,N_4057,N_4027);
nand U7973 (N_7973,N_4467,N_4658);
or U7974 (N_7974,N_5814,N_3088);
and U7975 (N_7975,N_5550,N_5654);
xor U7976 (N_7976,N_4921,N_4492);
and U7977 (N_7977,N_5534,N_5753);
and U7978 (N_7978,N_3908,N_4844);
and U7979 (N_7979,N_4865,N_5712);
nor U7980 (N_7980,N_5541,N_4631);
or U7981 (N_7981,N_3375,N_4451);
and U7982 (N_7982,N_3816,N_4443);
or U7983 (N_7983,N_5230,N_5017);
nand U7984 (N_7984,N_3243,N_3586);
or U7985 (N_7985,N_3128,N_3033);
nand U7986 (N_7986,N_4141,N_4295);
and U7987 (N_7987,N_3966,N_5797);
nor U7988 (N_7988,N_3030,N_4312);
or U7989 (N_7989,N_4324,N_4011);
or U7990 (N_7990,N_3411,N_3825);
and U7991 (N_7991,N_4895,N_3689);
and U7992 (N_7992,N_4056,N_3806);
nor U7993 (N_7993,N_5954,N_5202);
or U7994 (N_7994,N_4011,N_5201);
nor U7995 (N_7995,N_4997,N_4661);
or U7996 (N_7996,N_4652,N_5322);
nand U7997 (N_7997,N_4074,N_4992);
nand U7998 (N_7998,N_3759,N_5847);
nand U7999 (N_7999,N_5279,N_3738);
nand U8000 (N_8000,N_3557,N_3296);
or U8001 (N_8001,N_5713,N_5777);
nand U8002 (N_8002,N_4284,N_5779);
nor U8003 (N_8003,N_5342,N_5143);
or U8004 (N_8004,N_5243,N_5406);
or U8005 (N_8005,N_5433,N_4889);
and U8006 (N_8006,N_3142,N_5351);
nand U8007 (N_8007,N_4987,N_5342);
and U8008 (N_8008,N_3146,N_5876);
nand U8009 (N_8009,N_3493,N_3406);
nand U8010 (N_8010,N_5012,N_3200);
nor U8011 (N_8011,N_3068,N_4239);
and U8012 (N_8012,N_3170,N_5614);
and U8013 (N_8013,N_3474,N_4346);
nor U8014 (N_8014,N_4258,N_5286);
nor U8015 (N_8015,N_4033,N_3551);
and U8016 (N_8016,N_4999,N_5038);
nor U8017 (N_8017,N_5391,N_4358);
and U8018 (N_8018,N_5980,N_4546);
nor U8019 (N_8019,N_4086,N_3985);
and U8020 (N_8020,N_4649,N_4905);
and U8021 (N_8021,N_3952,N_4287);
or U8022 (N_8022,N_4250,N_4404);
nand U8023 (N_8023,N_4579,N_4267);
and U8024 (N_8024,N_3132,N_3150);
nand U8025 (N_8025,N_5192,N_4336);
nand U8026 (N_8026,N_4945,N_5163);
or U8027 (N_8027,N_4484,N_4308);
nor U8028 (N_8028,N_3440,N_3437);
nor U8029 (N_8029,N_5021,N_3588);
nor U8030 (N_8030,N_4018,N_3357);
nand U8031 (N_8031,N_5803,N_5271);
and U8032 (N_8032,N_3175,N_5660);
and U8033 (N_8033,N_4280,N_5092);
nor U8034 (N_8034,N_4939,N_4998);
and U8035 (N_8035,N_3717,N_3394);
and U8036 (N_8036,N_4152,N_3792);
nor U8037 (N_8037,N_4717,N_4496);
nor U8038 (N_8038,N_3084,N_3761);
nor U8039 (N_8039,N_4864,N_3764);
and U8040 (N_8040,N_5754,N_4842);
or U8041 (N_8041,N_3355,N_4660);
nand U8042 (N_8042,N_4199,N_3720);
and U8043 (N_8043,N_5681,N_3676);
nor U8044 (N_8044,N_5091,N_4563);
or U8045 (N_8045,N_5316,N_3722);
nand U8046 (N_8046,N_3118,N_5684);
or U8047 (N_8047,N_5646,N_4292);
and U8048 (N_8048,N_4708,N_5435);
nand U8049 (N_8049,N_5907,N_3173);
and U8050 (N_8050,N_5173,N_5697);
nand U8051 (N_8051,N_5396,N_3816);
or U8052 (N_8052,N_5862,N_3339);
and U8053 (N_8053,N_3498,N_3240);
and U8054 (N_8054,N_3122,N_5229);
or U8055 (N_8055,N_4500,N_3464);
nor U8056 (N_8056,N_4430,N_5566);
or U8057 (N_8057,N_3297,N_5548);
nand U8058 (N_8058,N_5271,N_4660);
and U8059 (N_8059,N_5468,N_5394);
nor U8060 (N_8060,N_3043,N_3768);
or U8061 (N_8061,N_4686,N_5455);
nor U8062 (N_8062,N_3393,N_5163);
or U8063 (N_8063,N_5501,N_4552);
nor U8064 (N_8064,N_3050,N_3936);
nand U8065 (N_8065,N_3283,N_4560);
nor U8066 (N_8066,N_4731,N_4499);
or U8067 (N_8067,N_3336,N_4757);
nor U8068 (N_8068,N_3918,N_4674);
or U8069 (N_8069,N_4594,N_5967);
xnor U8070 (N_8070,N_5062,N_3314);
nor U8071 (N_8071,N_4340,N_3234);
and U8072 (N_8072,N_3374,N_3936);
or U8073 (N_8073,N_4261,N_4196);
or U8074 (N_8074,N_4461,N_5851);
nand U8075 (N_8075,N_3422,N_5441);
or U8076 (N_8076,N_3577,N_4188);
nor U8077 (N_8077,N_3312,N_5748);
or U8078 (N_8078,N_5978,N_3913);
nand U8079 (N_8079,N_3278,N_4207);
and U8080 (N_8080,N_4904,N_4164);
nor U8081 (N_8081,N_5319,N_3260);
or U8082 (N_8082,N_4603,N_5080);
nor U8083 (N_8083,N_3193,N_4561);
and U8084 (N_8084,N_4530,N_3947);
nor U8085 (N_8085,N_4154,N_5763);
or U8086 (N_8086,N_4584,N_3444);
nor U8087 (N_8087,N_3202,N_5822);
or U8088 (N_8088,N_4611,N_4252);
nand U8089 (N_8089,N_4324,N_4185);
and U8090 (N_8090,N_5587,N_4503);
nor U8091 (N_8091,N_4466,N_4126);
and U8092 (N_8092,N_5690,N_5342);
nand U8093 (N_8093,N_5735,N_5134);
nor U8094 (N_8094,N_5206,N_4552);
nor U8095 (N_8095,N_4682,N_4151);
and U8096 (N_8096,N_4034,N_3993);
and U8097 (N_8097,N_5091,N_4639);
nor U8098 (N_8098,N_3328,N_5333);
or U8099 (N_8099,N_3133,N_5151);
or U8100 (N_8100,N_3358,N_4375);
nand U8101 (N_8101,N_4844,N_3423);
and U8102 (N_8102,N_3681,N_5502);
or U8103 (N_8103,N_3609,N_4356);
or U8104 (N_8104,N_5004,N_3411);
nor U8105 (N_8105,N_5199,N_3682);
nor U8106 (N_8106,N_3022,N_3190);
or U8107 (N_8107,N_5793,N_3395);
or U8108 (N_8108,N_5922,N_3409);
nor U8109 (N_8109,N_4170,N_4641);
and U8110 (N_8110,N_3693,N_4369);
nand U8111 (N_8111,N_4123,N_4581);
or U8112 (N_8112,N_4963,N_3589);
and U8113 (N_8113,N_3398,N_3770);
nor U8114 (N_8114,N_4808,N_5532);
or U8115 (N_8115,N_4627,N_3535);
and U8116 (N_8116,N_4802,N_3028);
and U8117 (N_8117,N_4480,N_5699);
xnor U8118 (N_8118,N_4979,N_3293);
nor U8119 (N_8119,N_4017,N_4948);
and U8120 (N_8120,N_4935,N_5876);
and U8121 (N_8121,N_3359,N_5862);
or U8122 (N_8122,N_3010,N_3006);
and U8123 (N_8123,N_3252,N_4879);
or U8124 (N_8124,N_5173,N_4963);
or U8125 (N_8125,N_3540,N_5485);
or U8126 (N_8126,N_3399,N_3041);
or U8127 (N_8127,N_4580,N_3069);
and U8128 (N_8128,N_5779,N_5550);
nand U8129 (N_8129,N_5176,N_3456);
nor U8130 (N_8130,N_4549,N_4194);
nor U8131 (N_8131,N_5642,N_5772);
or U8132 (N_8132,N_5352,N_3147);
and U8133 (N_8133,N_5627,N_4034);
and U8134 (N_8134,N_4925,N_5361);
and U8135 (N_8135,N_3208,N_3937);
nor U8136 (N_8136,N_4552,N_3495);
and U8137 (N_8137,N_4442,N_3707);
or U8138 (N_8138,N_3918,N_4744);
nand U8139 (N_8139,N_3838,N_4521);
nand U8140 (N_8140,N_4888,N_3071);
nand U8141 (N_8141,N_4121,N_4707);
nand U8142 (N_8142,N_5384,N_5495);
or U8143 (N_8143,N_3084,N_4471);
nor U8144 (N_8144,N_4689,N_5889);
nand U8145 (N_8145,N_4049,N_3153);
nand U8146 (N_8146,N_3171,N_3908);
and U8147 (N_8147,N_3587,N_3916);
nand U8148 (N_8148,N_5380,N_4242);
nand U8149 (N_8149,N_3363,N_3051);
and U8150 (N_8150,N_5265,N_4314);
nor U8151 (N_8151,N_3987,N_3959);
and U8152 (N_8152,N_4360,N_4246);
and U8153 (N_8153,N_5812,N_5179);
and U8154 (N_8154,N_5993,N_3475);
or U8155 (N_8155,N_4749,N_3514);
and U8156 (N_8156,N_3859,N_5290);
xnor U8157 (N_8157,N_5721,N_5791);
or U8158 (N_8158,N_3092,N_5147);
nor U8159 (N_8159,N_5440,N_4842);
or U8160 (N_8160,N_5510,N_4884);
nor U8161 (N_8161,N_5414,N_4803);
and U8162 (N_8162,N_4233,N_5718);
and U8163 (N_8163,N_3575,N_4087);
nand U8164 (N_8164,N_3926,N_3847);
or U8165 (N_8165,N_5894,N_3705);
and U8166 (N_8166,N_5796,N_5400);
or U8167 (N_8167,N_4223,N_5276);
or U8168 (N_8168,N_5744,N_3792);
and U8169 (N_8169,N_5205,N_3219);
and U8170 (N_8170,N_5015,N_4623);
or U8171 (N_8171,N_3508,N_5176);
nor U8172 (N_8172,N_3392,N_3860);
nor U8173 (N_8173,N_5039,N_3861);
or U8174 (N_8174,N_3609,N_4375);
nor U8175 (N_8175,N_3608,N_3851);
nand U8176 (N_8176,N_5761,N_5461);
or U8177 (N_8177,N_5062,N_3586);
nor U8178 (N_8178,N_4200,N_5998);
or U8179 (N_8179,N_3203,N_4345);
nand U8180 (N_8180,N_5138,N_3139);
and U8181 (N_8181,N_3589,N_5351);
and U8182 (N_8182,N_4549,N_3240);
and U8183 (N_8183,N_4778,N_4985);
and U8184 (N_8184,N_4924,N_5830);
and U8185 (N_8185,N_4085,N_3728);
nor U8186 (N_8186,N_3070,N_5555);
or U8187 (N_8187,N_5412,N_4161);
and U8188 (N_8188,N_5725,N_4130);
nor U8189 (N_8189,N_4816,N_5198);
nand U8190 (N_8190,N_5650,N_4480);
nor U8191 (N_8191,N_5550,N_4361);
nor U8192 (N_8192,N_4957,N_4191);
nand U8193 (N_8193,N_5451,N_5802);
nand U8194 (N_8194,N_5839,N_4838);
and U8195 (N_8195,N_5928,N_3409);
nor U8196 (N_8196,N_4147,N_3473);
and U8197 (N_8197,N_5677,N_3148);
or U8198 (N_8198,N_5888,N_4120);
nor U8199 (N_8199,N_4257,N_5380);
and U8200 (N_8200,N_5833,N_3347);
nor U8201 (N_8201,N_4286,N_5999);
nand U8202 (N_8202,N_4530,N_4509);
nor U8203 (N_8203,N_3214,N_3282);
and U8204 (N_8204,N_3710,N_4794);
or U8205 (N_8205,N_5829,N_5251);
nor U8206 (N_8206,N_3185,N_3208);
and U8207 (N_8207,N_3761,N_3615);
nand U8208 (N_8208,N_5525,N_5345);
and U8209 (N_8209,N_5678,N_3955);
nand U8210 (N_8210,N_5389,N_3873);
nor U8211 (N_8211,N_5875,N_4285);
and U8212 (N_8212,N_4231,N_4394);
nor U8213 (N_8213,N_5946,N_4749);
and U8214 (N_8214,N_5415,N_5725);
or U8215 (N_8215,N_5689,N_4411);
nor U8216 (N_8216,N_3521,N_3757);
nor U8217 (N_8217,N_4401,N_4086);
nor U8218 (N_8218,N_4259,N_3834);
nor U8219 (N_8219,N_4086,N_4777);
xnor U8220 (N_8220,N_4421,N_3320);
and U8221 (N_8221,N_4089,N_4259);
or U8222 (N_8222,N_5333,N_3634);
and U8223 (N_8223,N_4728,N_5804);
and U8224 (N_8224,N_4335,N_4443);
and U8225 (N_8225,N_3196,N_4236);
and U8226 (N_8226,N_5199,N_3254);
nand U8227 (N_8227,N_4423,N_4843);
nor U8228 (N_8228,N_5802,N_3510);
and U8229 (N_8229,N_3303,N_4060);
or U8230 (N_8230,N_5934,N_5115);
and U8231 (N_8231,N_3738,N_5417);
and U8232 (N_8232,N_4584,N_4189);
nor U8233 (N_8233,N_5392,N_3432);
nor U8234 (N_8234,N_3572,N_3069);
nand U8235 (N_8235,N_4916,N_3638);
nor U8236 (N_8236,N_4592,N_3611);
and U8237 (N_8237,N_4044,N_5614);
nor U8238 (N_8238,N_4750,N_5614);
nor U8239 (N_8239,N_5279,N_4252);
or U8240 (N_8240,N_3979,N_4404);
nand U8241 (N_8241,N_5789,N_3044);
and U8242 (N_8242,N_3764,N_5695);
nand U8243 (N_8243,N_5183,N_4049);
nand U8244 (N_8244,N_3217,N_5444);
nor U8245 (N_8245,N_3894,N_5150);
or U8246 (N_8246,N_4894,N_3062);
and U8247 (N_8247,N_3823,N_4093);
nor U8248 (N_8248,N_3918,N_4099);
nor U8249 (N_8249,N_3119,N_5224);
or U8250 (N_8250,N_4866,N_5380);
and U8251 (N_8251,N_3087,N_3470);
nor U8252 (N_8252,N_5367,N_4031);
or U8253 (N_8253,N_3983,N_4789);
nor U8254 (N_8254,N_3592,N_3247);
or U8255 (N_8255,N_3963,N_3918);
or U8256 (N_8256,N_3832,N_3200);
nand U8257 (N_8257,N_5339,N_5010);
nor U8258 (N_8258,N_5019,N_4372);
and U8259 (N_8259,N_4095,N_4269);
xnor U8260 (N_8260,N_3629,N_3726);
or U8261 (N_8261,N_5811,N_3569);
nor U8262 (N_8262,N_5078,N_5031);
or U8263 (N_8263,N_4748,N_3679);
nor U8264 (N_8264,N_4691,N_3962);
or U8265 (N_8265,N_5182,N_5551);
or U8266 (N_8266,N_5118,N_4502);
nor U8267 (N_8267,N_3333,N_4105);
nor U8268 (N_8268,N_5317,N_4191);
nand U8269 (N_8269,N_4437,N_3946);
or U8270 (N_8270,N_4470,N_5279);
and U8271 (N_8271,N_4007,N_3142);
or U8272 (N_8272,N_4968,N_3316);
nand U8273 (N_8273,N_5228,N_3117);
nor U8274 (N_8274,N_4875,N_5436);
or U8275 (N_8275,N_3792,N_5708);
nor U8276 (N_8276,N_4332,N_3189);
nand U8277 (N_8277,N_4564,N_3858);
nor U8278 (N_8278,N_3680,N_5060);
and U8279 (N_8279,N_5625,N_5419);
nand U8280 (N_8280,N_3548,N_4427);
or U8281 (N_8281,N_3275,N_4921);
or U8282 (N_8282,N_5002,N_4709);
nor U8283 (N_8283,N_3815,N_5279);
nor U8284 (N_8284,N_5309,N_5917);
or U8285 (N_8285,N_4286,N_5790);
nor U8286 (N_8286,N_3219,N_3476);
or U8287 (N_8287,N_3490,N_3172);
nor U8288 (N_8288,N_3458,N_4831);
nor U8289 (N_8289,N_4625,N_3793);
nor U8290 (N_8290,N_5438,N_5632);
nor U8291 (N_8291,N_5921,N_4958);
and U8292 (N_8292,N_4867,N_5877);
or U8293 (N_8293,N_5059,N_5018);
nor U8294 (N_8294,N_4393,N_5860);
nand U8295 (N_8295,N_3540,N_3462);
nand U8296 (N_8296,N_3462,N_3703);
nand U8297 (N_8297,N_3213,N_5495);
nor U8298 (N_8298,N_4877,N_5462);
or U8299 (N_8299,N_5994,N_4579);
nand U8300 (N_8300,N_4552,N_3194);
or U8301 (N_8301,N_5683,N_5936);
nor U8302 (N_8302,N_4617,N_5822);
nor U8303 (N_8303,N_3871,N_3118);
nand U8304 (N_8304,N_5237,N_5587);
and U8305 (N_8305,N_5196,N_3872);
or U8306 (N_8306,N_5673,N_5273);
and U8307 (N_8307,N_4934,N_4777);
and U8308 (N_8308,N_3632,N_3685);
nand U8309 (N_8309,N_4948,N_4489);
and U8310 (N_8310,N_5855,N_5612);
nand U8311 (N_8311,N_4663,N_4519);
nand U8312 (N_8312,N_5191,N_5526);
and U8313 (N_8313,N_4521,N_3515);
nand U8314 (N_8314,N_5669,N_4493);
nand U8315 (N_8315,N_3359,N_3248);
and U8316 (N_8316,N_4484,N_4536);
nor U8317 (N_8317,N_5214,N_5287);
nand U8318 (N_8318,N_5750,N_3736);
nor U8319 (N_8319,N_5068,N_3526);
nand U8320 (N_8320,N_3944,N_5310);
nor U8321 (N_8321,N_4862,N_4766);
or U8322 (N_8322,N_5402,N_4010);
nand U8323 (N_8323,N_5692,N_5027);
nand U8324 (N_8324,N_3772,N_3269);
nor U8325 (N_8325,N_5320,N_4598);
nor U8326 (N_8326,N_4617,N_5675);
nand U8327 (N_8327,N_3785,N_4579);
nand U8328 (N_8328,N_5611,N_4130);
and U8329 (N_8329,N_3830,N_4946);
nand U8330 (N_8330,N_3048,N_4768);
or U8331 (N_8331,N_5990,N_5105);
nor U8332 (N_8332,N_3192,N_3725);
nand U8333 (N_8333,N_4090,N_3188);
nand U8334 (N_8334,N_4000,N_5454);
and U8335 (N_8335,N_5113,N_5512);
or U8336 (N_8336,N_3401,N_4652);
nand U8337 (N_8337,N_4190,N_5122);
nand U8338 (N_8338,N_4785,N_3486);
or U8339 (N_8339,N_5035,N_3186);
nor U8340 (N_8340,N_5474,N_3670);
and U8341 (N_8341,N_4313,N_3888);
nand U8342 (N_8342,N_5953,N_5371);
nor U8343 (N_8343,N_3817,N_3518);
and U8344 (N_8344,N_5784,N_4006);
nand U8345 (N_8345,N_4485,N_3791);
nor U8346 (N_8346,N_5378,N_3267);
and U8347 (N_8347,N_3415,N_5338);
nor U8348 (N_8348,N_4445,N_3395);
or U8349 (N_8349,N_4311,N_3487);
and U8350 (N_8350,N_5788,N_5424);
nor U8351 (N_8351,N_4475,N_3610);
and U8352 (N_8352,N_5504,N_5203);
or U8353 (N_8353,N_3390,N_4143);
nand U8354 (N_8354,N_5714,N_3562);
or U8355 (N_8355,N_4506,N_5839);
nor U8356 (N_8356,N_4114,N_3568);
and U8357 (N_8357,N_4535,N_3010);
nand U8358 (N_8358,N_3775,N_5730);
nor U8359 (N_8359,N_5227,N_4392);
and U8360 (N_8360,N_4195,N_4423);
or U8361 (N_8361,N_5577,N_4921);
and U8362 (N_8362,N_5416,N_5423);
and U8363 (N_8363,N_3059,N_4486);
or U8364 (N_8364,N_5063,N_4347);
nor U8365 (N_8365,N_3687,N_3659);
or U8366 (N_8366,N_5015,N_5678);
nor U8367 (N_8367,N_3967,N_3464);
nand U8368 (N_8368,N_4610,N_4197);
nand U8369 (N_8369,N_5270,N_3941);
nand U8370 (N_8370,N_3568,N_5128);
or U8371 (N_8371,N_5996,N_3477);
nor U8372 (N_8372,N_5128,N_5118);
and U8373 (N_8373,N_4884,N_3031);
and U8374 (N_8374,N_4898,N_4603);
nor U8375 (N_8375,N_5015,N_4509);
nor U8376 (N_8376,N_5628,N_4547);
nor U8377 (N_8377,N_4011,N_5431);
nand U8378 (N_8378,N_4308,N_3330);
and U8379 (N_8379,N_3169,N_4870);
and U8380 (N_8380,N_5713,N_3184);
nand U8381 (N_8381,N_3098,N_3259);
and U8382 (N_8382,N_4085,N_5012);
or U8383 (N_8383,N_5230,N_3894);
or U8384 (N_8384,N_3154,N_3307);
nor U8385 (N_8385,N_5021,N_3701);
nor U8386 (N_8386,N_3472,N_3784);
nand U8387 (N_8387,N_3040,N_5826);
nor U8388 (N_8388,N_3789,N_4012);
nand U8389 (N_8389,N_4755,N_4358);
nor U8390 (N_8390,N_5341,N_5049);
or U8391 (N_8391,N_4675,N_5095);
nor U8392 (N_8392,N_3376,N_3508);
nand U8393 (N_8393,N_4503,N_3081);
and U8394 (N_8394,N_3495,N_4683);
nor U8395 (N_8395,N_5134,N_4789);
nor U8396 (N_8396,N_3648,N_5179);
and U8397 (N_8397,N_3264,N_5522);
or U8398 (N_8398,N_5601,N_3272);
and U8399 (N_8399,N_4112,N_5007);
or U8400 (N_8400,N_5080,N_4351);
or U8401 (N_8401,N_4187,N_4872);
and U8402 (N_8402,N_4232,N_3389);
nand U8403 (N_8403,N_5828,N_5429);
nor U8404 (N_8404,N_5041,N_5164);
and U8405 (N_8405,N_5036,N_3843);
and U8406 (N_8406,N_4769,N_3587);
and U8407 (N_8407,N_4616,N_3142);
and U8408 (N_8408,N_3797,N_5543);
or U8409 (N_8409,N_5479,N_4586);
nand U8410 (N_8410,N_5389,N_4575);
nand U8411 (N_8411,N_4613,N_3630);
or U8412 (N_8412,N_3712,N_3410);
nand U8413 (N_8413,N_3388,N_5057);
and U8414 (N_8414,N_5210,N_4982);
nand U8415 (N_8415,N_3985,N_5205);
nor U8416 (N_8416,N_3713,N_3356);
nand U8417 (N_8417,N_4079,N_4314);
or U8418 (N_8418,N_3474,N_4988);
and U8419 (N_8419,N_4803,N_3345);
and U8420 (N_8420,N_5223,N_3887);
xnor U8421 (N_8421,N_5573,N_4971);
and U8422 (N_8422,N_3781,N_5431);
nand U8423 (N_8423,N_3284,N_5786);
and U8424 (N_8424,N_5123,N_4344);
nor U8425 (N_8425,N_4771,N_3353);
nor U8426 (N_8426,N_3686,N_3278);
nand U8427 (N_8427,N_5297,N_5259);
or U8428 (N_8428,N_4172,N_5825);
nand U8429 (N_8429,N_5343,N_3606);
or U8430 (N_8430,N_5574,N_3687);
nand U8431 (N_8431,N_4334,N_4763);
and U8432 (N_8432,N_4849,N_3394);
nor U8433 (N_8433,N_5187,N_4429);
or U8434 (N_8434,N_5657,N_4212);
nor U8435 (N_8435,N_4489,N_4782);
or U8436 (N_8436,N_5371,N_4030);
nand U8437 (N_8437,N_4457,N_4391);
or U8438 (N_8438,N_4031,N_4193);
and U8439 (N_8439,N_3148,N_3721);
nor U8440 (N_8440,N_4119,N_4713);
or U8441 (N_8441,N_5201,N_3566);
and U8442 (N_8442,N_3791,N_4549);
nor U8443 (N_8443,N_3664,N_5265);
and U8444 (N_8444,N_5171,N_4759);
nand U8445 (N_8445,N_4395,N_4284);
nand U8446 (N_8446,N_5035,N_3954);
nor U8447 (N_8447,N_5950,N_4933);
or U8448 (N_8448,N_5259,N_4949);
or U8449 (N_8449,N_3498,N_3624);
nand U8450 (N_8450,N_5179,N_3831);
and U8451 (N_8451,N_5510,N_5671);
nand U8452 (N_8452,N_5956,N_3828);
nor U8453 (N_8453,N_5383,N_5727);
and U8454 (N_8454,N_5799,N_5138);
and U8455 (N_8455,N_5698,N_4060);
nand U8456 (N_8456,N_3941,N_4964);
nor U8457 (N_8457,N_5589,N_5323);
nand U8458 (N_8458,N_3077,N_4348);
or U8459 (N_8459,N_3561,N_3438);
nor U8460 (N_8460,N_4190,N_5757);
and U8461 (N_8461,N_3644,N_5010);
or U8462 (N_8462,N_5517,N_4140);
nand U8463 (N_8463,N_3534,N_4607);
and U8464 (N_8464,N_3769,N_3470);
nor U8465 (N_8465,N_3319,N_5150);
nand U8466 (N_8466,N_3169,N_3476);
nor U8467 (N_8467,N_3597,N_4852);
or U8468 (N_8468,N_5415,N_3295);
nor U8469 (N_8469,N_3274,N_4795);
and U8470 (N_8470,N_5641,N_3109);
nand U8471 (N_8471,N_5068,N_4483);
and U8472 (N_8472,N_4337,N_3901);
nand U8473 (N_8473,N_5554,N_3909);
or U8474 (N_8474,N_5535,N_5291);
and U8475 (N_8475,N_3127,N_4327);
or U8476 (N_8476,N_4071,N_3137);
and U8477 (N_8477,N_5854,N_5715);
or U8478 (N_8478,N_3096,N_4651);
nor U8479 (N_8479,N_3774,N_5678);
or U8480 (N_8480,N_3729,N_5089);
nand U8481 (N_8481,N_4940,N_3939);
and U8482 (N_8482,N_3112,N_4833);
nor U8483 (N_8483,N_5249,N_5187);
and U8484 (N_8484,N_4168,N_4373);
and U8485 (N_8485,N_5581,N_4693);
nand U8486 (N_8486,N_5798,N_3632);
nor U8487 (N_8487,N_4804,N_3391);
nand U8488 (N_8488,N_3834,N_5405);
and U8489 (N_8489,N_5928,N_5794);
nand U8490 (N_8490,N_5415,N_3299);
nand U8491 (N_8491,N_5978,N_4845);
nor U8492 (N_8492,N_3600,N_4700);
nor U8493 (N_8493,N_4120,N_4037);
nand U8494 (N_8494,N_3378,N_5839);
or U8495 (N_8495,N_4182,N_4870);
or U8496 (N_8496,N_3402,N_3608);
nand U8497 (N_8497,N_4358,N_4120);
or U8498 (N_8498,N_5551,N_3318);
or U8499 (N_8499,N_3287,N_4837);
nor U8500 (N_8500,N_4869,N_3344);
nand U8501 (N_8501,N_3588,N_4224);
nand U8502 (N_8502,N_4584,N_4359);
or U8503 (N_8503,N_5780,N_5039);
nor U8504 (N_8504,N_4083,N_4362);
nand U8505 (N_8505,N_4192,N_4847);
nand U8506 (N_8506,N_5045,N_4626);
nor U8507 (N_8507,N_3300,N_4778);
nor U8508 (N_8508,N_4453,N_3262);
and U8509 (N_8509,N_4153,N_3361);
nand U8510 (N_8510,N_3293,N_3624);
nand U8511 (N_8511,N_5240,N_5542);
and U8512 (N_8512,N_5530,N_3706);
or U8513 (N_8513,N_3882,N_4893);
and U8514 (N_8514,N_5266,N_5646);
nor U8515 (N_8515,N_4915,N_4299);
nor U8516 (N_8516,N_4456,N_4038);
and U8517 (N_8517,N_3899,N_3881);
nor U8518 (N_8518,N_3440,N_3291);
and U8519 (N_8519,N_5412,N_3660);
or U8520 (N_8520,N_3706,N_3478);
nor U8521 (N_8521,N_3539,N_3759);
or U8522 (N_8522,N_4971,N_5853);
nand U8523 (N_8523,N_5855,N_3247);
and U8524 (N_8524,N_5227,N_3015);
and U8525 (N_8525,N_3048,N_3657);
and U8526 (N_8526,N_4591,N_3388);
nor U8527 (N_8527,N_5792,N_5478);
nor U8528 (N_8528,N_3205,N_5381);
or U8529 (N_8529,N_3470,N_5962);
nor U8530 (N_8530,N_4152,N_5637);
nand U8531 (N_8531,N_4769,N_4141);
or U8532 (N_8532,N_3105,N_5648);
or U8533 (N_8533,N_4688,N_3133);
or U8534 (N_8534,N_4169,N_3725);
or U8535 (N_8535,N_3217,N_5562);
nand U8536 (N_8536,N_4021,N_5796);
nor U8537 (N_8537,N_3956,N_5124);
and U8538 (N_8538,N_4220,N_5543);
or U8539 (N_8539,N_5766,N_3327);
or U8540 (N_8540,N_3431,N_4280);
nor U8541 (N_8541,N_4556,N_5192);
nor U8542 (N_8542,N_3463,N_3163);
nand U8543 (N_8543,N_3495,N_5196);
or U8544 (N_8544,N_3925,N_4330);
or U8545 (N_8545,N_5626,N_3866);
or U8546 (N_8546,N_5572,N_3149);
nand U8547 (N_8547,N_3474,N_4765);
or U8548 (N_8548,N_4147,N_5511);
or U8549 (N_8549,N_3292,N_4029);
nand U8550 (N_8550,N_5800,N_4557);
and U8551 (N_8551,N_3085,N_3155);
and U8552 (N_8552,N_4371,N_3066);
nor U8553 (N_8553,N_5073,N_5746);
or U8554 (N_8554,N_5139,N_5754);
or U8555 (N_8555,N_5689,N_4976);
nor U8556 (N_8556,N_3482,N_4874);
or U8557 (N_8557,N_4097,N_4473);
nor U8558 (N_8558,N_3930,N_5324);
or U8559 (N_8559,N_4632,N_4652);
nand U8560 (N_8560,N_4995,N_5450);
nor U8561 (N_8561,N_5533,N_3278);
or U8562 (N_8562,N_5131,N_4128);
nand U8563 (N_8563,N_5886,N_5858);
or U8564 (N_8564,N_5825,N_5593);
nand U8565 (N_8565,N_5259,N_4631);
nand U8566 (N_8566,N_4064,N_3407);
nand U8567 (N_8567,N_3135,N_3837);
and U8568 (N_8568,N_3076,N_5044);
nor U8569 (N_8569,N_5461,N_5483);
or U8570 (N_8570,N_4214,N_4733);
nand U8571 (N_8571,N_4116,N_3678);
nor U8572 (N_8572,N_5474,N_5583);
nand U8573 (N_8573,N_3041,N_5393);
or U8574 (N_8574,N_4151,N_5122);
nand U8575 (N_8575,N_3889,N_5288);
and U8576 (N_8576,N_4550,N_4945);
xnor U8577 (N_8577,N_5634,N_5376);
or U8578 (N_8578,N_5006,N_3418);
xor U8579 (N_8579,N_4674,N_4739);
or U8580 (N_8580,N_4834,N_4094);
nand U8581 (N_8581,N_3170,N_4266);
or U8582 (N_8582,N_4044,N_3709);
nor U8583 (N_8583,N_4334,N_4908);
nor U8584 (N_8584,N_3064,N_4616);
nor U8585 (N_8585,N_5721,N_5261);
nor U8586 (N_8586,N_3664,N_4471);
or U8587 (N_8587,N_3856,N_4518);
and U8588 (N_8588,N_5147,N_4589);
nor U8589 (N_8589,N_5157,N_5310);
and U8590 (N_8590,N_5514,N_5010);
or U8591 (N_8591,N_4625,N_5412);
nand U8592 (N_8592,N_3713,N_3729);
and U8593 (N_8593,N_4811,N_3651);
nand U8594 (N_8594,N_3839,N_5843);
or U8595 (N_8595,N_3436,N_3076);
nand U8596 (N_8596,N_3694,N_4669);
nand U8597 (N_8597,N_5613,N_4914);
or U8598 (N_8598,N_3741,N_3436);
nor U8599 (N_8599,N_3809,N_4251);
nand U8600 (N_8600,N_4986,N_5185);
nand U8601 (N_8601,N_3167,N_3914);
nand U8602 (N_8602,N_4121,N_4111);
and U8603 (N_8603,N_5805,N_5943);
nor U8604 (N_8604,N_4925,N_4765);
and U8605 (N_8605,N_5943,N_3322);
or U8606 (N_8606,N_4555,N_5901);
nor U8607 (N_8607,N_4655,N_4616);
nand U8608 (N_8608,N_3522,N_5446);
and U8609 (N_8609,N_4483,N_3850);
and U8610 (N_8610,N_3754,N_3333);
and U8611 (N_8611,N_5246,N_5139);
and U8612 (N_8612,N_3242,N_4450);
and U8613 (N_8613,N_3148,N_5154);
or U8614 (N_8614,N_3925,N_3464);
or U8615 (N_8615,N_3785,N_3057);
nand U8616 (N_8616,N_5683,N_3780);
nand U8617 (N_8617,N_3271,N_3780);
nand U8618 (N_8618,N_4567,N_5856);
and U8619 (N_8619,N_4537,N_3570);
and U8620 (N_8620,N_5329,N_4709);
nor U8621 (N_8621,N_4249,N_4265);
and U8622 (N_8622,N_5568,N_3739);
or U8623 (N_8623,N_4669,N_3790);
and U8624 (N_8624,N_3317,N_3604);
nor U8625 (N_8625,N_5826,N_4640);
nor U8626 (N_8626,N_5092,N_3314);
nand U8627 (N_8627,N_3202,N_3373);
or U8628 (N_8628,N_5194,N_4603);
nand U8629 (N_8629,N_5933,N_5567);
nor U8630 (N_8630,N_4668,N_3491);
and U8631 (N_8631,N_4171,N_5128);
or U8632 (N_8632,N_5762,N_3127);
nor U8633 (N_8633,N_5689,N_4131);
nor U8634 (N_8634,N_3852,N_5508);
and U8635 (N_8635,N_3936,N_3702);
nor U8636 (N_8636,N_4419,N_5081);
or U8637 (N_8637,N_4491,N_3608);
xnor U8638 (N_8638,N_3436,N_5059);
or U8639 (N_8639,N_3490,N_4585);
nand U8640 (N_8640,N_4451,N_3325);
and U8641 (N_8641,N_3914,N_4186);
nor U8642 (N_8642,N_5733,N_5664);
nand U8643 (N_8643,N_4586,N_3112);
nor U8644 (N_8644,N_3215,N_5608);
nor U8645 (N_8645,N_5798,N_5176);
or U8646 (N_8646,N_4115,N_5000);
and U8647 (N_8647,N_5888,N_4397);
or U8648 (N_8648,N_3519,N_5361);
nand U8649 (N_8649,N_3944,N_5358);
and U8650 (N_8650,N_4924,N_4404);
and U8651 (N_8651,N_5434,N_4860);
nor U8652 (N_8652,N_4028,N_5047);
nor U8653 (N_8653,N_4287,N_3284);
and U8654 (N_8654,N_3312,N_3434);
nor U8655 (N_8655,N_3326,N_4501);
and U8656 (N_8656,N_3438,N_5123);
and U8657 (N_8657,N_4424,N_4913);
or U8658 (N_8658,N_3500,N_3578);
and U8659 (N_8659,N_4202,N_3169);
nor U8660 (N_8660,N_3914,N_4719);
and U8661 (N_8661,N_4355,N_3845);
and U8662 (N_8662,N_4602,N_5393);
and U8663 (N_8663,N_5848,N_5487);
and U8664 (N_8664,N_3763,N_5389);
nor U8665 (N_8665,N_4283,N_5127);
nand U8666 (N_8666,N_3381,N_5290);
nand U8667 (N_8667,N_5102,N_3079);
nor U8668 (N_8668,N_4918,N_5799);
nand U8669 (N_8669,N_3974,N_3961);
nor U8670 (N_8670,N_3830,N_4082);
nand U8671 (N_8671,N_4071,N_3236);
and U8672 (N_8672,N_5790,N_5408);
and U8673 (N_8673,N_5317,N_5762);
nand U8674 (N_8674,N_5637,N_5047);
nor U8675 (N_8675,N_4413,N_4072);
and U8676 (N_8676,N_3442,N_3757);
and U8677 (N_8677,N_4338,N_5689);
nand U8678 (N_8678,N_3863,N_5044);
or U8679 (N_8679,N_5626,N_4303);
nor U8680 (N_8680,N_4157,N_3450);
or U8681 (N_8681,N_5966,N_3765);
nor U8682 (N_8682,N_3192,N_5553);
nand U8683 (N_8683,N_5630,N_3205);
nor U8684 (N_8684,N_5103,N_4381);
nand U8685 (N_8685,N_5511,N_4671);
and U8686 (N_8686,N_4849,N_5538);
or U8687 (N_8687,N_3379,N_5253);
nand U8688 (N_8688,N_5393,N_3309);
or U8689 (N_8689,N_4638,N_4747);
nor U8690 (N_8690,N_4511,N_3023);
and U8691 (N_8691,N_4564,N_4886);
nand U8692 (N_8692,N_3542,N_3020);
or U8693 (N_8693,N_5224,N_4894);
or U8694 (N_8694,N_3839,N_5622);
nor U8695 (N_8695,N_4676,N_3479);
nor U8696 (N_8696,N_3510,N_3081);
nor U8697 (N_8697,N_3646,N_4485);
and U8698 (N_8698,N_3964,N_4284);
nand U8699 (N_8699,N_5088,N_5537);
nor U8700 (N_8700,N_3833,N_4594);
or U8701 (N_8701,N_4728,N_5977);
and U8702 (N_8702,N_4484,N_3550);
nand U8703 (N_8703,N_4686,N_3230);
and U8704 (N_8704,N_3827,N_3866);
nor U8705 (N_8705,N_3324,N_3578);
nand U8706 (N_8706,N_4861,N_3840);
nor U8707 (N_8707,N_5340,N_5151);
or U8708 (N_8708,N_3135,N_4117);
and U8709 (N_8709,N_5050,N_5039);
nor U8710 (N_8710,N_4865,N_4473);
nor U8711 (N_8711,N_4102,N_3493);
and U8712 (N_8712,N_5202,N_3960);
nand U8713 (N_8713,N_5695,N_3169);
and U8714 (N_8714,N_4088,N_5450);
or U8715 (N_8715,N_4558,N_5963);
nand U8716 (N_8716,N_4806,N_4634);
or U8717 (N_8717,N_4938,N_3114);
or U8718 (N_8718,N_4807,N_4167);
or U8719 (N_8719,N_3772,N_4635);
nor U8720 (N_8720,N_5283,N_5903);
and U8721 (N_8721,N_5749,N_3227);
or U8722 (N_8722,N_5690,N_4084);
nand U8723 (N_8723,N_3651,N_5349);
nand U8724 (N_8724,N_3196,N_3552);
and U8725 (N_8725,N_4728,N_3863);
nor U8726 (N_8726,N_5820,N_5557);
or U8727 (N_8727,N_3731,N_5628);
and U8728 (N_8728,N_5248,N_4708);
and U8729 (N_8729,N_5457,N_3632);
and U8730 (N_8730,N_4872,N_3780);
xor U8731 (N_8731,N_3473,N_3386);
xnor U8732 (N_8732,N_4223,N_4729);
xor U8733 (N_8733,N_5672,N_3428);
or U8734 (N_8734,N_5322,N_3654);
nor U8735 (N_8735,N_3242,N_4296);
or U8736 (N_8736,N_5872,N_5267);
and U8737 (N_8737,N_3507,N_3606);
or U8738 (N_8738,N_3088,N_5088);
or U8739 (N_8739,N_4308,N_3474);
nor U8740 (N_8740,N_4849,N_5065);
nand U8741 (N_8741,N_3935,N_4488);
nor U8742 (N_8742,N_4448,N_4265);
or U8743 (N_8743,N_5067,N_3874);
nand U8744 (N_8744,N_4001,N_5114);
and U8745 (N_8745,N_4539,N_5725);
nor U8746 (N_8746,N_5630,N_4764);
or U8747 (N_8747,N_3502,N_4033);
nand U8748 (N_8748,N_5775,N_4075);
nor U8749 (N_8749,N_3430,N_3659);
nand U8750 (N_8750,N_5157,N_5491);
nand U8751 (N_8751,N_5061,N_5294);
or U8752 (N_8752,N_5785,N_4182);
or U8753 (N_8753,N_3341,N_5212);
or U8754 (N_8754,N_3084,N_3039);
and U8755 (N_8755,N_3338,N_4038);
and U8756 (N_8756,N_5916,N_4434);
and U8757 (N_8757,N_4137,N_5873);
nor U8758 (N_8758,N_5080,N_4977);
nor U8759 (N_8759,N_5656,N_3535);
or U8760 (N_8760,N_3338,N_4208);
or U8761 (N_8761,N_5305,N_4116);
or U8762 (N_8762,N_4470,N_5096);
nand U8763 (N_8763,N_3059,N_4981);
or U8764 (N_8764,N_3132,N_3780);
or U8765 (N_8765,N_5261,N_5292);
and U8766 (N_8766,N_4050,N_5683);
nor U8767 (N_8767,N_5562,N_3784);
and U8768 (N_8768,N_5133,N_5298);
nor U8769 (N_8769,N_3691,N_3814);
or U8770 (N_8770,N_4657,N_5779);
and U8771 (N_8771,N_3920,N_3090);
or U8772 (N_8772,N_3359,N_5040);
nand U8773 (N_8773,N_4797,N_4773);
or U8774 (N_8774,N_5880,N_3623);
nand U8775 (N_8775,N_4943,N_4045);
and U8776 (N_8776,N_4819,N_4987);
or U8777 (N_8777,N_5150,N_3016);
nand U8778 (N_8778,N_4729,N_3269);
and U8779 (N_8779,N_3933,N_4718);
or U8780 (N_8780,N_5428,N_3949);
nand U8781 (N_8781,N_3160,N_3047);
nor U8782 (N_8782,N_4848,N_3332);
nand U8783 (N_8783,N_3996,N_4029);
and U8784 (N_8784,N_3726,N_4864);
or U8785 (N_8785,N_3915,N_3176);
nor U8786 (N_8786,N_3176,N_3405);
and U8787 (N_8787,N_5667,N_5970);
or U8788 (N_8788,N_4622,N_4591);
and U8789 (N_8789,N_5884,N_5499);
and U8790 (N_8790,N_3362,N_3455);
or U8791 (N_8791,N_5729,N_5553);
and U8792 (N_8792,N_5028,N_3246);
and U8793 (N_8793,N_4416,N_5192);
or U8794 (N_8794,N_3224,N_3262);
and U8795 (N_8795,N_4704,N_3064);
or U8796 (N_8796,N_5470,N_4355);
nor U8797 (N_8797,N_3640,N_5830);
nor U8798 (N_8798,N_4233,N_5160);
and U8799 (N_8799,N_5900,N_3513);
or U8800 (N_8800,N_4260,N_4919);
or U8801 (N_8801,N_3760,N_5287);
nand U8802 (N_8802,N_4538,N_4742);
and U8803 (N_8803,N_3585,N_3430);
and U8804 (N_8804,N_5317,N_5841);
nand U8805 (N_8805,N_3350,N_3429);
or U8806 (N_8806,N_3373,N_5486);
nor U8807 (N_8807,N_5880,N_3173);
nor U8808 (N_8808,N_3277,N_3942);
and U8809 (N_8809,N_3936,N_3758);
and U8810 (N_8810,N_3954,N_5504);
nand U8811 (N_8811,N_5035,N_4438);
and U8812 (N_8812,N_4935,N_4194);
and U8813 (N_8813,N_3916,N_3017);
nor U8814 (N_8814,N_4431,N_3030);
and U8815 (N_8815,N_4795,N_5362);
nor U8816 (N_8816,N_3668,N_3178);
nor U8817 (N_8817,N_3294,N_4045);
or U8818 (N_8818,N_4794,N_4059);
nor U8819 (N_8819,N_4667,N_5515);
and U8820 (N_8820,N_5402,N_5816);
or U8821 (N_8821,N_5581,N_3910);
nand U8822 (N_8822,N_4443,N_3581);
or U8823 (N_8823,N_3251,N_3819);
or U8824 (N_8824,N_4608,N_3045);
nor U8825 (N_8825,N_4141,N_4005);
nor U8826 (N_8826,N_3280,N_4443);
or U8827 (N_8827,N_3534,N_4325);
nand U8828 (N_8828,N_4274,N_3201);
nor U8829 (N_8829,N_5696,N_3415);
nand U8830 (N_8830,N_5342,N_4886);
or U8831 (N_8831,N_4259,N_5419);
nor U8832 (N_8832,N_4240,N_4349);
and U8833 (N_8833,N_4686,N_5180);
nor U8834 (N_8834,N_3099,N_3345);
or U8835 (N_8835,N_3067,N_4699);
nor U8836 (N_8836,N_4213,N_4940);
nor U8837 (N_8837,N_4551,N_4969);
nand U8838 (N_8838,N_5198,N_4248);
nor U8839 (N_8839,N_4194,N_3792);
nor U8840 (N_8840,N_4485,N_4619);
or U8841 (N_8841,N_4268,N_4465);
or U8842 (N_8842,N_3537,N_5196);
nand U8843 (N_8843,N_5641,N_4820);
nand U8844 (N_8844,N_3428,N_3728);
and U8845 (N_8845,N_4130,N_4401);
or U8846 (N_8846,N_4350,N_5614);
nor U8847 (N_8847,N_5466,N_3058);
nor U8848 (N_8848,N_4492,N_5724);
nand U8849 (N_8849,N_5373,N_5525);
or U8850 (N_8850,N_3845,N_3345);
nor U8851 (N_8851,N_3383,N_3357);
nor U8852 (N_8852,N_3055,N_4167);
or U8853 (N_8853,N_4036,N_5375);
or U8854 (N_8854,N_4529,N_3628);
nor U8855 (N_8855,N_3720,N_4187);
or U8856 (N_8856,N_4479,N_5988);
nand U8857 (N_8857,N_5772,N_3024);
and U8858 (N_8858,N_3313,N_4356);
or U8859 (N_8859,N_4871,N_5276);
or U8860 (N_8860,N_4391,N_3581);
and U8861 (N_8861,N_4201,N_4806);
xor U8862 (N_8862,N_3089,N_4078);
and U8863 (N_8863,N_3292,N_4841);
and U8864 (N_8864,N_3578,N_3698);
nand U8865 (N_8865,N_4877,N_3717);
nand U8866 (N_8866,N_3416,N_4863);
nand U8867 (N_8867,N_3551,N_5996);
and U8868 (N_8868,N_5304,N_5678);
and U8869 (N_8869,N_5317,N_5898);
or U8870 (N_8870,N_4936,N_3817);
nand U8871 (N_8871,N_3894,N_4757);
nor U8872 (N_8872,N_5445,N_5604);
and U8873 (N_8873,N_3938,N_3054);
and U8874 (N_8874,N_3287,N_3736);
nand U8875 (N_8875,N_4477,N_4022);
and U8876 (N_8876,N_5497,N_4929);
nand U8877 (N_8877,N_3437,N_5191);
nand U8878 (N_8878,N_5148,N_3683);
nand U8879 (N_8879,N_3215,N_3074);
nand U8880 (N_8880,N_3423,N_3864);
nor U8881 (N_8881,N_4613,N_4041);
and U8882 (N_8882,N_5806,N_3404);
nor U8883 (N_8883,N_4605,N_5959);
xnor U8884 (N_8884,N_3068,N_4183);
and U8885 (N_8885,N_5484,N_5829);
or U8886 (N_8886,N_3865,N_5028);
nand U8887 (N_8887,N_3630,N_5346);
and U8888 (N_8888,N_3287,N_5647);
nor U8889 (N_8889,N_3669,N_3270);
and U8890 (N_8890,N_3416,N_5442);
nand U8891 (N_8891,N_4448,N_5746);
and U8892 (N_8892,N_5133,N_5851);
and U8893 (N_8893,N_5015,N_4782);
nand U8894 (N_8894,N_3639,N_3293);
nand U8895 (N_8895,N_3107,N_4990);
or U8896 (N_8896,N_5720,N_3583);
nor U8897 (N_8897,N_3922,N_5070);
and U8898 (N_8898,N_3026,N_3382);
or U8899 (N_8899,N_5679,N_4803);
nand U8900 (N_8900,N_4254,N_4299);
nand U8901 (N_8901,N_3910,N_5673);
nand U8902 (N_8902,N_4674,N_4599);
and U8903 (N_8903,N_3851,N_3834);
nor U8904 (N_8904,N_3065,N_3967);
nand U8905 (N_8905,N_3988,N_3112);
nand U8906 (N_8906,N_5361,N_5547);
nor U8907 (N_8907,N_5567,N_4524);
nor U8908 (N_8908,N_3435,N_3750);
and U8909 (N_8909,N_3480,N_3677);
nand U8910 (N_8910,N_5344,N_5510);
nor U8911 (N_8911,N_4845,N_3483);
nand U8912 (N_8912,N_5560,N_5595);
and U8913 (N_8913,N_3840,N_4329);
nor U8914 (N_8914,N_5202,N_4465);
nor U8915 (N_8915,N_4791,N_4743);
nor U8916 (N_8916,N_5905,N_5650);
nor U8917 (N_8917,N_4110,N_4118);
nand U8918 (N_8918,N_4339,N_5560);
and U8919 (N_8919,N_4820,N_5603);
nor U8920 (N_8920,N_4814,N_3947);
nor U8921 (N_8921,N_5675,N_5763);
or U8922 (N_8922,N_5586,N_5628);
and U8923 (N_8923,N_3397,N_5805);
or U8924 (N_8924,N_5348,N_3324);
nor U8925 (N_8925,N_5854,N_4940);
or U8926 (N_8926,N_5739,N_4076);
nor U8927 (N_8927,N_5566,N_5981);
nand U8928 (N_8928,N_3007,N_3998);
nor U8929 (N_8929,N_3695,N_4684);
nand U8930 (N_8930,N_3995,N_4478);
nand U8931 (N_8931,N_3917,N_5495);
and U8932 (N_8932,N_5760,N_5274);
nand U8933 (N_8933,N_3741,N_4341);
nand U8934 (N_8934,N_5560,N_5240);
and U8935 (N_8935,N_5459,N_3786);
nand U8936 (N_8936,N_3622,N_4149);
or U8937 (N_8937,N_3136,N_4512);
and U8938 (N_8938,N_4319,N_3403);
and U8939 (N_8939,N_4437,N_5266);
and U8940 (N_8940,N_4911,N_5044);
or U8941 (N_8941,N_3741,N_5075);
nand U8942 (N_8942,N_5817,N_5974);
nand U8943 (N_8943,N_3964,N_5309);
nor U8944 (N_8944,N_3559,N_4730);
nor U8945 (N_8945,N_5571,N_4214);
nor U8946 (N_8946,N_3485,N_3820);
or U8947 (N_8947,N_3706,N_4237);
nand U8948 (N_8948,N_5661,N_5415);
nand U8949 (N_8949,N_3635,N_4231);
xor U8950 (N_8950,N_4437,N_4325);
or U8951 (N_8951,N_3916,N_4552);
nor U8952 (N_8952,N_4333,N_4448);
or U8953 (N_8953,N_3105,N_5744);
nand U8954 (N_8954,N_5447,N_3022);
nand U8955 (N_8955,N_4985,N_5559);
and U8956 (N_8956,N_3794,N_5280);
and U8957 (N_8957,N_4874,N_3105);
nand U8958 (N_8958,N_4480,N_3357);
or U8959 (N_8959,N_4947,N_4710);
and U8960 (N_8960,N_4807,N_5741);
and U8961 (N_8961,N_4653,N_4821);
and U8962 (N_8962,N_4234,N_5224);
nand U8963 (N_8963,N_4158,N_3903);
nand U8964 (N_8964,N_4593,N_5400);
nand U8965 (N_8965,N_3113,N_3195);
and U8966 (N_8966,N_3804,N_5878);
nor U8967 (N_8967,N_3113,N_3144);
nand U8968 (N_8968,N_3115,N_3934);
or U8969 (N_8969,N_5468,N_3251);
and U8970 (N_8970,N_3634,N_5845);
nor U8971 (N_8971,N_5689,N_3812);
nor U8972 (N_8972,N_5146,N_3651);
nor U8973 (N_8973,N_3603,N_4811);
nand U8974 (N_8974,N_3363,N_5855);
and U8975 (N_8975,N_4842,N_4729);
or U8976 (N_8976,N_3336,N_3525);
and U8977 (N_8977,N_4106,N_5210);
nor U8978 (N_8978,N_5927,N_4282);
and U8979 (N_8979,N_4484,N_4249);
and U8980 (N_8980,N_4483,N_3129);
and U8981 (N_8981,N_3509,N_5673);
nand U8982 (N_8982,N_4417,N_3085);
nor U8983 (N_8983,N_3262,N_4894);
nand U8984 (N_8984,N_4002,N_5776);
or U8985 (N_8985,N_4882,N_3548);
nor U8986 (N_8986,N_3898,N_4997);
nand U8987 (N_8987,N_3358,N_3504);
or U8988 (N_8988,N_5977,N_4799);
nand U8989 (N_8989,N_5877,N_4060);
nand U8990 (N_8990,N_5275,N_3632);
or U8991 (N_8991,N_4447,N_3076);
nand U8992 (N_8992,N_3672,N_4713);
and U8993 (N_8993,N_3684,N_5007);
nand U8994 (N_8994,N_3408,N_4882);
or U8995 (N_8995,N_5394,N_3449);
nor U8996 (N_8996,N_3742,N_5353);
nand U8997 (N_8997,N_3968,N_4973);
nor U8998 (N_8998,N_4741,N_4780);
nor U8999 (N_8999,N_5694,N_4317);
or U9000 (N_9000,N_8301,N_8452);
or U9001 (N_9001,N_7857,N_7191);
or U9002 (N_9002,N_6462,N_6585);
nor U9003 (N_9003,N_8095,N_7248);
nand U9004 (N_9004,N_8345,N_6946);
or U9005 (N_9005,N_8417,N_7873);
and U9006 (N_9006,N_6651,N_6716);
and U9007 (N_9007,N_8473,N_7382);
nand U9008 (N_9008,N_6980,N_6380);
nor U9009 (N_9009,N_7696,N_7299);
or U9010 (N_9010,N_8629,N_7179);
or U9011 (N_9011,N_7917,N_6315);
nand U9012 (N_9012,N_6618,N_7199);
nand U9013 (N_9013,N_7748,N_8216);
nor U9014 (N_9014,N_7300,N_8268);
or U9015 (N_9015,N_8371,N_7358);
or U9016 (N_9016,N_7131,N_6898);
or U9017 (N_9017,N_8506,N_7979);
nor U9018 (N_9018,N_7818,N_7619);
nand U9019 (N_9019,N_8315,N_8894);
nand U9020 (N_9020,N_6525,N_8622);
nand U9021 (N_9021,N_7853,N_6699);
nand U9022 (N_9022,N_6105,N_8702);
and U9023 (N_9023,N_6912,N_8669);
nor U9024 (N_9024,N_6993,N_6026);
nor U9025 (N_9025,N_8842,N_6162);
or U9026 (N_9026,N_8377,N_8246);
nand U9027 (N_9027,N_7942,N_8289);
nor U9028 (N_9028,N_8500,N_8888);
nand U9029 (N_9029,N_7760,N_8010);
nand U9030 (N_9030,N_6337,N_6413);
nor U9031 (N_9031,N_7690,N_8620);
nand U9032 (N_9032,N_8633,N_6244);
nor U9033 (N_9033,N_7269,N_7765);
and U9034 (N_9034,N_7871,N_7812);
and U9035 (N_9035,N_7801,N_8775);
nor U9036 (N_9036,N_8762,N_7699);
nand U9037 (N_9037,N_8146,N_6101);
or U9038 (N_9038,N_6919,N_7065);
nand U9039 (N_9039,N_7270,N_6705);
or U9040 (N_9040,N_7354,N_8140);
or U9041 (N_9041,N_8038,N_7557);
nand U9042 (N_9042,N_7249,N_8687);
nor U9043 (N_9043,N_6146,N_8061);
nand U9044 (N_9044,N_8237,N_8162);
nor U9045 (N_9045,N_8919,N_6369);
or U9046 (N_9046,N_8461,N_7414);
and U9047 (N_9047,N_8256,N_6995);
and U9048 (N_9048,N_6990,N_6886);
or U9049 (N_9049,N_6043,N_6550);
and U9050 (N_9050,N_6098,N_8652);
nor U9051 (N_9051,N_7866,N_6677);
or U9052 (N_9052,N_8899,N_6269);
or U9053 (N_9053,N_8437,N_6516);
and U9054 (N_9054,N_6675,N_8610);
nor U9055 (N_9055,N_6108,N_7044);
nor U9056 (N_9056,N_6356,N_8576);
nand U9057 (N_9057,N_8259,N_8456);
and U9058 (N_9058,N_8395,N_6349);
nor U9059 (N_9059,N_7473,N_8589);
and U9060 (N_9060,N_7291,N_6834);
and U9061 (N_9061,N_7701,N_8340);
nor U9062 (N_9062,N_7892,N_7413);
and U9063 (N_9063,N_8243,N_8333);
nand U9064 (N_9064,N_7355,N_8644);
nor U9065 (N_9065,N_8878,N_8201);
nor U9066 (N_9066,N_6727,N_7235);
nand U9067 (N_9067,N_6933,N_7284);
nand U9068 (N_9068,N_7626,N_6346);
nor U9069 (N_9069,N_6156,N_7539);
nor U9070 (N_9070,N_6366,N_7273);
or U9071 (N_9071,N_8580,N_6936);
or U9072 (N_9072,N_7947,N_7729);
nand U9073 (N_9073,N_6647,N_6323);
or U9074 (N_9074,N_8968,N_7884);
and U9075 (N_9075,N_8106,N_8877);
or U9076 (N_9076,N_8701,N_6505);
nor U9077 (N_9077,N_8936,N_6720);
and U9078 (N_9078,N_6318,N_8334);
and U9079 (N_9079,N_8360,N_8659);
or U9080 (N_9080,N_6560,N_6010);
nand U9081 (N_9081,N_8169,N_6908);
nand U9082 (N_9082,N_8786,N_6594);
nor U9083 (N_9083,N_6818,N_8002);
nor U9084 (N_9084,N_7608,N_7802);
or U9085 (N_9085,N_6351,N_6648);
nor U9086 (N_9086,N_6313,N_7566);
or U9087 (N_9087,N_8895,N_8076);
nand U9088 (N_9088,N_7776,N_6592);
nor U9089 (N_9089,N_8611,N_8553);
or U9090 (N_9090,N_7939,N_6778);
nor U9091 (N_9091,N_6041,N_8770);
or U9092 (N_9092,N_6330,N_7813);
or U9093 (N_9093,N_8047,N_8678);
and U9094 (N_9094,N_7037,N_6111);
nor U9095 (N_9095,N_7401,N_8616);
nor U9096 (N_9096,N_6000,N_6379);
and U9097 (N_9097,N_7773,N_6093);
nor U9098 (N_9098,N_7604,N_6414);
nand U9099 (N_9099,N_6674,N_7767);
or U9100 (N_9100,N_8107,N_6023);
nand U9101 (N_9101,N_8472,N_6407);
or U9102 (N_9102,N_8781,N_8517);
and U9103 (N_9103,N_7797,N_7987);
and U9104 (N_9104,N_8865,N_8828);
nor U9105 (N_9105,N_7181,N_6521);
and U9106 (N_9106,N_7847,N_7999);
and U9107 (N_9107,N_7005,N_7930);
nand U9108 (N_9108,N_7313,N_7811);
nor U9109 (N_9109,N_8675,N_8866);
or U9110 (N_9110,N_6861,N_7250);
nand U9111 (N_9111,N_6166,N_7303);
nand U9112 (N_9112,N_8411,N_7097);
nor U9113 (N_9113,N_6582,N_7558);
and U9114 (N_9114,N_6080,N_6728);
or U9115 (N_9115,N_6416,N_7860);
nand U9116 (N_9116,N_8011,N_8640);
or U9117 (N_9117,N_7334,N_6203);
nor U9118 (N_9118,N_6611,N_6391);
nand U9119 (N_9119,N_6520,N_6220);
nand U9120 (N_9120,N_7470,N_7571);
or U9121 (N_9121,N_6737,N_6623);
nand U9122 (N_9122,N_8392,N_6446);
nor U9123 (N_9123,N_7443,N_6374);
nand U9124 (N_9124,N_8822,N_8588);
nand U9125 (N_9125,N_8292,N_6045);
and U9126 (N_9126,N_8338,N_6364);
and U9127 (N_9127,N_6562,N_6254);
or U9128 (N_9128,N_7200,N_8223);
or U9129 (N_9129,N_7777,N_6642);
nand U9130 (N_9130,N_6875,N_7074);
and U9131 (N_9131,N_6548,N_8367);
or U9132 (N_9132,N_8432,N_8440);
nand U9133 (N_9133,N_6841,N_7996);
nor U9134 (N_9134,N_7563,N_8348);
nor U9135 (N_9135,N_7839,N_8030);
nand U9136 (N_9136,N_8829,N_6665);
nor U9137 (N_9137,N_8721,N_7896);
nor U9138 (N_9138,N_8302,N_8487);
and U9139 (N_9139,N_8914,N_8141);
nand U9140 (N_9140,N_8881,N_7075);
xnor U9141 (N_9141,N_6989,N_7721);
or U9142 (N_9142,N_8695,N_6773);
nor U9143 (N_9143,N_7038,N_6281);
and U9144 (N_9144,N_6290,N_6267);
or U9145 (N_9145,N_6653,N_8833);
and U9146 (N_9146,N_6533,N_7895);
nand U9147 (N_9147,N_8189,N_8904);
nand U9148 (N_9148,N_7057,N_8855);
or U9149 (N_9149,N_6634,N_7011);
nor U9150 (N_9150,N_7416,N_8564);
or U9151 (N_9151,N_6478,N_6873);
nor U9152 (N_9152,N_7345,N_7309);
and U9153 (N_9153,N_8118,N_6866);
nor U9154 (N_9154,N_8160,N_7444);
nand U9155 (N_9155,N_6113,N_8072);
or U9156 (N_9156,N_6803,N_7157);
or U9157 (N_9157,N_8778,N_8493);
nand U9158 (N_9158,N_7310,N_8510);
and U9159 (N_9159,N_7140,N_8849);
nand U9160 (N_9160,N_7955,N_8804);
or U9161 (N_9161,N_7295,N_6388);
nand U9162 (N_9162,N_7020,N_8998);
and U9163 (N_9163,N_6030,N_8668);
nor U9164 (N_9164,N_7753,N_6325);
or U9165 (N_9165,N_7043,N_8747);
nand U9166 (N_9166,N_6524,N_7676);
and U9167 (N_9167,N_8327,N_7500);
nand U9168 (N_9168,N_8089,N_7596);
or U9169 (N_9169,N_8884,N_6020);
nor U9170 (N_9170,N_6445,N_8671);
nor U9171 (N_9171,N_8399,N_7610);
nand U9172 (N_9172,N_8516,N_6810);
nor U9173 (N_9173,N_8502,N_6401);
or U9174 (N_9174,N_6477,N_7185);
or U9175 (N_9175,N_8730,N_8000);
and U9176 (N_9176,N_7297,N_8518);
or U9177 (N_9177,N_7953,N_7228);
nand U9178 (N_9178,N_7646,N_8606);
nand U9179 (N_9179,N_6174,N_7899);
nand U9180 (N_9180,N_7377,N_8422);
and U9181 (N_9181,N_8260,N_7808);
nor U9182 (N_9182,N_8304,N_6792);
or U9183 (N_9183,N_7513,N_7920);
and U9184 (N_9184,N_8347,N_6876);
nor U9185 (N_9185,N_7872,N_7318);
or U9186 (N_9186,N_7775,N_6535);
or U9187 (N_9187,N_6495,N_6259);
nand U9188 (N_9188,N_6321,N_8492);
nor U9189 (N_9189,N_7287,N_7417);
nand U9190 (N_9190,N_7991,N_6539);
and U9191 (N_9191,N_7912,N_7536);
or U9192 (N_9192,N_7360,N_6055);
nand U9193 (N_9193,N_6126,N_8218);
or U9194 (N_9194,N_7886,N_6037);
nor U9195 (N_9195,N_6285,N_8803);
nand U9196 (N_9196,N_7576,N_6785);
and U9197 (N_9197,N_7176,N_8264);
nor U9198 (N_9198,N_8841,N_8285);
nor U9199 (N_9199,N_7010,N_7496);
and U9200 (N_9200,N_7363,N_7954);
nand U9201 (N_9201,N_6581,N_7386);
and U9202 (N_9202,N_6280,N_7552);
and U9203 (N_9203,N_6250,N_8320);
nand U9204 (N_9204,N_8635,N_8966);
nand U9205 (N_9205,N_8646,N_8688);
or U9206 (N_9206,N_7819,N_8079);
and U9207 (N_9207,N_6722,N_6942);
nand U9208 (N_9208,N_7509,N_6887);
or U9209 (N_9209,N_7754,N_8390);
or U9210 (N_9210,N_7915,N_8749);
or U9211 (N_9211,N_6129,N_6862);
nand U9212 (N_9212,N_6421,N_8382);
nand U9213 (N_9213,N_6506,N_7072);
nand U9214 (N_9214,N_7630,N_7829);
nand U9215 (N_9215,N_8810,N_6572);
or U9216 (N_9216,N_7901,N_7550);
or U9217 (N_9217,N_6344,N_6249);
nand U9218 (N_9218,N_8044,N_7830);
or U9219 (N_9219,N_8806,N_6965);
or U9220 (N_9220,N_8240,N_7451);
and U9221 (N_9221,N_7590,N_7961);
nand U9222 (N_9222,N_8293,N_8125);
xnor U9223 (N_9223,N_8273,N_7675);
or U9224 (N_9224,N_8167,N_7832);
nor U9225 (N_9225,N_7547,N_8637);
or U9226 (N_9226,N_7893,N_7631);
nand U9227 (N_9227,N_6226,N_6317);
nand U9228 (N_9228,N_8159,N_8134);
nand U9229 (N_9229,N_6135,N_6089);
nor U9230 (N_9230,N_8607,N_6694);
nand U9231 (N_9231,N_6133,N_7421);
nand U9232 (N_9232,N_7101,N_8941);
and U9233 (N_9233,N_7929,N_8761);
or U9234 (N_9234,N_6595,N_7361);
nand U9235 (N_9235,N_6956,N_8288);
nand U9236 (N_9236,N_8060,N_6002);
and U9237 (N_9237,N_8186,N_8976);
or U9238 (N_9238,N_8631,N_7335);
and U9239 (N_9239,N_6381,N_7396);
nor U9240 (N_9240,N_8501,N_6710);
or U9241 (N_9241,N_6179,N_7843);
or U9242 (N_9242,N_7528,N_6920);
nand U9243 (N_9243,N_8183,N_6409);
nand U9244 (N_9244,N_6408,N_7257);
nor U9245 (N_9245,N_7183,N_7123);
and U9246 (N_9246,N_8766,N_7628);
nand U9247 (N_9247,N_6760,N_6776);
xnor U9248 (N_9248,N_8485,N_8253);
and U9249 (N_9249,N_7491,N_8950);
and U9250 (N_9250,N_6540,N_8997);
nor U9251 (N_9251,N_8051,N_8021);
nand U9252 (N_9252,N_8867,N_7804);
nand U9253 (N_9253,N_7856,N_8241);
and U9254 (N_9254,N_8312,N_8498);
and U9255 (N_9255,N_8341,N_6609);
or U9256 (N_9256,N_7711,N_6922);
nand U9257 (N_9257,N_6260,N_7218);
nand U9258 (N_9258,N_6114,N_7054);
nor U9259 (N_9259,N_8691,N_8729);
or U9260 (N_9260,N_7007,N_7095);
or U9261 (N_9261,N_7809,N_8715);
nand U9262 (N_9262,N_6470,N_7651);
and U9263 (N_9263,N_6221,N_7837);
or U9264 (N_9264,N_8918,N_8109);
nand U9265 (N_9265,N_8636,N_7454);
and U9266 (N_9266,N_7616,N_8322);
nand U9267 (N_9267,N_6498,N_8336);
or U9268 (N_9268,N_8959,N_8540);
nand U9269 (N_9269,N_7261,N_6522);
and U9270 (N_9270,N_6650,N_7375);
or U9271 (N_9271,N_7092,N_8057);
xor U9272 (N_9272,N_6513,N_6452);
nand U9273 (N_9273,N_8660,N_8156);
nand U9274 (N_9274,N_8880,N_8429);
nor U9275 (N_9275,N_6970,N_8228);
nand U9276 (N_9276,N_8433,N_6112);
or U9277 (N_9277,N_7861,N_8284);
nand U9278 (N_9278,N_8590,N_7120);
or U9279 (N_9279,N_6177,N_7378);
or U9280 (N_9280,N_8554,N_7112);
nor U9281 (N_9281,N_7073,N_8670);
nor U9282 (N_9282,N_7784,N_7436);
or U9283 (N_9283,N_7679,N_6011);
and U9284 (N_9284,N_6211,N_6399);
and U9285 (N_9285,N_7541,N_7677);
or U9286 (N_9286,N_8446,N_8266);
and U9287 (N_9287,N_6499,N_6868);
and U9288 (N_9288,N_8490,N_7125);
and U9289 (N_9289,N_6935,N_7420);
or U9290 (N_9290,N_8605,N_8062);
and U9291 (N_9291,N_6631,N_7122);
nor U9292 (N_9292,N_8555,N_6729);
nor U9293 (N_9293,N_8591,N_6939);
or U9294 (N_9294,N_7602,N_6361);
and U9295 (N_9295,N_6555,N_8978);
and U9296 (N_9296,N_7133,N_8848);
or U9297 (N_9297,N_6237,N_6863);
and U9298 (N_9298,N_8296,N_8545);
and U9299 (N_9299,N_8113,N_8132);
and U9300 (N_9300,N_6613,N_6219);
and U9301 (N_9301,N_7343,N_6941);
nand U9302 (N_9302,N_7973,N_6423);
nand U9303 (N_9303,N_7068,N_7669);
or U9304 (N_9304,N_8108,N_6756);
nand U9305 (N_9305,N_8984,N_8386);
and U9306 (N_9306,N_8722,N_6894);
and U9307 (N_9307,N_8650,N_7408);
nor U9308 (N_9308,N_6823,N_6116);
and U9309 (N_9309,N_6475,N_7988);
and U9310 (N_9310,N_8584,N_8835);
nor U9311 (N_9311,N_7707,N_7222);
or U9312 (N_9312,N_7495,N_7494);
nand U9313 (N_9313,N_7186,N_7277);
and U9314 (N_9314,N_6564,N_8898);
nand U9315 (N_9315,N_8357,N_7722);
nor U9316 (N_9316,N_7168,N_8704);
and U9317 (N_9317,N_7138,N_7689);
nor U9318 (N_9318,N_6947,N_6487);
nor U9319 (N_9319,N_6489,N_6807);
or U9320 (N_9320,N_8102,N_8346);
nand U9321 (N_9321,N_7993,N_6441);
nor U9322 (N_9322,N_7772,N_8585);
nor U9323 (N_9323,N_8641,N_6718);
nand U9324 (N_9324,N_6025,N_6316);
nand U9325 (N_9325,N_8211,N_7152);
nor U9326 (N_9326,N_7709,N_6557);
nand U9327 (N_9327,N_8449,N_6804);
or U9328 (N_9328,N_7803,N_7134);
and U9329 (N_9329,N_6725,N_8040);
nor U9330 (N_9330,N_7145,N_7527);
or U9331 (N_9331,N_7461,N_6012);
nor U9332 (N_9332,N_6256,N_8155);
and U9333 (N_9333,N_8020,N_8627);
and U9334 (N_9334,N_8619,N_7650);
and U9335 (N_9335,N_6552,N_8931);
nand U9336 (N_9336,N_6273,N_6230);
nor U9337 (N_9337,N_6232,N_7844);
or U9338 (N_9338,N_6436,N_8909);
nor U9339 (N_9339,N_7990,N_6405);
nor U9340 (N_9340,N_8519,N_6734);
or U9341 (N_9341,N_7022,N_7487);
nor U9342 (N_9342,N_8582,N_8488);
nor U9343 (N_9343,N_7742,N_7735);
nor U9344 (N_9344,N_7219,N_6295);
xnor U9345 (N_9345,N_7202,N_6537);
nor U9346 (N_9346,N_6668,N_6235);
and U9347 (N_9347,N_7763,N_8401);
nand U9348 (N_9348,N_7237,N_8892);
nor U9349 (N_9349,N_6197,N_7166);
and U9350 (N_9350,N_7066,N_7644);
nor U9351 (N_9351,N_7919,N_8406);
and U9352 (N_9352,N_8496,N_7366);
nor U9353 (N_9353,N_8489,N_8009);
nor U9354 (N_9354,N_6530,N_8421);
or U9355 (N_9355,N_8317,N_6578);
nand U9356 (N_9356,N_8066,N_8311);
nor U9357 (N_9357,N_7666,N_8850);
nor U9358 (N_9358,N_6526,N_7967);
nor U9359 (N_9359,N_6629,N_8073);
nand U9360 (N_9360,N_8734,N_7210);
nor U9361 (N_9361,N_6385,N_8269);
nor U9362 (N_9362,N_7150,N_7595);
or U9363 (N_9363,N_6271,N_8407);
nand U9364 (N_9364,N_8732,N_7964);
xor U9365 (N_9365,N_8091,N_8475);
nor U9366 (N_9366,N_6345,N_8235);
nor U9367 (N_9367,N_7041,N_6107);
nand U9368 (N_9368,N_7067,N_6155);
nand U9369 (N_9369,N_7908,N_7732);
nor U9370 (N_9370,N_7474,N_6590);
and U9371 (N_9371,N_6851,N_6044);
nand U9372 (N_9372,N_6144,N_6967);
and U9373 (N_9373,N_7614,N_6897);
nor U9374 (N_9374,N_6556,N_7681);
or U9375 (N_9375,N_7958,N_7922);
or U9376 (N_9376,N_7718,N_7293);
nand U9377 (N_9377,N_6063,N_7174);
nand U9378 (N_9378,N_8710,N_6865);
nand U9379 (N_9379,N_8552,N_6453);
nand U9380 (N_9380,N_8335,N_8932);
nor U9381 (N_9381,N_6263,N_6902);
or U9382 (N_9382,N_8905,N_7759);
and U9383 (N_9383,N_6895,N_8165);
or U9384 (N_9384,N_6683,N_8686);
nand U9385 (N_9385,N_7121,N_8250);
and U9386 (N_9386,N_6333,N_7523);
nor U9387 (N_9387,N_7082,N_6504);
or U9388 (N_9388,N_7537,N_8275);
nor U9389 (N_9389,N_8960,N_6422);
or U9390 (N_9390,N_6264,N_6850);
or U9391 (N_9391,N_8801,N_8546);
nand U9392 (N_9392,N_7726,N_6471);
nor U9393 (N_9393,N_7684,N_6950);
and U9394 (N_9394,N_7466,N_6047);
or U9395 (N_9395,N_7560,N_6960);
or U9396 (N_9396,N_6066,N_7221);
nor U9397 (N_9397,N_6547,N_8426);
nand U9398 (N_9398,N_7464,N_6322);
nand U9399 (N_9399,N_7731,N_8025);
and U9400 (N_9400,N_8001,N_7647);
nor U9401 (N_9401,N_8768,N_8059);
and U9402 (N_9402,N_7457,N_8916);
and U9403 (N_9403,N_8839,N_8019);
nand U9404 (N_9404,N_7836,N_6899);
nor U9405 (N_9405,N_8436,N_6529);
or U9406 (N_9406,N_7822,N_6809);
nand U9407 (N_9407,N_8098,N_6128);
and U9408 (N_9408,N_6619,N_6884);
nor U9409 (N_9409,N_8054,N_8906);
nand U9410 (N_9410,N_8365,N_8511);
nand U9411 (N_9411,N_8874,N_6064);
and U9412 (N_9412,N_7260,N_8719);
and U9413 (N_9413,N_6222,N_8043);
nand U9414 (N_9414,N_8035,N_6469);
and U9415 (N_9415,N_8813,N_6309);
nand U9416 (N_9416,N_8093,N_6549);
and U9417 (N_9417,N_8832,N_7910);
nand U9418 (N_9418,N_6509,N_7409);
nor U9419 (N_9419,N_8225,N_7438);
nor U9420 (N_9420,N_7551,N_8114);
nor U9421 (N_9421,N_6510,N_8415);
nor U9422 (N_9422,N_7136,N_6885);
nor U9423 (N_9423,N_8128,N_7555);
nand U9424 (N_9424,N_6743,N_6343);
nor U9425 (N_9425,N_7924,N_8369);
nor U9426 (N_9426,N_7490,N_6274);
and U9427 (N_9427,N_6764,N_8547);
or U9428 (N_9428,N_7580,N_7637);
nand U9429 (N_9429,N_7327,N_8090);
nor U9430 (N_9430,N_6874,N_6654);
nand U9431 (N_9431,N_6352,N_7290);
nand U9432 (N_9432,N_6186,N_7518);
and U9433 (N_9433,N_7109,N_7499);
or U9434 (N_9434,N_7691,N_7880);
nand U9435 (N_9435,N_6419,N_7468);
nor U9436 (N_9436,N_8970,N_8864);
nand U9437 (N_9437,N_8767,N_8278);
and U9438 (N_9438,N_6007,N_6410);
and U9439 (N_9439,N_7139,N_8934);
nor U9440 (N_9440,N_8129,N_7959);
or U9441 (N_9441,N_6224,N_6740);
nor U9442 (N_9442,N_7662,N_6151);
or U9443 (N_9443,N_6437,N_7592);
nand U9444 (N_9444,N_6217,N_7411);
nor U9445 (N_9445,N_7493,N_7683);
or U9446 (N_9446,N_7531,N_7578);
and U9447 (N_9447,N_6953,N_7639);
nor U9448 (N_9448,N_6328,N_6104);
or U9449 (N_9449,N_6003,N_8205);
nor U9450 (N_9450,N_8824,N_7053);
nor U9451 (N_9451,N_6781,N_6958);
nor U9452 (N_9452,N_8318,N_6209);
nand U9453 (N_9453,N_8007,N_6790);
nor U9454 (N_9454,N_6234,N_8330);
nor U9455 (N_9455,N_8651,N_7437);
nor U9456 (N_9456,N_8769,N_6327);
and U9457 (N_9457,N_8818,N_8696);
nand U9458 (N_9458,N_8151,N_8823);
and U9459 (N_9459,N_7846,N_7342);
nand U9460 (N_9460,N_7562,N_7589);
nand U9461 (N_9461,N_7976,N_8736);
and U9462 (N_9462,N_6216,N_8963);
nor U9463 (N_9463,N_6977,N_6466);
nand U9464 (N_9464,N_8570,N_7745);
nand U9465 (N_9465,N_6753,N_6551);
or U9466 (N_9466,N_7027,N_7026);
nand U9467 (N_9467,N_6854,N_7577);
or U9468 (N_9468,N_8996,N_6703);
and U9469 (N_9469,N_7201,N_7340);
and U9470 (N_9470,N_7814,N_6201);
and U9471 (N_9471,N_7405,N_6424);
nor U9472 (N_9472,N_7716,N_7758);
and U9473 (N_9473,N_7175,N_8396);
or U9474 (N_9474,N_8470,N_8513);
or U9475 (N_9475,N_7061,N_8374);
or U9476 (N_9476,N_6719,N_7648);
and U9477 (N_9477,N_6392,N_8210);
nor U9478 (N_9478,N_6485,N_6614);
nor U9479 (N_9479,N_8003,N_6434);
and U9480 (N_9480,N_6279,N_6181);
nor U9481 (N_9481,N_8886,N_7278);
nor U9482 (N_9482,N_6759,N_7105);
or U9483 (N_9483,N_7586,N_7935);
nand U9484 (N_9484,N_6981,N_6971);
and U9485 (N_9485,N_7720,N_6831);
nand U9486 (N_9486,N_8331,N_6354);
nor U9487 (N_9487,N_6029,N_7806);
nor U9488 (N_9488,N_6350,N_6238);
or U9489 (N_9489,N_7661,N_7481);
or U9490 (N_9490,N_6692,N_7522);
nor U9491 (N_9491,N_8692,N_7376);
or U9492 (N_9492,N_8463,N_6120);
and U9493 (N_9493,N_7713,N_6763);
and U9494 (N_9494,N_7130,N_6680);
nor U9495 (N_9495,N_8935,N_7515);
or U9496 (N_9496,N_8940,N_6915);
or U9497 (N_9497,N_8574,N_7399);
nand U9498 (N_9498,N_6507,N_8049);
and U9499 (N_9499,N_6033,N_8703);
or U9500 (N_9500,N_7158,N_7769);
or U9501 (N_9501,N_6934,N_7505);
nand U9502 (N_9502,N_7267,N_6888);
or U9503 (N_9503,N_6893,N_7243);
and U9504 (N_9504,N_6463,N_7710);
nor U9505 (N_9505,N_8840,N_6094);
or U9506 (N_9506,N_6117,N_8466);
or U9507 (N_9507,N_8653,N_6494);
or U9508 (N_9508,N_8634,N_8939);
and U9509 (N_9509,N_8920,N_7205);
and U9510 (N_9510,N_7956,N_6869);
or U9511 (N_9511,N_8388,N_7172);
and U9512 (N_9512,N_8063,N_6660);
or U9513 (N_9513,N_6242,N_8116);
or U9514 (N_9514,N_8987,N_7282);
nand U9515 (N_9515,N_6571,N_8359);
or U9516 (N_9516,N_8977,N_7756);
nor U9517 (N_9517,N_6802,N_7632);
xor U9518 (N_9518,N_7216,N_7259);
or U9519 (N_9519,N_8682,N_6472);
nand U9520 (N_9520,N_8363,N_6534);
or U9521 (N_9521,N_8708,N_8742);
nor U9522 (N_9522,N_7909,N_6797);
nand U9523 (N_9523,N_6468,N_6298);
nor U9524 (N_9524,N_7059,N_8676);
or U9525 (N_9525,N_8927,N_8161);
or U9526 (N_9526,N_8414,N_6262);
and U9527 (N_9527,N_6567,N_8814);
nor U9528 (N_9528,N_7142,N_6481);
or U9529 (N_9529,N_8989,N_6974);
and U9530 (N_9530,N_6954,N_8529);
nor U9531 (N_9531,N_8229,N_8004);
nor U9532 (N_9532,N_7167,N_7739);
nor U9533 (N_9533,N_8845,N_6754);
or U9534 (N_9534,N_8563,N_6766);
and U9535 (N_9535,N_8131,N_8756);
nor U9536 (N_9536,N_8673,N_7271);
and U9537 (N_9537,N_6844,N_6696);
nand U9538 (N_9538,N_8725,N_6086);
nand U9539 (N_9539,N_8664,N_7159);
nand U9540 (N_9540,N_6786,N_7923);
and U9541 (N_9541,N_8716,N_8561);
nor U9542 (N_9542,N_6568,N_8297);
or U9543 (N_9543,N_8087,N_8027);
and U9544 (N_9544,N_7606,N_6929);
nand U9545 (N_9545,N_7406,N_8618);
nor U9546 (N_9546,N_6655,N_6430);
or U9547 (N_9547,N_6576,N_8022);
and U9548 (N_9548,N_8457,N_7519);
nor U9549 (N_9549,N_7102,N_7231);
and U9550 (N_9550,N_8568,N_8577);
and U9551 (N_9551,N_8967,N_8046);
or U9552 (N_9552,N_7203,N_8792);
and U9553 (N_9553,N_7826,N_8202);
and U9554 (N_9554,N_7362,N_6545);
and U9555 (N_9555,N_7565,N_8364);
or U9556 (N_9556,N_7538,N_6758);
nor U9557 (N_9557,N_6021,N_7244);
and U9558 (N_9558,N_7728,N_7317);
or U9559 (N_9559,N_6910,N_7934);
or U9560 (N_9560,N_6951,N_6656);
nand U9561 (N_9561,N_6752,N_8565);
or U9562 (N_9562,N_8053,N_8709);
and U9563 (N_9563,N_7863,N_6355);
nor U9564 (N_9564,N_8339,N_7877);
or U9565 (N_9565,N_6948,N_7864);
and U9566 (N_9566,N_7050,N_6474);
or U9567 (N_9567,N_6788,N_7835);
or U9568 (N_9568,N_8082,N_8139);
or U9569 (N_9569,N_7391,N_6907);
or U9570 (N_9570,N_7107,N_6903);
or U9571 (N_9571,N_7693,N_6768);
or U9572 (N_9572,N_6396,N_8227);
or U9573 (N_9573,N_8314,N_7501);
nand U9574 (N_9574,N_8649,N_7963);
or U9575 (N_9575,N_7768,N_6016);
or U9576 (N_9576,N_8300,N_6079);
and U9577 (N_9577,N_6577,N_8104);
nor U9578 (N_9578,N_7948,N_7636);
and U9579 (N_9579,N_8219,N_8366);
nor U9580 (N_9580,N_8424,N_7032);
or U9581 (N_9581,N_7642,N_6060);
and U9582 (N_9582,N_8790,N_6736);
nor U9583 (N_9583,N_8844,N_7793);
and U9584 (N_9584,N_7104,N_6964);
and U9585 (N_9585,N_6852,N_7352);
and U9586 (N_9586,N_6573,N_8748);
or U9587 (N_9587,N_8924,N_6730);
nor U9588 (N_9588,N_6353,N_7780);
or U9589 (N_9589,N_6652,N_6305);
and U9590 (N_9590,N_7198,N_8524);
nor U9591 (N_9591,N_8638,N_8525);
and U9592 (N_9592,N_6687,N_6372);
and U9593 (N_9593,N_6672,N_6492);
xor U9594 (N_9594,N_6048,N_8913);
or U9595 (N_9595,N_8887,N_6531);
nor U9596 (N_9596,N_8103,N_7333);
or U9597 (N_9597,N_7482,N_8763);
nor U9598 (N_9598,N_6825,N_7600);
nor U9599 (N_9599,N_8777,N_6982);
nand U9600 (N_9600,N_6214,N_6600);
or U9601 (N_9601,N_6812,N_7572);
nand U9602 (N_9602,N_6225,N_7449);
nand U9603 (N_9603,N_7276,N_6090);
or U9604 (N_9604,N_7874,N_8538);
nor U9605 (N_9605,N_7048,N_6775);
nand U9606 (N_9606,N_7674,N_8014);
or U9607 (N_9607,N_7534,N_8858);
nand U9608 (N_9608,N_8903,N_7283);
and U9609 (N_9609,N_7144,N_6180);
nand U9610 (N_9610,N_6403,N_8549);
and U9611 (N_9611,N_8600,N_7274);
and U9612 (N_9612,N_8922,N_7903);
nand U9613 (N_9613,N_6099,N_6627);
nand U9614 (N_9614,N_7926,N_7365);
nor U9615 (N_9615,N_6796,N_6544);
nand U9616 (N_9616,N_7845,N_8055);
and U9617 (N_9617,N_8680,N_6054);
or U9618 (N_9618,N_7478,N_7514);
nor U9619 (N_9619,N_7380,N_8410);
xnor U9620 (N_9620,N_7236,N_7155);
nor U9621 (N_9621,N_8071,N_6691);
or U9622 (N_9622,N_6735,N_7452);
nand U9623 (N_9623,N_6569,N_7087);
nor U9624 (N_9624,N_6957,N_6191);
and U9625 (N_9625,N_7952,N_6676);
or U9626 (N_9626,N_6076,N_7664);
or U9627 (N_9627,N_6817,N_6190);
and U9628 (N_9628,N_7217,N_7504);
and U9629 (N_9629,N_7162,N_7770);
or U9630 (N_9630,N_7370,N_8194);
or U9631 (N_9631,N_6515,N_8954);
nand U9632 (N_9632,N_7442,N_6360);
and U9633 (N_9633,N_6561,N_6943);
nand U9634 (N_9634,N_7000,N_8290);
or U9635 (N_9635,N_8232,N_8316);
nand U9636 (N_9636,N_7189,N_6639);
and U9637 (N_9637,N_7878,N_6476);
or U9638 (N_9638,N_8361,N_8667);
or U9639 (N_9639,N_7063,N_7292);
nor U9640 (N_9640,N_6726,N_7447);
nand U9641 (N_9641,N_7932,N_6169);
or U9642 (N_9642,N_7965,N_7392);
and U9643 (N_9643,N_8689,N_7727);
nand U9644 (N_9644,N_7532,N_6307);
nor U9645 (N_9645,N_8326,N_6959);
nor U9646 (N_9646,N_8875,N_8755);
nor U9647 (N_9647,N_7114,N_6832);
nand U9648 (N_9648,N_8249,N_7573);
nand U9649 (N_9649,N_8528,N_8765);
nor U9650 (N_9650,N_6966,N_8893);
and U9651 (N_9651,N_8994,N_6883);
nor U9652 (N_9652,N_8558,N_7213);
nand U9653 (N_9653,N_6389,N_8973);
nor U9654 (N_9654,N_8203,N_8562);
nor U9655 (N_9655,N_8608,N_8130);
nand U9656 (N_9656,N_7254,N_8008);
nor U9657 (N_9657,N_7981,N_6840);
nor U9658 (N_9658,N_8945,N_6877);
and U9659 (N_9659,N_8230,N_8137);
xnor U9660 (N_9660,N_6284,N_6748);
and U9661 (N_9661,N_6579,N_6387);
and U9662 (N_9662,N_7264,N_8423);
and U9663 (N_9663,N_6926,N_8930);
and U9664 (N_9664,N_8896,N_7798);
or U9665 (N_9665,N_7400,N_6664);
nand U9666 (N_9666,N_8975,N_8707);
nor U9667 (N_9667,N_7398,N_6955);
nand U9668 (N_9668,N_8609,N_6925);
nor U9669 (N_9669,N_6272,N_6163);
nor U9670 (N_9670,N_6543,N_6152);
or U9671 (N_9671,N_6574,N_6787);
nand U9672 (N_9672,N_7127,N_8482);
and U9673 (N_9673,N_6188,N_8902);
nor U9674 (N_9674,N_8809,N_6258);
or U9675 (N_9675,N_7698,N_6062);
or U9676 (N_9676,N_6923,N_6377);
or U9677 (N_9677,N_8221,N_6292);
and U9678 (N_9678,N_6164,N_7058);
nor U9679 (N_9679,N_7624,N_7663);
nand U9680 (N_9680,N_7229,N_6136);
and U9681 (N_9681,N_8827,N_6384);
nor U9682 (N_9682,N_6293,N_6398);
nor U9683 (N_9683,N_6386,N_7762);
nor U9684 (N_9684,N_8979,N_7164);
nor U9685 (N_9685,N_6227,N_7298);
or U9686 (N_9686,N_7374,N_7719);
and U9687 (N_9687,N_7972,N_8154);
nand U9688 (N_9688,N_7384,N_7385);
and U9689 (N_9689,N_8425,N_6824);
or U9690 (N_9690,N_8307,N_7099);
and U9691 (N_9691,N_8750,N_6442);
nand U9692 (N_9692,N_7906,N_6124);
or U9693 (N_9693,N_7975,N_6559);
nand U9694 (N_9694,N_6075,N_8962);
nand U9695 (N_9695,N_6334,N_6493);
or U9696 (N_9696,N_7325,N_7211);
nand U9697 (N_9697,N_7791,N_8274);
or U9698 (N_9698,N_8484,N_6833);
and U9699 (N_9699,N_8387,N_7275);
nor U9700 (N_9700,N_7089,N_7206);
nand U9701 (N_9701,N_7692,N_7882);
nand U9702 (N_9702,N_6771,N_7412);
or U9703 (N_9703,N_7062,N_6314);
nor U9704 (N_9704,N_8535,N_7842);
or U9705 (N_9705,N_8964,N_6921);
nor U9706 (N_9706,N_8384,N_7561);
or U9707 (N_9707,N_6014,N_8681);
and U9708 (N_9708,N_7194,N_7230);
and U9709 (N_9709,N_7480,N_6774);
or U9710 (N_9710,N_8006,N_7623);
nand U9711 (N_9711,N_8915,N_8586);
nand U9712 (N_9712,N_6239,N_6945);
nor U9713 (N_9713,N_7995,N_7840);
nor U9714 (N_9714,N_8404,N_7285);
or U9715 (N_9715,N_6878,N_8911);
nor U9716 (N_9716,N_7078,N_6828);
and U9717 (N_9717,N_7730,N_8291);
or U9718 (N_9718,N_6288,N_7950);
nor U9719 (N_9719,N_8873,N_8085);
and U9720 (N_9720,N_8526,N_7143);
nand U9721 (N_9721,N_6496,N_7315);
nor U9722 (N_9722,N_8075,N_6411);
or U9723 (N_9723,N_7778,N_7258);
and U9724 (N_9724,N_6265,N_7238);
nor U9725 (N_9725,N_7004,N_8551);
nand U9726 (N_9726,N_6906,N_8295);
and U9727 (N_9727,N_6022,N_7738);
and U9728 (N_9728,N_7700,N_8251);
nand U9729 (N_9729,N_6072,N_6100);
and U9730 (N_9730,N_7289,N_8891);
or U9731 (N_9731,N_8569,N_8117);
or U9732 (N_9732,N_6085,N_8907);
nor U9733 (N_9733,N_6371,N_8193);
and U9734 (N_9734,N_6448,N_7655);
nand U9735 (N_9735,N_7106,N_8207);
nand U9736 (N_9736,N_6130,N_7982);
or U9737 (N_9737,N_7914,N_6900);
or U9738 (N_9738,N_7855,N_6213);
xor U9739 (N_9739,N_6514,N_6928);
nor U9740 (N_9740,N_6808,N_7656);
or U9741 (N_9741,N_8971,N_7098);
nand U9742 (N_9742,N_7907,N_7706);
nor U9743 (N_9743,N_8153,N_6248);
nand U9744 (N_9744,N_6142,N_7321);
or U9745 (N_9745,N_8099,N_6171);
and U9746 (N_9746,N_8897,N_7171);
nor U9747 (N_9747,N_8697,N_6711);
and U9748 (N_9748,N_8148,N_7369);
and U9749 (N_9749,N_8258,N_7314);
and U9750 (N_9750,N_8744,N_8263);
and U9751 (N_9751,N_7820,N_7331);
and U9752 (N_9752,N_8069,N_7697);
nor U9753 (N_9753,N_6373,N_8949);
and U9754 (N_9754,N_7233,N_7512);
or U9755 (N_9755,N_8505,N_8509);
or U9756 (N_9756,N_7585,N_6005);
xor U9757 (N_9757,N_6765,N_7649);
nor U9758 (N_9758,N_6645,N_8621);
nor U9759 (N_9759,N_6207,N_8579);
nor U9760 (N_9760,N_7240,N_7851);
nor U9761 (N_9761,N_8349,N_7091);
and U9762 (N_9762,N_6603,N_6949);
nand U9763 (N_9763,N_6121,N_6909);
or U9764 (N_9764,N_7025,N_6836);
or U9765 (N_9765,N_6110,N_7766);
nor U9766 (N_9766,N_6431,N_6363);
or U9767 (N_9767,N_6546,N_6501);
nand U9768 (N_9768,N_6750,N_6616);
or U9769 (N_9769,N_6092,N_8376);
and U9770 (N_9770,N_8441,N_7476);
nor U9771 (N_9771,N_6731,N_6523);
nor U9772 (N_9772,N_8628,N_8133);
and U9773 (N_9773,N_7251,N_6704);
and U9774 (N_9774,N_6706,N_6641);
or U9775 (N_9775,N_8596,N_7633);
nor U9776 (N_9776,N_6202,N_6986);
or U9777 (N_9777,N_7463,N_8448);
and U9778 (N_9778,N_7774,N_8879);
and U9779 (N_9779,N_8872,N_6622);
or U9780 (N_9780,N_8726,N_7288);
or U9781 (N_9781,N_7428,N_7615);
and U9782 (N_9782,N_6517,N_6311);
or U9783 (N_9783,N_7838,N_6739);
or U9784 (N_9784,N_7749,N_6938);
nor U9785 (N_9785,N_7440,N_7553);
and U9786 (N_9786,N_7418,N_7823);
nand U9787 (N_9787,N_7262,N_6077);
nor U9788 (N_9788,N_6701,N_6053);
and U9789 (N_9789,N_7301,N_7296);
and U9790 (N_9790,N_8412,N_8192);
and U9791 (N_9791,N_8805,N_7093);
nand U9792 (N_9792,N_7944,N_6320);
xnor U9793 (N_9793,N_8969,N_6102);
or U9794 (N_9794,N_7387,N_8270);
nand U9795 (N_9795,N_8068,N_7779);
or U9796 (N_9796,N_7665,N_6669);
and U9797 (N_9797,N_8871,N_6795);
or U9798 (N_9798,N_6761,N_8852);
and U9799 (N_9799,N_6630,N_7554);
nor U9800 (N_9800,N_8995,N_6198);
nand U9801 (N_9801,N_6519,N_8029);
nand U9802 (N_9802,N_7936,N_6801);
and U9803 (N_9803,N_6204,N_7071);
nor U9804 (N_9804,N_6640,N_7868);
nor U9805 (N_9805,N_7389,N_7214);
nand U9806 (N_9806,N_6607,N_6826);
nand U9807 (N_9807,N_6329,N_6732);
xnor U9808 (N_9808,N_7404,N_6218);
nand U9809 (N_9809,N_8052,N_7497);
or U9810 (N_9810,N_6013,N_6712);
nor U9811 (N_9811,N_7351,N_8276);
nor U9812 (N_9812,N_8536,N_6362);
xor U9813 (N_9813,N_7195,N_8795);
nand U9814 (N_9814,N_6390,N_6192);
nor U9815 (N_9815,N_7761,N_8587);
nor U9816 (N_9816,N_8900,N_6261);
or U9817 (N_9817,N_7364,N_7227);
and U9818 (N_9818,N_6588,N_8626);
and U9819 (N_9819,N_7245,N_7962);
and U9820 (N_9820,N_7305,N_6615);
nor U9821 (N_9821,N_6583,N_8356);
or U9822 (N_9822,N_6843,N_6924);
or U9823 (N_9823,N_8937,N_7088);
and U9824 (N_9824,N_7548,N_7347);
nor U9825 (N_9825,N_6429,N_7927);
nor U9826 (N_9826,N_8758,N_8743);
or U9827 (N_9827,N_8084,N_6842);
nor U9828 (N_9828,N_7492,N_8252);
or U9829 (N_9829,N_7717,N_6870);
and U9830 (N_9830,N_7110,N_7373);
nand U9831 (N_9831,N_8663,N_6268);
or U9832 (N_9832,N_8853,N_6697);
or U9833 (N_9833,N_8797,N_8514);
and U9834 (N_9834,N_7597,N_6395);
or U9835 (N_9835,N_7241,N_7862);
nand U9836 (N_9836,N_6347,N_8630);
nor U9837 (N_9837,N_6185,N_8603);
nand U9838 (N_9838,N_8497,N_8857);
nand U9839 (N_9839,N_7643,N_6464);
and U9840 (N_9840,N_7569,N_7450);
nand U9841 (N_9841,N_8149,N_8244);
and U9842 (N_9842,N_7545,N_7521);
nor U9843 (N_9843,N_6433,N_6916);
nand U9844 (N_9844,N_6291,N_7584);
nor U9845 (N_9845,N_8974,N_6253);
nand U9846 (N_9846,N_7725,N_7799);
nor U9847 (N_9847,N_6438,N_6194);
or U9848 (N_9848,N_8791,N_7115);
nand U9849 (N_9849,N_7371,N_6241);
nand U9850 (N_9850,N_7682,N_8811);
nand U9851 (N_9851,N_8281,N_6626);
nand U9852 (N_9852,N_8321,N_6638);
or U9853 (N_9853,N_8479,N_7137);
and U9854 (N_9854,N_8544,N_6502);
nor U9855 (N_9855,N_7510,N_7714);
nand U9856 (N_9856,N_6088,N_8282);
or U9857 (N_9857,N_6017,N_6231);
nor U9858 (N_9858,N_7704,N_8550);
and U9859 (N_9859,N_7272,N_8224);
and U9860 (N_9860,N_8860,N_8353);
or U9861 (N_9861,N_6751,N_6158);
nand U9862 (N_9862,N_8720,N_8168);
or U9863 (N_9863,N_8615,N_6173);
nor U9864 (N_9864,N_8738,N_8843);
or U9865 (N_9865,N_6443,N_6846);
and U9866 (N_9866,N_6335,N_6518);
and U9867 (N_9867,N_6604,N_6979);
nand U9868 (N_9868,N_8398,N_8126);
nand U9869 (N_9869,N_8533,N_6927);
or U9870 (N_9870,N_7827,N_8245);
and U9871 (N_9871,N_7641,N_8471);
nor U9872 (N_9872,N_6406,N_6083);
nand U9873 (N_9873,N_8459,N_7117);
and U9874 (N_9874,N_6657,N_7108);
nor U9875 (N_9875,N_6755,N_6901);
nand U9876 (N_9876,N_7750,N_8947);
or U9877 (N_9877,N_8521,N_7156);
nor U9878 (N_9878,N_7407,N_6837);
nand U9879 (N_9879,N_7170,N_7888);
or U9880 (N_9880,N_8993,N_8416);
and U9881 (N_9881,N_7094,N_8328);
and U9882 (N_9882,N_7997,N_7266);
and U9883 (N_9883,N_6963,N_7395);
nand U9884 (N_9884,N_7594,N_6644);
nor U9885 (N_9885,N_8350,N_7989);
and U9886 (N_9886,N_8705,N_7070);
or U9887 (N_9887,N_8101,N_7429);
or U9888 (N_9888,N_8745,N_8419);
nor U9889 (N_9889,N_7311,N_8121);
nand U9890 (N_9890,N_6154,N_7036);
nand U9891 (N_9891,N_7867,N_7006);
nand U9892 (N_9892,N_6565,N_7224);
nand U9893 (N_9893,N_7379,N_6039);
or U9894 (N_9894,N_8788,N_8889);
or U9895 (N_9895,N_8015,N_8503);
or U9896 (N_9896,N_6798,N_7702);
nand U9897 (N_9897,N_8654,N_6015);
nor U9898 (N_9898,N_7030,N_7543);
and U9899 (N_9899,N_8789,N_8303);
nand U9900 (N_9900,N_7879,N_7256);
nor U9901 (N_9901,N_6229,N_8236);
and U9902 (N_9902,N_8890,N_7056);
and U9903 (N_9903,N_8921,N_7567);
and U9904 (N_9904,N_7787,N_6714);
or U9905 (N_9905,N_7530,N_8272);
or U9906 (N_9906,N_8393,N_8123);
nand U9907 (N_9907,N_6891,N_7430);
and U9908 (N_9908,N_7265,N_8982);
or U9909 (N_9909,N_7671,N_7308);
or U9910 (N_9910,N_6415,N_6393);
nor U9911 (N_9911,N_7344,N_6772);
nor U9912 (N_9912,N_8176,N_7326);
nor U9913 (N_9913,N_7517,N_6137);
or U9914 (N_9914,N_8557,N_6427);
nor U9915 (N_9915,N_7484,N_6770);
or U9916 (N_9916,N_8812,N_6038);
and U9917 (N_9917,N_8859,N_8277);
and U9918 (N_9918,N_7187,N_8368);
nand U9919 (N_9919,N_7883,N_7076);
or U9920 (N_9920,N_6208,N_6597);
or U9921 (N_9921,N_6338,N_8821);
nor U9922 (N_9922,N_8370,N_8173);
and U9923 (N_9923,N_7980,N_8815);
or U9924 (N_9924,N_8170,N_8271);
nor U9925 (N_9925,N_6490,N_7079);
nor U9926 (N_9926,N_6860,N_8953);
nor U9927 (N_9927,N_6051,N_6150);
or U9928 (N_9928,N_7225,N_8380);
and U9929 (N_9929,N_8556,N_6435);
or U9930 (N_9930,N_8023,N_7746);
nand U9931 (N_9931,N_6176,N_6690);
nand U9932 (N_9932,N_7786,N_7042);
nor U9933 (N_9933,N_8494,N_8257);
nand U9934 (N_9934,N_8760,N_7357);
nor U9935 (N_9935,N_7173,N_6073);
and U9936 (N_9936,N_7028,N_7905);
and U9937 (N_9937,N_6845,N_8468);
or U9938 (N_9938,N_7977,N_6527);
nand U9939 (N_9939,N_8991,N_7338);
nor U9940 (N_9940,N_6589,N_7118);
and U9941 (N_9941,N_6175,N_8474);
and U9942 (N_9942,N_6969,N_8986);
nand U9943 (N_9943,N_8442,N_8142);
or U9944 (N_9944,N_8508,N_8830);
xnor U9945 (N_9945,N_8507,N_6301);
and U9946 (N_9946,N_8265,N_6294);
nor U9947 (N_9947,N_8771,N_7086);
or U9948 (N_9948,N_8174,N_8706);
or U9949 (N_9949,N_6918,N_6061);
and U9950 (N_9950,N_7232,N_7190);
nor U9951 (N_9951,N_8443,N_6983);
nor U9952 (N_9952,N_6252,N_7833);
or U9953 (N_9953,N_7207,N_7782);
and U9954 (N_9954,N_6637,N_8166);
nor U9955 (N_9955,N_6822,N_7322);
nor U9956 (N_9956,N_8787,N_6465);
nor U9957 (N_9957,N_8379,N_7992);
nand U9958 (N_9958,N_6440,N_8643);
nand U9959 (N_9959,N_8764,N_7582);
or U9960 (N_9960,N_8105,N_6008);
or U9961 (N_9961,N_6042,N_8753);
or U9962 (N_9962,N_7852,N_6367);
or U9963 (N_9963,N_6459,N_8802);
and U9964 (N_9964,N_8152,N_6821);
nor U9965 (N_9965,N_6246,N_7966);
and U9966 (N_9966,N_7703,N_8467);
or U9967 (N_9967,N_8096,N_8713);
or U9968 (N_9968,N_7575,N_7568);
and U9969 (N_9969,N_6632,N_8693);
nand U9970 (N_9970,N_7477,N_7858);
nand U9971 (N_9971,N_7785,N_6240);
or U9972 (N_9972,N_6805,N_6819);
or U9973 (N_9973,N_6458,N_8785);
nand U9974 (N_9974,N_6681,N_6161);
and U9975 (N_9975,N_6746,N_6339);
nor U9976 (N_9976,N_8163,N_6799);
nor U9977 (N_9977,N_8598,N_6460);
nor U9978 (N_9978,N_7925,N_7715);
or U9979 (N_9979,N_6892,N_6662);
nor U9980 (N_9980,N_8445,N_6078);
nor U9981 (N_9981,N_7359,N_6591);
nor U9982 (N_9982,N_8354,N_6598);
and U9983 (N_9983,N_8352,N_6376);
nand U9984 (N_9984,N_8248,N_7593);
nand U9985 (N_9985,N_6744,N_8005);
nand U9986 (N_9986,N_8834,N_6247);
nor U9987 (N_9987,N_7549,N_7077);
nor U9988 (N_9988,N_8480,N_7184);
or U9989 (N_9989,N_8267,N_8150);
and U9990 (N_9990,N_6605,N_8581);
nor U9991 (N_9991,N_8751,N_7503);
nor U9992 (N_9992,N_6663,N_6069);
nor U9993 (N_9993,N_7535,N_7601);
or U9994 (N_9994,N_8727,N_8929);
nand U9995 (N_9995,N_6784,N_6497);
nor U9996 (N_9996,N_7946,N_7587);
and U9997 (N_9997,N_6684,N_7014);
nand U9998 (N_9998,N_7998,N_7794);
nor U9999 (N_9999,N_7546,N_8213);
xnor U10000 (N_10000,N_6184,N_8796);
and U10001 (N_10001,N_6858,N_7629);
nand U10002 (N_10002,N_7850,N_7419);
or U10003 (N_10003,N_8124,N_7618);
nand U10004 (N_10004,N_7859,N_8784);
nand U10005 (N_10005,N_7462,N_6829);
nor U10006 (N_10006,N_6741,N_7938);
nor U10007 (N_10007,N_7239,N_7312);
nand U10008 (N_10008,N_7393,N_7752);
nand U10009 (N_10009,N_7329,N_6695);
nand U10010 (N_10010,N_6118,N_8773);
nand U10011 (N_10011,N_7581,N_7402);
and U10012 (N_10012,N_8214,N_8119);
or U10013 (N_10013,N_7060,N_6304);
or U10014 (N_10014,N_7286,N_8031);
nor U10015 (N_10015,N_8067,N_8306);
nor U10016 (N_10016,N_8397,N_7747);
or U10017 (N_10017,N_6417,N_7002);
or U10018 (N_10018,N_6276,N_6331);
nand U10019 (N_10019,N_6153,N_8658);
or U10020 (N_10020,N_6308,N_8575);
nand U10021 (N_10021,N_8531,N_6125);
and U10022 (N_10022,N_8212,N_6779);
or U10023 (N_10023,N_8342,N_6006);
or U10024 (N_10024,N_7533,N_8120);
nor U10025 (N_10025,N_8476,N_8958);
or U10026 (N_10026,N_8583,N_6794);
nor U10027 (N_10027,N_8542,N_7453);
nor U10028 (N_10028,N_8665,N_6457);
nand U10029 (N_10029,N_8016,N_8122);
and U10030 (N_10030,N_8595,N_6811);
and U10031 (N_10031,N_8195,N_7141);
or U10032 (N_10032,N_8981,N_7783);
nand U10033 (N_10033,N_6067,N_8612);
and U10034 (N_10034,N_6500,N_6932);
nor U10035 (N_10035,N_8413,N_6649);
nand U10036 (N_10036,N_6911,N_7021);
nor U10037 (N_10037,N_6976,N_6300);
or U10038 (N_10038,N_8798,N_7817);
or U10039 (N_10039,N_7016,N_8869);
and U10040 (N_10040,N_7805,N_8418);
nand U10041 (N_10041,N_8454,N_8741);
and U10042 (N_10042,N_8614,N_7940);
xnor U10043 (N_10043,N_8280,N_7128);
or U10044 (N_10044,N_6071,N_8319);
nor U10045 (N_10045,N_6867,N_8794);
nand U10046 (N_10046,N_6606,N_8846);
or U10047 (N_10047,N_7069,N_6486);
or U10048 (N_10048,N_7403,N_8746);
nand U10049 (N_10049,N_6123,N_7426);
nor U10050 (N_10050,N_7196,N_8222);
or U10051 (N_10051,N_8018,N_6070);
nand U10052 (N_10052,N_8728,N_8405);
nand U10053 (N_10053,N_7605,N_7435);
nand U10054 (N_10054,N_8677,N_7734);
and U10055 (N_10055,N_8933,N_7090);
and U10056 (N_10056,N_6621,N_7645);
or U10057 (N_10057,N_6196,N_8283);
and U10058 (N_10058,N_8013,N_6383);
nor U10059 (N_10059,N_8391,N_8825);
nor U10060 (N_10060,N_6074,N_7223);
and U10061 (N_10061,N_6643,N_6447);
and U10062 (N_10062,N_6587,N_8883);
nand U10063 (N_10063,N_6052,N_8543);
or U10064 (N_10064,N_7129,N_7017);
and U10065 (N_10065,N_6115,N_8329);
or U10066 (N_10066,N_7668,N_8375);
nand U10067 (N_10067,N_7751,N_7741);
and U10068 (N_10068,N_6001,N_8144);
or U10069 (N_10069,N_7891,N_7986);
and U10070 (N_10070,N_6454,N_6299);
nand U10071 (N_10071,N_8733,N_6997);
nand U10072 (N_10072,N_8672,N_7163);
nor U10073 (N_10073,N_6103,N_6871);
or U10074 (N_10074,N_7328,N_8807);
or U10075 (N_10075,N_6782,N_8988);
nor U10076 (N_10076,N_7889,N_8772);
nor U10077 (N_10077,N_7755,N_7897);
nand U10078 (N_10078,N_7841,N_7051);
or U10079 (N_10079,N_6332,N_8532);
nand U10080 (N_10080,N_8209,N_6835);
or U10081 (N_10081,N_8080,N_8648);
and U10082 (N_10082,N_6783,N_7100);
or U10083 (N_10083,N_8774,N_6145);
nand U10084 (N_10084,N_7336,N_6087);
and U10085 (N_10085,N_6019,N_8188);
nor U10086 (N_10086,N_7540,N_8381);
and U10087 (N_10087,N_8180,N_7035);
nand U10088 (N_10088,N_7724,N_7653);
nand U10089 (N_10089,N_8826,N_6095);
nor U10090 (N_10090,N_6097,N_7433);
and U10091 (N_10091,N_7529,N_7096);
nor U10092 (N_10092,N_8233,N_6302);
nand U10093 (N_10093,N_6451,N_7970);
or U10094 (N_10094,N_8373,N_8185);
nor U10095 (N_10095,N_8078,N_8199);
nor U10096 (N_10096,N_8039,N_7031);
nand U10097 (N_10097,N_6456,N_8625);
nor U10098 (N_10098,N_7471,N_7612);
nor U10099 (N_10099,N_7670,N_7712);
or U10100 (N_10100,N_8145,N_8685);
and U10101 (N_10101,N_6999,N_8045);
nand U10102 (N_10102,N_6141,N_7916);
and U10103 (N_10103,N_6402,N_7943);
and U10104 (N_10104,N_6686,N_7165);
nand U10105 (N_10105,N_6789,N_6439);
xnor U10106 (N_10106,N_6806,N_8602);
nand U10107 (N_10107,N_8537,N_7733);
nand U10108 (N_10108,N_6491,N_6815);
nor U10109 (N_10109,N_8838,N_8037);
and U10110 (N_10110,N_7455,N_8861);
nor U10111 (N_10111,N_8816,N_7434);
or U10112 (N_10112,N_6420,N_7294);
nor U10113 (N_10113,N_7445,N_6206);
or U10114 (N_10114,N_7694,N_7367);
nor U10115 (N_10115,N_7015,N_8187);
or U10116 (N_10116,N_6287,N_6689);
and U10117 (N_10117,N_6961,N_6172);
and U10118 (N_10118,N_7467,N_7064);
and U10119 (N_10119,N_7045,N_8196);
nand U10120 (N_10120,N_6882,N_6988);
and U10121 (N_10121,N_7825,N_8050);
nand U10122 (N_10122,N_8836,N_8083);
or U10123 (N_10123,N_8572,N_6896);
nand U10124 (N_10124,N_6131,N_8028);
or U10125 (N_10125,N_6245,N_6512);
and U10126 (N_10126,N_7498,N_7446);
nand U10127 (N_10127,N_6312,N_8548);
nor U10128 (N_10128,N_7667,N_8923);
and U10129 (N_10129,N_7388,N_7951);
nor U10130 (N_10130,N_7588,N_6673);
nor U10131 (N_10131,N_6049,N_6266);
and U10132 (N_10132,N_7771,N_7599);
or U10133 (N_10133,N_7460,N_8956);
nand U10134 (N_10134,N_7009,N_7609);
and U10135 (N_10135,N_8420,N_6940);
and U10136 (N_10136,N_8298,N_7029);
nor U10137 (N_10137,N_7348,N_7255);
or U10138 (N_10138,N_6432,N_8567);
and U10139 (N_10139,N_8520,N_6917);
and U10140 (N_10140,N_8495,N_7885);
and U10141 (N_10141,N_7024,N_8985);
nor U10142 (N_10142,N_7472,N_8573);
nor U10143 (N_10143,N_8599,N_8428);
or U10144 (N_10144,N_7246,N_7744);
or U10145 (N_10145,N_8863,N_7686);
or U10146 (N_10146,N_8081,N_7620);
nand U10147 (N_10147,N_8723,N_6791);
nand U10148 (N_10148,N_6709,N_6488);
and U10149 (N_10149,N_6134,N_6056);
or U10150 (N_10150,N_6503,N_7084);
nand U10151 (N_10151,N_6306,N_6511);
and U10152 (N_10152,N_7193,N_7816);
nand U10153 (N_10153,N_8980,N_8431);
and U10154 (N_10154,N_6009,N_8655);
or U10155 (N_10155,N_8048,N_6058);
or U10156 (N_10156,N_8372,N_8094);
nor U10157 (N_10157,N_8190,N_6479);
and U10158 (N_10158,N_6282,N_6081);
and U10159 (N_10159,N_7019,N_8731);
and U10160 (N_10160,N_8478,N_8070);
nor U10161 (N_10161,N_8324,N_6168);
and U10162 (N_10162,N_6864,N_7372);
or U10163 (N_10163,N_6636,N_6659);
and U10164 (N_10164,N_6713,N_6119);
and U10165 (N_10165,N_8946,N_6658);
nor U10166 (N_10166,N_6998,N_8385);
nand U10167 (N_10167,N_7356,N_6536);
and U10168 (N_10168,N_7579,N_6359);
nor U10169 (N_10169,N_7969,N_6195);
nor U10170 (N_10170,N_8402,N_8110);
or U10171 (N_10171,N_7304,N_7876);
or U10172 (N_10172,N_6586,N_8444);
nand U10173 (N_10173,N_6624,N_6160);
or U10174 (N_10174,N_7949,N_7350);
and U10175 (N_10175,N_6178,N_8666);
xnor U10176 (N_10176,N_7621,N_8639);
and U10177 (N_10177,N_8624,N_6157);
and U10178 (N_10178,N_6678,N_6599);
and U10179 (N_10179,N_8972,N_8512);
or U10180 (N_10180,N_6814,N_7945);
or U10181 (N_10181,N_7617,N_7678);
or U10182 (N_10182,N_6357,N_8115);
nor U10183 (N_10183,N_7415,N_8279);
nor U10184 (N_10184,N_6702,N_6889);
nand U10185 (N_10185,N_8656,N_6397);
or U10186 (N_10186,N_7933,N_8912);
nand U10187 (N_10187,N_8559,N_8305);
or U10188 (N_10188,N_8486,N_6972);
and U10189 (N_10189,N_7898,N_6461);
nor U10190 (N_10190,N_6212,N_6140);
nor U10191 (N_10191,N_8847,N_7502);
nor U10192 (N_10192,N_7339,N_8308);
and U10193 (N_10193,N_7252,N_8092);
and U10194 (N_10194,N_8462,N_6994);
or U10195 (N_10195,N_7657,N_6319);
or U10196 (N_10196,N_7306,N_7737);
nand U10197 (N_10197,N_6473,N_7796);
or U10198 (N_10198,N_8679,N_8530);
nor U10199 (N_10199,N_7394,N_7431);
nor U10200 (N_10200,N_6872,N_7913);
nand U10201 (N_10201,N_6880,N_7013);
nor U10202 (N_10202,N_7425,N_6394);
or U10203 (N_10203,N_7381,N_6904);
or U10204 (N_10204,N_6879,N_6324);
and U10205 (N_10205,N_7410,N_7640);
nor U10206 (N_10206,N_8012,N_8204);
nor U10207 (N_10207,N_7113,N_8724);
or U10208 (N_10208,N_8310,N_8592);
and U10209 (N_10209,N_7685,N_6757);
and U10210 (N_10210,N_7208,N_8566);
and U10211 (N_10211,N_6050,N_8632);
and U10212 (N_10212,N_6620,N_7346);
or U10213 (N_10213,N_7169,N_6289);
nor U10214 (N_10214,N_7638,N_8657);
nor U10215 (N_10215,N_6303,N_7180);
nor U10216 (N_10216,N_8481,N_8438);
nor U10217 (N_10217,N_6189,N_6996);
nor U10218 (N_10218,N_7475,N_8323);
and U10219 (N_10219,N_6816,N_6820);
nor U10220 (N_10220,N_7215,N_7652);
and U10221 (N_10221,N_7324,N_8097);
and U10222 (N_10222,N_7659,N_8534);
nor U10223 (N_10223,N_6091,N_8033);
nor U10224 (N_10224,N_7489,N_7220);
and U10225 (N_10225,N_8217,N_7397);
or U10226 (N_10226,N_8220,N_8699);
nor U10227 (N_10227,N_8718,N_8578);
and U10228 (N_10228,N_7469,N_6057);
nor U10229 (N_10229,N_6856,N_7524);
and U10230 (N_10230,N_6426,N_8694);
nand U10231 (N_10231,N_6418,N_7008);
or U10232 (N_10232,N_7148,N_7984);
nand U10233 (N_10233,N_6024,N_6721);
nand U10234 (N_10234,N_7119,N_8042);
nor U10235 (N_10235,N_8286,N_6028);
or U10236 (N_10236,N_8571,N_6257);
nor U10237 (N_10237,N_8135,N_7598);
and U10238 (N_10238,N_6275,N_8036);
nand U10239 (N_10239,N_7622,N_8460);
nor U10240 (N_10240,N_7281,N_7800);
or U10241 (N_10241,N_8242,N_6973);
or U10242 (N_10242,N_7544,N_7918);
nor U10243 (N_10243,N_8740,N_7427);
or U10244 (N_10244,N_6027,N_8351);
or U10245 (N_10245,N_7887,N_8901);
and U10246 (N_10246,N_8820,N_6601);
and U10247 (N_10247,N_7831,N_8464);
or U10248 (N_10248,N_6688,N_6575);
nand U10249 (N_10249,N_8337,N_6480);
or U10250 (N_10250,N_6149,N_7985);
and U10251 (N_10251,N_8074,N_7253);
nand U10252 (N_10252,N_7928,N_6742);
or U10253 (N_10253,N_7790,N_7740);
and U10254 (N_10254,N_8928,N_6612);
nor U10255 (N_10255,N_7126,N_8647);
nor U10256 (N_10256,N_6193,N_7869);
or U10257 (N_10257,N_7516,N_6286);
and U10258 (N_10258,N_7153,N_7828);
nor U10259 (N_10259,N_7319,N_7080);
nor U10260 (N_10260,N_8783,N_6827);
or U10261 (N_10261,N_7506,N_8147);
nand U10262 (N_10262,N_7900,N_7723);
nand U10263 (N_10263,N_8817,N_6554);
nor U10264 (N_10264,N_8439,N_7789);
and U10265 (N_10265,N_7047,N_7848);
and U10266 (N_10266,N_6148,N_7161);
or U10267 (N_10267,N_8182,N_7559);
or U10268 (N_10268,N_8455,N_6914);
and U10269 (N_10269,N_7263,N_8198);
and U10270 (N_10270,N_8434,N_7383);
or U10271 (N_10271,N_8754,N_7353);
nand U10272 (N_10272,N_7247,N_8943);
or U10273 (N_10273,N_6767,N_8714);
or U10274 (N_10274,N_6147,N_6849);
and U10275 (N_10275,N_6167,N_8735);
and U10276 (N_10276,N_8674,N_6205);
or U10277 (N_10277,N_6707,N_8451);
nor U10278 (N_10278,N_6170,N_6800);
nand U10279 (N_10279,N_7688,N_6084);
nor U10280 (N_10280,N_8197,N_6139);
nand U10281 (N_10281,N_7033,N_6187);
nor U10282 (N_10282,N_8782,N_7116);
or U10283 (N_10283,N_8862,N_8112);
and U10284 (N_10284,N_6183,N_6200);
nand U10285 (N_10285,N_7439,N_8819);
and U10286 (N_10286,N_8206,N_7083);
and U10287 (N_10287,N_6685,N_7212);
and U10288 (N_10288,N_6348,N_8851);
or U10289 (N_10289,N_7349,N_6270);
nand U10290 (N_10290,N_8504,N_6215);
nor U10291 (N_10291,N_6370,N_7705);
nand U10292 (N_10292,N_8458,N_7881);
and U10293 (N_10293,N_7921,N_7556);
nor U10294 (N_10294,N_7736,N_7607);
and U10295 (N_10295,N_8779,N_6542);
nand U10296 (N_10296,N_7052,N_8925);
or U10297 (N_10297,N_6570,N_6859);
and U10298 (N_10298,N_8870,N_8992);
or U10299 (N_10299,N_7695,N_7978);
and U10300 (N_10300,N_8983,N_7583);
xnor U10301 (N_10301,N_6985,N_8158);
or U10302 (N_10302,N_7870,N_6670);
nand U10303 (N_10303,N_6633,N_8717);
nand U10304 (N_10304,N_8700,N_7849);
or U10305 (N_10305,N_8181,N_6944);
nand U10306 (N_10306,N_7875,N_8064);
or U10307 (N_10307,N_7423,N_8961);
nand U10308 (N_10308,N_6004,N_6278);
or U10309 (N_10309,N_7974,N_6780);
nor U10310 (N_10310,N_7432,N_6793);
and U10311 (N_10311,N_8942,N_7234);
and U10312 (N_10312,N_8613,N_7625);
nand U10313 (N_10313,N_7570,N_6968);
nand U10314 (N_10314,N_8910,N_8739);
or U10315 (N_10315,N_6937,N_6310);
nor U10316 (N_10316,N_7815,N_7307);
nand U10317 (N_10317,N_7834,N_6717);
nor U10318 (N_10318,N_7994,N_6625);
nand U10319 (N_10319,N_6584,N_8034);
or U10320 (N_10320,N_7441,N_8856);
and U10321 (N_10321,N_7795,N_7757);
and U10322 (N_10322,N_7390,N_6031);
and U10323 (N_10323,N_8944,N_7937);
or U10324 (N_10324,N_8171,N_6138);
and U10325 (N_10325,N_8831,N_6608);
nand U10326 (N_10326,N_7613,N_7941);
or U10327 (N_10327,N_6400,N_8127);
or U10328 (N_10328,N_6848,N_8837);
or U10329 (N_10329,N_7894,N_6455);
or U10330 (N_10330,N_6159,N_6553);
and U10331 (N_10331,N_6747,N_6830);
and U10332 (N_10332,N_7983,N_6068);
or U10333 (N_10333,N_8175,N_7627);
and U10334 (N_10334,N_8294,N_7635);
nand U10335 (N_10335,N_6566,N_8254);
nor U10336 (N_10336,N_7154,N_8200);
and U10337 (N_10337,N_7465,N_8593);
nor U10338 (N_10338,N_7660,N_6593);
or U10339 (N_10339,N_8313,N_6962);
nand U10340 (N_10340,N_8876,N_6182);
nand U10341 (N_10341,N_6723,N_8759);
and U10342 (N_10342,N_8711,N_7003);
or U10343 (N_10343,N_8617,N_7865);
or U10344 (N_10344,N_8086,N_6375);
or U10345 (N_10345,N_8400,N_6342);
nand U10346 (N_10346,N_6666,N_6528);
nor U10347 (N_10347,N_6646,N_8157);
nand U10348 (N_10348,N_7049,N_8332);
or U10349 (N_10349,N_7458,N_8287);
and U10350 (N_10350,N_7902,N_7111);
and U10351 (N_10351,N_6855,N_7673);
and U10352 (N_10352,N_6813,N_8024);
or U10353 (N_10353,N_6036,N_6745);
or U10354 (N_10354,N_8362,N_8215);
nand U10355 (N_10355,N_7242,N_7708);
nor U10356 (N_10356,N_6853,N_7603);
nand U10357 (N_10357,N_6881,N_8435);
and U10358 (N_10358,N_6223,N_8032);
nand U10359 (N_10359,N_6236,N_8683);
nand U10360 (N_10360,N_8854,N_8757);
and U10361 (N_10361,N_8100,N_6769);
and U10362 (N_10362,N_6358,N_6404);
nor U10363 (N_10363,N_7911,N_6449);
or U10364 (N_10364,N_8299,N_7957);
and U10365 (N_10365,N_7279,N_8208);
nor U10366 (N_10366,N_6444,N_7743);
or U10367 (N_10367,N_6890,N_6749);
and U10368 (N_10368,N_8065,N_8908);
nand U10369 (N_10369,N_7764,N_8483);
or U10370 (N_10370,N_8965,N_8469);
nand U10371 (N_10371,N_8138,N_6482);
xnor U10372 (N_10372,N_6132,N_6952);
or U10373 (N_10373,N_7146,N_8325);
nand U10374 (N_10374,N_7520,N_8164);
or U10375 (N_10375,N_6661,N_7135);
nor U10376 (N_10376,N_8358,N_6035);
and U10377 (N_10377,N_6724,N_8800);
nor U10378 (N_10378,N_6715,N_6368);
nand U10379 (N_10379,N_8999,N_7316);
nand U10380 (N_10380,N_8661,N_7204);
nor U10381 (N_10381,N_6034,N_7781);
nor U10382 (N_10382,N_8179,N_6467);
or U10383 (N_10383,N_6580,N_7178);
nand U10384 (N_10384,N_6297,N_7368);
nand U10385 (N_10385,N_8239,N_8642);
nor U10386 (N_10386,N_7507,N_8184);
and U10387 (N_10387,N_8383,N_6857);
or U10388 (N_10388,N_8560,N_6484);
nor U10389 (N_10389,N_6987,N_6733);
and U10390 (N_10390,N_6340,N_8926);
nand U10391 (N_10391,N_6040,N_7968);
nand U10392 (N_10392,N_8515,N_8955);
or U10393 (N_10393,N_8752,N_6283);
nor U10394 (N_10394,N_8389,N_8938);
or U10395 (N_10395,N_6382,N_7807);
or U10396 (N_10396,N_8394,N_6777);
nand U10397 (N_10397,N_8527,N_8948);
and U10398 (N_10398,N_7197,N_6336);
nand U10399 (N_10399,N_7323,N_6378);
nand U10400 (N_10400,N_8868,N_6847);
nand U10401 (N_10401,N_6365,N_7040);
and U10402 (N_10402,N_8594,N_6984);
and U10403 (N_10403,N_8136,N_6538);
nor U10404 (N_10404,N_7854,N_8343);
or U10405 (N_10405,N_8491,N_7055);
and U10406 (N_10406,N_8238,N_8378);
or U10407 (N_10407,N_7424,N_6667);
nand U10408 (N_10408,N_6693,N_8522);
nand U10409 (N_10409,N_7788,N_6199);
or U10410 (N_10410,N_6082,N_7485);
or U10411 (N_10411,N_8409,N_6602);
nand U10412 (N_10412,N_8231,N_6483);
nand U10413 (N_10413,N_7302,N_8698);
nand U10414 (N_10414,N_7821,N_8226);
and U10415 (N_10415,N_7488,N_6975);
nor U10416 (N_10416,N_8355,N_6563);
nand U10417 (N_10417,N_6991,N_8523);
and U10418 (N_10418,N_7337,N_6428);
nor U10419 (N_10419,N_8088,N_8427);
or U10420 (N_10420,N_8477,N_6931);
nand U10421 (N_10421,N_6296,N_6930);
nand U10422 (N_10422,N_7459,N_7526);
or U10423 (N_10423,N_6096,N_7151);
and U10424 (N_10424,N_7511,N_8951);
or U10425 (N_10425,N_6635,N_7448);
nand U10426 (N_10426,N_8191,N_6341);
nor U10427 (N_10427,N_6913,N_7226);
or U10428 (N_10428,N_6412,N_7147);
nor U10429 (N_10429,N_6018,N_7209);
nand U10430 (N_10430,N_7611,N_7085);
nor U10431 (N_10431,N_7268,N_8247);
nand U10432 (N_10432,N_7479,N_8403);
nand U10433 (N_10433,N_8712,N_8882);
and U10434 (N_10434,N_7023,N_8261);
and U10435 (N_10435,N_6046,N_8539);
or U10436 (N_10436,N_8234,N_8780);
nand U10437 (N_10437,N_7188,N_7486);
nor U10438 (N_10438,N_7039,N_7018);
or U10439 (N_10439,N_7330,N_8408);
and U10440 (N_10440,N_8604,N_6558);
nor U10441 (N_10441,N_7792,N_8262);
nand U10442 (N_10442,N_7931,N_7810);
nor U10443 (N_10443,N_6243,N_8450);
or U10444 (N_10444,N_6065,N_8344);
or U10445 (N_10445,N_7542,N_8499);
and U10446 (N_10446,N_7132,N_8597);
and U10447 (N_10447,N_6628,N_7456);
nand U10448 (N_10448,N_7824,N_8885);
or U10449 (N_10449,N_7332,N_8541);
nand U10450 (N_10450,N_8737,N_8957);
or U10451 (N_10451,N_6106,N_6450);
or U10452 (N_10452,N_7320,N_7182);
nand U10453 (N_10453,N_6210,N_8453);
nor U10454 (N_10454,N_7483,N_7149);
nand U10455 (N_10455,N_6059,N_8017);
or U10456 (N_10456,N_8684,N_6508);
nand U10457 (N_10457,N_6425,N_8026);
and U10458 (N_10458,N_7124,N_8447);
or U10459 (N_10459,N_8056,N_8111);
nand U10460 (N_10460,N_6682,N_6617);
or U10461 (N_10461,N_6708,N_7525);
or U10462 (N_10462,N_7904,N_8799);
nor U10463 (N_10463,N_8917,N_8178);
or U10464 (N_10464,N_7654,N_7046);
nand U10465 (N_10465,N_6143,N_6905);
and U10466 (N_10466,N_7680,N_6228);
nand U10467 (N_10467,N_7103,N_8645);
nor U10468 (N_10468,N_7574,N_8041);
and U10469 (N_10469,N_6541,N_6032);
xor U10470 (N_10470,N_6838,N_8465);
or U10471 (N_10471,N_6532,N_6109);
and U10472 (N_10472,N_6255,N_8662);
nand U10473 (N_10473,N_8690,N_6992);
and U10474 (N_10474,N_7034,N_7280);
nand U10475 (N_10475,N_8309,N_8172);
nand U10476 (N_10476,N_6671,N_8601);
and U10477 (N_10477,N_7160,N_6839);
nand U10478 (N_10478,N_7591,N_7634);
or U10479 (N_10479,N_7508,N_7192);
or U10480 (N_10480,N_7001,N_7177);
or U10481 (N_10481,N_8077,N_6700);
nand U10482 (N_10482,N_6122,N_7081);
nand U10483 (N_10483,N_8430,N_6610);
nor U10484 (N_10484,N_8776,N_6277);
or U10485 (N_10485,N_8793,N_7012);
nand U10486 (N_10486,N_7890,N_6165);
nor U10487 (N_10487,N_8623,N_7687);
or U10488 (N_10488,N_6326,N_8952);
or U10489 (N_10489,N_6978,N_8143);
nor U10490 (N_10490,N_7960,N_7658);
xnor U10491 (N_10491,N_6596,N_7564);
or U10492 (N_10492,N_8255,N_6679);
nor U10493 (N_10493,N_8058,N_7422);
nor U10494 (N_10494,N_6127,N_6698);
xor U10495 (N_10495,N_6251,N_7341);
nand U10496 (N_10496,N_8990,N_6738);
and U10497 (N_10497,N_6762,N_8808);
nor U10498 (N_10498,N_6233,N_8177);
nor U10499 (N_10499,N_7672,N_7971);
or U10500 (N_10500,N_6682,N_7075);
nand U10501 (N_10501,N_8210,N_6552);
and U10502 (N_10502,N_8913,N_6461);
nor U10503 (N_10503,N_8645,N_8300);
nand U10504 (N_10504,N_6814,N_8124);
nand U10505 (N_10505,N_8755,N_8499);
nor U10506 (N_10506,N_8801,N_7515);
or U10507 (N_10507,N_8551,N_8651);
nand U10508 (N_10508,N_6084,N_8734);
and U10509 (N_10509,N_6137,N_8815);
nand U10510 (N_10510,N_7670,N_6835);
and U10511 (N_10511,N_7151,N_6460);
or U10512 (N_10512,N_6977,N_7894);
and U10513 (N_10513,N_8346,N_8106);
and U10514 (N_10514,N_6365,N_8140);
nand U10515 (N_10515,N_8691,N_8114);
nor U10516 (N_10516,N_7212,N_7494);
nor U10517 (N_10517,N_7890,N_6613);
or U10518 (N_10518,N_7535,N_8957);
nor U10519 (N_10519,N_6615,N_7957);
and U10520 (N_10520,N_7820,N_6944);
or U10521 (N_10521,N_6591,N_8717);
and U10522 (N_10522,N_7675,N_6328);
and U10523 (N_10523,N_8603,N_8069);
nand U10524 (N_10524,N_7754,N_6241);
and U10525 (N_10525,N_7437,N_8113);
nand U10526 (N_10526,N_8334,N_6887);
nor U10527 (N_10527,N_7934,N_6170);
and U10528 (N_10528,N_6013,N_6140);
and U10529 (N_10529,N_6339,N_6808);
or U10530 (N_10530,N_6577,N_6990);
nor U10531 (N_10531,N_8312,N_6912);
nor U10532 (N_10532,N_7236,N_6498);
nor U10533 (N_10533,N_8363,N_7006);
nor U10534 (N_10534,N_6594,N_8435);
and U10535 (N_10535,N_6234,N_6168);
nand U10536 (N_10536,N_6228,N_8101);
nor U10537 (N_10537,N_6899,N_7158);
nand U10538 (N_10538,N_7635,N_6868);
and U10539 (N_10539,N_7674,N_6904);
or U10540 (N_10540,N_8602,N_6264);
nand U10541 (N_10541,N_7818,N_7563);
and U10542 (N_10542,N_8057,N_8947);
or U10543 (N_10543,N_8713,N_7530);
and U10544 (N_10544,N_8153,N_6572);
or U10545 (N_10545,N_8382,N_8393);
nor U10546 (N_10546,N_7896,N_7279);
nand U10547 (N_10547,N_6629,N_8486);
nand U10548 (N_10548,N_7070,N_6432);
nand U10549 (N_10549,N_8195,N_8688);
nor U10550 (N_10550,N_7640,N_8257);
or U10551 (N_10551,N_7224,N_6473);
nand U10552 (N_10552,N_8825,N_6454);
nor U10553 (N_10553,N_6615,N_6868);
nand U10554 (N_10554,N_8662,N_8656);
and U10555 (N_10555,N_6282,N_8758);
or U10556 (N_10556,N_7383,N_6422);
nor U10557 (N_10557,N_7223,N_7540);
and U10558 (N_10558,N_8325,N_6487);
or U10559 (N_10559,N_8542,N_6850);
nor U10560 (N_10560,N_6682,N_8219);
and U10561 (N_10561,N_7119,N_6078);
nor U10562 (N_10562,N_8018,N_8812);
nor U10563 (N_10563,N_7619,N_8427);
nor U10564 (N_10564,N_8876,N_7508);
nor U10565 (N_10565,N_8206,N_8799);
or U10566 (N_10566,N_6739,N_6170);
nor U10567 (N_10567,N_8730,N_7225);
and U10568 (N_10568,N_8644,N_7943);
and U10569 (N_10569,N_6604,N_8272);
and U10570 (N_10570,N_7752,N_7064);
nor U10571 (N_10571,N_8938,N_7867);
nand U10572 (N_10572,N_8762,N_6326);
nand U10573 (N_10573,N_7692,N_8997);
and U10574 (N_10574,N_6609,N_6310);
or U10575 (N_10575,N_7062,N_6360);
nand U10576 (N_10576,N_7001,N_7927);
and U10577 (N_10577,N_7964,N_7075);
nor U10578 (N_10578,N_7995,N_7468);
nand U10579 (N_10579,N_7127,N_8446);
or U10580 (N_10580,N_6093,N_7935);
nor U10581 (N_10581,N_7507,N_8260);
nor U10582 (N_10582,N_7593,N_8564);
or U10583 (N_10583,N_8110,N_8504);
or U10584 (N_10584,N_6932,N_6139);
nand U10585 (N_10585,N_7594,N_7961);
nor U10586 (N_10586,N_8899,N_7582);
or U10587 (N_10587,N_6597,N_7030);
nor U10588 (N_10588,N_6265,N_7759);
and U10589 (N_10589,N_6457,N_8235);
and U10590 (N_10590,N_8913,N_7629);
nand U10591 (N_10591,N_8571,N_8761);
or U10592 (N_10592,N_8457,N_7138);
nor U10593 (N_10593,N_6695,N_6827);
and U10594 (N_10594,N_6388,N_7529);
or U10595 (N_10595,N_7535,N_6883);
nand U10596 (N_10596,N_7384,N_8861);
nand U10597 (N_10597,N_6650,N_8448);
nor U10598 (N_10598,N_8068,N_6273);
nor U10599 (N_10599,N_7763,N_8382);
nor U10600 (N_10600,N_8559,N_6670);
nand U10601 (N_10601,N_7496,N_8864);
or U10602 (N_10602,N_8469,N_8299);
nand U10603 (N_10603,N_6997,N_6577);
or U10604 (N_10604,N_8962,N_7936);
nor U10605 (N_10605,N_8244,N_7092);
nand U10606 (N_10606,N_6896,N_7155);
xor U10607 (N_10607,N_7874,N_8906);
nor U10608 (N_10608,N_6123,N_7523);
or U10609 (N_10609,N_8898,N_7372);
and U10610 (N_10610,N_6689,N_7744);
and U10611 (N_10611,N_8447,N_6845);
or U10612 (N_10612,N_6561,N_7032);
nand U10613 (N_10613,N_6183,N_8090);
nand U10614 (N_10614,N_8533,N_6811);
xnor U10615 (N_10615,N_6253,N_7235);
nor U10616 (N_10616,N_8877,N_6622);
and U10617 (N_10617,N_7148,N_6281);
and U10618 (N_10618,N_6940,N_6484);
nand U10619 (N_10619,N_6903,N_8765);
nand U10620 (N_10620,N_8999,N_6430);
nor U10621 (N_10621,N_6696,N_8521);
and U10622 (N_10622,N_7074,N_7979);
nor U10623 (N_10623,N_8715,N_7405);
or U10624 (N_10624,N_7606,N_8898);
and U10625 (N_10625,N_6273,N_8058);
and U10626 (N_10626,N_6474,N_8695);
nand U10627 (N_10627,N_6277,N_7751);
and U10628 (N_10628,N_8679,N_6878);
nand U10629 (N_10629,N_6168,N_7953);
nand U10630 (N_10630,N_6621,N_7220);
nor U10631 (N_10631,N_6421,N_7114);
nor U10632 (N_10632,N_7895,N_7985);
and U10633 (N_10633,N_8713,N_7337);
nor U10634 (N_10634,N_6370,N_8500);
nand U10635 (N_10635,N_6480,N_8067);
or U10636 (N_10636,N_7474,N_7005);
nand U10637 (N_10637,N_7108,N_6742);
nor U10638 (N_10638,N_7556,N_8530);
nor U10639 (N_10639,N_7556,N_6741);
or U10640 (N_10640,N_8247,N_7663);
and U10641 (N_10641,N_6758,N_7725);
and U10642 (N_10642,N_6895,N_6512);
or U10643 (N_10643,N_6666,N_8659);
nand U10644 (N_10644,N_8113,N_8680);
or U10645 (N_10645,N_8444,N_8461);
nor U10646 (N_10646,N_6626,N_7771);
nand U10647 (N_10647,N_7707,N_8775);
or U10648 (N_10648,N_8104,N_8651);
and U10649 (N_10649,N_8510,N_7384);
nand U10650 (N_10650,N_6740,N_7067);
or U10651 (N_10651,N_8036,N_7722);
nor U10652 (N_10652,N_8936,N_7189);
and U10653 (N_10653,N_7133,N_6351);
nor U10654 (N_10654,N_7774,N_6053);
nor U10655 (N_10655,N_7662,N_7510);
nor U10656 (N_10656,N_6540,N_8529);
nand U10657 (N_10657,N_7465,N_7067);
or U10658 (N_10658,N_8323,N_8553);
nor U10659 (N_10659,N_7062,N_8364);
and U10660 (N_10660,N_6989,N_7803);
and U10661 (N_10661,N_8080,N_8561);
nand U10662 (N_10662,N_6652,N_8476);
or U10663 (N_10663,N_7814,N_8834);
nand U10664 (N_10664,N_6477,N_7527);
nand U10665 (N_10665,N_7020,N_8812);
nor U10666 (N_10666,N_6641,N_6311);
nor U10667 (N_10667,N_6022,N_6676);
or U10668 (N_10668,N_6215,N_6968);
or U10669 (N_10669,N_7736,N_6703);
nand U10670 (N_10670,N_8921,N_6800);
nor U10671 (N_10671,N_7670,N_8584);
nand U10672 (N_10672,N_7818,N_8631);
nor U10673 (N_10673,N_8137,N_7501);
nor U10674 (N_10674,N_7348,N_8022);
nand U10675 (N_10675,N_8285,N_8047);
and U10676 (N_10676,N_7970,N_7769);
or U10677 (N_10677,N_8020,N_7007);
nand U10678 (N_10678,N_7700,N_6530);
nor U10679 (N_10679,N_8868,N_6237);
and U10680 (N_10680,N_6707,N_6207);
nand U10681 (N_10681,N_8180,N_7418);
or U10682 (N_10682,N_6321,N_7261);
or U10683 (N_10683,N_8598,N_8331);
nand U10684 (N_10684,N_6342,N_7152);
and U10685 (N_10685,N_8907,N_6797);
nor U10686 (N_10686,N_7821,N_8470);
and U10687 (N_10687,N_8962,N_6591);
nor U10688 (N_10688,N_8954,N_7226);
nand U10689 (N_10689,N_6100,N_7781);
or U10690 (N_10690,N_7713,N_6067);
or U10691 (N_10691,N_6853,N_8984);
or U10692 (N_10692,N_7125,N_6109);
nor U10693 (N_10693,N_7049,N_6810);
or U10694 (N_10694,N_7673,N_8436);
or U10695 (N_10695,N_6897,N_8051);
nor U10696 (N_10696,N_8867,N_7569);
nand U10697 (N_10697,N_6401,N_6593);
or U10698 (N_10698,N_8358,N_6191);
nand U10699 (N_10699,N_8268,N_8123);
and U10700 (N_10700,N_7368,N_6350);
or U10701 (N_10701,N_7628,N_8269);
nor U10702 (N_10702,N_7057,N_8872);
or U10703 (N_10703,N_7926,N_6366);
nor U10704 (N_10704,N_8126,N_8452);
or U10705 (N_10705,N_8358,N_8943);
nor U10706 (N_10706,N_7504,N_7553);
and U10707 (N_10707,N_6995,N_6251);
nand U10708 (N_10708,N_7911,N_6991);
and U10709 (N_10709,N_6839,N_6633);
nor U10710 (N_10710,N_8998,N_7531);
or U10711 (N_10711,N_8337,N_7098);
nor U10712 (N_10712,N_6193,N_7180);
and U10713 (N_10713,N_8531,N_6831);
and U10714 (N_10714,N_6840,N_8450);
or U10715 (N_10715,N_8851,N_6296);
nand U10716 (N_10716,N_6581,N_7963);
nor U10717 (N_10717,N_6557,N_8760);
and U10718 (N_10718,N_6727,N_7293);
nor U10719 (N_10719,N_7646,N_8447);
and U10720 (N_10720,N_8622,N_8209);
or U10721 (N_10721,N_6529,N_7704);
and U10722 (N_10722,N_6876,N_6564);
or U10723 (N_10723,N_7436,N_7656);
nand U10724 (N_10724,N_7412,N_6582);
xor U10725 (N_10725,N_7339,N_7397);
and U10726 (N_10726,N_6527,N_6746);
nand U10727 (N_10727,N_6106,N_6330);
nor U10728 (N_10728,N_8113,N_8105);
and U10729 (N_10729,N_6535,N_8511);
or U10730 (N_10730,N_6260,N_7228);
or U10731 (N_10731,N_7995,N_8649);
and U10732 (N_10732,N_6177,N_6890);
nor U10733 (N_10733,N_7054,N_6267);
nand U10734 (N_10734,N_7221,N_7207);
nor U10735 (N_10735,N_7723,N_7172);
nand U10736 (N_10736,N_6327,N_6383);
nor U10737 (N_10737,N_7455,N_7425);
nor U10738 (N_10738,N_8522,N_6249);
or U10739 (N_10739,N_8537,N_7929);
nand U10740 (N_10740,N_6609,N_8957);
and U10741 (N_10741,N_6395,N_7807);
and U10742 (N_10742,N_8688,N_6510);
nor U10743 (N_10743,N_8827,N_6577);
nor U10744 (N_10744,N_6790,N_7302);
nor U10745 (N_10745,N_8414,N_6203);
nand U10746 (N_10746,N_6991,N_8999);
nand U10747 (N_10747,N_7963,N_7658);
nand U10748 (N_10748,N_6055,N_6904);
nor U10749 (N_10749,N_6154,N_7659);
nand U10750 (N_10750,N_7905,N_6936);
xor U10751 (N_10751,N_7474,N_7455);
or U10752 (N_10752,N_6154,N_7519);
and U10753 (N_10753,N_6392,N_6201);
nand U10754 (N_10754,N_7258,N_7326);
nand U10755 (N_10755,N_6200,N_7864);
nand U10756 (N_10756,N_8632,N_7489);
nand U10757 (N_10757,N_6382,N_8013);
and U10758 (N_10758,N_8492,N_6747);
and U10759 (N_10759,N_6790,N_6487);
or U10760 (N_10760,N_8308,N_8763);
nand U10761 (N_10761,N_8622,N_8103);
nand U10762 (N_10762,N_7609,N_7272);
or U10763 (N_10763,N_6341,N_7331);
or U10764 (N_10764,N_8102,N_8863);
and U10765 (N_10765,N_6675,N_8277);
or U10766 (N_10766,N_6686,N_7324);
and U10767 (N_10767,N_6044,N_7219);
and U10768 (N_10768,N_8094,N_8921);
or U10769 (N_10769,N_7388,N_8468);
and U10770 (N_10770,N_7588,N_7207);
nor U10771 (N_10771,N_8177,N_8652);
nor U10772 (N_10772,N_7264,N_7048);
or U10773 (N_10773,N_7482,N_7666);
and U10774 (N_10774,N_8502,N_6996);
and U10775 (N_10775,N_6787,N_8085);
and U10776 (N_10776,N_7381,N_7309);
or U10777 (N_10777,N_6651,N_7706);
or U10778 (N_10778,N_7320,N_7321);
nand U10779 (N_10779,N_8179,N_6565);
nand U10780 (N_10780,N_8711,N_6848);
nor U10781 (N_10781,N_7544,N_6024);
nand U10782 (N_10782,N_8051,N_8926);
or U10783 (N_10783,N_7414,N_7135);
nor U10784 (N_10784,N_7301,N_7266);
and U10785 (N_10785,N_8833,N_6621);
and U10786 (N_10786,N_7875,N_6397);
nand U10787 (N_10787,N_8674,N_6416);
or U10788 (N_10788,N_7479,N_6646);
or U10789 (N_10789,N_8488,N_6649);
or U10790 (N_10790,N_6306,N_8547);
nor U10791 (N_10791,N_6190,N_6554);
and U10792 (N_10792,N_8813,N_7769);
nand U10793 (N_10793,N_8424,N_6974);
nand U10794 (N_10794,N_7673,N_7215);
nor U10795 (N_10795,N_8548,N_8514);
or U10796 (N_10796,N_8571,N_8701);
or U10797 (N_10797,N_7295,N_8784);
nand U10798 (N_10798,N_8457,N_6477);
and U10799 (N_10799,N_7359,N_8863);
nor U10800 (N_10800,N_6376,N_6936);
nand U10801 (N_10801,N_6173,N_6118);
nand U10802 (N_10802,N_6861,N_7982);
and U10803 (N_10803,N_8166,N_6791);
nand U10804 (N_10804,N_6486,N_8360);
and U10805 (N_10805,N_6825,N_7198);
or U10806 (N_10806,N_7551,N_7081);
and U10807 (N_10807,N_6267,N_7937);
and U10808 (N_10808,N_6972,N_6009);
nand U10809 (N_10809,N_7138,N_8223);
nor U10810 (N_10810,N_6523,N_7815);
or U10811 (N_10811,N_6063,N_6301);
nor U10812 (N_10812,N_8929,N_7707);
and U10813 (N_10813,N_7221,N_6933);
or U10814 (N_10814,N_8070,N_8316);
nand U10815 (N_10815,N_7683,N_8047);
and U10816 (N_10816,N_7369,N_8980);
nand U10817 (N_10817,N_7303,N_7364);
nor U10818 (N_10818,N_7519,N_7046);
or U10819 (N_10819,N_7802,N_6388);
nand U10820 (N_10820,N_8278,N_6717);
nor U10821 (N_10821,N_8061,N_7670);
or U10822 (N_10822,N_7595,N_6147);
and U10823 (N_10823,N_7865,N_7505);
nor U10824 (N_10824,N_8004,N_7813);
or U10825 (N_10825,N_8470,N_6907);
nor U10826 (N_10826,N_6256,N_6942);
or U10827 (N_10827,N_8470,N_7092);
nand U10828 (N_10828,N_8471,N_6323);
nand U10829 (N_10829,N_8400,N_7681);
and U10830 (N_10830,N_7601,N_7325);
and U10831 (N_10831,N_6012,N_8972);
nand U10832 (N_10832,N_7953,N_8524);
or U10833 (N_10833,N_7539,N_7796);
or U10834 (N_10834,N_6385,N_7425);
nand U10835 (N_10835,N_6288,N_6255);
nand U10836 (N_10836,N_6374,N_7140);
or U10837 (N_10837,N_8517,N_6723);
and U10838 (N_10838,N_6689,N_6449);
and U10839 (N_10839,N_6699,N_8128);
nand U10840 (N_10840,N_8208,N_8133);
or U10841 (N_10841,N_7421,N_8724);
and U10842 (N_10842,N_8790,N_6703);
or U10843 (N_10843,N_8812,N_8503);
or U10844 (N_10844,N_7870,N_8484);
nor U10845 (N_10845,N_6352,N_8687);
nand U10846 (N_10846,N_8001,N_6511);
and U10847 (N_10847,N_6389,N_8947);
and U10848 (N_10848,N_8488,N_7018);
or U10849 (N_10849,N_8178,N_6438);
nand U10850 (N_10850,N_8940,N_8218);
or U10851 (N_10851,N_8429,N_8728);
nand U10852 (N_10852,N_7355,N_7927);
nand U10853 (N_10853,N_7075,N_6132);
nand U10854 (N_10854,N_6046,N_6340);
and U10855 (N_10855,N_6217,N_6924);
or U10856 (N_10856,N_7002,N_6428);
nor U10857 (N_10857,N_6937,N_8802);
nand U10858 (N_10858,N_6858,N_6682);
or U10859 (N_10859,N_8502,N_6732);
and U10860 (N_10860,N_7453,N_7372);
nand U10861 (N_10861,N_6686,N_6346);
nor U10862 (N_10862,N_8186,N_7039);
or U10863 (N_10863,N_7473,N_6593);
nand U10864 (N_10864,N_8584,N_6561);
or U10865 (N_10865,N_7138,N_7532);
nor U10866 (N_10866,N_8223,N_7184);
or U10867 (N_10867,N_8638,N_7844);
and U10868 (N_10868,N_8307,N_8708);
and U10869 (N_10869,N_6404,N_6622);
nor U10870 (N_10870,N_6188,N_7759);
nor U10871 (N_10871,N_6392,N_8622);
nor U10872 (N_10872,N_8331,N_6698);
or U10873 (N_10873,N_8048,N_7892);
nor U10874 (N_10874,N_7181,N_6896);
and U10875 (N_10875,N_8522,N_8240);
nor U10876 (N_10876,N_6499,N_8477);
nor U10877 (N_10877,N_8641,N_7735);
and U10878 (N_10878,N_7960,N_7844);
nor U10879 (N_10879,N_7869,N_6689);
nand U10880 (N_10880,N_7326,N_8026);
and U10881 (N_10881,N_6433,N_7183);
and U10882 (N_10882,N_8856,N_7274);
nand U10883 (N_10883,N_7997,N_7607);
nor U10884 (N_10884,N_7358,N_7444);
nor U10885 (N_10885,N_6282,N_6456);
or U10886 (N_10886,N_8627,N_6897);
and U10887 (N_10887,N_8652,N_6380);
or U10888 (N_10888,N_6052,N_7591);
nand U10889 (N_10889,N_8507,N_7734);
nand U10890 (N_10890,N_7649,N_8675);
or U10891 (N_10891,N_6648,N_7291);
nor U10892 (N_10892,N_7798,N_7545);
nor U10893 (N_10893,N_8265,N_8077);
nor U10894 (N_10894,N_6015,N_6362);
or U10895 (N_10895,N_8227,N_7988);
or U10896 (N_10896,N_7554,N_6151);
or U10897 (N_10897,N_8248,N_8343);
or U10898 (N_10898,N_8409,N_7630);
nand U10899 (N_10899,N_7885,N_6990);
nor U10900 (N_10900,N_8973,N_7787);
and U10901 (N_10901,N_7290,N_6590);
nor U10902 (N_10902,N_7012,N_6038);
xor U10903 (N_10903,N_7664,N_7044);
nand U10904 (N_10904,N_7256,N_6041);
nor U10905 (N_10905,N_6556,N_6943);
or U10906 (N_10906,N_6427,N_7865);
nor U10907 (N_10907,N_6280,N_8650);
nand U10908 (N_10908,N_6460,N_6861);
nand U10909 (N_10909,N_6548,N_8781);
nand U10910 (N_10910,N_7013,N_7723);
nand U10911 (N_10911,N_6638,N_6884);
or U10912 (N_10912,N_8739,N_8038);
and U10913 (N_10913,N_6686,N_7828);
or U10914 (N_10914,N_8708,N_8880);
nand U10915 (N_10915,N_8450,N_6505);
or U10916 (N_10916,N_7898,N_7874);
or U10917 (N_10917,N_8041,N_8239);
nor U10918 (N_10918,N_8498,N_8690);
nor U10919 (N_10919,N_8005,N_6757);
and U10920 (N_10920,N_6920,N_8615);
nor U10921 (N_10921,N_8443,N_6130);
or U10922 (N_10922,N_6123,N_8961);
nor U10923 (N_10923,N_8945,N_6333);
and U10924 (N_10924,N_7082,N_6735);
nor U10925 (N_10925,N_8438,N_7493);
nor U10926 (N_10926,N_7542,N_6993);
or U10927 (N_10927,N_8525,N_6516);
and U10928 (N_10928,N_7929,N_6506);
or U10929 (N_10929,N_8378,N_7781);
or U10930 (N_10930,N_7996,N_8091);
or U10931 (N_10931,N_8916,N_7199);
and U10932 (N_10932,N_7918,N_6661);
or U10933 (N_10933,N_7474,N_7288);
or U10934 (N_10934,N_7744,N_7442);
or U10935 (N_10935,N_6494,N_7376);
nor U10936 (N_10936,N_6418,N_7052);
nor U10937 (N_10937,N_8457,N_8731);
nor U10938 (N_10938,N_8111,N_6159);
or U10939 (N_10939,N_8376,N_7145);
and U10940 (N_10940,N_6620,N_7829);
or U10941 (N_10941,N_6920,N_7380);
nand U10942 (N_10942,N_6101,N_8992);
or U10943 (N_10943,N_8487,N_7520);
nor U10944 (N_10944,N_6634,N_6637);
nand U10945 (N_10945,N_7423,N_7258);
or U10946 (N_10946,N_6819,N_8960);
nor U10947 (N_10947,N_7078,N_8159);
nor U10948 (N_10948,N_6118,N_8672);
or U10949 (N_10949,N_8360,N_8596);
or U10950 (N_10950,N_8606,N_7541);
nand U10951 (N_10951,N_6888,N_7702);
nor U10952 (N_10952,N_8510,N_7818);
and U10953 (N_10953,N_6391,N_8883);
nand U10954 (N_10954,N_6941,N_8095);
and U10955 (N_10955,N_8627,N_7937);
or U10956 (N_10956,N_7640,N_8161);
nor U10957 (N_10957,N_6003,N_8519);
or U10958 (N_10958,N_7583,N_8151);
and U10959 (N_10959,N_8116,N_8062);
nor U10960 (N_10960,N_7944,N_8215);
or U10961 (N_10961,N_6469,N_8362);
nor U10962 (N_10962,N_6380,N_8514);
nor U10963 (N_10963,N_6307,N_7339);
and U10964 (N_10964,N_8584,N_7506);
nor U10965 (N_10965,N_8655,N_7155);
nor U10966 (N_10966,N_8343,N_7764);
or U10967 (N_10967,N_7863,N_6539);
nor U10968 (N_10968,N_7756,N_7353);
nand U10969 (N_10969,N_7382,N_6242);
and U10970 (N_10970,N_8521,N_6755);
and U10971 (N_10971,N_6726,N_6214);
and U10972 (N_10972,N_6717,N_7414);
nor U10973 (N_10973,N_8420,N_8189);
nand U10974 (N_10974,N_8976,N_7098);
nor U10975 (N_10975,N_8117,N_8427);
nand U10976 (N_10976,N_8423,N_6771);
nor U10977 (N_10977,N_6710,N_8812);
and U10978 (N_10978,N_7001,N_7278);
or U10979 (N_10979,N_8736,N_7080);
nor U10980 (N_10980,N_6033,N_6439);
nor U10981 (N_10981,N_6442,N_7528);
and U10982 (N_10982,N_6405,N_6580);
xnor U10983 (N_10983,N_8375,N_7744);
nor U10984 (N_10984,N_8665,N_8563);
nand U10985 (N_10985,N_7385,N_7178);
and U10986 (N_10986,N_7502,N_6042);
or U10987 (N_10987,N_6777,N_6926);
nand U10988 (N_10988,N_8964,N_6770);
and U10989 (N_10989,N_8159,N_6838);
nor U10990 (N_10990,N_7430,N_8624);
or U10991 (N_10991,N_7713,N_6221);
and U10992 (N_10992,N_7361,N_8426);
and U10993 (N_10993,N_8359,N_8782);
nand U10994 (N_10994,N_8961,N_8630);
nand U10995 (N_10995,N_8220,N_7067);
or U10996 (N_10996,N_6455,N_7152);
or U10997 (N_10997,N_7017,N_7294);
or U10998 (N_10998,N_8308,N_6810);
and U10999 (N_10999,N_8087,N_6995);
or U11000 (N_11000,N_7537,N_6268);
and U11001 (N_11001,N_7572,N_7251);
nand U11002 (N_11002,N_6317,N_6931);
and U11003 (N_11003,N_8716,N_6338);
nand U11004 (N_11004,N_7180,N_6587);
nand U11005 (N_11005,N_7597,N_7110);
and U11006 (N_11006,N_6429,N_7893);
nor U11007 (N_11007,N_6090,N_6416);
and U11008 (N_11008,N_7597,N_8398);
or U11009 (N_11009,N_8160,N_6802);
and U11010 (N_11010,N_7495,N_6355);
nand U11011 (N_11011,N_7294,N_8415);
or U11012 (N_11012,N_7706,N_8053);
nand U11013 (N_11013,N_8711,N_7505);
nand U11014 (N_11014,N_8317,N_8080);
nor U11015 (N_11015,N_8287,N_8297);
and U11016 (N_11016,N_8328,N_6131);
or U11017 (N_11017,N_6066,N_6343);
nor U11018 (N_11018,N_6257,N_6683);
and U11019 (N_11019,N_6378,N_6702);
nand U11020 (N_11020,N_6652,N_7729);
or U11021 (N_11021,N_6098,N_7812);
or U11022 (N_11022,N_6998,N_8459);
and U11023 (N_11023,N_6944,N_6789);
and U11024 (N_11024,N_8517,N_8956);
nor U11025 (N_11025,N_6509,N_7883);
nor U11026 (N_11026,N_6529,N_6689);
nand U11027 (N_11027,N_6412,N_7271);
xnor U11028 (N_11028,N_8453,N_8048);
nand U11029 (N_11029,N_8119,N_8768);
or U11030 (N_11030,N_6647,N_8791);
nor U11031 (N_11031,N_7882,N_8943);
and U11032 (N_11032,N_7405,N_6609);
nor U11033 (N_11033,N_8929,N_8270);
and U11034 (N_11034,N_7232,N_8559);
nand U11035 (N_11035,N_7448,N_6499);
and U11036 (N_11036,N_7680,N_6899);
nor U11037 (N_11037,N_6308,N_6417);
nand U11038 (N_11038,N_7862,N_8471);
nor U11039 (N_11039,N_6619,N_7881);
and U11040 (N_11040,N_7287,N_7119);
or U11041 (N_11041,N_8312,N_7218);
nor U11042 (N_11042,N_7039,N_6665);
or U11043 (N_11043,N_7574,N_8835);
nor U11044 (N_11044,N_6201,N_6961);
nand U11045 (N_11045,N_6093,N_7416);
and U11046 (N_11046,N_8176,N_8608);
nor U11047 (N_11047,N_6325,N_7248);
nand U11048 (N_11048,N_8187,N_7720);
and U11049 (N_11049,N_7978,N_6481);
or U11050 (N_11050,N_8129,N_7508);
nand U11051 (N_11051,N_8822,N_7757);
or U11052 (N_11052,N_6568,N_8242);
nor U11053 (N_11053,N_8540,N_7035);
nand U11054 (N_11054,N_6956,N_8210);
nor U11055 (N_11055,N_6522,N_7805);
nor U11056 (N_11056,N_8190,N_6636);
and U11057 (N_11057,N_7087,N_8968);
or U11058 (N_11058,N_8510,N_8091);
nor U11059 (N_11059,N_7026,N_7128);
nor U11060 (N_11060,N_7557,N_7128);
and U11061 (N_11061,N_6549,N_7384);
nor U11062 (N_11062,N_7923,N_8273);
and U11063 (N_11063,N_8332,N_8519);
nor U11064 (N_11064,N_6098,N_6331);
and U11065 (N_11065,N_6364,N_6590);
or U11066 (N_11066,N_7879,N_7765);
nor U11067 (N_11067,N_7484,N_6941);
or U11068 (N_11068,N_6857,N_8821);
or U11069 (N_11069,N_6750,N_7674);
or U11070 (N_11070,N_6911,N_6418);
and U11071 (N_11071,N_8567,N_8945);
nand U11072 (N_11072,N_8455,N_8148);
nand U11073 (N_11073,N_6905,N_7113);
nor U11074 (N_11074,N_7883,N_7927);
nand U11075 (N_11075,N_8630,N_6904);
nand U11076 (N_11076,N_8668,N_8681);
nor U11077 (N_11077,N_6672,N_6221);
nand U11078 (N_11078,N_8983,N_8626);
nor U11079 (N_11079,N_6349,N_7769);
xnor U11080 (N_11080,N_7929,N_7955);
nand U11081 (N_11081,N_6356,N_6280);
and U11082 (N_11082,N_6735,N_8932);
nand U11083 (N_11083,N_6017,N_7319);
or U11084 (N_11084,N_8428,N_7678);
nand U11085 (N_11085,N_7952,N_8096);
nor U11086 (N_11086,N_6399,N_8874);
and U11087 (N_11087,N_7570,N_6515);
nand U11088 (N_11088,N_8178,N_7397);
nand U11089 (N_11089,N_7305,N_6721);
nand U11090 (N_11090,N_7533,N_6054);
nand U11091 (N_11091,N_8169,N_6119);
or U11092 (N_11092,N_8515,N_8507);
nand U11093 (N_11093,N_7744,N_6361);
and U11094 (N_11094,N_8188,N_6926);
nor U11095 (N_11095,N_8444,N_6537);
nor U11096 (N_11096,N_6160,N_6284);
nand U11097 (N_11097,N_7564,N_8452);
or U11098 (N_11098,N_7008,N_6885);
nor U11099 (N_11099,N_6174,N_7454);
or U11100 (N_11100,N_6770,N_7669);
and U11101 (N_11101,N_7504,N_7468);
nor U11102 (N_11102,N_7116,N_7590);
and U11103 (N_11103,N_7779,N_6231);
or U11104 (N_11104,N_7959,N_6951);
and U11105 (N_11105,N_7051,N_7794);
nor U11106 (N_11106,N_6630,N_8571);
nand U11107 (N_11107,N_7320,N_7634);
and U11108 (N_11108,N_8245,N_8889);
nor U11109 (N_11109,N_7724,N_8518);
or U11110 (N_11110,N_8992,N_6679);
nor U11111 (N_11111,N_6393,N_8028);
or U11112 (N_11112,N_7275,N_8567);
or U11113 (N_11113,N_6677,N_7482);
nand U11114 (N_11114,N_8968,N_8212);
nand U11115 (N_11115,N_6087,N_8057);
nor U11116 (N_11116,N_6022,N_8757);
nand U11117 (N_11117,N_8594,N_6004);
or U11118 (N_11118,N_8913,N_6621);
nor U11119 (N_11119,N_8320,N_6009);
nand U11120 (N_11120,N_7686,N_6617);
nand U11121 (N_11121,N_7884,N_8724);
or U11122 (N_11122,N_7562,N_8495);
nor U11123 (N_11123,N_6477,N_6369);
nand U11124 (N_11124,N_8147,N_6155);
or U11125 (N_11125,N_7183,N_8821);
and U11126 (N_11126,N_6042,N_6297);
or U11127 (N_11127,N_6947,N_6407);
nand U11128 (N_11128,N_6947,N_6249);
nor U11129 (N_11129,N_6636,N_7383);
nand U11130 (N_11130,N_7408,N_8632);
nor U11131 (N_11131,N_6418,N_6133);
and U11132 (N_11132,N_7596,N_7353);
nor U11133 (N_11133,N_8401,N_6488);
nand U11134 (N_11134,N_6791,N_6720);
or U11135 (N_11135,N_6222,N_8647);
and U11136 (N_11136,N_7026,N_8176);
nor U11137 (N_11137,N_8576,N_8799);
or U11138 (N_11138,N_6058,N_6147);
and U11139 (N_11139,N_6716,N_6213);
nor U11140 (N_11140,N_7636,N_8808);
or U11141 (N_11141,N_8415,N_6600);
or U11142 (N_11142,N_6483,N_7199);
or U11143 (N_11143,N_7212,N_7819);
nor U11144 (N_11144,N_7070,N_7300);
nor U11145 (N_11145,N_7584,N_8910);
or U11146 (N_11146,N_8996,N_7747);
nand U11147 (N_11147,N_7020,N_7034);
and U11148 (N_11148,N_7255,N_8150);
nor U11149 (N_11149,N_8135,N_8239);
or U11150 (N_11150,N_7471,N_6503);
and U11151 (N_11151,N_8869,N_7298);
nand U11152 (N_11152,N_8713,N_8339);
nor U11153 (N_11153,N_7180,N_8000);
or U11154 (N_11154,N_7805,N_8380);
nor U11155 (N_11155,N_8836,N_6705);
or U11156 (N_11156,N_6383,N_7033);
or U11157 (N_11157,N_6570,N_8279);
nor U11158 (N_11158,N_7364,N_8316);
nor U11159 (N_11159,N_6936,N_7457);
nand U11160 (N_11160,N_6577,N_7237);
and U11161 (N_11161,N_6718,N_8789);
nor U11162 (N_11162,N_8342,N_8454);
and U11163 (N_11163,N_6307,N_6453);
nand U11164 (N_11164,N_6037,N_8453);
nor U11165 (N_11165,N_7274,N_8900);
nor U11166 (N_11166,N_7535,N_8894);
nand U11167 (N_11167,N_8190,N_6008);
and U11168 (N_11168,N_6402,N_8074);
and U11169 (N_11169,N_6034,N_8012);
nand U11170 (N_11170,N_8129,N_8840);
and U11171 (N_11171,N_8616,N_6968);
or U11172 (N_11172,N_8015,N_7586);
nand U11173 (N_11173,N_8628,N_7253);
nand U11174 (N_11174,N_6521,N_7165);
and U11175 (N_11175,N_6087,N_7612);
nor U11176 (N_11176,N_7507,N_7837);
nand U11177 (N_11177,N_6469,N_8376);
nor U11178 (N_11178,N_6125,N_7777);
and U11179 (N_11179,N_7596,N_7148);
or U11180 (N_11180,N_8637,N_8973);
nor U11181 (N_11181,N_6944,N_7004);
or U11182 (N_11182,N_6233,N_7379);
nor U11183 (N_11183,N_7143,N_6546);
nor U11184 (N_11184,N_7763,N_8669);
and U11185 (N_11185,N_7705,N_6485);
nor U11186 (N_11186,N_7524,N_6446);
or U11187 (N_11187,N_6755,N_7796);
nor U11188 (N_11188,N_8178,N_6237);
nand U11189 (N_11189,N_6647,N_8333);
and U11190 (N_11190,N_6781,N_8228);
nand U11191 (N_11191,N_6947,N_6199);
nand U11192 (N_11192,N_8403,N_6962);
nand U11193 (N_11193,N_8665,N_7328);
nor U11194 (N_11194,N_6747,N_7141);
or U11195 (N_11195,N_8342,N_6553);
nor U11196 (N_11196,N_7087,N_8135);
xor U11197 (N_11197,N_6298,N_6129);
or U11198 (N_11198,N_7219,N_7037);
nor U11199 (N_11199,N_6330,N_6020);
nand U11200 (N_11200,N_7425,N_7209);
or U11201 (N_11201,N_8650,N_6592);
and U11202 (N_11202,N_8251,N_8815);
or U11203 (N_11203,N_7450,N_6934);
nand U11204 (N_11204,N_7979,N_7376);
nand U11205 (N_11205,N_7760,N_6029);
and U11206 (N_11206,N_8660,N_6206);
and U11207 (N_11207,N_8828,N_8631);
and U11208 (N_11208,N_6824,N_6356);
nor U11209 (N_11209,N_7358,N_8680);
nand U11210 (N_11210,N_6903,N_6590);
nand U11211 (N_11211,N_6388,N_8181);
and U11212 (N_11212,N_7506,N_8259);
nand U11213 (N_11213,N_6941,N_6376);
and U11214 (N_11214,N_8601,N_7505);
and U11215 (N_11215,N_8163,N_7243);
nor U11216 (N_11216,N_7874,N_8077);
nand U11217 (N_11217,N_6563,N_7493);
or U11218 (N_11218,N_7837,N_6003);
and U11219 (N_11219,N_7340,N_6160);
and U11220 (N_11220,N_7525,N_7388);
nand U11221 (N_11221,N_8021,N_7583);
or U11222 (N_11222,N_8656,N_7069);
nor U11223 (N_11223,N_8657,N_8588);
and U11224 (N_11224,N_6299,N_7567);
nand U11225 (N_11225,N_7602,N_6000);
or U11226 (N_11226,N_7247,N_6972);
nor U11227 (N_11227,N_8932,N_6135);
nor U11228 (N_11228,N_8871,N_7144);
nand U11229 (N_11229,N_7383,N_6224);
nand U11230 (N_11230,N_7020,N_7019);
xor U11231 (N_11231,N_8062,N_7916);
nor U11232 (N_11232,N_6184,N_8848);
and U11233 (N_11233,N_7775,N_8286);
nand U11234 (N_11234,N_6829,N_8027);
nand U11235 (N_11235,N_8285,N_6186);
nand U11236 (N_11236,N_8800,N_8877);
or U11237 (N_11237,N_7967,N_7707);
or U11238 (N_11238,N_8723,N_8138);
and U11239 (N_11239,N_6774,N_7554);
nand U11240 (N_11240,N_7066,N_7232);
and U11241 (N_11241,N_7115,N_7258);
nand U11242 (N_11242,N_6992,N_6836);
nor U11243 (N_11243,N_8684,N_7387);
nand U11244 (N_11244,N_7784,N_8641);
nor U11245 (N_11245,N_6438,N_6716);
nor U11246 (N_11246,N_8888,N_8143);
nor U11247 (N_11247,N_6156,N_7258);
or U11248 (N_11248,N_7388,N_7731);
nand U11249 (N_11249,N_6474,N_7259);
xor U11250 (N_11250,N_7205,N_6101);
or U11251 (N_11251,N_7516,N_7145);
and U11252 (N_11252,N_6137,N_7587);
nand U11253 (N_11253,N_8131,N_8414);
or U11254 (N_11254,N_6485,N_6349);
and U11255 (N_11255,N_7004,N_7390);
and U11256 (N_11256,N_8742,N_7236);
nand U11257 (N_11257,N_7806,N_8764);
nand U11258 (N_11258,N_6616,N_6624);
or U11259 (N_11259,N_7462,N_7833);
or U11260 (N_11260,N_8656,N_6868);
nand U11261 (N_11261,N_8538,N_6844);
or U11262 (N_11262,N_6901,N_7367);
and U11263 (N_11263,N_7879,N_7188);
nor U11264 (N_11264,N_8204,N_8254);
and U11265 (N_11265,N_8535,N_6808);
nand U11266 (N_11266,N_8592,N_6593);
and U11267 (N_11267,N_6018,N_8459);
nand U11268 (N_11268,N_8742,N_6530);
or U11269 (N_11269,N_7199,N_6654);
or U11270 (N_11270,N_8548,N_6018);
or U11271 (N_11271,N_8368,N_6435);
nand U11272 (N_11272,N_8813,N_7067);
nor U11273 (N_11273,N_8291,N_8482);
and U11274 (N_11274,N_6463,N_6143);
nor U11275 (N_11275,N_7079,N_6406);
nor U11276 (N_11276,N_7728,N_7888);
and U11277 (N_11277,N_8280,N_6942);
nor U11278 (N_11278,N_7634,N_8125);
nor U11279 (N_11279,N_7472,N_7903);
nor U11280 (N_11280,N_8470,N_8293);
nor U11281 (N_11281,N_8564,N_7838);
nor U11282 (N_11282,N_8019,N_6867);
or U11283 (N_11283,N_7901,N_7753);
or U11284 (N_11284,N_6895,N_7474);
and U11285 (N_11285,N_8265,N_7097);
and U11286 (N_11286,N_7281,N_7870);
and U11287 (N_11287,N_7766,N_8833);
or U11288 (N_11288,N_8320,N_7928);
or U11289 (N_11289,N_6508,N_6319);
nand U11290 (N_11290,N_6376,N_8533);
and U11291 (N_11291,N_6629,N_8626);
nand U11292 (N_11292,N_7449,N_7826);
nand U11293 (N_11293,N_8014,N_7364);
and U11294 (N_11294,N_7499,N_8231);
and U11295 (N_11295,N_6517,N_6131);
or U11296 (N_11296,N_7841,N_8150);
and U11297 (N_11297,N_7838,N_8897);
nand U11298 (N_11298,N_6416,N_7497);
nor U11299 (N_11299,N_8075,N_8855);
or U11300 (N_11300,N_6545,N_7145);
nand U11301 (N_11301,N_7100,N_6432);
or U11302 (N_11302,N_7596,N_8530);
nand U11303 (N_11303,N_6463,N_8053);
and U11304 (N_11304,N_7390,N_8718);
and U11305 (N_11305,N_7472,N_8544);
nor U11306 (N_11306,N_6703,N_7396);
nand U11307 (N_11307,N_6414,N_7816);
nor U11308 (N_11308,N_8718,N_8214);
and U11309 (N_11309,N_8218,N_7164);
and U11310 (N_11310,N_8943,N_7419);
nor U11311 (N_11311,N_8767,N_6330);
nor U11312 (N_11312,N_8546,N_6955);
nor U11313 (N_11313,N_6232,N_7546);
or U11314 (N_11314,N_6090,N_8142);
and U11315 (N_11315,N_8416,N_8748);
nor U11316 (N_11316,N_8334,N_6534);
or U11317 (N_11317,N_6405,N_8032);
nor U11318 (N_11318,N_8230,N_6331);
nand U11319 (N_11319,N_6098,N_6970);
or U11320 (N_11320,N_6626,N_7808);
nand U11321 (N_11321,N_6190,N_7571);
or U11322 (N_11322,N_7486,N_6337);
or U11323 (N_11323,N_6682,N_8151);
nor U11324 (N_11324,N_8475,N_7880);
or U11325 (N_11325,N_6826,N_7695);
and U11326 (N_11326,N_8110,N_8411);
or U11327 (N_11327,N_8691,N_8073);
nor U11328 (N_11328,N_7836,N_8070);
and U11329 (N_11329,N_7146,N_7871);
nand U11330 (N_11330,N_8161,N_7869);
and U11331 (N_11331,N_8796,N_6444);
and U11332 (N_11332,N_8328,N_6581);
and U11333 (N_11333,N_6137,N_8078);
or U11334 (N_11334,N_7039,N_6138);
nand U11335 (N_11335,N_6770,N_6500);
or U11336 (N_11336,N_6628,N_8228);
or U11337 (N_11337,N_7723,N_8965);
or U11338 (N_11338,N_8703,N_8507);
or U11339 (N_11339,N_6713,N_7481);
xnor U11340 (N_11340,N_6640,N_7939);
or U11341 (N_11341,N_8792,N_6322);
or U11342 (N_11342,N_8734,N_6132);
and U11343 (N_11343,N_8084,N_8144);
and U11344 (N_11344,N_7831,N_8696);
nor U11345 (N_11345,N_7709,N_8931);
nor U11346 (N_11346,N_7644,N_8017);
or U11347 (N_11347,N_7535,N_8976);
and U11348 (N_11348,N_8033,N_6277);
nor U11349 (N_11349,N_8449,N_6728);
or U11350 (N_11350,N_6180,N_6241);
and U11351 (N_11351,N_7543,N_8315);
nor U11352 (N_11352,N_7080,N_6623);
nand U11353 (N_11353,N_8175,N_7383);
nor U11354 (N_11354,N_8389,N_8457);
nor U11355 (N_11355,N_8371,N_8661);
or U11356 (N_11356,N_6093,N_6169);
or U11357 (N_11357,N_8181,N_6294);
nand U11358 (N_11358,N_6960,N_8110);
nand U11359 (N_11359,N_8021,N_7965);
or U11360 (N_11360,N_7936,N_7780);
nor U11361 (N_11361,N_7279,N_6556);
nand U11362 (N_11362,N_7678,N_7762);
and U11363 (N_11363,N_8429,N_7515);
nor U11364 (N_11364,N_8554,N_6149);
nor U11365 (N_11365,N_7414,N_7465);
nand U11366 (N_11366,N_6898,N_7941);
and U11367 (N_11367,N_7827,N_7322);
nand U11368 (N_11368,N_7793,N_6919);
and U11369 (N_11369,N_8751,N_7936);
and U11370 (N_11370,N_6353,N_6681);
nor U11371 (N_11371,N_6535,N_6558);
and U11372 (N_11372,N_7737,N_8874);
nor U11373 (N_11373,N_8567,N_6692);
nor U11374 (N_11374,N_8182,N_7060);
and U11375 (N_11375,N_6164,N_7383);
and U11376 (N_11376,N_7092,N_6561);
nor U11377 (N_11377,N_8724,N_8548);
and U11378 (N_11378,N_7263,N_6298);
or U11379 (N_11379,N_8863,N_6137);
or U11380 (N_11380,N_7411,N_6904);
or U11381 (N_11381,N_6683,N_8451);
nand U11382 (N_11382,N_7410,N_8246);
nor U11383 (N_11383,N_8450,N_8479);
or U11384 (N_11384,N_6470,N_7027);
or U11385 (N_11385,N_6287,N_6941);
nor U11386 (N_11386,N_7385,N_8447);
or U11387 (N_11387,N_8526,N_6553);
nor U11388 (N_11388,N_8345,N_8482);
nor U11389 (N_11389,N_6331,N_6975);
nand U11390 (N_11390,N_8329,N_6256);
nor U11391 (N_11391,N_8946,N_6290);
nor U11392 (N_11392,N_8207,N_7199);
nor U11393 (N_11393,N_8798,N_7407);
and U11394 (N_11394,N_7169,N_6640);
or U11395 (N_11395,N_8367,N_6651);
nor U11396 (N_11396,N_7450,N_7264);
or U11397 (N_11397,N_6587,N_7395);
or U11398 (N_11398,N_8162,N_7131);
nor U11399 (N_11399,N_8230,N_7063);
or U11400 (N_11400,N_8642,N_7909);
nand U11401 (N_11401,N_7996,N_8189);
and U11402 (N_11402,N_7850,N_7900);
and U11403 (N_11403,N_7288,N_7872);
and U11404 (N_11404,N_7970,N_6513);
and U11405 (N_11405,N_7366,N_6777);
nor U11406 (N_11406,N_6258,N_6875);
or U11407 (N_11407,N_6321,N_7543);
nand U11408 (N_11408,N_7624,N_6697);
nor U11409 (N_11409,N_8827,N_7637);
and U11410 (N_11410,N_7309,N_8704);
nand U11411 (N_11411,N_6058,N_8870);
nand U11412 (N_11412,N_6182,N_8254);
nor U11413 (N_11413,N_6243,N_6904);
or U11414 (N_11414,N_8238,N_7722);
nor U11415 (N_11415,N_6315,N_6432);
and U11416 (N_11416,N_8071,N_7768);
and U11417 (N_11417,N_7601,N_7845);
or U11418 (N_11418,N_8482,N_6581);
nand U11419 (N_11419,N_7952,N_6825);
or U11420 (N_11420,N_6328,N_7699);
nand U11421 (N_11421,N_8261,N_7104);
or U11422 (N_11422,N_7602,N_6421);
nand U11423 (N_11423,N_8091,N_8137);
nor U11424 (N_11424,N_7010,N_8771);
nand U11425 (N_11425,N_8705,N_8458);
nand U11426 (N_11426,N_7250,N_6349);
or U11427 (N_11427,N_8392,N_8438);
or U11428 (N_11428,N_7121,N_8089);
or U11429 (N_11429,N_6569,N_8034);
or U11430 (N_11430,N_7175,N_7582);
nor U11431 (N_11431,N_8445,N_8648);
or U11432 (N_11432,N_8621,N_7113);
and U11433 (N_11433,N_7560,N_7625);
and U11434 (N_11434,N_8906,N_8087);
or U11435 (N_11435,N_7359,N_6433);
or U11436 (N_11436,N_8651,N_8918);
nand U11437 (N_11437,N_7012,N_6078);
and U11438 (N_11438,N_7475,N_7891);
nand U11439 (N_11439,N_8246,N_7671);
and U11440 (N_11440,N_8004,N_8024);
nor U11441 (N_11441,N_7857,N_6846);
nor U11442 (N_11442,N_6523,N_8343);
or U11443 (N_11443,N_8745,N_7894);
and U11444 (N_11444,N_7675,N_6407);
nor U11445 (N_11445,N_8301,N_6731);
nor U11446 (N_11446,N_6978,N_6832);
and U11447 (N_11447,N_7989,N_8146);
and U11448 (N_11448,N_7558,N_7225);
nand U11449 (N_11449,N_6874,N_7332);
or U11450 (N_11450,N_8335,N_8809);
nand U11451 (N_11451,N_6401,N_7093);
nor U11452 (N_11452,N_6697,N_7114);
or U11453 (N_11453,N_7985,N_6858);
or U11454 (N_11454,N_7729,N_7943);
nor U11455 (N_11455,N_7684,N_6997);
nand U11456 (N_11456,N_7334,N_6378);
or U11457 (N_11457,N_7126,N_7878);
or U11458 (N_11458,N_8511,N_8467);
and U11459 (N_11459,N_6218,N_7274);
or U11460 (N_11460,N_7800,N_7578);
or U11461 (N_11461,N_8048,N_8060);
or U11462 (N_11462,N_6204,N_6427);
and U11463 (N_11463,N_6453,N_6140);
or U11464 (N_11464,N_8869,N_6965);
nand U11465 (N_11465,N_8807,N_8462);
nand U11466 (N_11466,N_8621,N_6333);
or U11467 (N_11467,N_7940,N_6886);
nand U11468 (N_11468,N_6068,N_7660);
or U11469 (N_11469,N_8813,N_7191);
or U11470 (N_11470,N_7989,N_7164);
nor U11471 (N_11471,N_7584,N_6578);
nor U11472 (N_11472,N_7935,N_6779);
nor U11473 (N_11473,N_8813,N_8265);
nand U11474 (N_11474,N_8276,N_6122);
xor U11475 (N_11475,N_7707,N_8039);
and U11476 (N_11476,N_6060,N_8505);
nand U11477 (N_11477,N_8139,N_6131);
nand U11478 (N_11478,N_8509,N_8176);
or U11479 (N_11479,N_6286,N_8690);
nor U11480 (N_11480,N_7194,N_7459);
nor U11481 (N_11481,N_7148,N_6834);
and U11482 (N_11482,N_8905,N_6075);
nor U11483 (N_11483,N_6946,N_6630);
nor U11484 (N_11484,N_6706,N_6796);
nand U11485 (N_11485,N_6887,N_7333);
and U11486 (N_11486,N_7846,N_7309);
and U11487 (N_11487,N_8127,N_6174);
and U11488 (N_11488,N_7857,N_8536);
and U11489 (N_11489,N_8835,N_7428);
nand U11490 (N_11490,N_8540,N_8196);
nand U11491 (N_11491,N_6068,N_7512);
nand U11492 (N_11492,N_8010,N_8982);
or U11493 (N_11493,N_7830,N_6752);
or U11494 (N_11494,N_6429,N_8832);
or U11495 (N_11495,N_6289,N_6651);
nand U11496 (N_11496,N_8296,N_6771);
nor U11497 (N_11497,N_7250,N_8285);
nor U11498 (N_11498,N_8104,N_7209);
xor U11499 (N_11499,N_8032,N_8501);
and U11500 (N_11500,N_6157,N_6132);
or U11501 (N_11501,N_6318,N_6691);
and U11502 (N_11502,N_6331,N_8708);
and U11503 (N_11503,N_7467,N_6900);
nand U11504 (N_11504,N_6687,N_7606);
and U11505 (N_11505,N_8147,N_7668);
nand U11506 (N_11506,N_7566,N_7920);
and U11507 (N_11507,N_8366,N_8229);
and U11508 (N_11508,N_8586,N_7832);
nand U11509 (N_11509,N_7709,N_6725);
and U11510 (N_11510,N_8040,N_7878);
nor U11511 (N_11511,N_7795,N_7181);
and U11512 (N_11512,N_8114,N_7247);
nor U11513 (N_11513,N_7530,N_8489);
nand U11514 (N_11514,N_6101,N_7754);
or U11515 (N_11515,N_7099,N_7671);
or U11516 (N_11516,N_8971,N_6033);
or U11517 (N_11517,N_7066,N_6058);
and U11518 (N_11518,N_6703,N_8191);
xor U11519 (N_11519,N_7365,N_7769);
and U11520 (N_11520,N_6937,N_7835);
and U11521 (N_11521,N_7604,N_8769);
nor U11522 (N_11522,N_8538,N_8839);
nor U11523 (N_11523,N_6365,N_7079);
and U11524 (N_11524,N_8634,N_8096);
nor U11525 (N_11525,N_7833,N_7134);
nand U11526 (N_11526,N_6471,N_6948);
and U11527 (N_11527,N_6933,N_8886);
nor U11528 (N_11528,N_8500,N_6691);
nor U11529 (N_11529,N_6627,N_8370);
nand U11530 (N_11530,N_6166,N_6868);
nor U11531 (N_11531,N_8547,N_8288);
or U11532 (N_11532,N_7002,N_7510);
xor U11533 (N_11533,N_7152,N_7113);
or U11534 (N_11534,N_7853,N_6142);
nand U11535 (N_11535,N_8634,N_7538);
or U11536 (N_11536,N_6017,N_7154);
and U11537 (N_11537,N_7313,N_6973);
or U11538 (N_11538,N_8523,N_8772);
nand U11539 (N_11539,N_8333,N_6574);
nand U11540 (N_11540,N_8901,N_8292);
and U11541 (N_11541,N_8755,N_8235);
nand U11542 (N_11542,N_6543,N_7863);
nor U11543 (N_11543,N_8504,N_8432);
and U11544 (N_11544,N_6036,N_8757);
nor U11545 (N_11545,N_6408,N_7601);
or U11546 (N_11546,N_8617,N_7708);
or U11547 (N_11547,N_7783,N_7801);
and U11548 (N_11548,N_6898,N_8233);
or U11549 (N_11549,N_8069,N_6566);
nor U11550 (N_11550,N_6967,N_7953);
nor U11551 (N_11551,N_6396,N_7566);
or U11552 (N_11552,N_6715,N_8209);
and U11553 (N_11553,N_8289,N_7434);
nor U11554 (N_11554,N_6037,N_6965);
or U11555 (N_11555,N_6773,N_6252);
nand U11556 (N_11556,N_6977,N_8501);
nor U11557 (N_11557,N_6932,N_7831);
and U11558 (N_11558,N_7263,N_6167);
nor U11559 (N_11559,N_8399,N_8203);
and U11560 (N_11560,N_6166,N_8296);
nor U11561 (N_11561,N_6186,N_6511);
nor U11562 (N_11562,N_8268,N_8157);
nor U11563 (N_11563,N_7011,N_7360);
and U11564 (N_11564,N_8066,N_6929);
nor U11565 (N_11565,N_8389,N_7761);
nor U11566 (N_11566,N_8189,N_7549);
nand U11567 (N_11567,N_8519,N_7834);
or U11568 (N_11568,N_6159,N_8341);
or U11569 (N_11569,N_6354,N_7500);
and U11570 (N_11570,N_7750,N_6872);
or U11571 (N_11571,N_8006,N_7776);
nand U11572 (N_11572,N_7500,N_7609);
nand U11573 (N_11573,N_6355,N_6091);
nor U11574 (N_11574,N_8603,N_6625);
and U11575 (N_11575,N_8348,N_8862);
or U11576 (N_11576,N_8514,N_6750);
or U11577 (N_11577,N_8111,N_7831);
or U11578 (N_11578,N_6940,N_7297);
and U11579 (N_11579,N_7133,N_6133);
and U11580 (N_11580,N_6915,N_8939);
nand U11581 (N_11581,N_8922,N_8023);
nor U11582 (N_11582,N_6445,N_7199);
xor U11583 (N_11583,N_8930,N_6023);
nand U11584 (N_11584,N_7617,N_7592);
nor U11585 (N_11585,N_6720,N_7866);
nor U11586 (N_11586,N_8955,N_8754);
nand U11587 (N_11587,N_8566,N_8896);
and U11588 (N_11588,N_6961,N_8498);
and U11589 (N_11589,N_7507,N_7868);
nand U11590 (N_11590,N_7412,N_8123);
nor U11591 (N_11591,N_8167,N_6536);
nand U11592 (N_11592,N_8758,N_6876);
and U11593 (N_11593,N_8818,N_7008);
nand U11594 (N_11594,N_6038,N_6711);
nor U11595 (N_11595,N_8153,N_7339);
nor U11596 (N_11596,N_7328,N_7231);
or U11597 (N_11597,N_8777,N_7918);
and U11598 (N_11598,N_6143,N_6507);
or U11599 (N_11599,N_6047,N_7787);
and U11600 (N_11600,N_6209,N_7803);
and U11601 (N_11601,N_8888,N_6652);
and U11602 (N_11602,N_7736,N_8866);
or U11603 (N_11603,N_8131,N_6946);
nor U11604 (N_11604,N_8652,N_6991);
or U11605 (N_11605,N_6196,N_8230);
or U11606 (N_11606,N_8784,N_6321);
nor U11607 (N_11607,N_8160,N_6449);
nand U11608 (N_11608,N_8857,N_7464);
or U11609 (N_11609,N_7804,N_8305);
nand U11610 (N_11610,N_6807,N_6826);
xor U11611 (N_11611,N_8519,N_8817);
and U11612 (N_11612,N_6313,N_8849);
or U11613 (N_11613,N_7830,N_7385);
and U11614 (N_11614,N_8812,N_6199);
nor U11615 (N_11615,N_7887,N_7192);
and U11616 (N_11616,N_8419,N_6708);
or U11617 (N_11617,N_6831,N_6929);
nor U11618 (N_11618,N_8816,N_6604);
nand U11619 (N_11619,N_7678,N_8214);
nor U11620 (N_11620,N_6075,N_6905);
nor U11621 (N_11621,N_7243,N_8132);
or U11622 (N_11622,N_6843,N_7167);
nor U11623 (N_11623,N_6303,N_8588);
nor U11624 (N_11624,N_6092,N_7632);
or U11625 (N_11625,N_8159,N_6162);
and U11626 (N_11626,N_6947,N_6023);
and U11627 (N_11627,N_7569,N_7008);
or U11628 (N_11628,N_6164,N_6716);
nor U11629 (N_11629,N_7883,N_6240);
and U11630 (N_11630,N_7900,N_7937);
and U11631 (N_11631,N_8678,N_8221);
nor U11632 (N_11632,N_8040,N_6227);
or U11633 (N_11633,N_8356,N_8371);
or U11634 (N_11634,N_6106,N_6793);
and U11635 (N_11635,N_8514,N_8637);
nand U11636 (N_11636,N_7353,N_7483);
nand U11637 (N_11637,N_6465,N_6658);
and U11638 (N_11638,N_7617,N_8504);
and U11639 (N_11639,N_6188,N_6656);
nand U11640 (N_11640,N_6639,N_8271);
nor U11641 (N_11641,N_8574,N_8322);
nor U11642 (N_11642,N_8536,N_7145);
nor U11643 (N_11643,N_7274,N_7808);
nand U11644 (N_11644,N_8253,N_6869);
nand U11645 (N_11645,N_8303,N_7909);
and U11646 (N_11646,N_6911,N_8795);
nor U11647 (N_11647,N_7397,N_8594);
and U11648 (N_11648,N_6445,N_7779);
nand U11649 (N_11649,N_7736,N_6305);
nor U11650 (N_11650,N_7305,N_7757);
nand U11651 (N_11651,N_6561,N_7105);
nor U11652 (N_11652,N_7103,N_8611);
nor U11653 (N_11653,N_7741,N_6259);
and U11654 (N_11654,N_7387,N_8718);
nor U11655 (N_11655,N_8446,N_8756);
nor U11656 (N_11656,N_7210,N_8085);
or U11657 (N_11657,N_6155,N_7272);
nor U11658 (N_11658,N_6151,N_7866);
and U11659 (N_11659,N_8491,N_6145);
nand U11660 (N_11660,N_7051,N_7673);
nand U11661 (N_11661,N_8617,N_6213);
or U11662 (N_11662,N_7820,N_7737);
nand U11663 (N_11663,N_8846,N_8460);
and U11664 (N_11664,N_7900,N_8713);
nand U11665 (N_11665,N_6030,N_8686);
nor U11666 (N_11666,N_6072,N_6843);
or U11667 (N_11667,N_8785,N_8141);
nand U11668 (N_11668,N_6119,N_6224);
nor U11669 (N_11669,N_8702,N_7387);
nor U11670 (N_11670,N_6583,N_7290);
nand U11671 (N_11671,N_7236,N_8203);
or U11672 (N_11672,N_8064,N_6079);
nor U11673 (N_11673,N_8822,N_6257);
nor U11674 (N_11674,N_7137,N_8689);
nand U11675 (N_11675,N_8420,N_7786);
and U11676 (N_11676,N_7944,N_7859);
and U11677 (N_11677,N_8682,N_8923);
nand U11678 (N_11678,N_7189,N_7231);
nor U11679 (N_11679,N_8336,N_6540);
and U11680 (N_11680,N_8077,N_7510);
nand U11681 (N_11681,N_7359,N_6070);
or U11682 (N_11682,N_6933,N_6581);
and U11683 (N_11683,N_6949,N_8122);
or U11684 (N_11684,N_7496,N_8523);
and U11685 (N_11685,N_6280,N_7577);
nor U11686 (N_11686,N_8582,N_6942);
and U11687 (N_11687,N_8136,N_7613);
and U11688 (N_11688,N_6233,N_6054);
nor U11689 (N_11689,N_7242,N_8705);
and U11690 (N_11690,N_8398,N_7771);
and U11691 (N_11691,N_7072,N_6866);
nor U11692 (N_11692,N_8956,N_8593);
nor U11693 (N_11693,N_7020,N_8301);
and U11694 (N_11694,N_8679,N_6871);
nand U11695 (N_11695,N_7644,N_6869);
and U11696 (N_11696,N_6028,N_7446);
nor U11697 (N_11697,N_6283,N_7743);
or U11698 (N_11698,N_8817,N_6674);
nand U11699 (N_11699,N_7969,N_8238);
and U11700 (N_11700,N_8892,N_7876);
or U11701 (N_11701,N_8467,N_7754);
and U11702 (N_11702,N_8070,N_8756);
and U11703 (N_11703,N_7840,N_7493);
and U11704 (N_11704,N_8960,N_8740);
nand U11705 (N_11705,N_8138,N_6370);
and U11706 (N_11706,N_6171,N_6576);
or U11707 (N_11707,N_8906,N_7135);
nand U11708 (N_11708,N_7344,N_6383);
nor U11709 (N_11709,N_7853,N_7740);
nor U11710 (N_11710,N_8010,N_6280);
or U11711 (N_11711,N_7948,N_8625);
or U11712 (N_11712,N_8081,N_8524);
nor U11713 (N_11713,N_8238,N_6883);
or U11714 (N_11714,N_7647,N_8558);
or U11715 (N_11715,N_8737,N_7671);
or U11716 (N_11716,N_7579,N_8096);
and U11717 (N_11717,N_8419,N_7761);
or U11718 (N_11718,N_6692,N_8710);
nor U11719 (N_11719,N_7229,N_6000);
and U11720 (N_11720,N_8754,N_7178);
and U11721 (N_11721,N_8971,N_8486);
nor U11722 (N_11722,N_6831,N_8685);
and U11723 (N_11723,N_8734,N_8486);
or U11724 (N_11724,N_7661,N_6961);
or U11725 (N_11725,N_8993,N_8601);
and U11726 (N_11726,N_6372,N_7172);
and U11727 (N_11727,N_8871,N_7190);
or U11728 (N_11728,N_8590,N_6758);
or U11729 (N_11729,N_8279,N_7761);
nor U11730 (N_11730,N_7957,N_8155);
nor U11731 (N_11731,N_8558,N_6831);
nand U11732 (N_11732,N_8054,N_6582);
nand U11733 (N_11733,N_8684,N_8165);
and U11734 (N_11734,N_6488,N_8053);
nor U11735 (N_11735,N_6891,N_7667);
nor U11736 (N_11736,N_7544,N_7518);
and U11737 (N_11737,N_7364,N_7812);
nor U11738 (N_11738,N_8864,N_7083);
and U11739 (N_11739,N_7076,N_6031);
nand U11740 (N_11740,N_8517,N_8259);
or U11741 (N_11741,N_6420,N_7110);
and U11742 (N_11742,N_7997,N_8463);
nand U11743 (N_11743,N_7661,N_6073);
xnor U11744 (N_11744,N_7292,N_8674);
and U11745 (N_11745,N_7325,N_6461);
or U11746 (N_11746,N_7907,N_8197);
and U11747 (N_11747,N_6862,N_8736);
or U11748 (N_11748,N_8831,N_8402);
or U11749 (N_11749,N_7121,N_6916);
and U11750 (N_11750,N_6262,N_8058);
nor U11751 (N_11751,N_6277,N_7131);
nor U11752 (N_11752,N_7050,N_6520);
and U11753 (N_11753,N_8600,N_8896);
and U11754 (N_11754,N_6626,N_7553);
nor U11755 (N_11755,N_6018,N_6187);
nor U11756 (N_11756,N_7279,N_8119);
nand U11757 (N_11757,N_7120,N_6932);
and U11758 (N_11758,N_7562,N_6053);
or U11759 (N_11759,N_7484,N_8234);
nor U11760 (N_11760,N_8791,N_7779);
nor U11761 (N_11761,N_7893,N_6809);
and U11762 (N_11762,N_6037,N_7481);
or U11763 (N_11763,N_6019,N_6210);
nor U11764 (N_11764,N_6024,N_8285);
or U11765 (N_11765,N_7343,N_7805);
or U11766 (N_11766,N_8003,N_7245);
or U11767 (N_11767,N_8819,N_6353);
nand U11768 (N_11768,N_7932,N_7410);
or U11769 (N_11769,N_7620,N_8318);
nand U11770 (N_11770,N_6907,N_6860);
nor U11771 (N_11771,N_8200,N_8265);
and U11772 (N_11772,N_8464,N_6622);
or U11773 (N_11773,N_8037,N_7130);
or U11774 (N_11774,N_7049,N_6307);
and U11775 (N_11775,N_6374,N_7633);
and U11776 (N_11776,N_6248,N_8102);
or U11777 (N_11777,N_8485,N_8503);
and U11778 (N_11778,N_7607,N_8309);
and U11779 (N_11779,N_7980,N_6333);
nand U11780 (N_11780,N_8127,N_6863);
and U11781 (N_11781,N_7402,N_7728);
or U11782 (N_11782,N_8406,N_8305);
nand U11783 (N_11783,N_6721,N_7170);
nand U11784 (N_11784,N_7712,N_8312);
or U11785 (N_11785,N_6889,N_6040);
nor U11786 (N_11786,N_6093,N_6039);
nand U11787 (N_11787,N_7924,N_8697);
or U11788 (N_11788,N_8814,N_8744);
and U11789 (N_11789,N_8972,N_7426);
nor U11790 (N_11790,N_8782,N_6102);
nand U11791 (N_11791,N_7948,N_7960);
nand U11792 (N_11792,N_6348,N_7154);
nand U11793 (N_11793,N_8599,N_7112);
nor U11794 (N_11794,N_6559,N_6463);
xor U11795 (N_11795,N_7798,N_7614);
and U11796 (N_11796,N_8341,N_7409);
and U11797 (N_11797,N_8744,N_6132);
nor U11798 (N_11798,N_6423,N_6586);
or U11799 (N_11799,N_7949,N_7616);
nor U11800 (N_11800,N_7025,N_6363);
and U11801 (N_11801,N_8734,N_6819);
or U11802 (N_11802,N_6727,N_8545);
and U11803 (N_11803,N_6385,N_6196);
nor U11804 (N_11804,N_8557,N_8878);
nor U11805 (N_11805,N_8726,N_8845);
nand U11806 (N_11806,N_7502,N_7428);
nor U11807 (N_11807,N_6374,N_7594);
xor U11808 (N_11808,N_7187,N_8998);
and U11809 (N_11809,N_8454,N_8035);
nand U11810 (N_11810,N_6183,N_6158);
nand U11811 (N_11811,N_7920,N_8503);
and U11812 (N_11812,N_7059,N_6502);
nand U11813 (N_11813,N_8561,N_6808);
and U11814 (N_11814,N_6911,N_7992);
nand U11815 (N_11815,N_7323,N_8770);
and U11816 (N_11816,N_6538,N_7537);
or U11817 (N_11817,N_8964,N_7637);
nor U11818 (N_11818,N_7360,N_7671);
nor U11819 (N_11819,N_6608,N_8305);
or U11820 (N_11820,N_8307,N_6411);
or U11821 (N_11821,N_7044,N_8564);
nor U11822 (N_11822,N_8542,N_8581);
nor U11823 (N_11823,N_8929,N_8199);
nor U11824 (N_11824,N_6991,N_8207);
or U11825 (N_11825,N_7088,N_8598);
nand U11826 (N_11826,N_7378,N_6538);
nor U11827 (N_11827,N_7600,N_6507);
nand U11828 (N_11828,N_8971,N_8968);
nor U11829 (N_11829,N_8791,N_8884);
nand U11830 (N_11830,N_8314,N_7236);
and U11831 (N_11831,N_8529,N_8708);
and U11832 (N_11832,N_6787,N_7295);
nor U11833 (N_11833,N_6960,N_7130);
nor U11834 (N_11834,N_7862,N_7348);
nand U11835 (N_11835,N_8088,N_6742);
nand U11836 (N_11836,N_7242,N_8014);
and U11837 (N_11837,N_8334,N_8732);
or U11838 (N_11838,N_6446,N_7226);
and U11839 (N_11839,N_8800,N_8246);
nand U11840 (N_11840,N_7644,N_7581);
and U11841 (N_11841,N_6376,N_6840);
nor U11842 (N_11842,N_6918,N_8379);
or U11843 (N_11843,N_6390,N_8112);
nand U11844 (N_11844,N_7718,N_7016);
nand U11845 (N_11845,N_6212,N_8357);
or U11846 (N_11846,N_7066,N_8555);
or U11847 (N_11847,N_6050,N_8706);
or U11848 (N_11848,N_8714,N_8577);
and U11849 (N_11849,N_6610,N_7047);
nand U11850 (N_11850,N_7272,N_8599);
or U11851 (N_11851,N_7629,N_6456);
or U11852 (N_11852,N_6836,N_8481);
or U11853 (N_11853,N_8716,N_8114);
nand U11854 (N_11854,N_8460,N_6270);
nor U11855 (N_11855,N_8390,N_8093);
or U11856 (N_11856,N_6086,N_8298);
or U11857 (N_11857,N_8389,N_8154);
or U11858 (N_11858,N_8550,N_6578);
nand U11859 (N_11859,N_8632,N_8140);
or U11860 (N_11860,N_6918,N_6646);
nor U11861 (N_11861,N_7964,N_7335);
nor U11862 (N_11862,N_7597,N_8171);
or U11863 (N_11863,N_7997,N_8740);
and U11864 (N_11864,N_6687,N_8733);
nor U11865 (N_11865,N_7918,N_6487);
nand U11866 (N_11866,N_6449,N_6918);
nor U11867 (N_11867,N_7573,N_7605);
nor U11868 (N_11868,N_8131,N_8174);
or U11869 (N_11869,N_6913,N_8369);
nand U11870 (N_11870,N_8392,N_8650);
nand U11871 (N_11871,N_8271,N_6194);
or U11872 (N_11872,N_7894,N_6620);
or U11873 (N_11873,N_6572,N_8384);
nor U11874 (N_11874,N_7138,N_6278);
nor U11875 (N_11875,N_6663,N_7472);
nor U11876 (N_11876,N_8075,N_6303);
nor U11877 (N_11877,N_7345,N_8872);
nor U11878 (N_11878,N_8369,N_7953);
nor U11879 (N_11879,N_6502,N_6621);
nand U11880 (N_11880,N_6483,N_8637);
and U11881 (N_11881,N_6421,N_6341);
and U11882 (N_11882,N_7656,N_7351);
or U11883 (N_11883,N_7583,N_6408);
or U11884 (N_11884,N_6430,N_7171);
nand U11885 (N_11885,N_8560,N_7260);
nand U11886 (N_11886,N_6905,N_7573);
nor U11887 (N_11887,N_7443,N_7936);
nor U11888 (N_11888,N_6374,N_7105);
nand U11889 (N_11889,N_7469,N_7542);
and U11890 (N_11890,N_8456,N_6308);
nand U11891 (N_11891,N_6854,N_7486);
nor U11892 (N_11892,N_7033,N_6824);
nor U11893 (N_11893,N_6419,N_7940);
and U11894 (N_11894,N_7954,N_8492);
and U11895 (N_11895,N_6998,N_7128);
nand U11896 (N_11896,N_6047,N_7328);
nand U11897 (N_11897,N_8960,N_6106);
nor U11898 (N_11898,N_6118,N_7266);
or U11899 (N_11899,N_8876,N_8573);
nand U11900 (N_11900,N_8873,N_7202);
nand U11901 (N_11901,N_7465,N_8469);
nor U11902 (N_11902,N_7648,N_7001);
and U11903 (N_11903,N_7256,N_6864);
nor U11904 (N_11904,N_8641,N_8700);
or U11905 (N_11905,N_7296,N_8814);
or U11906 (N_11906,N_7942,N_6168);
or U11907 (N_11907,N_7745,N_6186);
or U11908 (N_11908,N_8300,N_7550);
or U11909 (N_11909,N_7069,N_8009);
nor U11910 (N_11910,N_8153,N_6004);
nand U11911 (N_11911,N_8343,N_8599);
and U11912 (N_11912,N_6149,N_6645);
nor U11913 (N_11913,N_7979,N_6913);
nand U11914 (N_11914,N_6461,N_8797);
or U11915 (N_11915,N_8200,N_8927);
and U11916 (N_11916,N_7405,N_6077);
or U11917 (N_11917,N_7602,N_6255);
or U11918 (N_11918,N_6357,N_8426);
and U11919 (N_11919,N_7884,N_6309);
or U11920 (N_11920,N_8125,N_8677);
nand U11921 (N_11921,N_8043,N_7788);
or U11922 (N_11922,N_6953,N_7388);
or U11923 (N_11923,N_8877,N_6848);
or U11924 (N_11924,N_6686,N_8195);
nand U11925 (N_11925,N_8358,N_6234);
and U11926 (N_11926,N_8670,N_8003);
nor U11927 (N_11927,N_6150,N_6077);
nand U11928 (N_11928,N_7251,N_7753);
nand U11929 (N_11929,N_7114,N_6842);
and U11930 (N_11930,N_8689,N_7904);
or U11931 (N_11931,N_8903,N_6945);
nor U11932 (N_11932,N_8866,N_6675);
and U11933 (N_11933,N_8900,N_8514);
or U11934 (N_11934,N_7686,N_8223);
and U11935 (N_11935,N_6298,N_6102);
nor U11936 (N_11936,N_8745,N_8348);
nor U11937 (N_11937,N_8101,N_6093);
nand U11938 (N_11938,N_6411,N_7113);
or U11939 (N_11939,N_8961,N_6970);
nor U11940 (N_11940,N_6972,N_6613);
or U11941 (N_11941,N_7692,N_8247);
nor U11942 (N_11942,N_7463,N_7715);
nor U11943 (N_11943,N_6390,N_7667);
and U11944 (N_11944,N_6988,N_6713);
or U11945 (N_11945,N_8683,N_6726);
and U11946 (N_11946,N_7156,N_8433);
and U11947 (N_11947,N_8842,N_7718);
and U11948 (N_11948,N_8750,N_6534);
or U11949 (N_11949,N_8708,N_6048);
nand U11950 (N_11950,N_7235,N_8246);
nand U11951 (N_11951,N_6517,N_6453);
or U11952 (N_11952,N_7476,N_7597);
nand U11953 (N_11953,N_7447,N_7118);
nor U11954 (N_11954,N_6782,N_7934);
or U11955 (N_11955,N_7642,N_6763);
nand U11956 (N_11956,N_8859,N_7843);
nor U11957 (N_11957,N_6700,N_8803);
or U11958 (N_11958,N_7854,N_7447);
or U11959 (N_11959,N_8696,N_6809);
xnor U11960 (N_11960,N_6750,N_6493);
or U11961 (N_11961,N_8998,N_6588);
and U11962 (N_11962,N_8893,N_7968);
nor U11963 (N_11963,N_8809,N_6591);
nor U11964 (N_11964,N_7946,N_8054);
or U11965 (N_11965,N_6614,N_7980);
or U11966 (N_11966,N_7963,N_6546);
or U11967 (N_11967,N_8049,N_8417);
nor U11968 (N_11968,N_7592,N_8186);
or U11969 (N_11969,N_7645,N_8639);
nand U11970 (N_11970,N_6509,N_7932);
and U11971 (N_11971,N_6716,N_6033);
nor U11972 (N_11972,N_6436,N_8869);
and U11973 (N_11973,N_6551,N_8755);
or U11974 (N_11974,N_8137,N_6803);
or U11975 (N_11975,N_6429,N_8206);
nor U11976 (N_11976,N_8222,N_6293);
nand U11977 (N_11977,N_8872,N_6734);
nor U11978 (N_11978,N_7308,N_6550);
nor U11979 (N_11979,N_7239,N_7142);
nand U11980 (N_11980,N_7531,N_6237);
or U11981 (N_11981,N_8933,N_6488);
or U11982 (N_11982,N_7552,N_6201);
nor U11983 (N_11983,N_6155,N_6311);
nand U11984 (N_11984,N_8735,N_7195);
nand U11985 (N_11985,N_6863,N_7914);
nand U11986 (N_11986,N_6629,N_7108);
nor U11987 (N_11987,N_7210,N_6040);
nor U11988 (N_11988,N_6321,N_6166);
nand U11989 (N_11989,N_7061,N_6418);
nand U11990 (N_11990,N_7486,N_6570);
xor U11991 (N_11991,N_7699,N_8837);
nor U11992 (N_11992,N_7388,N_8027);
nand U11993 (N_11993,N_7152,N_7535);
or U11994 (N_11994,N_8190,N_6969);
or U11995 (N_11995,N_8468,N_7719);
and U11996 (N_11996,N_6094,N_6771);
and U11997 (N_11997,N_8457,N_7800);
nor U11998 (N_11998,N_6998,N_7093);
nor U11999 (N_11999,N_6723,N_6540);
nand U12000 (N_12000,N_10428,N_11767);
and U12001 (N_12001,N_10868,N_11772);
xor U12002 (N_12002,N_11400,N_10431);
nand U12003 (N_12003,N_10682,N_9914);
nand U12004 (N_12004,N_10328,N_9534);
and U12005 (N_12005,N_10308,N_11221);
nor U12006 (N_12006,N_9748,N_9184);
nand U12007 (N_12007,N_10147,N_10375);
nand U12008 (N_12008,N_10944,N_11074);
nand U12009 (N_12009,N_9578,N_9747);
nor U12010 (N_12010,N_11028,N_9478);
or U12011 (N_12011,N_9252,N_11473);
and U12012 (N_12012,N_11693,N_9244);
nor U12013 (N_12013,N_11387,N_11618);
nor U12014 (N_12014,N_11493,N_9028);
or U12015 (N_12015,N_9528,N_9506);
nor U12016 (N_12016,N_9736,N_11427);
and U12017 (N_12017,N_11231,N_9020);
or U12018 (N_12018,N_10137,N_9925);
nand U12019 (N_12019,N_9492,N_9554);
nor U12020 (N_12020,N_9809,N_9339);
and U12021 (N_12021,N_9574,N_11858);
and U12022 (N_12022,N_10794,N_11513);
or U12023 (N_12023,N_10237,N_10288);
and U12024 (N_12024,N_10277,N_10098);
and U12025 (N_12025,N_10012,N_9246);
or U12026 (N_12026,N_11334,N_10313);
nand U12027 (N_12027,N_11616,N_9209);
nand U12028 (N_12028,N_11453,N_9963);
nand U12029 (N_12029,N_11316,N_9344);
nor U12030 (N_12030,N_11025,N_10932);
and U12031 (N_12031,N_9536,N_10786);
and U12032 (N_12032,N_11429,N_11771);
nand U12033 (N_12033,N_10481,N_9620);
or U12034 (N_12034,N_11588,N_9843);
and U12035 (N_12035,N_9277,N_9178);
nor U12036 (N_12036,N_11175,N_10565);
or U12037 (N_12037,N_9547,N_11019);
or U12038 (N_12038,N_11509,N_9597);
or U12039 (N_12039,N_11105,N_9684);
or U12040 (N_12040,N_10606,N_9776);
xor U12041 (N_12041,N_9972,N_9657);
or U12042 (N_12042,N_10728,N_10394);
and U12043 (N_12043,N_10739,N_9069);
nor U12044 (N_12044,N_9258,N_11361);
nand U12045 (N_12045,N_11350,N_10229);
or U12046 (N_12046,N_9458,N_10222);
nand U12047 (N_12047,N_9543,N_11174);
nand U12048 (N_12048,N_11783,N_11814);
nor U12049 (N_12049,N_10245,N_9402);
xor U12050 (N_12050,N_10262,N_9175);
nor U12051 (N_12051,N_10272,N_10675);
and U12052 (N_12052,N_9874,N_10840);
and U12053 (N_12053,N_10287,N_10472);
xnor U12054 (N_12054,N_9978,N_9881);
xor U12055 (N_12055,N_11474,N_10990);
or U12056 (N_12056,N_10065,N_10710);
nand U12057 (N_12057,N_10030,N_11714);
nor U12058 (N_12058,N_11343,N_9135);
nand U12059 (N_12059,N_11785,N_11776);
and U12060 (N_12060,N_9380,N_11058);
nand U12061 (N_12061,N_10215,N_11866);
nand U12062 (N_12062,N_11533,N_9349);
nand U12063 (N_12063,N_9969,N_11116);
and U12064 (N_12064,N_9987,N_11907);
nor U12065 (N_12065,N_10669,N_10418);
nand U12066 (N_12066,N_11452,N_11271);
and U12067 (N_12067,N_9529,N_9230);
nor U12068 (N_12068,N_11345,N_10782);
nor U12069 (N_12069,N_11071,N_11634);
and U12070 (N_12070,N_9188,N_10841);
nor U12071 (N_12071,N_11979,N_9318);
nand U12072 (N_12072,N_10749,N_10956);
or U12073 (N_12073,N_9703,N_11485);
nand U12074 (N_12074,N_9455,N_11086);
nor U12075 (N_12075,N_9082,N_10372);
nor U12076 (N_12076,N_11152,N_9954);
nor U12077 (N_12077,N_10358,N_10874);
or U12078 (N_12078,N_9428,N_10570);
nand U12079 (N_12079,N_11134,N_9770);
nand U12080 (N_12080,N_9565,N_9783);
nand U12081 (N_12081,N_11365,N_9389);
nor U12082 (N_12082,N_9051,N_10359);
nand U12083 (N_12083,N_9701,N_9757);
and U12084 (N_12084,N_10371,N_10656);
or U12085 (N_12085,N_10620,N_10459);
and U12086 (N_12086,N_11463,N_10397);
nand U12087 (N_12087,N_10491,N_9032);
or U12088 (N_12088,N_10479,N_10083);
or U12089 (N_12089,N_10631,N_10989);
nor U12090 (N_12090,N_9731,N_9625);
or U12091 (N_12091,N_10536,N_11690);
nand U12092 (N_12092,N_11909,N_11812);
nor U12093 (N_12093,N_10953,N_11667);
or U12094 (N_12094,N_10158,N_10842);
nand U12095 (N_12095,N_10997,N_10090);
or U12096 (N_12096,N_10453,N_9553);
or U12097 (N_12097,N_10760,N_9544);
or U12098 (N_12098,N_11506,N_10929);
and U12099 (N_12099,N_9837,N_11855);
nand U12100 (N_12100,N_10048,N_9950);
and U12101 (N_12101,N_10216,N_10547);
nor U12102 (N_12102,N_9559,N_10100);
and U12103 (N_12103,N_11575,N_10720);
nand U12104 (N_12104,N_10876,N_9900);
nand U12105 (N_12105,N_9326,N_10689);
or U12106 (N_12106,N_11272,N_9222);
and U12107 (N_12107,N_11965,N_10124);
and U12108 (N_12108,N_10066,N_11311);
nand U12109 (N_12109,N_11120,N_9599);
or U12110 (N_12110,N_9399,N_11442);
and U12111 (N_12111,N_10832,N_10688);
and U12112 (N_12112,N_11516,N_9269);
and U12113 (N_12113,N_10044,N_9871);
nand U12114 (N_12114,N_10591,N_9280);
or U12115 (N_12115,N_9310,N_10343);
and U12116 (N_12116,N_9114,N_11494);
or U12117 (N_12117,N_9345,N_9424);
and U12118 (N_12118,N_11613,N_10817);
and U12119 (N_12119,N_9745,N_11821);
and U12120 (N_12120,N_9921,N_11695);
or U12121 (N_12121,N_11004,N_11021);
nor U12122 (N_12122,N_9005,N_11180);
nand U12123 (N_12123,N_10278,N_10869);
or U12124 (N_12124,N_9159,N_11067);
or U12125 (N_12125,N_10896,N_9132);
and U12126 (N_12126,N_9287,N_11947);
nand U12127 (N_12127,N_10807,N_11097);
nor U12128 (N_12128,N_10562,N_11655);
and U12129 (N_12129,N_10121,N_9686);
nand U12130 (N_12130,N_11203,N_11209);
or U12131 (N_12131,N_11728,N_9491);
nor U12132 (N_12132,N_9439,N_10823);
or U12133 (N_12133,N_11628,N_11054);
nor U12134 (N_12134,N_11883,N_9728);
nand U12135 (N_12135,N_11531,N_11041);
or U12136 (N_12136,N_10027,N_9739);
and U12137 (N_12137,N_9434,N_11782);
nand U12138 (N_12138,N_11731,N_9756);
or U12139 (N_12139,N_10858,N_10680);
or U12140 (N_12140,N_9884,N_10438);
or U12141 (N_12141,N_11087,N_11591);
nor U12142 (N_12142,N_11050,N_10612);
and U12143 (N_12143,N_11060,N_9066);
or U12144 (N_12144,N_9680,N_10092);
nor U12145 (N_12145,N_9859,N_10169);
nor U12146 (N_12146,N_11636,N_10724);
nand U12147 (N_12147,N_11301,N_9250);
nor U12148 (N_12148,N_9569,N_9303);
nand U12149 (N_12149,N_11184,N_11286);
nor U12150 (N_12150,N_11872,N_11355);
and U12151 (N_12151,N_9294,N_10805);
nor U12152 (N_12152,N_9595,N_9168);
nand U12153 (N_12153,N_9790,N_9635);
or U12154 (N_12154,N_10487,N_10081);
nand U12155 (N_12155,N_11946,N_9946);
nor U12156 (N_12156,N_11341,N_9170);
and U12157 (N_12157,N_11002,N_10762);
nor U12158 (N_12158,N_9527,N_10392);
nand U12159 (N_12159,N_10164,N_10069);
nand U12160 (N_12160,N_10273,N_10243);
nor U12161 (N_12161,N_11709,N_11626);
nand U12162 (N_12162,N_9503,N_9512);
xnor U12163 (N_12163,N_10527,N_11479);
and U12164 (N_12164,N_9834,N_10150);
or U12165 (N_12165,N_10902,N_9140);
or U12166 (N_12166,N_9289,N_9470);
nor U12167 (N_12167,N_10563,N_11265);
nand U12168 (N_12168,N_10240,N_10152);
and U12169 (N_12169,N_11455,N_10155);
and U12170 (N_12170,N_10727,N_10787);
and U12171 (N_12171,N_11213,N_9496);
or U12172 (N_12172,N_10391,N_11331);
and U12173 (N_12173,N_11088,N_11358);
nand U12174 (N_12174,N_9000,N_9733);
nor U12175 (N_12175,N_11015,N_9202);
and U12176 (N_12176,N_11980,N_9760);
nand U12177 (N_12177,N_9511,N_11718);
and U12178 (N_12178,N_11149,N_9227);
nor U12179 (N_12179,N_11698,N_11929);
and U12180 (N_12180,N_9562,N_11310);
or U12181 (N_12181,N_11754,N_11692);
or U12182 (N_12182,N_9600,N_9690);
or U12183 (N_12183,N_9379,N_10629);
and U12184 (N_12184,N_10653,N_10063);
nand U12185 (N_12185,N_11110,N_9011);
nand U12186 (N_12186,N_9290,N_10758);
nor U12187 (N_12187,N_9273,N_10156);
nor U12188 (N_12188,N_9989,N_9457);
nor U12189 (N_12189,N_11870,N_9922);
or U12190 (N_12190,N_9221,N_10381);
nand U12191 (N_12191,N_10951,N_10552);
nand U12192 (N_12192,N_11235,N_11916);
or U12193 (N_12193,N_11344,N_11022);
and U12194 (N_12194,N_9846,N_10139);
and U12195 (N_12195,N_10828,N_10555);
nand U12196 (N_12196,N_11918,N_9327);
and U12197 (N_12197,N_9466,N_11986);
xnor U12198 (N_12198,N_9358,N_10023);
and U12199 (N_12199,N_11746,N_9644);
and U12200 (N_12200,N_11079,N_11156);
and U12201 (N_12201,N_10336,N_11863);
and U12202 (N_12202,N_9813,N_9915);
and U12203 (N_12203,N_9134,N_10184);
nand U12204 (N_12204,N_10289,N_10441);
or U12205 (N_12205,N_11046,N_11416);
nand U12206 (N_12206,N_9866,N_10839);
and U12207 (N_12207,N_11961,N_10910);
nand U12208 (N_12208,N_11837,N_9452);
nand U12209 (N_12209,N_11321,N_11859);
nand U12210 (N_12210,N_9473,N_11619);
and U12211 (N_12211,N_9072,N_11244);
or U12212 (N_12212,N_10042,N_9019);
and U12213 (N_12213,N_10293,N_10159);
nand U12214 (N_12214,N_11445,N_11633);
and U12215 (N_12215,N_10978,N_11124);
nor U12216 (N_12216,N_9422,N_10909);
and U12217 (N_12217,N_10779,N_11700);
nand U12218 (N_12218,N_9984,N_10276);
and U12219 (N_12219,N_10578,N_9870);
or U12220 (N_12220,N_11987,N_11642);
nor U12221 (N_12221,N_9461,N_10761);
nor U12222 (N_12222,N_9023,N_10489);
nor U12223 (N_12223,N_11262,N_11585);
nand U12224 (N_12224,N_9568,N_11538);
or U12225 (N_12225,N_11127,N_10880);
nand U12226 (N_12226,N_10300,N_10338);
nor U12227 (N_12227,N_11838,N_9228);
and U12228 (N_12228,N_9026,N_10434);
nand U12229 (N_12229,N_9676,N_11254);
and U12230 (N_12230,N_9828,N_10693);
and U12231 (N_12231,N_11238,N_10040);
and U12232 (N_12232,N_11297,N_11291);
or U12233 (N_12233,N_11791,N_9668);
nand U12234 (N_12234,N_11792,N_11083);
nand U12235 (N_12235,N_10440,N_9566);
xor U12236 (N_12236,N_10493,N_9329);
or U12237 (N_12237,N_9715,N_9615);
or U12238 (N_12238,N_10622,N_9173);
nand U12239 (N_12239,N_10502,N_11414);
nor U12240 (N_12240,N_11958,N_11336);
and U12241 (N_12241,N_10490,N_9588);
or U12242 (N_12242,N_11101,N_11832);
and U12243 (N_12243,N_11666,N_10845);
nor U12244 (N_12244,N_11080,N_10878);
and U12245 (N_12245,N_11926,N_11972);
xor U12246 (N_12246,N_9365,N_11402);
and U12247 (N_12247,N_10099,N_9335);
nand U12248 (N_12248,N_9386,N_11373);
and U12249 (N_12249,N_11182,N_9800);
or U12250 (N_12250,N_11397,N_9719);
or U12251 (N_12251,N_10926,N_10463);
nand U12252 (N_12252,N_11486,N_11500);
nor U12253 (N_12253,N_10192,N_11664);
and U12254 (N_12254,N_11062,N_10347);
or U12255 (N_12255,N_9893,N_9133);
nor U12256 (N_12256,N_9479,N_11749);
nand U12257 (N_12257,N_10865,N_11830);
nor U12258 (N_12258,N_9139,N_10549);
or U12259 (N_12259,N_11614,N_11813);
or U12260 (N_12260,N_11118,N_10447);
or U12261 (N_12261,N_11172,N_11534);
nand U12262 (N_12262,N_10002,N_11912);
and U12263 (N_12263,N_10651,N_9048);
nand U12264 (N_12264,N_9275,N_10960);
or U12265 (N_12265,N_10464,N_11132);
nand U12266 (N_12266,N_9862,N_10970);
nor U12267 (N_12267,N_10324,N_9674);
nand U12268 (N_12268,N_9361,N_9714);
nand U12269 (N_12269,N_10905,N_11662);
nor U12270 (N_12270,N_11976,N_11276);
or U12271 (N_12271,N_10444,N_10473);
nand U12272 (N_12272,N_10542,N_11045);
nand U12273 (N_12273,N_9817,N_9502);
nand U12274 (N_12274,N_11153,N_11809);
and U12275 (N_12275,N_11242,N_11535);
and U12276 (N_12276,N_9899,N_10888);
nand U12277 (N_12277,N_10275,N_9419);
or U12278 (N_12278,N_11611,N_10683);
or U12279 (N_12279,N_9158,N_10475);
nor U12280 (N_12280,N_10574,N_10129);
or U12281 (N_12281,N_9769,N_9414);
and U12282 (N_12282,N_10889,N_10251);
and U12283 (N_12283,N_11927,N_10711);
nor U12284 (N_12284,N_10561,N_9537);
or U12285 (N_12285,N_10016,N_11465);
nor U12286 (N_12286,N_9805,N_10666);
and U12287 (N_12287,N_9086,N_9876);
and U12288 (N_12288,N_11314,N_10526);
nor U12289 (N_12289,N_10247,N_9027);
nor U12290 (N_12290,N_11181,N_10064);
nand U12291 (N_12291,N_10532,N_10480);
nand U12292 (N_12292,N_10142,N_11368);
nand U12293 (N_12293,N_10748,N_11775);
nand U12294 (N_12294,N_11970,N_9779);
or U12295 (N_12295,N_9360,N_10531);
nand U12296 (N_12296,N_9117,N_9602);
and U12297 (N_12297,N_11454,N_10914);
or U12298 (N_12298,N_9049,N_9410);
nand U12299 (N_12299,N_9396,N_9163);
and U12300 (N_12300,N_11135,N_9631);
nor U12301 (N_12301,N_11320,N_10763);
and U12302 (N_12302,N_9123,N_9610);
and U12303 (N_12303,N_11154,N_9796);
or U12304 (N_12304,N_9157,N_9183);
nor U12305 (N_12305,N_9970,N_10166);
nand U12306 (N_12306,N_11803,N_11128);
and U12307 (N_12307,N_9591,N_11997);
nor U12308 (N_12308,N_11293,N_10678);
and U12309 (N_12309,N_11846,N_9627);
or U12310 (N_12310,N_9695,N_9663);
xor U12311 (N_12311,N_9832,N_11865);
or U12312 (N_12312,N_10604,N_10936);
or U12313 (N_12313,N_11953,N_10344);
and U12314 (N_12314,N_11186,N_11777);
or U12315 (N_12315,N_10311,N_10274);
nand U12316 (N_12316,N_9219,N_9076);
nand U12317 (N_12317,N_11439,N_11201);
and U12318 (N_12318,N_10639,N_9116);
or U12319 (N_12319,N_11527,N_9030);
nor U12320 (N_12320,N_11969,N_10122);
and U12321 (N_12321,N_9482,N_10316);
nand U12322 (N_12322,N_9764,N_10173);
nor U12323 (N_12323,N_9791,N_9308);
and U12324 (N_12324,N_10716,N_9077);
nand U12325 (N_12325,N_9882,N_11507);
nor U12326 (N_12326,N_9823,N_10518);
nor U12327 (N_12327,N_9018,N_11547);
or U12328 (N_12328,N_9357,N_10827);
and U12329 (N_12329,N_9751,N_10172);
xor U12330 (N_12330,N_11715,N_11652);
and U12331 (N_12331,N_11112,N_9249);
nand U12332 (N_12332,N_11084,N_9603);
or U12333 (N_12333,N_11993,N_10177);
or U12334 (N_12334,N_9265,N_9679);
or U12335 (N_12335,N_10577,N_10759);
nand U12336 (N_12336,N_9678,N_9609);
or U12337 (N_12337,N_9993,N_11359);
nor U12338 (N_12338,N_10408,N_10259);
nand U12339 (N_12339,N_11716,N_10354);
nor U12340 (N_12340,N_10681,N_9645);
nand U12341 (N_12341,N_9067,N_11263);
nand U12342 (N_12342,N_11512,N_10253);
or U12343 (N_12343,N_10234,N_10947);
and U12344 (N_12344,N_9863,N_10373);
nor U12345 (N_12345,N_10553,N_11475);
or U12346 (N_12346,N_11099,N_11299);
and U12347 (N_12347,N_10690,N_11708);
nand U12348 (N_12348,N_9895,N_11085);
nor U12349 (N_12349,N_11415,N_10742);
or U12350 (N_12350,N_11146,N_11874);
nor U12351 (N_12351,N_11784,N_10449);
nand U12352 (N_12352,N_10568,N_11957);
nand U12353 (N_12353,N_9400,N_11300);
and U12354 (N_12354,N_9641,N_9858);
nand U12355 (N_12355,N_9237,N_10927);
nand U12356 (N_12356,N_11401,N_9824);
or U12357 (N_12357,N_10377,N_9592);
nand U12358 (N_12358,N_11339,N_11963);
nor U12359 (N_12359,N_9854,N_10744);
and U12360 (N_12360,N_11755,N_9376);
nor U12361 (N_12361,N_11082,N_9351);
and U12362 (N_12362,N_11810,N_10813);
nor U12363 (N_12363,N_10705,N_9853);
and U12364 (N_12364,N_11047,N_9078);
or U12365 (N_12365,N_11375,N_11757);
nor U12366 (N_12366,N_9912,N_10333);
nand U12367 (N_12367,N_11206,N_11974);
or U12368 (N_12368,N_9943,N_9507);
nand U12369 (N_12369,N_9847,N_10265);
nand U12370 (N_12370,N_10556,N_11943);
nor U12371 (N_12371,N_9035,N_11337);
or U12372 (N_12372,N_10427,N_11230);
or U12373 (N_12373,N_9421,N_10646);
nor U12374 (N_12374,N_11018,N_10168);
or U12375 (N_12375,N_11717,N_9029);
nand U12376 (N_12376,N_9299,N_11624);
nor U12377 (N_12377,N_11839,N_10700);
nand U12378 (N_12378,N_10596,N_11308);
nor U12379 (N_12379,N_11685,N_11761);
and U12380 (N_12380,N_11504,N_9064);
nand U12381 (N_12381,N_9391,N_11956);
nand U12382 (N_12382,N_9702,N_9453);
or U12383 (N_12383,N_11228,N_9334);
and U12384 (N_12384,N_11012,N_10189);
nor U12385 (N_12385,N_9236,N_10741);
and U12386 (N_12386,N_11584,N_10478);
and U12387 (N_12387,N_9883,N_11207);
or U12388 (N_12388,N_10721,N_11579);
and U12389 (N_12389,N_10691,N_10406);
and U12390 (N_12390,N_11497,N_9949);
and U12391 (N_12391,N_9677,N_11143);
nand U12392 (N_12392,N_9047,N_11638);
and U12393 (N_12393,N_11917,N_11119);
and U12394 (N_12394,N_10178,N_10032);
nand U12395 (N_12395,N_9688,N_9742);
xor U12396 (N_12396,N_10113,N_11468);
nand U12397 (N_12397,N_11225,N_11223);
nand U12398 (N_12398,N_11699,N_10497);
nand U12399 (N_12399,N_10022,N_9836);
nand U12400 (N_12400,N_9724,N_10923);
or U12401 (N_12401,N_10196,N_10645);
or U12402 (N_12402,N_11496,N_11061);
or U12403 (N_12403,N_11501,N_11278);
nand U12404 (N_12404,N_11735,N_9643);
or U12405 (N_12405,N_9190,N_9730);
nand U12406 (N_12406,N_11179,N_10210);
or U12407 (N_12407,N_9350,N_9520);
nand U12408 (N_12408,N_9122,N_11519);
nand U12409 (N_12409,N_10860,N_10625);
nand U12410 (N_12410,N_10414,N_11878);
nor U12411 (N_12411,N_11081,N_9095);
or U12412 (N_12412,N_9792,N_10600);
or U12413 (N_12413,N_10988,N_9939);
or U12414 (N_12414,N_9555,N_9979);
nand U12415 (N_12415,N_11729,N_9533);
or U12416 (N_12416,N_10423,N_10161);
nor U12417 (N_12417,N_11736,N_11815);
nand U12418 (N_12418,N_10389,N_10894);
nor U12419 (N_12419,N_11014,N_10571);
nand U12420 (N_12420,N_9842,N_10241);
nand U12421 (N_12421,N_10881,N_9260);
nand U12422 (N_12422,N_10933,N_9024);
nand U12423 (N_12423,N_10831,N_11913);
and U12424 (N_12424,N_11612,N_11191);
or U12425 (N_12425,N_10851,N_10004);
xnor U12426 (N_12426,N_10437,N_11756);
and U12427 (N_12427,N_9761,N_9903);
and U12428 (N_12428,N_11131,N_9877);
nor U12429 (N_12429,N_11890,N_11332);
nand U12430 (N_12430,N_10321,N_10714);
and U12431 (N_12431,N_11871,N_9998);
nand U12432 (N_12432,N_10572,N_11437);
or U12433 (N_12433,N_9074,N_9567);
or U12434 (N_12434,N_11901,N_11428);
or U12435 (N_12435,N_9061,N_9613);
and U12436 (N_12436,N_10558,N_10117);
and U12437 (N_12437,N_9655,N_11532);
nor U12438 (N_12438,N_10977,N_9211);
nor U12439 (N_12439,N_11139,N_11945);
xor U12440 (N_12440,N_10655,N_11650);
and U12441 (N_12441,N_11670,N_9623);
nand U12442 (N_12442,N_10110,N_11819);
and U12443 (N_12443,N_9541,N_9103);
nand U12444 (N_12444,N_9772,N_10985);
nand U12445 (N_12445,N_9012,N_11834);
nand U12446 (N_12446,N_9112,N_9759);
or U12447 (N_12447,N_10291,N_11727);
and U12448 (N_12448,N_9068,N_10393);
or U12449 (N_12449,N_10154,N_11920);
nand U12450 (N_12450,N_11395,N_11418);
and U12451 (N_12451,N_10384,N_9879);
or U12452 (N_12452,N_11704,N_10746);
nand U12453 (N_12453,N_10550,N_11936);
and U12454 (N_12454,N_10329,N_11349);
or U12455 (N_12455,N_9716,N_10587);
nand U12456 (N_12456,N_11456,N_9266);
nor U12457 (N_12457,N_11933,N_10738);
and U12458 (N_12458,N_10367,N_11217);
and U12459 (N_12459,N_10310,N_9229);
nor U12460 (N_12460,N_11040,N_10454);
and U12461 (N_12461,N_11555,N_9581);
nor U12462 (N_12462,N_9377,N_9660);
or U12463 (N_12463,N_10000,N_11677);
and U12464 (N_12464,N_9021,N_11204);
and U12465 (N_12465,N_10452,N_9448);
and U12466 (N_12466,N_9206,N_9463);
nand U12467 (N_12467,N_9505,N_9632);
nor U12468 (N_12468,N_11564,N_11919);
and U12469 (N_12469,N_10987,N_9161);
nand U12470 (N_12470,N_9951,N_10709);
or U12471 (N_12471,N_9333,N_11366);
nor U12472 (N_12472,N_9902,N_11466);
nand U12473 (N_12473,N_11033,N_11380);
nand U12474 (N_12474,N_9160,N_11686);
and U12475 (N_12475,N_9241,N_11171);
and U12476 (N_12476,N_10118,N_11657);
nor U12477 (N_12477,N_9167,N_10641);
nor U12478 (N_12478,N_9297,N_10426);
or U12479 (N_12479,N_10699,N_9446);
and U12480 (N_12480,N_10026,N_11115);
and U12481 (N_12481,N_9097,N_10084);
nor U12482 (N_12482,N_10846,N_9734);
nand U12483 (N_12483,N_11769,N_11362);
and U12484 (N_12484,N_10593,N_9750);
or U12485 (N_12485,N_10077,N_11867);
nor U12486 (N_12486,N_9711,N_10116);
and U12487 (N_12487,N_11899,N_10921);
nor U12488 (N_12488,N_10140,N_11672);
or U12489 (N_12489,N_11446,N_9570);
or U12490 (N_12490,N_11290,N_11357);
or U12491 (N_12491,N_9187,N_11266);
or U12492 (N_12492,N_10912,N_10269);
or U12493 (N_12493,N_10486,N_9392);
nand U12494 (N_12494,N_10753,N_9826);
nor U12495 (N_12495,N_10143,N_9671);
nor U12496 (N_12496,N_10070,N_11848);
nand U12497 (N_12497,N_11603,N_10341);
nor U12498 (N_12498,N_9004,N_11881);
and U12499 (N_12499,N_9687,N_11093);
nor U12500 (N_12500,N_11369,N_11106);
nor U12501 (N_12501,N_10105,N_10633);
nor U12502 (N_12502,N_11583,N_11719);
and U12503 (N_12503,N_11739,N_9493);
and U12504 (N_12504,N_11944,N_10660);
nand U12505 (N_12505,N_10370,N_9062);
nor U12506 (N_12506,N_10356,N_10864);
nor U12507 (N_12507,N_11306,N_10543);
and U12508 (N_12508,N_11663,N_9885);
and U12509 (N_12509,N_10857,N_9189);
xnor U12510 (N_12510,N_11549,N_11637);
nor U12511 (N_12511,N_9582,N_11352);
and U12512 (N_12512,N_10019,N_10835);
nand U12513 (N_12513,N_10174,N_11137);
nor U12514 (N_12514,N_10213,N_10580);
nand U12515 (N_12515,N_10330,N_10435);
nor U12516 (N_12516,N_9002,N_11932);
nand U12517 (N_12517,N_9444,N_10569);
nor U12518 (N_12518,N_10795,N_9234);
nand U12519 (N_12519,N_10797,N_11168);
nor U12520 (N_12520,N_10506,N_9065);
and U12521 (N_12521,N_11440,N_10713);
nor U12522 (N_12522,N_9320,N_11595);
or U12523 (N_12523,N_11602,N_11406);
nand U12524 (N_12524,N_11741,N_11471);
nand U12525 (N_12525,N_9649,N_10443);
nor U12526 (N_12526,N_11537,N_11324);
nor U12527 (N_12527,N_10496,N_10975);
and U12528 (N_12528,N_9775,N_10862);
or U12529 (N_12529,N_11481,N_9046);
and U12530 (N_12530,N_10733,N_9359);
nand U12531 (N_12531,N_11107,N_9563);
nand U12532 (N_12532,N_10602,N_10607);
nor U12533 (N_12533,N_10627,N_10072);
or U12534 (N_12534,N_10867,N_10884);
nor U12535 (N_12535,N_11539,N_11831);
nor U12536 (N_12536,N_10319,N_9872);
or U12537 (N_12537,N_9477,N_11882);
or U12538 (N_12538,N_9120,N_11632);
nor U12539 (N_12539,N_11811,N_9852);
nor U12540 (N_12540,N_10590,N_10186);
nand U12541 (N_12541,N_10640,N_10494);
nand U12542 (N_12542,N_11759,N_9749);
and U12543 (N_12543,N_11720,N_10764);
nor U12544 (N_12544,N_9406,N_11333);
nand U12545 (N_12545,N_10296,N_9364);
or U12546 (N_12546,N_9991,N_11451);
or U12547 (N_12547,N_11029,N_9407);
nor U12548 (N_12548,N_10694,N_11896);
or U12549 (N_12549,N_9149,N_10332);
or U12550 (N_12550,N_10270,N_11762);
nand U12551 (N_12551,N_10672,N_11627);
and U12552 (N_12552,N_10209,N_11178);
nor U12553 (N_12553,N_10123,N_9789);
or U12554 (N_12554,N_10939,N_9741);
or U12555 (N_12555,N_9540,N_10946);
nand U12556 (N_12556,N_10503,N_11296);
or U12557 (N_12557,N_11732,N_10352);
nand U12558 (N_12558,N_9841,N_11669);
nand U12559 (N_12559,N_9683,N_11210);
and U12560 (N_12560,N_10855,N_10938);
nand U12561 (N_12561,N_10650,N_9415);
and U12562 (N_12562,N_9521,N_10548);
or U12563 (N_12563,N_10996,N_11450);
and U12564 (N_12564,N_11222,N_9732);
nor U12565 (N_12565,N_9777,N_10232);
or U12566 (N_12566,N_10608,N_11610);
and U12567 (N_12567,N_9692,N_9031);
nand U12568 (N_12568,N_9586,N_9517);
or U12569 (N_12569,N_9015,N_9363);
or U12570 (N_12570,N_11781,N_10195);
nor U12571 (N_12571,N_10226,N_10621);
and U12572 (N_12572,N_10974,N_9651);
nand U12573 (N_12573,N_10965,N_11804);
nand U12574 (N_12574,N_11470,N_10616);
and U12575 (N_12575,N_9058,N_9601);
nor U12576 (N_12576,N_10501,N_9705);
nor U12577 (N_12577,N_10357,N_10292);
or U12578 (N_12578,N_10219,N_9224);
or U12579 (N_12579,N_9235,N_11457);
or U12580 (N_12580,N_10952,N_9934);
or U12581 (N_12581,N_10962,N_11284);
nand U12582 (N_12582,N_11954,N_11219);
nor U12583 (N_12583,N_10696,N_9799);
and U12584 (N_12584,N_11458,N_11802);
or U12585 (N_12585,N_9580,N_11794);
or U12586 (N_12586,N_10236,N_9291);
and U12587 (N_12587,N_11653,N_10318);
or U12588 (N_12588,N_10734,N_11680);
or U12589 (N_12589,N_10998,N_10266);
or U12590 (N_12590,N_10246,N_9485);
and U12591 (N_12591,N_11598,N_11129);
or U12592 (N_12592,N_11476,N_9718);
nor U12593 (N_12593,N_9171,N_11706);
nor U12594 (N_12594,N_9059,N_11150);
or U12595 (N_12595,N_10589,N_9382);
and U12596 (N_12596,N_11576,N_10185);
nor U12597 (N_12597,N_10132,N_10723);
nand U12598 (N_12598,N_11173,N_10767);
nand U12599 (N_12599,N_11582,N_9650);
nand U12600 (N_12600,N_11003,N_10575);
nand U12601 (N_12601,N_11267,N_11676);
nor U12602 (N_12602,N_9328,N_11646);
or U12603 (N_12603,N_11200,N_11930);
nor U12604 (N_12604,N_11169,N_9825);
and U12605 (N_12605,N_9101,N_9944);
nor U12606 (N_12606,N_9956,N_9214);
and U12607 (N_12607,N_11302,N_10821);
nand U12608 (N_12608,N_11654,N_9181);
and U12609 (N_12609,N_9626,N_9367);
nor U12610 (N_12610,N_9640,N_10365);
and U12611 (N_12611,N_11623,N_10942);
or U12612 (N_12612,N_10630,N_10204);
or U12613 (N_12613,N_10958,N_10521);
or U12614 (N_12614,N_11318,N_11556);
and U12615 (N_12615,N_11508,N_10260);
nand U12616 (N_12616,N_10366,N_10006);
or U12617 (N_12617,N_9940,N_11006);
and U12618 (N_12618,N_11960,N_10120);
and U12619 (N_12619,N_11144,N_10882);
or U12620 (N_12620,N_11967,N_9488);
xor U12621 (N_12621,N_11467,N_11660);
or U12622 (N_12622,N_9475,N_11572);
nand U12623 (N_12623,N_9152,N_9707);
nand U12624 (N_12624,N_9413,N_10829);
nand U12625 (N_12625,N_9199,N_9127);
nand U12626 (N_12626,N_10702,N_9590);
nor U12627 (N_12627,N_11688,N_11411);
or U12628 (N_12628,N_11023,N_10810);
and U12629 (N_12629,N_11381,N_10535);
nor U12630 (N_12630,N_9585,N_9185);
nor U12631 (N_12631,N_10055,N_10395);
and U12632 (N_12632,N_11779,N_11856);
or U12633 (N_12633,N_11273,N_11522);
or U12634 (N_12634,N_10583,N_11705);
and U12635 (N_12635,N_11910,N_9911);
and U12636 (N_12636,N_9390,N_9906);
xnor U12637 (N_12637,N_9661,N_11780);
or U12638 (N_12638,N_11066,N_11900);
and U12639 (N_12639,N_9829,N_10299);
or U12640 (N_12640,N_11971,N_9316);
nand U12641 (N_12641,N_10754,N_10080);
nor U12642 (N_12642,N_10849,N_10648);
nor U12643 (N_12643,N_9604,N_9111);
nand U12644 (N_12644,N_10770,N_11239);
or U12645 (N_12645,N_11111,N_9830);
or U12646 (N_12646,N_10848,N_9194);
nand U12647 (N_12647,N_10752,N_10637);
and U12648 (N_12648,N_10020,N_10007);
or U12649 (N_12649,N_9932,N_11240);
or U12650 (N_12650,N_11973,N_9384);
or U12651 (N_12651,N_11261,N_10339);
nor U12652 (N_12652,N_10980,N_11224);
nand U12653 (N_12653,N_9803,N_10180);
xnor U12654 (N_12654,N_9835,N_9892);
nand U12655 (N_12655,N_10825,N_11915);
or U12656 (N_12656,N_9948,N_9648);
and U12657 (N_12657,N_9038,N_9322);
nor U12658 (N_12658,N_10386,N_10778);
nand U12659 (N_12659,N_10153,N_10410);
and U12660 (N_12660,N_9727,N_10991);
nor U12661 (N_12661,N_11188,N_11448);
nand U12662 (N_12662,N_10467,N_9125);
nand U12663 (N_12663,N_9106,N_9524);
or U12664 (N_12664,N_10183,N_10802);
or U12665 (N_12665,N_11280,N_9217);
nor U12666 (N_12666,N_10170,N_11922);
nand U12667 (N_12667,N_10029,N_10919);
and U12668 (N_12668,N_10233,N_10875);
nand U12669 (N_12669,N_10483,N_11030);
nand U12670 (N_12670,N_10628,N_10928);
nand U12671 (N_12671,N_9037,N_9370);
or U12672 (N_12672,N_10976,N_10895);
nor U12673 (N_12673,N_11557,N_11409);
or U12674 (N_12674,N_9408,N_10907);
or U12675 (N_12675,N_11032,N_10211);
nand U12676 (N_12676,N_10041,N_11275);
nand U12677 (N_12677,N_9990,N_9454);
or U12678 (N_12678,N_10791,N_9247);
and U12679 (N_12679,N_10039,N_11382);
and U12680 (N_12680,N_11248,N_10731);
nor U12681 (N_12681,N_11104,N_11712);
and U12682 (N_12682,N_9735,N_10028);
nor U12683 (N_12683,N_9223,N_10018);
or U12684 (N_12684,N_9460,N_10199);
nand U12685 (N_12685,N_10126,N_9926);
or U12686 (N_12686,N_11599,N_9420);
nand U12687 (N_12687,N_10320,N_9418);
or U12688 (N_12688,N_11952,N_10515);
nand U12689 (N_12689,N_9725,N_11298);
and U12690 (N_12690,N_11133,N_10157);
nor U12691 (N_12691,N_10144,N_11063);
or U12692 (N_12692,N_11020,N_11911);
nor U12693 (N_12693,N_11577,N_11229);
and U12694 (N_12694,N_9288,N_11499);
or U12695 (N_12695,N_10450,N_11013);
or U12696 (N_12696,N_11938,N_9781);
or U12697 (N_12697,N_10239,N_10446);
nor U12698 (N_12698,N_9464,N_11256);
and U12699 (N_12699,N_11026,N_11198);
nor U12700 (N_12700,N_10283,N_10335);
nand U12701 (N_12701,N_9137,N_9498);
nor U12702 (N_12702,N_11567,N_9743);
or U12703 (N_12703,N_10451,N_11553);
nor U12704 (N_12704,N_9240,N_9923);
nand U12705 (N_12705,N_11561,N_10538);
and U12706 (N_12706,N_10820,N_10230);
and U12707 (N_12707,N_9412,N_11966);
nand U12708 (N_12708,N_10911,N_11902);
and U12709 (N_12709,N_11158,N_9740);
nand U12710 (N_12710,N_10362,N_9094);
nor U12711 (N_12711,N_9374,N_11743);
or U12712 (N_12712,N_11885,N_10145);
and U12713 (N_12713,N_10286,N_11243);
or U12714 (N_12714,N_10403,N_9664);
or U12715 (N_12715,N_11304,N_11836);
nand U12716 (N_12716,N_10814,N_10220);
nor U12717 (N_12717,N_10057,N_10046);
nor U12718 (N_12718,N_9195,N_10419);
nor U12719 (N_12719,N_9976,N_9353);
nand U12720 (N_12720,N_11315,N_11363);
or U12721 (N_12721,N_9484,N_10819);
and U12722 (N_12722,N_9093,N_11130);
nand U12723 (N_12723,N_11981,N_11528);
nand U12724 (N_12724,N_10257,N_9089);
or U12725 (N_12725,N_11114,N_9387);
nor U12726 (N_12726,N_9807,N_10227);
and U12727 (N_12727,N_9633,N_10109);
or U12728 (N_12728,N_10516,N_10967);
and U12729 (N_12729,N_11196,N_9481);
or U12730 (N_12730,N_10133,N_9840);
nand U12731 (N_12731,N_11713,N_11007);
nor U12732 (N_12732,N_11580,N_11123);
and U12733 (N_12733,N_11620,N_10088);
nand U12734 (N_12734,N_9279,N_9274);
or U12735 (N_12735,N_11649,N_11625);
nand U12736 (N_12736,N_11027,N_9036);
or U12737 (N_12737,N_11723,N_10053);
nand U12738 (N_12738,N_11822,N_11897);
xnor U12739 (N_12739,N_10350,N_10866);
nor U12740 (N_12740,N_10726,N_11593);
or U12741 (N_12741,N_11095,N_10217);
nor U12742 (N_12742,N_10416,N_9710);
nor U12743 (N_12743,N_9788,N_11682);
and U12744 (N_12744,N_11826,N_11742);
and U12745 (N_12745,N_9887,N_10130);
or U12746 (N_12746,N_11992,N_9416);
nand U12747 (N_12747,N_10388,N_11805);
and U12748 (N_12748,N_11586,N_9196);
or U12749 (N_12749,N_10033,N_11648);
and U12750 (N_12750,N_11701,N_9681);
and U12751 (N_12751,N_11227,N_9022);
nand U12752 (N_12752,N_9430,N_11542);
nor U12753 (N_12753,N_10225,N_10708);
nand U12754 (N_12754,N_9313,N_10013);
nor U12755 (N_12755,N_9208,N_9981);
nor U12756 (N_12756,N_9126,N_10112);
and U12757 (N_12757,N_9973,N_11404);
and U12758 (N_12758,N_10457,N_9472);
and U12759 (N_12759,N_11108,N_11077);
and U12760 (N_12760,N_11420,N_9694);
nand U12761 (N_12761,N_9480,N_11430);
nor U12762 (N_12762,N_11668,N_9774);
or U12763 (N_12763,N_10038,N_10551);
and U12764 (N_12764,N_11277,N_11484);
nand U12765 (N_12765,N_10765,N_10775);
and U12766 (N_12766,N_11996,N_10883);
nor U12767 (N_12767,N_10104,N_10203);
nand U12768 (N_12768,N_10474,N_11069);
and U12769 (N_12769,N_10729,N_10722);
nand U12770 (N_12770,N_11573,N_10737);
or U12771 (N_12771,N_9584,N_10348);
and U12772 (N_12772,N_10193,N_9073);
or U12773 (N_12773,N_9302,N_9839);
nor U12774 (N_12774,N_9436,N_10799);
and U12775 (N_12775,N_9780,N_11905);
and U12776 (N_12776,N_10188,N_9352);
nand U12777 (N_12777,N_10353,N_11820);
nand U12778 (N_12778,N_10465,N_11990);
nand U12779 (N_12779,N_9025,N_11844);
nor U12780 (N_12780,N_9873,N_11991);
nand U12781 (N_12781,N_9706,N_9820);
or U12782 (N_12782,N_11257,N_11740);
nand U12783 (N_12783,N_9251,N_10662);
nor U12784 (N_12784,N_9545,N_11737);
nand U12785 (N_12785,N_11630,N_11631);
or U12786 (N_12786,N_9284,N_10698);
and U12787 (N_12787,N_11396,N_9624);
or U12788 (N_12788,N_9109,N_10559);
or U12789 (N_12789,N_9486,N_11478);
or U12790 (N_12790,N_11941,N_11383);
or U12791 (N_12791,N_9889,N_9332);
or U12792 (N_12792,N_9523,N_11778);
nor U12793 (N_12793,N_9945,N_11236);
and U12794 (N_12794,N_9426,N_10379);
and U12795 (N_12795,N_11661,N_9268);
or U12796 (N_12796,N_11389,N_11226);
and U12797 (N_12797,N_9787,N_9177);
nand U12798 (N_12798,N_9220,N_11808);
nand U12799 (N_12799,N_9752,N_11730);
nand U12800 (N_12800,N_9154,N_10665);
nor U12801 (N_12801,N_11214,N_11554);
nor U12802 (N_12802,N_10331,N_11841);
nand U12803 (N_12803,N_11563,N_11328);
nor U12804 (N_12804,N_9083,N_9869);
and U12805 (N_12805,N_11148,N_9658);
or U12806 (N_12806,N_11994,N_10115);
or U12807 (N_12807,N_10636,N_10498);
and U12808 (N_12808,N_9737,N_11059);
and U12809 (N_12809,N_10009,N_9346);
or U12810 (N_12810,N_11807,N_9652);
nand U12811 (N_12811,N_9856,N_11109);
and U12812 (N_12812,N_10959,N_10982);
and U12813 (N_12813,N_10424,N_9239);
or U12814 (N_12814,N_11068,N_9530);
xor U12815 (N_12815,N_9713,N_11908);
or U12816 (N_12816,N_9438,N_11758);
xor U12817 (N_12817,N_9385,N_9314);
nand U12818 (N_12818,N_11353,N_11853);
nand U12819 (N_12819,N_11658,N_10968);
and U12820 (N_12820,N_9729,N_9798);
and U12821 (N_12821,N_11869,N_9811);
nand U12822 (N_12822,N_11895,N_10468);
or U12823 (N_12823,N_10429,N_10146);
or U12824 (N_12824,N_11860,N_9292);
nor U12825 (N_12825,N_10345,N_9670);
and U12826 (N_12826,N_11982,N_11574);
nand U12827 (N_12827,N_9875,N_9155);
nor U12828 (N_12828,N_9849,N_10374);
or U12829 (N_12829,N_11892,N_9151);
nand U12830 (N_12830,N_11875,N_9685);
nand U12831 (N_12831,N_11391,N_11589);
or U12832 (N_12832,N_9953,N_9401);
nand U12833 (N_12833,N_11745,N_9336);
nor U12834 (N_12834,N_10852,N_9369);
or U12835 (N_12835,N_10190,N_11205);
or U12836 (N_12836,N_11386,N_11951);
nand U12837 (N_12837,N_9372,N_9855);
nand U12838 (N_12838,N_11211,N_9445);
and U12839 (N_12839,N_11935,N_10201);
nor U12840 (N_12840,N_10284,N_10160);
or U12841 (N_12841,N_10812,N_11565);
and U12842 (N_12842,N_11829,N_11053);
or U12843 (N_12843,N_9682,N_9102);
or U12844 (N_12844,N_10854,N_11438);
or U12845 (N_12845,N_9901,N_11921);
nand U12846 (N_12846,N_10837,N_9317);
or U12847 (N_12847,N_11995,N_10079);
or U12848 (N_12848,N_10873,N_10605);
or U12849 (N_12849,N_10268,N_10214);
and U12850 (N_12850,N_11823,N_9539);
and U12851 (N_12851,N_9462,N_10207);
nor U12852 (N_12852,N_11959,N_10771);
or U12853 (N_12853,N_9232,N_10294);
nor U12854 (N_12854,N_11570,N_10337);
xor U12855 (N_12855,N_10898,N_11998);
nand U12856 (N_12856,N_9145,N_9306);
nand U12857 (N_12857,N_9459,N_11218);
or U12858 (N_12858,N_10049,N_9767);
or U12859 (N_12859,N_10512,N_11558);
nor U12860 (N_12860,N_9198,N_10635);
or U12861 (N_12861,N_11008,N_10134);
or U12862 (N_12862,N_9886,N_9699);
and U12863 (N_12863,N_10302,N_9556);
or U12864 (N_12864,N_10413,N_10103);
and U12865 (N_12865,N_11766,N_10400);
nor U12866 (N_12866,N_11295,N_9935);
nand U12867 (N_12867,N_11928,N_10613);
nor U12868 (N_12868,N_9927,N_11733);
and U12869 (N_12869,N_11233,N_10539);
nor U12870 (N_12870,N_9704,N_9778);
nand U12871 (N_12871,N_10307,N_10390);
and U12872 (N_12872,N_9043,N_9952);
or U12873 (N_12873,N_11529,N_9007);
nor U12874 (N_12874,N_10052,N_9766);
or U12875 (N_12875,N_11798,N_10686);
nor U12876 (N_12876,N_10244,N_11566);
or U12877 (N_12877,N_11237,N_9606);
and U12878 (N_12878,N_9992,N_10477);
nor U12879 (N_12879,N_11126,N_10138);
or U12880 (N_12880,N_11056,N_11170);
or U12881 (N_12881,N_9100,N_11459);
and U12882 (N_12882,N_9551,N_11421);
nor U12883 (N_12883,N_10261,N_11873);
and U12884 (N_12884,N_10279,N_9618);
nor U12885 (N_12885,N_11644,N_9443);
or U12886 (N_12886,N_10712,N_10981);
or U12887 (N_12887,N_10511,N_10545);
nand U12888 (N_12888,N_9063,N_9071);
or U12889 (N_12889,N_10582,N_9816);
and U12890 (N_12890,N_11977,N_10643);
nor U12891 (N_12891,N_9215,N_11888);
nor U12892 (N_12892,N_11403,N_9253);
nand U12893 (N_12893,N_9243,N_9471);
and U12894 (N_12894,N_9558,N_9197);
nor U12895 (N_12895,N_10872,N_11691);
nor U12896 (N_12896,N_11984,N_11313);
nor U12897 (N_12897,N_9994,N_9142);
nand U12898 (N_12898,N_11287,N_10087);
nand U12899 (N_12899,N_11360,N_9343);
or U12900 (N_12900,N_11955,N_10461);
or U12901 (N_12901,N_9340,N_10836);
or U12902 (N_12902,N_10455,N_10025);
or U12903 (N_12903,N_11392,N_11923);
or U12904 (N_12904,N_11495,N_11825);
nor U12905 (N_12905,N_10396,N_10290);
or U12906 (N_12906,N_10383,N_9868);
or U12907 (N_12907,N_9216,N_9042);
nor U12908 (N_12908,N_9959,N_11894);
nor U12909 (N_12909,N_9003,N_10445);
nor U12910 (N_12910,N_9331,N_10530);
and U12911 (N_12911,N_11525,N_9616);
nor U12912 (N_12912,N_10010,N_9867);
and U12913 (N_12913,N_9726,N_10061);
or U12914 (N_12914,N_11281,N_11884);
and U12915 (N_12915,N_10508,N_10769);
nor U12916 (N_12916,N_11569,N_11724);
and U12917 (N_12917,N_10417,N_11039);
nor U12918 (N_12918,N_9500,N_11678);
xnor U12919 (N_12919,N_10306,N_9085);
nor U12920 (N_12920,N_11164,N_10972);
nand U12921 (N_12921,N_10663,N_10504);
nor U12922 (N_12922,N_9342,N_9325);
or U12923 (N_12923,N_10718,N_9810);
nand U12924 (N_12924,N_9404,N_10517);
nand U12925 (N_12925,N_10937,N_11818);
nor U12926 (N_12926,N_11514,N_11751);
nor U12927 (N_12927,N_9433,N_9281);
nand U12928 (N_12928,N_10740,N_11195);
and U12929 (N_12929,N_11490,N_11245);
and U12930 (N_12930,N_9535,N_11405);
or U12931 (N_12931,N_10037,N_11121);
and U12932 (N_12932,N_9947,N_11376);
or U12933 (N_12933,N_11162,N_10584);
and U12934 (N_12934,N_11354,N_10796);
nand U12935 (N_12935,N_9977,N_11346);
or U12936 (N_12936,N_11806,N_10271);
nor U12937 (N_12937,N_10719,N_11530);
and U12938 (N_12938,N_10460,N_11444);
or U12939 (N_12939,N_11787,N_11629);
and U12940 (N_12940,N_11090,N_9205);
nand U12941 (N_12941,N_10524,N_10351);
nand U12942 (N_12942,N_11517,N_10317);
nand U12943 (N_12943,N_10094,N_10223);
nor U12944 (N_12944,N_10228,N_10913);
and U12945 (N_12945,N_10466,N_11594);
or U12946 (N_12946,N_10179,N_10623);
and U12947 (N_12947,N_10024,N_11388);
or U12948 (N_12948,N_10212,N_9238);
nor U12949 (N_12949,N_11434,N_11796);
nor U12950 (N_12950,N_10175,N_9587);
or U12951 (N_12951,N_11544,N_11734);
nand U12952 (N_12952,N_9878,N_11232);
or U12953 (N_12953,N_9115,N_11432);
nand U12954 (N_12954,N_11964,N_9278);
or U12955 (N_12955,N_11710,N_11103);
or U12956 (N_12956,N_10404,N_9165);
xnor U12957 (N_12957,N_10412,N_11931);
nand U12958 (N_12958,N_10482,N_9666);
or U12959 (N_12959,N_9162,N_10182);
nand U12960 (N_12960,N_11876,N_9309);
nor U12961 (N_12961,N_10385,N_10401);
and U12962 (N_12962,N_9305,N_10008);
xnor U12963 (N_12963,N_10948,N_10697);
or U12964 (N_12964,N_9936,N_9845);
nand U12965 (N_12965,N_9179,N_10254);
or U12966 (N_12966,N_9347,N_9300);
and U12967 (N_12967,N_10181,N_9315);
or U12968 (N_12968,N_9647,N_10755);
and U12969 (N_12969,N_9296,N_11398);
nand U12970 (N_12970,N_11122,N_11988);
or U12971 (N_12971,N_9098,N_11145);
nand U12972 (N_12972,N_11165,N_10824);
and U12973 (N_12973,N_9411,N_10005);
and U12974 (N_12974,N_11840,N_9006);
nor U12975 (N_12975,N_10045,N_10626);
nor U12976 (N_12976,N_9113,N_9397);
or U12977 (N_12977,N_11999,N_10971);
and U12978 (N_12978,N_10058,N_11592);
nand U12979 (N_12979,N_9617,N_10901);
or U12980 (N_12980,N_10963,N_10595);
nor U12981 (N_12981,N_9967,N_9440);
nand U12982 (N_12982,N_10541,N_10102);
nand U12983 (N_12983,N_10334,N_11893);
or U12984 (N_12984,N_11985,N_11850);
nor U12985 (N_12985,N_11510,N_10800);
nor U12986 (N_12986,N_11939,N_10492);
nand U12987 (N_12987,N_9815,N_9450);
nand U12988 (N_12988,N_10887,N_9794);
or U12989 (N_12989,N_11645,N_10745);
and U12990 (N_12990,N_11303,N_11279);
or U12991 (N_12991,N_9129,N_9508);
and U12992 (N_12992,N_10792,N_10904);
and U12993 (N_12993,N_11753,N_11335);
and U12994 (N_12994,N_9958,N_10931);
nand U12995 (N_12995,N_10916,N_11562);
and U12996 (N_12996,N_11760,N_9909);
nand U12997 (N_12997,N_9483,N_10448);
or U12998 (N_12998,N_10941,N_11622);
nand U12999 (N_12999,N_11689,N_9612);
nand U13000 (N_13000,N_9009,N_10657);
nor U13001 (N_13001,N_10068,N_10847);
nor U13002 (N_13002,N_10597,N_9980);
nand U13003 (N_13003,N_9225,N_9793);
or U13004 (N_13004,N_10774,N_10485);
nor U13005 (N_13005,N_9561,N_9538);
nor U13006 (N_13006,N_10659,N_9354);
and U13007 (N_13007,N_9518,N_9896);
nor U13008 (N_13008,N_10523,N_11234);
nor U13009 (N_13009,N_10658,N_9201);
or U13010 (N_13010,N_10955,N_10804);
nor U13011 (N_13011,N_9546,N_10528);
or U13012 (N_13012,N_9282,N_9639);
and U13013 (N_13013,N_11447,N_10111);
and U13014 (N_13014,N_9689,N_10349);
or U13015 (N_13015,N_11511,N_10692);
nor U13016 (N_13016,N_11502,N_10036);
or U13017 (N_13017,N_9468,N_11764);
or U13018 (N_13018,N_10281,N_10415);
nand U13019 (N_13019,N_9822,N_9465);
nand U13020 (N_13020,N_11949,N_11422);
nand U13021 (N_13021,N_9804,N_10964);
nor U13022 (N_13022,N_9929,N_10202);
nor U13023 (N_13023,N_10499,N_9293);
or U13024 (N_13024,N_11789,N_9398);
and U13025 (N_13025,N_11413,N_10879);
and U13026 (N_13026,N_11089,N_10644);
or U13027 (N_13027,N_10264,N_9338);
and U13028 (N_13028,N_10520,N_9819);
or U13029 (N_13029,N_11370,N_9040);
xor U13030 (N_13030,N_9960,N_10001);
nand U13031 (N_13031,N_10073,N_11659);
nand U13032 (N_13032,N_10677,N_11433);
and U13033 (N_13033,N_11774,N_10031);
and U13034 (N_13034,N_10834,N_9773);
or U13035 (N_13035,N_10056,N_10886);
and U13036 (N_13036,N_10255,N_10267);
nor U13037 (N_13037,N_11925,N_9937);
or U13038 (N_13038,N_10076,N_9393);
nor U13039 (N_13039,N_9088,N_11177);
nor U13040 (N_13040,N_9107,N_10218);
nand U13041 (N_13041,N_9985,N_10534);
or U13042 (N_13042,N_11587,N_10101);
and U13043 (N_13043,N_9053,N_10766);
nor U13044 (N_13044,N_11091,N_10830);
or U13045 (N_13045,N_9974,N_9427);
and U13046 (N_13046,N_9758,N_11608);
nand U13047 (N_13047,N_11009,N_11160);
and U13048 (N_13048,N_9786,N_9908);
and U13049 (N_13049,N_11725,N_11868);
or U13050 (N_13050,N_11722,N_11898);
or U13051 (N_13051,N_11551,N_9768);
nor U13052 (N_13052,N_10085,N_9593);
and U13053 (N_13053,N_11138,N_9261);
or U13054 (N_13054,N_10409,N_9001);
nor U13055 (N_13055,N_9611,N_10432);
or U13056 (N_13056,N_9166,N_10091);
and U13057 (N_13057,N_9801,N_10934);
nand U13058 (N_13058,N_11251,N_9607);
and U13059 (N_13059,N_10149,N_9110);
nor U13060 (N_13060,N_11016,N_9432);
nor U13061 (N_13061,N_10730,N_11249);
nand U13062 (N_13062,N_10695,N_10816);
nor U13063 (N_13063,N_10194,N_10421);
and U13064 (N_13064,N_11671,N_9942);
nand U13065 (N_13065,N_11472,N_9851);
or U13066 (N_13066,N_10674,N_9904);
and U13067 (N_13067,N_10634,N_9233);
and U13068 (N_13068,N_9355,N_10125);
and U13069 (N_13069,N_10992,N_11364);
or U13070 (N_13070,N_11449,N_9860);
nand U13071 (N_13071,N_9108,N_9662);
and U13072 (N_13072,N_10986,N_10346);
nor U13073 (N_13073,N_9833,N_10235);
or U13074 (N_13074,N_11187,N_9802);
nand U13075 (N_13075,N_10471,N_11469);
and U13076 (N_13076,N_11797,N_9785);
and U13077 (N_13077,N_11904,N_11312);
nor U13078 (N_13078,N_11167,N_9080);
and U13079 (N_13079,N_9857,N_11055);
nand U13080 (N_13080,N_11384,N_9099);
and U13081 (N_13081,N_10811,N_9104);
or U13082 (N_13082,N_10844,N_10863);
nand U13083 (N_13083,N_10973,N_9550);
nor U13084 (N_13084,N_11480,N_11590);
nand U13085 (N_13085,N_9575,N_9267);
nand U13086 (N_13086,N_9081,N_9144);
nor U13087 (N_13087,N_10533,N_9366);
nor U13088 (N_13088,N_10768,N_10249);
and U13089 (N_13089,N_11356,N_11498);
nand U13090 (N_13090,N_11377,N_10314);
and U13091 (N_13091,N_11425,N_9207);
nor U13092 (N_13092,N_10312,N_10994);
or U13093 (N_13093,N_11034,N_9193);
nor U13094 (N_13094,N_9200,N_9495);
nor U13095 (N_13095,N_11694,N_10436);
nor U13096 (N_13096,N_10035,N_10197);
nor U13097 (N_13097,N_9673,N_10983);
and U13098 (N_13098,N_9653,N_11117);
nand U13099 (N_13099,N_10743,N_11326);
or U13100 (N_13100,N_11163,N_9146);
nand U13101 (N_13101,N_10784,N_9797);
and U13102 (N_13102,N_10684,N_11711);
and U13103 (N_13103,N_9571,N_11568);
or U13104 (N_13104,N_10495,N_10305);
nand U13105 (N_13105,N_9169,N_11864);
and U13106 (N_13106,N_11877,N_11288);
nor U13107 (N_13107,N_10838,N_11436);
nor U13108 (N_13108,N_10043,N_11903);
and U13109 (N_13109,N_9552,N_10297);
and U13110 (N_13110,N_11560,N_11379);
nor U13111 (N_13111,N_9675,N_9373);
nand U13112 (N_13112,N_9494,N_9070);
nor U13113 (N_13113,N_9721,N_9696);
nor U13114 (N_13114,N_10315,N_10430);
and U13115 (N_13115,N_9449,N_9514);
and U13116 (N_13116,N_9079,N_10050);
nor U13117 (N_13117,N_9256,N_9248);
nor U13118 (N_13118,N_11348,N_9646);
and U13119 (N_13119,N_9753,N_10798);
or U13120 (N_13120,N_11371,N_10422);
nand U13121 (N_13121,N_10208,N_10224);
nor U13122 (N_13122,N_10322,N_11543);
nand U13123 (N_13123,N_9880,N_10624);
or U13124 (N_13124,N_10411,N_11887);
and U13125 (N_13125,N_11748,N_10871);
nand U13126 (N_13126,N_10925,N_11559);
nand U13127 (N_13127,N_9368,N_10420);
nand U13128 (N_13128,N_10906,N_9153);
nor U13129 (N_13129,N_11518,N_10507);
nand U13130 (N_13130,N_11541,N_11721);
or U13131 (N_13131,N_9573,N_11393);
and U13132 (N_13132,N_10544,N_10918);
nor U13133 (N_13133,N_11697,N_11857);
nor U13134 (N_13134,N_11978,N_10141);
and U13135 (N_13135,N_10285,N_11258);
or U13136 (N_13136,N_11000,N_10304);
nor U13137 (N_13137,N_10706,N_10340);
or U13138 (N_13138,N_11609,N_9806);
nand U13139 (N_13139,N_9405,N_10573);
nand U13140 (N_13140,N_10586,N_9245);
nand U13141 (N_13141,N_11816,N_10668);
and U13142 (N_13142,N_10309,N_10850);
or U13143 (N_13143,N_11399,N_11043);
and U13144 (N_13144,N_10176,N_11524);
and U13145 (N_13145,N_10060,N_11269);
nor U13146 (N_13146,N_9557,N_9812);
and U13147 (N_13147,N_9182,N_10529);
nor U13148 (N_13148,N_10047,N_10704);
and U13149 (N_13149,N_9119,N_9628);
and U13150 (N_13150,N_11942,N_11651);
or U13151 (N_13151,N_9619,N_11526);
and U13152 (N_13152,N_11673,N_9017);
nor U13153 (N_13153,N_9672,N_11880);
and U13154 (N_13154,N_11283,N_10148);
and U13155 (N_13155,N_11906,N_9148);
nor U13156 (N_13156,N_11801,N_9084);
and U13157 (N_13157,N_9409,N_10062);
nand U13158 (N_13158,N_9596,N_9966);
and U13159 (N_13159,N_10783,N_10368);
and U13160 (N_13160,N_9519,N_11036);
nor U13161 (N_13161,N_10592,N_10870);
or U13162 (N_13162,N_11889,N_10685);
or U13163 (N_13163,N_11424,N_9717);
nand U13164 (N_13164,N_10979,N_11051);
nand U13165 (N_13165,N_10505,N_11322);
and U13166 (N_13166,N_11540,N_10756);
or U13167 (N_13167,N_10917,N_9982);
or U13168 (N_13168,N_10900,N_9917);
nor U13169 (N_13169,N_9150,N_9489);
nand U13170 (N_13170,N_11319,N_10950);
nor U13171 (N_13171,N_10363,N_9096);
xnor U13172 (N_13172,N_9988,N_10818);
nand U13173 (N_13173,N_10585,N_10603);
and U13174 (N_13174,N_9838,N_10679);
nor U13175 (N_13175,N_10715,N_9499);
or U13176 (N_13176,N_11419,N_10011);
nand U13177 (N_13177,N_11851,N_11462);
or U13178 (N_13178,N_10525,N_9041);
nor U13179 (N_13179,N_11378,N_11763);
nand U13180 (N_13180,N_9765,N_10642);
and U13181 (N_13181,N_9964,N_10510);
and U13182 (N_13182,N_11192,N_11435);
nor U13183 (N_13183,N_9054,N_9467);
nor U13184 (N_13184,N_9045,N_9861);
nor U13185 (N_13185,N_10361,N_10200);
nor U13186 (N_13186,N_10034,N_9920);
and U13187 (N_13187,N_10405,N_9995);
nor U13188 (N_13188,N_9056,N_9515);
and U13189 (N_13189,N_11010,N_10097);
and U13190 (N_13190,N_10167,N_9034);
nand U13191 (N_13191,N_9180,N_10803);
or U13192 (N_13192,N_9986,N_10119);
and U13193 (N_13193,N_11048,N_11548);
nor U13194 (N_13194,N_9532,N_10136);
or U13195 (N_13195,N_9283,N_11703);
and U13196 (N_13196,N_9131,N_10861);
or U13197 (N_13197,N_10893,N_11989);
and U13198 (N_13198,N_9272,N_11255);
or U13199 (N_13199,N_11461,N_9850);
nand U13200 (N_13200,N_9898,N_10387);
xnor U13201 (N_13201,N_10323,N_10484);
xnor U13202 (N_13202,N_10935,N_10833);
nor U13203 (N_13203,N_11505,N_11076);
and U13204 (N_13204,N_9864,N_9656);
and U13205 (N_13205,N_10131,N_9356);
and U13206 (N_13206,N_9091,N_9905);
and U13207 (N_13207,N_10890,N_11151);
nor U13208 (N_13208,N_10632,N_10576);
nor U13209 (N_13209,N_9513,N_10903);
and U13210 (N_13210,N_10187,N_9827);
nor U13211 (N_13211,N_11488,N_11049);
nand U13212 (N_13212,N_11294,N_11477);
or U13213 (N_13213,N_10750,N_9755);
nor U13214 (N_13214,N_10899,N_10707);
xor U13215 (N_13215,N_9118,N_10082);
or U13216 (N_13216,N_9771,N_11270);
and U13217 (N_13217,N_11489,N_10915);
or U13218 (N_13218,N_10071,N_10557);
or U13219 (N_13219,N_10509,N_9665);
nand U13220 (N_13220,N_11788,N_11656);
or U13221 (N_13221,N_10922,N_9894);
nor U13222 (N_13222,N_9324,N_11417);
or U13223 (N_13223,N_10703,N_9192);
or U13224 (N_13224,N_11828,N_11268);
or U13225 (N_13225,N_10908,N_11600);
nand U13226 (N_13226,N_9522,N_10250);
or U13227 (N_13227,N_9092,N_10258);
and U13228 (N_13228,N_10513,N_11487);
or U13229 (N_13229,N_9888,N_10095);
nor U13230 (N_13230,N_11426,N_10611);
and U13231 (N_13231,N_10221,N_11216);
and U13232 (N_13232,N_9913,N_11601);
nand U13233 (N_13233,N_9594,N_10252);
and U13234 (N_13234,N_10500,N_11197);
nor U13235 (N_13235,N_11770,N_10067);
or U13236 (N_13236,N_9531,N_9700);
and U13237 (N_13237,N_9975,N_10280);
nor U13238 (N_13238,N_9697,N_9075);
nand U13239 (N_13239,N_11962,N_11702);
nor U13240 (N_13240,N_11289,N_9897);
nand U13241 (N_13241,N_10943,N_10295);
nor U13242 (N_13242,N_11190,N_10949);
nand U13243 (N_13243,N_11250,N_10789);
and U13244 (N_13244,N_10128,N_10198);
and U13245 (N_13245,N_11675,N_10021);
or U13246 (N_13246,N_9255,N_10380);
nand U13247 (N_13247,N_9709,N_11795);
or U13248 (N_13248,N_9204,N_9298);
and U13249 (N_13249,N_9128,N_11879);
nand U13250 (N_13250,N_9996,N_9955);
xor U13251 (N_13251,N_10376,N_9712);
or U13252 (N_13252,N_11674,N_10015);
or U13253 (N_13253,N_9212,N_10303);
nand U13254 (N_13254,N_9330,N_9583);
nor U13255 (N_13255,N_10355,N_9997);
and U13256 (N_13256,N_11824,N_9744);
or U13257 (N_13257,N_11157,N_11523);
nand U13258 (N_13258,N_10652,N_11305);
nand U13259 (N_13259,N_10609,N_9638);
nand U13260 (N_13260,N_9691,N_9254);
and U13261 (N_13261,N_9050,N_11604);
or U13262 (N_13262,N_9605,N_10135);
xnor U13263 (N_13263,N_10892,N_9576);
nor U13264 (N_13264,N_11193,N_11017);
nor U13265 (N_13265,N_11431,N_11323);
nand U13266 (N_13266,N_9311,N_9542);
nor U13267 (N_13267,N_10790,N_9723);
nor U13268 (N_13268,N_11264,N_11597);
nand U13269 (N_13269,N_11073,N_11641);
nor U13270 (N_13270,N_11024,N_9844);
or U13271 (N_13271,N_11078,N_9388);
nor U13272 (N_13272,N_9371,N_9501);
and U13273 (N_13273,N_11292,N_10736);
or U13274 (N_13274,N_10127,N_9307);
or U13275 (N_13275,N_10442,N_9164);
nand U13276 (N_13276,N_9469,N_11327);
nor U13277 (N_13277,N_10954,N_9509);
nand U13278 (N_13278,N_10930,N_9423);
nand U13279 (N_13279,N_9105,N_10378);
and U13280 (N_13280,N_9052,N_11687);
and U13281 (N_13281,N_10282,N_9435);
or U13282 (N_13282,N_11001,N_10425);
or U13283 (N_13283,N_10407,N_11241);
or U13284 (N_13284,N_11545,N_11817);
or U13285 (N_13285,N_11679,N_10205);
or U13286 (N_13286,N_11408,N_10456);
or U13287 (N_13287,N_9572,N_9654);
nor U13288 (N_13288,N_10788,N_10751);
or U13289 (N_13289,N_11464,N_11035);
nand U13290 (N_13290,N_11924,N_9451);
or U13291 (N_13291,N_11854,N_11102);
nand U13292 (N_13292,N_10614,N_10369);
and U13293 (N_13293,N_9141,N_9226);
and U13294 (N_13294,N_9560,N_11259);
or U13295 (N_13295,N_11793,N_10263);
nor U13296 (N_13296,N_9490,N_9381);
or U13297 (N_13297,N_11307,N_9983);
nand U13298 (N_13298,N_10519,N_10439);
or U13299 (N_13299,N_9456,N_9630);
and U13300 (N_13300,N_11940,N_9431);
or U13301 (N_13301,N_11338,N_11786);
and U13302 (N_13302,N_11665,N_10326);
and U13303 (N_13303,N_11546,N_9754);
nand U13304 (N_13304,N_10206,N_9138);
nor U13305 (N_13305,N_11738,N_11166);
nor U13306 (N_13306,N_11194,N_10661);
or U13307 (N_13307,N_11246,N_10093);
and U13308 (N_13308,N_9263,N_9971);
and U13309 (N_13309,N_10231,N_10619);
or U13310 (N_13310,N_9564,N_9337);
nand U13311 (N_13311,N_10003,N_11847);
nor U13312 (N_13312,N_11845,N_9634);
nor U13313 (N_13313,N_9147,N_10801);
nand U13314 (N_13314,N_10059,N_9060);
xnor U13315 (N_13315,N_11536,N_10673);
and U13316 (N_13316,N_9476,N_11492);
nand U13317 (N_13317,N_9487,N_10560);
nand U13318 (N_13318,N_9667,N_11385);
and U13319 (N_13319,N_10248,N_9348);
nand U13320 (N_13320,N_9383,N_11460);
nand U13321 (N_13321,N_9931,N_10398);
or U13322 (N_13322,N_10114,N_10165);
nor U13323 (N_13323,N_10969,N_9013);
nand U13324 (N_13324,N_9548,N_11765);
nor U13325 (N_13325,N_11861,N_9784);
nand U13326 (N_13326,N_11220,N_10924);
xor U13327 (N_13327,N_11140,N_10325);
nor U13328 (N_13328,N_11064,N_11726);
or U13329 (N_13329,N_10687,N_10757);
nand U13330 (N_13330,N_9930,N_10171);
or U13331 (N_13331,N_9285,N_11044);
nor U13332 (N_13332,N_10567,N_10540);
nor U13333 (N_13333,N_9210,N_11072);
or U13334 (N_13334,N_11578,N_10618);
or U13335 (N_13335,N_10075,N_11070);
nor U13336 (N_13336,N_9999,N_10327);
and U13337 (N_13337,N_11410,N_11640);
xnor U13338 (N_13338,N_9941,N_9782);
nor U13339 (N_13339,N_9965,N_10945);
nor U13340 (N_13340,N_9016,N_10089);
nor U13341 (N_13341,N_10647,N_9708);
and U13342 (N_13342,N_9417,N_10999);
and U13343 (N_13343,N_11983,N_9698);
nor U13344 (N_13344,N_11968,N_9821);
and U13345 (N_13345,N_10402,N_9818);
or U13346 (N_13346,N_11552,N_11423);
and U13347 (N_13347,N_11849,N_11094);
nor U13348 (N_13348,N_9271,N_10785);
nor U13349 (N_13349,N_11605,N_11483);
nor U13350 (N_13350,N_11596,N_11199);
or U13351 (N_13351,N_11937,N_10676);
nor U13352 (N_13352,N_11707,N_11390);
nor U13353 (N_13353,N_11948,N_9341);
or U13354 (N_13354,N_10732,N_9362);
nand U13355 (N_13355,N_10617,N_11325);
and U13356 (N_13356,N_9916,N_9938);
or U13357 (N_13357,N_10610,N_10017);
nand U13358 (N_13358,N_11744,N_9795);
or U13359 (N_13359,N_11768,N_10238);
nor U13360 (N_13360,N_11253,N_9589);
or U13361 (N_13361,N_10470,N_10601);
nand U13362 (N_13362,N_11520,N_10701);
and U13363 (N_13363,N_11752,N_11161);
and U13364 (N_13364,N_9323,N_10462);
and U13365 (N_13365,N_9516,N_11155);
or U13366 (N_13366,N_11571,N_11639);
nor U13367 (N_13367,N_9762,N_10806);
or U13368 (N_13368,N_9746,N_9174);
or U13369 (N_13369,N_10163,N_10433);
and U13370 (N_13370,N_10891,N_9526);
nor U13371 (N_13371,N_9172,N_11934);
and U13372 (N_13372,N_9242,N_10537);
xnor U13373 (N_13373,N_10086,N_9375);
and U13374 (N_13374,N_9621,N_10793);
or U13375 (N_13375,N_11862,N_11342);
or U13376 (N_13376,N_9738,N_9044);
or U13377 (N_13377,N_9441,N_9504);
nand U13378 (N_13378,N_9130,N_9218);
nand U13379 (N_13379,N_11347,N_9629);
nand U13380 (N_13380,N_10581,N_9814);
nand U13381 (N_13381,N_9928,N_9919);
nand U13382 (N_13382,N_11683,N_9312);
or U13383 (N_13383,N_11443,N_11052);
nor U13384 (N_13384,N_10014,N_10773);
or U13385 (N_13385,N_9319,N_11125);
or U13386 (N_13386,N_9231,N_11005);
and U13387 (N_13387,N_11647,N_9286);
nor U13388 (N_13388,N_10096,N_10476);
nand U13389 (N_13389,N_9008,N_11412);
or U13390 (N_13390,N_11330,N_10843);
nand U13391 (N_13391,N_11914,N_10074);
and U13392 (N_13392,N_10671,N_11247);
and U13393 (N_13393,N_9301,N_11252);
nand U13394 (N_13394,N_11833,N_9962);
or U13395 (N_13395,N_9933,N_9425);
nand U13396 (N_13396,N_10920,N_10717);
and U13397 (N_13397,N_9598,N_10078);
nor U13398 (N_13398,N_9033,N_9865);
nor U13399 (N_13399,N_10885,N_11185);
nor U13400 (N_13400,N_10877,N_9295);
nor U13401 (N_13401,N_11282,N_11037);
or U13402 (N_13402,N_11843,N_9321);
and U13403 (N_13403,N_10107,N_11159);
or U13404 (N_13404,N_10522,N_9010);
nor U13405 (N_13405,N_11057,N_10301);
and U13406 (N_13406,N_11503,N_9203);
and U13407 (N_13407,N_10822,N_11750);
or U13408 (N_13408,N_11950,N_11491);
or U13409 (N_13409,N_10670,N_10780);
nor U13410 (N_13410,N_11065,N_11521);
or U13411 (N_13411,N_10776,N_9039);
and U13412 (N_13412,N_9614,N_9525);
nand U13413 (N_13413,N_10859,N_11827);
nand U13414 (N_13414,N_10588,N_9156);
nor U13415 (N_13415,N_9378,N_11367);
and U13416 (N_13416,N_10151,N_10654);
and U13417 (N_13417,N_10382,N_9579);
and U13418 (N_13418,N_10594,N_11607);
nand U13419 (N_13419,N_11147,N_9442);
nand U13420 (N_13420,N_11615,N_11096);
nand U13421 (N_13421,N_11113,N_11351);
nor U13422 (N_13422,N_9143,N_10995);
and U13423 (N_13423,N_11852,N_10897);
or U13424 (N_13424,N_9270,N_11038);
nand U13425 (N_13425,N_11183,N_10772);
or U13426 (N_13426,N_10815,N_11100);
or U13427 (N_13427,N_11891,N_10242);
nor U13428 (N_13428,N_9055,N_9474);
nor U13429 (N_13429,N_11142,N_10993);
nand U13430 (N_13430,N_9693,N_10256);
and U13431 (N_13431,N_11441,N_9090);
and U13432 (N_13432,N_10735,N_10162);
nor U13433 (N_13433,N_9262,N_11581);
or U13434 (N_13434,N_11317,N_10808);
or U13435 (N_13435,N_9642,N_10638);
and U13436 (N_13436,N_11260,N_9510);
nand U13437 (N_13437,N_11799,N_11136);
or U13438 (N_13438,N_9437,N_11309);
nand U13439 (N_13439,N_11975,N_10469);
and U13440 (N_13440,N_9808,N_10564);
and U13441 (N_13441,N_11340,N_11274);
and U13442 (N_13442,N_10856,N_11617);
and U13443 (N_13443,N_9669,N_9659);
and U13444 (N_13444,N_11684,N_10360);
nor U13445 (N_13445,N_9257,N_11189);
nand U13446 (N_13446,N_11372,N_10599);
nor U13447 (N_13447,N_11747,N_9608);
nand U13448 (N_13448,N_9191,N_11042);
and U13449 (N_13449,N_11075,N_10054);
or U13450 (N_13450,N_11141,N_11643);
nand U13451 (N_13451,N_11790,N_10809);
nand U13452 (N_13452,N_10106,N_9549);
or U13453 (N_13453,N_9124,N_10826);
or U13454 (N_13454,N_9429,N_10488);
nor U13455 (N_13455,N_10546,N_10298);
nor U13456 (N_13456,N_9848,N_11773);
and U13457 (N_13457,N_10579,N_9259);
nor U13458 (N_13458,N_11515,N_11285);
and U13459 (N_13459,N_9891,N_10940);
nor U13460 (N_13460,N_10966,N_11835);
and U13461 (N_13461,N_11681,N_11098);
and U13462 (N_13462,N_9577,N_9890);
nand U13463 (N_13463,N_9924,N_11374);
nor U13464 (N_13464,N_10664,N_10747);
or U13465 (N_13465,N_11621,N_9622);
and U13466 (N_13466,N_11031,N_11606);
or U13467 (N_13467,N_11635,N_11202);
and U13468 (N_13468,N_11208,N_10554);
and U13469 (N_13469,N_10781,N_10615);
nor U13470 (N_13470,N_9497,N_10725);
and U13471 (N_13471,N_11011,N_9831);
and U13472 (N_13472,N_10108,N_9910);
nor U13473 (N_13473,N_9957,N_9720);
and U13474 (N_13474,N_9014,N_10566);
nand U13475 (N_13475,N_11092,N_9057);
nand U13476 (N_13476,N_9121,N_11329);
or U13477 (N_13477,N_9276,N_10649);
or U13478 (N_13478,N_11886,N_10853);
or U13479 (N_13479,N_9176,N_10957);
nor U13480 (N_13480,N_10051,N_9968);
nor U13481 (N_13481,N_9961,N_9264);
nand U13482 (N_13482,N_11407,N_11800);
nand U13483 (N_13483,N_10399,N_11212);
or U13484 (N_13484,N_9395,N_11394);
or U13485 (N_13485,N_9636,N_9637);
nor U13486 (N_13486,N_9447,N_9763);
or U13487 (N_13487,N_10984,N_9918);
nand U13488 (N_13488,N_11176,N_10191);
and U13489 (N_13489,N_11215,N_10961);
or U13490 (N_13490,N_10364,N_9403);
or U13491 (N_13491,N_10598,N_9136);
or U13492 (N_13492,N_11696,N_10667);
or U13493 (N_13493,N_9087,N_10342);
and U13494 (N_13494,N_10458,N_11842);
nor U13495 (N_13495,N_9304,N_9907);
nand U13496 (N_13496,N_11482,N_9722);
or U13497 (N_13497,N_10514,N_9186);
nand U13498 (N_13498,N_9394,N_10777);
and U13499 (N_13499,N_11550,N_9213);
nand U13500 (N_13500,N_11300,N_11954);
nor U13501 (N_13501,N_10192,N_11131);
nor U13502 (N_13502,N_11509,N_10544);
nand U13503 (N_13503,N_10445,N_9506);
nand U13504 (N_13504,N_10506,N_10791);
and U13505 (N_13505,N_11001,N_9080);
nand U13506 (N_13506,N_10459,N_11104);
and U13507 (N_13507,N_10637,N_11775);
xor U13508 (N_13508,N_10912,N_11354);
or U13509 (N_13509,N_10738,N_9360);
and U13510 (N_13510,N_10197,N_11955);
nand U13511 (N_13511,N_9204,N_9908);
nor U13512 (N_13512,N_11423,N_10692);
or U13513 (N_13513,N_9906,N_11373);
or U13514 (N_13514,N_9156,N_9839);
nand U13515 (N_13515,N_11605,N_10058);
and U13516 (N_13516,N_9451,N_9587);
nand U13517 (N_13517,N_10527,N_9865);
nor U13518 (N_13518,N_11506,N_11638);
or U13519 (N_13519,N_9304,N_11225);
or U13520 (N_13520,N_11656,N_10563);
and U13521 (N_13521,N_11268,N_11250);
nor U13522 (N_13522,N_9120,N_10778);
or U13523 (N_13523,N_9378,N_10746);
xor U13524 (N_13524,N_11535,N_11065);
and U13525 (N_13525,N_9858,N_10276);
nand U13526 (N_13526,N_11248,N_11863);
nand U13527 (N_13527,N_11523,N_11167);
nand U13528 (N_13528,N_10712,N_10059);
nor U13529 (N_13529,N_9481,N_9170);
nor U13530 (N_13530,N_11770,N_11386);
nand U13531 (N_13531,N_10337,N_9574);
and U13532 (N_13532,N_10013,N_11135);
or U13533 (N_13533,N_9997,N_9370);
nand U13534 (N_13534,N_11723,N_9270);
nand U13535 (N_13535,N_10361,N_11270);
nor U13536 (N_13536,N_11184,N_10902);
and U13537 (N_13537,N_11855,N_9023);
and U13538 (N_13538,N_9781,N_11475);
or U13539 (N_13539,N_10749,N_10298);
or U13540 (N_13540,N_9435,N_9665);
or U13541 (N_13541,N_9379,N_9283);
and U13542 (N_13542,N_10673,N_11957);
nor U13543 (N_13543,N_9099,N_11467);
nor U13544 (N_13544,N_10821,N_11553);
and U13545 (N_13545,N_9103,N_9323);
nand U13546 (N_13546,N_10632,N_11240);
nor U13547 (N_13547,N_11264,N_9192);
and U13548 (N_13548,N_9870,N_9961);
and U13549 (N_13549,N_11126,N_9596);
nor U13550 (N_13550,N_11779,N_10779);
nand U13551 (N_13551,N_9635,N_10987);
and U13552 (N_13552,N_10470,N_10353);
and U13553 (N_13553,N_10013,N_9352);
and U13554 (N_13554,N_9204,N_9143);
nor U13555 (N_13555,N_9985,N_9510);
and U13556 (N_13556,N_9923,N_10106);
and U13557 (N_13557,N_9261,N_10317);
nand U13558 (N_13558,N_10924,N_10468);
nor U13559 (N_13559,N_11081,N_9174);
or U13560 (N_13560,N_9906,N_10179);
or U13561 (N_13561,N_10840,N_9527);
or U13562 (N_13562,N_11128,N_9777);
nor U13563 (N_13563,N_9486,N_9872);
or U13564 (N_13564,N_9979,N_10405);
nor U13565 (N_13565,N_10410,N_11649);
or U13566 (N_13566,N_10703,N_11687);
nand U13567 (N_13567,N_11119,N_10732);
nor U13568 (N_13568,N_11590,N_9494);
nor U13569 (N_13569,N_11960,N_11643);
or U13570 (N_13570,N_9385,N_10267);
nand U13571 (N_13571,N_11897,N_9707);
nor U13572 (N_13572,N_9208,N_9843);
nor U13573 (N_13573,N_11927,N_11571);
nand U13574 (N_13574,N_11141,N_9484);
and U13575 (N_13575,N_9529,N_11145);
and U13576 (N_13576,N_11782,N_9002);
nand U13577 (N_13577,N_10704,N_11987);
nand U13578 (N_13578,N_9804,N_10711);
or U13579 (N_13579,N_10017,N_11953);
nand U13580 (N_13580,N_11559,N_10056);
and U13581 (N_13581,N_11896,N_11265);
and U13582 (N_13582,N_10606,N_9463);
or U13583 (N_13583,N_10630,N_9761);
nor U13584 (N_13584,N_11045,N_10383);
or U13585 (N_13585,N_11124,N_11572);
nand U13586 (N_13586,N_9487,N_10506);
or U13587 (N_13587,N_9231,N_9202);
nand U13588 (N_13588,N_11436,N_11364);
and U13589 (N_13589,N_10156,N_10059);
nand U13590 (N_13590,N_11629,N_10512);
nand U13591 (N_13591,N_9756,N_11982);
or U13592 (N_13592,N_11054,N_11472);
nor U13593 (N_13593,N_10453,N_9087);
or U13594 (N_13594,N_11377,N_9109);
and U13595 (N_13595,N_11273,N_9143);
xnor U13596 (N_13596,N_11462,N_11397);
and U13597 (N_13597,N_9704,N_10863);
and U13598 (N_13598,N_9254,N_9031);
and U13599 (N_13599,N_9760,N_9846);
nor U13600 (N_13600,N_9598,N_11839);
or U13601 (N_13601,N_11993,N_10211);
or U13602 (N_13602,N_9116,N_10885);
nand U13603 (N_13603,N_11934,N_10368);
and U13604 (N_13604,N_11571,N_9361);
xnor U13605 (N_13605,N_11975,N_9848);
or U13606 (N_13606,N_11466,N_9847);
or U13607 (N_13607,N_9897,N_9403);
nor U13608 (N_13608,N_9331,N_11983);
and U13609 (N_13609,N_10972,N_9616);
and U13610 (N_13610,N_10792,N_10417);
and U13611 (N_13611,N_9946,N_10791);
nor U13612 (N_13612,N_9196,N_9428);
and U13613 (N_13613,N_10263,N_11983);
and U13614 (N_13614,N_9961,N_9513);
nand U13615 (N_13615,N_10675,N_9136);
and U13616 (N_13616,N_11707,N_11021);
nand U13617 (N_13617,N_11252,N_9405);
nand U13618 (N_13618,N_11287,N_10927);
nor U13619 (N_13619,N_9543,N_10320);
nand U13620 (N_13620,N_11297,N_10082);
nor U13621 (N_13621,N_11096,N_11398);
nor U13622 (N_13622,N_10359,N_11833);
or U13623 (N_13623,N_9296,N_11067);
nor U13624 (N_13624,N_11357,N_10118);
nor U13625 (N_13625,N_10206,N_11580);
and U13626 (N_13626,N_10009,N_10341);
nand U13627 (N_13627,N_10680,N_11149);
nand U13628 (N_13628,N_9063,N_9235);
and U13629 (N_13629,N_11652,N_9575);
and U13630 (N_13630,N_10319,N_9203);
or U13631 (N_13631,N_10360,N_11407);
or U13632 (N_13632,N_11129,N_11603);
nand U13633 (N_13633,N_9220,N_9684);
and U13634 (N_13634,N_11865,N_9568);
nor U13635 (N_13635,N_11199,N_9536);
nor U13636 (N_13636,N_10929,N_11250);
nor U13637 (N_13637,N_10708,N_10943);
nand U13638 (N_13638,N_11247,N_10073);
nor U13639 (N_13639,N_11586,N_10859);
or U13640 (N_13640,N_11735,N_11405);
nor U13641 (N_13641,N_10177,N_9592);
and U13642 (N_13642,N_9687,N_10693);
nor U13643 (N_13643,N_9284,N_9901);
and U13644 (N_13644,N_10615,N_10771);
nand U13645 (N_13645,N_9592,N_9417);
or U13646 (N_13646,N_10882,N_9577);
and U13647 (N_13647,N_11883,N_11089);
and U13648 (N_13648,N_10078,N_11879);
nand U13649 (N_13649,N_11408,N_9749);
nand U13650 (N_13650,N_10770,N_10492);
nor U13651 (N_13651,N_11420,N_9119);
nor U13652 (N_13652,N_11889,N_9544);
or U13653 (N_13653,N_9227,N_11719);
nand U13654 (N_13654,N_9299,N_9729);
nand U13655 (N_13655,N_10162,N_10230);
nand U13656 (N_13656,N_11068,N_9375);
or U13657 (N_13657,N_11478,N_9345);
nor U13658 (N_13658,N_9940,N_10073);
and U13659 (N_13659,N_10001,N_11594);
nor U13660 (N_13660,N_10620,N_10605);
or U13661 (N_13661,N_10332,N_9158);
nand U13662 (N_13662,N_11394,N_9418);
and U13663 (N_13663,N_10894,N_9956);
or U13664 (N_13664,N_11435,N_11908);
and U13665 (N_13665,N_9184,N_11362);
or U13666 (N_13666,N_9673,N_11153);
nand U13667 (N_13667,N_9454,N_9376);
or U13668 (N_13668,N_10034,N_10079);
nand U13669 (N_13669,N_11982,N_10259);
nor U13670 (N_13670,N_11567,N_10887);
nand U13671 (N_13671,N_9877,N_11467);
or U13672 (N_13672,N_10865,N_11382);
and U13673 (N_13673,N_10792,N_11571);
and U13674 (N_13674,N_9320,N_9065);
nand U13675 (N_13675,N_10272,N_10726);
or U13676 (N_13676,N_10528,N_9138);
and U13677 (N_13677,N_11338,N_10301);
nand U13678 (N_13678,N_10660,N_10468);
nand U13679 (N_13679,N_9819,N_9666);
and U13680 (N_13680,N_11761,N_10803);
nand U13681 (N_13681,N_10310,N_10391);
and U13682 (N_13682,N_9120,N_11374);
nor U13683 (N_13683,N_10041,N_11123);
or U13684 (N_13684,N_11156,N_11271);
nor U13685 (N_13685,N_9538,N_9374);
and U13686 (N_13686,N_9205,N_9707);
nand U13687 (N_13687,N_11952,N_11279);
and U13688 (N_13688,N_11792,N_11399);
nand U13689 (N_13689,N_11470,N_10811);
and U13690 (N_13690,N_9857,N_11782);
nor U13691 (N_13691,N_9807,N_10656);
nand U13692 (N_13692,N_9077,N_9626);
nand U13693 (N_13693,N_11767,N_11569);
and U13694 (N_13694,N_11205,N_10874);
nand U13695 (N_13695,N_11164,N_10730);
or U13696 (N_13696,N_11772,N_10359);
and U13697 (N_13697,N_11575,N_10231);
nor U13698 (N_13698,N_11085,N_9145);
nand U13699 (N_13699,N_9091,N_10435);
nor U13700 (N_13700,N_11398,N_10533);
or U13701 (N_13701,N_11981,N_10171);
nor U13702 (N_13702,N_10346,N_9485);
nor U13703 (N_13703,N_10512,N_9473);
nor U13704 (N_13704,N_11821,N_9703);
and U13705 (N_13705,N_11511,N_9512);
or U13706 (N_13706,N_11629,N_9829);
nand U13707 (N_13707,N_11457,N_10404);
nand U13708 (N_13708,N_10000,N_10334);
nor U13709 (N_13709,N_10095,N_10696);
nand U13710 (N_13710,N_11781,N_10101);
nor U13711 (N_13711,N_11533,N_11606);
nand U13712 (N_13712,N_11655,N_11326);
or U13713 (N_13713,N_10688,N_9179);
and U13714 (N_13714,N_11943,N_11269);
and U13715 (N_13715,N_11343,N_11678);
and U13716 (N_13716,N_9214,N_9991);
or U13717 (N_13717,N_10406,N_11677);
and U13718 (N_13718,N_11364,N_9936);
nand U13719 (N_13719,N_9359,N_11738);
nor U13720 (N_13720,N_9023,N_9111);
nor U13721 (N_13721,N_10892,N_10404);
and U13722 (N_13722,N_11010,N_11790);
nand U13723 (N_13723,N_11003,N_11448);
nand U13724 (N_13724,N_10059,N_9673);
or U13725 (N_13725,N_10855,N_10074);
nand U13726 (N_13726,N_9453,N_9082);
nand U13727 (N_13727,N_10895,N_9651);
xnor U13728 (N_13728,N_10100,N_11426);
nand U13729 (N_13729,N_11583,N_9688);
or U13730 (N_13730,N_9213,N_11314);
nand U13731 (N_13731,N_10922,N_9704);
or U13732 (N_13732,N_10058,N_10168);
and U13733 (N_13733,N_9817,N_11620);
nand U13734 (N_13734,N_10886,N_9691);
xor U13735 (N_13735,N_10229,N_9918);
nand U13736 (N_13736,N_10269,N_11404);
nor U13737 (N_13737,N_11963,N_10607);
and U13738 (N_13738,N_10770,N_10995);
nand U13739 (N_13739,N_9979,N_10685);
or U13740 (N_13740,N_10767,N_11135);
and U13741 (N_13741,N_9223,N_9972);
and U13742 (N_13742,N_10950,N_11004);
or U13743 (N_13743,N_10688,N_9519);
and U13744 (N_13744,N_11178,N_11848);
nor U13745 (N_13745,N_9350,N_9258);
and U13746 (N_13746,N_9957,N_10495);
nand U13747 (N_13747,N_11992,N_10963);
or U13748 (N_13748,N_9292,N_9427);
nand U13749 (N_13749,N_9780,N_9579);
and U13750 (N_13750,N_10942,N_11052);
nand U13751 (N_13751,N_10219,N_11392);
or U13752 (N_13752,N_9600,N_10530);
nor U13753 (N_13753,N_9423,N_9277);
or U13754 (N_13754,N_11384,N_9715);
nand U13755 (N_13755,N_9740,N_10460);
or U13756 (N_13756,N_11014,N_11067);
nor U13757 (N_13757,N_11823,N_9354);
or U13758 (N_13758,N_10186,N_10518);
nor U13759 (N_13759,N_11322,N_11368);
nand U13760 (N_13760,N_11367,N_10654);
and U13761 (N_13761,N_9677,N_11946);
nand U13762 (N_13762,N_9356,N_9067);
nor U13763 (N_13763,N_11920,N_10551);
nand U13764 (N_13764,N_10821,N_11255);
and U13765 (N_13765,N_9272,N_9249);
xnor U13766 (N_13766,N_9585,N_10228);
and U13767 (N_13767,N_10113,N_9097);
or U13768 (N_13768,N_10106,N_9742);
and U13769 (N_13769,N_9755,N_10140);
nand U13770 (N_13770,N_11351,N_10541);
and U13771 (N_13771,N_9765,N_11458);
nand U13772 (N_13772,N_9573,N_11261);
nor U13773 (N_13773,N_10201,N_11245);
nor U13774 (N_13774,N_11333,N_11688);
and U13775 (N_13775,N_11215,N_11764);
nand U13776 (N_13776,N_11002,N_10945);
or U13777 (N_13777,N_9342,N_11199);
nand U13778 (N_13778,N_11877,N_11071);
and U13779 (N_13779,N_11696,N_11007);
nor U13780 (N_13780,N_10816,N_9558);
nand U13781 (N_13781,N_9066,N_11772);
nand U13782 (N_13782,N_11116,N_9370);
and U13783 (N_13783,N_9624,N_9369);
nand U13784 (N_13784,N_10975,N_11537);
nor U13785 (N_13785,N_10958,N_11518);
nand U13786 (N_13786,N_9033,N_11724);
nor U13787 (N_13787,N_9161,N_11009);
or U13788 (N_13788,N_10160,N_11595);
and U13789 (N_13789,N_11379,N_11223);
nor U13790 (N_13790,N_10109,N_11652);
nand U13791 (N_13791,N_11009,N_10762);
and U13792 (N_13792,N_10035,N_10264);
nor U13793 (N_13793,N_9202,N_10461);
nor U13794 (N_13794,N_9166,N_10439);
nor U13795 (N_13795,N_9181,N_11655);
and U13796 (N_13796,N_9942,N_10408);
nand U13797 (N_13797,N_10598,N_10709);
or U13798 (N_13798,N_10312,N_10454);
and U13799 (N_13799,N_10601,N_11281);
and U13800 (N_13800,N_10817,N_10564);
and U13801 (N_13801,N_10908,N_10630);
and U13802 (N_13802,N_11068,N_9037);
and U13803 (N_13803,N_9550,N_10098);
and U13804 (N_13804,N_9791,N_11310);
or U13805 (N_13805,N_10420,N_9181);
nand U13806 (N_13806,N_10490,N_10456);
nand U13807 (N_13807,N_10562,N_10389);
and U13808 (N_13808,N_11826,N_10968);
nand U13809 (N_13809,N_10861,N_9940);
or U13810 (N_13810,N_11615,N_10945);
nand U13811 (N_13811,N_11798,N_9107);
nand U13812 (N_13812,N_9509,N_11023);
and U13813 (N_13813,N_11032,N_10036);
and U13814 (N_13814,N_11295,N_11114);
nor U13815 (N_13815,N_11350,N_11829);
or U13816 (N_13816,N_11920,N_10328);
or U13817 (N_13817,N_10710,N_9818);
or U13818 (N_13818,N_9994,N_11657);
and U13819 (N_13819,N_11285,N_11756);
nand U13820 (N_13820,N_10645,N_10307);
and U13821 (N_13821,N_11025,N_10941);
nor U13822 (N_13822,N_11292,N_11133);
and U13823 (N_13823,N_11094,N_9190);
or U13824 (N_13824,N_10755,N_10128);
and U13825 (N_13825,N_11571,N_11975);
or U13826 (N_13826,N_9106,N_10568);
and U13827 (N_13827,N_11588,N_11381);
or U13828 (N_13828,N_9205,N_11630);
and U13829 (N_13829,N_11471,N_11366);
or U13830 (N_13830,N_11872,N_10085);
and U13831 (N_13831,N_9648,N_9639);
or U13832 (N_13832,N_11804,N_9196);
nor U13833 (N_13833,N_9538,N_11824);
and U13834 (N_13834,N_11192,N_9140);
nand U13835 (N_13835,N_9535,N_11334);
and U13836 (N_13836,N_9813,N_9270);
or U13837 (N_13837,N_11707,N_9530);
or U13838 (N_13838,N_9473,N_11037);
and U13839 (N_13839,N_11596,N_9840);
nor U13840 (N_13840,N_11844,N_9062);
nand U13841 (N_13841,N_10691,N_10496);
nand U13842 (N_13842,N_10401,N_11209);
xor U13843 (N_13843,N_9788,N_10551);
or U13844 (N_13844,N_9960,N_11421);
or U13845 (N_13845,N_11505,N_10571);
and U13846 (N_13846,N_10256,N_9291);
nor U13847 (N_13847,N_9201,N_11503);
nor U13848 (N_13848,N_11595,N_9119);
or U13849 (N_13849,N_9299,N_9519);
or U13850 (N_13850,N_11242,N_11183);
nor U13851 (N_13851,N_9298,N_10805);
or U13852 (N_13852,N_11134,N_11173);
nor U13853 (N_13853,N_11623,N_11526);
and U13854 (N_13854,N_9952,N_11240);
nand U13855 (N_13855,N_9770,N_10456);
nor U13856 (N_13856,N_9755,N_9006);
and U13857 (N_13857,N_9458,N_9646);
or U13858 (N_13858,N_9201,N_9682);
or U13859 (N_13859,N_9264,N_9319);
nand U13860 (N_13860,N_9982,N_11112);
nor U13861 (N_13861,N_9821,N_11941);
nor U13862 (N_13862,N_11795,N_10790);
or U13863 (N_13863,N_10452,N_10576);
or U13864 (N_13864,N_11684,N_9165);
nor U13865 (N_13865,N_11341,N_9052);
nand U13866 (N_13866,N_11120,N_10287);
nand U13867 (N_13867,N_10371,N_9158);
and U13868 (N_13868,N_9876,N_10092);
or U13869 (N_13869,N_10453,N_9045);
and U13870 (N_13870,N_10103,N_10106);
nand U13871 (N_13871,N_11765,N_10787);
nand U13872 (N_13872,N_10407,N_9391);
or U13873 (N_13873,N_10046,N_9420);
nand U13874 (N_13874,N_11893,N_9134);
or U13875 (N_13875,N_11902,N_11671);
or U13876 (N_13876,N_10593,N_11341);
nor U13877 (N_13877,N_11668,N_10054);
nor U13878 (N_13878,N_11434,N_11930);
nor U13879 (N_13879,N_11439,N_11284);
and U13880 (N_13880,N_9076,N_9554);
or U13881 (N_13881,N_10708,N_11140);
xnor U13882 (N_13882,N_11172,N_9672);
and U13883 (N_13883,N_10093,N_9584);
or U13884 (N_13884,N_11097,N_10018);
nor U13885 (N_13885,N_10114,N_11777);
nand U13886 (N_13886,N_9453,N_11866);
nor U13887 (N_13887,N_9930,N_11776);
or U13888 (N_13888,N_10266,N_9873);
and U13889 (N_13889,N_11665,N_10085);
nor U13890 (N_13890,N_10038,N_9531);
or U13891 (N_13891,N_9431,N_11713);
or U13892 (N_13892,N_10339,N_11111);
xor U13893 (N_13893,N_9364,N_9548);
or U13894 (N_13894,N_9635,N_11120);
and U13895 (N_13895,N_10095,N_10712);
nor U13896 (N_13896,N_10410,N_9471);
or U13897 (N_13897,N_10406,N_11514);
nor U13898 (N_13898,N_9793,N_10758);
and U13899 (N_13899,N_9274,N_9734);
and U13900 (N_13900,N_10431,N_10101);
nand U13901 (N_13901,N_9304,N_11882);
or U13902 (N_13902,N_10408,N_11961);
and U13903 (N_13903,N_11530,N_9530);
and U13904 (N_13904,N_9790,N_9810);
nor U13905 (N_13905,N_9511,N_10552);
nand U13906 (N_13906,N_11652,N_11292);
nand U13907 (N_13907,N_9503,N_11174);
and U13908 (N_13908,N_9763,N_9446);
or U13909 (N_13909,N_11134,N_11023);
or U13910 (N_13910,N_9909,N_10899);
or U13911 (N_13911,N_9830,N_11809);
nor U13912 (N_13912,N_10867,N_9900);
nor U13913 (N_13913,N_10535,N_11887);
and U13914 (N_13914,N_9642,N_9539);
or U13915 (N_13915,N_11306,N_9231);
and U13916 (N_13916,N_11951,N_11665);
and U13917 (N_13917,N_11983,N_9100);
nor U13918 (N_13918,N_9188,N_10123);
or U13919 (N_13919,N_11718,N_9706);
nand U13920 (N_13920,N_10495,N_9745);
xor U13921 (N_13921,N_10887,N_10938);
or U13922 (N_13922,N_11485,N_9940);
and U13923 (N_13923,N_9724,N_11914);
nor U13924 (N_13924,N_11423,N_11990);
nand U13925 (N_13925,N_9534,N_9478);
nor U13926 (N_13926,N_9958,N_9870);
nor U13927 (N_13927,N_9013,N_10254);
and U13928 (N_13928,N_9462,N_9113);
nand U13929 (N_13929,N_10341,N_10036);
nor U13930 (N_13930,N_9533,N_10779);
and U13931 (N_13931,N_9654,N_10229);
nor U13932 (N_13932,N_10275,N_10135);
nor U13933 (N_13933,N_11372,N_9856);
nor U13934 (N_13934,N_9779,N_9198);
nand U13935 (N_13935,N_11598,N_9379);
nand U13936 (N_13936,N_11374,N_10446);
and U13937 (N_13937,N_11057,N_10115);
nand U13938 (N_13938,N_9549,N_10698);
nor U13939 (N_13939,N_9780,N_10088);
nand U13940 (N_13940,N_9627,N_10185);
nor U13941 (N_13941,N_11740,N_9812);
and U13942 (N_13942,N_11537,N_11607);
nor U13943 (N_13943,N_10070,N_10584);
and U13944 (N_13944,N_10888,N_10232);
nand U13945 (N_13945,N_10013,N_9856);
or U13946 (N_13946,N_10464,N_11066);
and U13947 (N_13947,N_9515,N_10917);
or U13948 (N_13948,N_10733,N_10185);
nand U13949 (N_13949,N_11835,N_11137);
nor U13950 (N_13950,N_9989,N_11002);
xor U13951 (N_13951,N_11689,N_9748);
and U13952 (N_13952,N_9571,N_11677);
and U13953 (N_13953,N_11452,N_9731);
nor U13954 (N_13954,N_10552,N_11188);
nand U13955 (N_13955,N_11800,N_10499);
nor U13956 (N_13956,N_9689,N_9834);
nor U13957 (N_13957,N_9857,N_11788);
or U13958 (N_13958,N_10067,N_10061);
nand U13959 (N_13959,N_11910,N_10083);
nand U13960 (N_13960,N_11645,N_10242);
and U13961 (N_13961,N_11593,N_11710);
nand U13962 (N_13962,N_9442,N_9180);
nor U13963 (N_13963,N_11118,N_9427);
nor U13964 (N_13964,N_11104,N_9915);
nor U13965 (N_13965,N_11966,N_10949);
or U13966 (N_13966,N_10091,N_10392);
xor U13967 (N_13967,N_9781,N_10515);
and U13968 (N_13968,N_9643,N_11970);
nor U13969 (N_13969,N_11505,N_10596);
nor U13970 (N_13970,N_9963,N_10278);
nand U13971 (N_13971,N_9417,N_11923);
or U13972 (N_13972,N_9352,N_11638);
nor U13973 (N_13973,N_10835,N_9523);
nand U13974 (N_13974,N_11505,N_10653);
and U13975 (N_13975,N_11308,N_11502);
nand U13976 (N_13976,N_9967,N_10917);
or U13977 (N_13977,N_9301,N_10971);
and U13978 (N_13978,N_10542,N_9818);
or U13979 (N_13979,N_10613,N_9938);
nand U13980 (N_13980,N_10319,N_9498);
nor U13981 (N_13981,N_9018,N_10952);
or U13982 (N_13982,N_10694,N_11639);
and U13983 (N_13983,N_9222,N_10859);
nor U13984 (N_13984,N_11232,N_11970);
or U13985 (N_13985,N_11456,N_9838);
or U13986 (N_13986,N_9989,N_9505);
nand U13987 (N_13987,N_11646,N_9255);
or U13988 (N_13988,N_10006,N_11916);
nor U13989 (N_13989,N_10832,N_9387);
and U13990 (N_13990,N_10032,N_10069);
or U13991 (N_13991,N_11706,N_10616);
or U13992 (N_13992,N_9413,N_9484);
nand U13993 (N_13993,N_9292,N_9436);
and U13994 (N_13994,N_9529,N_10987);
or U13995 (N_13995,N_9191,N_10074);
and U13996 (N_13996,N_10783,N_11222);
and U13997 (N_13997,N_11738,N_10275);
nand U13998 (N_13998,N_9193,N_11467);
and U13999 (N_13999,N_11604,N_10018);
nand U14000 (N_14000,N_11458,N_10270);
nand U14001 (N_14001,N_11121,N_9022);
or U14002 (N_14002,N_10435,N_9467);
or U14003 (N_14003,N_11400,N_9663);
nand U14004 (N_14004,N_11974,N_9997);
and U14005 (N_14005,N_10567,N_10897);
and U14006 (N_14006,N_11109,N_11759);
or U14007 (N_14007,N_11707,N_9249);
or U14008 (N_14008,N_9417,N_9204);
and U14009 (N_14009,N_10702,N_10903);
nor U14010 (N_14010,N_9551,N_9074);
and U14011 (N_14011,N_9690,N_10859);
or U14012 (N_14012,N_10022,N_9447);
nor U14013 (N_14013,N_10655,N_9386);
nand U14014 (N_14014,N_9589,N_11170);
nand U14015 (N_14015,N_9406,N_9899);
nand U14016 (N_14016,N_9736,N_10206);
nor U14017 (N_14017,N_10764,N_10225);
nor U14018 (N_14018,N_10711,N_9270);
and U14019 (N_14019,N_11648,N_11516);
and U14020 (N_14020,N_10450,N_9426);
xnor U14021 (N_14021,N_11841,N_9241);
nand U14022 (N_14022,N_10232,N_9363);
or U14023 (N_14023,N_11223,N_9404);
nor U14024 (N_14024,N_9503,N_9120);
nand U14025 (N_14025,N_10671,N_9699);
nor U14026 (N_14026,N_10484,N_11217);
and U14027 (N_14027,N_9607,N_11444);
and U14028 (N_14028,N_9843,N_11942);
nor U14029 (N_14029,N_11697,N_10671);
nand U14030 (N_14030,N_10544,N_9035);
and U14031 (N_14031,N_9434,N_11585);
nand U14032 (N_14032,N_9730,N_9307);
nand U14033 (N_14033,N_9162,N_9642);
or U14034 (N_14034,N_9940,N_11451);
or U14035 (N_14035,N_11945,N_10197);
nor U14036 (N_14036,N_10122,N_11991);
and U14037 (N_14037,N_9153,N_11758);
nand U14038 (N_14038,N_10851,N_11314);
and U14039 (N_14039,N_11373,N_9431);
and U14040 (N_14040,N_10404,N_11021);
or U14041 (N_14041,N_10105,N_10498);
nor U14042 (N_14042,N_9858,N_9007);
nor U14043 (N_14043,N_9836,N_10665);
nand U14044 (N_14044,N_10773,N_9638);
nand U14045 (N_14045,N_11228,N_10325);
nand U14046 (N_14046,N_10858,N_9227);
and U14047 (N_14047,N_9628,N_11677);
nand U14048 (N_14048,N_11316,N_10856);
nor U14049 (N_14049,N_9345,N_11848);
nand U14050 (N_14050,N_11852,N_11755);
and U14051 (N_14051,N_9091,N_9551);
and U14052 (N_14052,N_11501,N_11728);
nand U14053 (N_14053,N_9830,N_9514);
and U14054 (N_14054,N_11006,N_10802);
and U14055 (N_14055,N_10531,N_10650);
or U14056 (N_14056,N_11929,N_11194);
xnor U14057 (N_14057,N_10904,N_9866);
nor U14058 (N_14058,N_11880,N_11957);
nand U14059 (N_14059,N_11154,N_10742);
or U14060 (N_14060,N_9939,N_9815);
or U14061 (N_14061,N_11965,N_9781);
and U14062 (N_14062,N_9277,N_11482);
and U14063 (N_14063,N_10184,N_10075);
nand U14064 (N_14064,N_11080,N_9297);
or U14065 (N_14065,N_9609,N_11484);
nor U14066 (N_14066,N_10417,N_10928);
and U14067 (N_14067,N_9564,N_11699);
xnor U14068 (N_14068,N_10530,N_11299);
nor U14069 (N_14069,N_10601,N_9209);
nand U14070 (N_14070,N_9415,N_10063);
and U14071 (N_14071,N_11990,N_10612);
nor U14072 (N_14072,N_10115,N_11268);
or U14073 (N_14073,N_10651,N_10773);
nand U14074 (N_14074,N_9320,N_9177);
and U14075 (N_14075,N_10419,N_11560);
or U14076 (N_14076,N_11209,N_10412);
nand U14077 (N_14077,N_9682,N_11622);
or U14078 (N_14078,N_10796,N_10250);
and U14079 (N_14079,N_10782,N_9290);
and U14080 (N_14080,N_9645,N_11954);
and U14081 (N_14081,N_11738,N_11759);
nor U14082 (N_14082,N_10925,N_9584);
nand U14083 (N_14083,N_10803,N_10893);
nor U14084 (N_14084,N_10026,N_11738);
nand U14085 (N_14085,N_9573,N_10627);
and U14086 (N_14086,N_9662,N_9407);
and U14087 (N_14087,N_9759,N_11269);
nand U14088 (N_14088,N_11583,N_10152);
and U14089 (N_14089,N_9611,N_9784);
and U14090 (N_14090,N_9778,N_10159);
and U14091 (N_14091,N_9761,N_11359);
or U14092 (N_14092,N_10591,N_9159);
nand U14093 (N_14093,N_11295,N_9118);
nand U14094 (N_14094,N_9656,N_10624);
or U14095 (N_14095,N_11758,N_10430);
and U14096 (N_14096,N_10626,N_9497);
or U14097 (N_14097,N_10780,N_9385);
nor U14098 (N_14098,N_10575,N_11115);
or U14099 (N_14099,N_11660,N_11647);
xnor U14100 (N_14100,N_9425,N_10088);
or U14101 (N_14101,N_9944,N_9932);
and U14102 (N_14102,N_9027,N_9894);
or U14103 (N_14103,N_11004,N_11140);
nor U14104 (N_14104,N_11138,N_9325);
and U14105 (N_14105,N_9172,N_10373);
nand U14106 (N_14106,N_9792,N_11503);
or U14107 (N_14107,N_10701,N_9389);
nor U14108 (N_14108,N_9887,N_9403);
nand U14109 (N_14109,N_11294,N_9170);
nand U14110 (N_14110,N_11647,N_10156);
and U14111 (N_14111,N_9689,N_9824);
nand U14112 (N_14112,N_10071,N_11909);
nor U14113 (N_14113,N_10673,N_11592);
nand U14114 (N_14114,N_10391,N_10337);
nor U14115 (N_14115,N_11347,N_9736);
or U14116 (N_14116,N_9740,N_9008);
and U14117 (N_14117,N_9724,N_10637);
nand U14118 (N_14118,N_9461,N_9522);
or U14119 (N_14119,N_10038,N_11488);
nor U14120 (N_14120,N_11471,N_11543);
or U14121 (N_14121,N_11571,N_11038);
or U14122 (N_14122,N_11029,N_11194);
and U14123 (N_14123,N_11131,N_11922);
nand U14124 (N_14124,N_9286,N_10017);
nand U14125 (N_14125,N_9028,N_10518);
or U14126 (N_14126,N_9375,N_11608);
nor U14127 (N_14127,N_10567,N_10454);
nand U14128 (N_14128,N_10251,N_10843);
nor U14129 (N_14129,N_9645,N_11129);
nor U14130 (N_14130,N_10708,N_11877);
nor U14131 (N_14131,N_11259,N_11731);
or U14132 (N_14132,N_10931,N_9257);
or U14133 (N_14133,N_9175,N_10684);
or U14134 (N_14134,N_9636,N_9164);
nor U14135 (N_14135,N_9672,N_9118);
nor U14136 (N_14136,N_11327,N_9224);
and U14137 (N_14137,N_11293,N_10759);
nand U14138 (N_14138,N_11620,N_9197);
or U14139 (N_14139,N_9951,N_10979);
nor U14140 (N_14140,N_11433,N_10466);
nand U14141 (N_14141,N_10419,N_9410);
nor U14142 (N_14142,N_11044,N_10958);
and U14143 (N_14143,N_9844,N_10754);
nand U14144 (N_14144,N_11782,N_9560);
or U14145 (N_14145,N_10910,N_9381);
nand U14146 (N_14146,N_11666,N_11191);
or U14147 (N_14147,N_11311,N_9507);
nand U14148 (N_14148,N_10062,N_10691);
nand U14149 (N_14149,N_9740,N_11494);
and U14150 (N_14150,N_11905,N_9813);
nor U14151 (N_14151,N_9756,N_11668);
nor U14152 (N_14152,N_9138,N_9353);
nand U14153 (N_14153,N_9212,N_11553);
and U14154 (N_14154,N_9596,N_11733);
nand U14155 (N_14155,N_10889,N_10691);
and U14156 (N_14156,N_11890,N_10118);
or U14157 (N_14157,N_10291,N_10083);
nor U14158 (N_14158,N_9917,N_11885);
nand U14159 (N_14159,N_11379,N_10771);
or U14160 (N_14160,N_10888,N_9416);
or U14161 (N_14161,N_10701,N_9754);
xor U14162 (N_14162,N_10323,N_11101);
or U14163 (N_14163,N_10670,N_11811);
xnor U14164 (N_14164,N_9523,N_10172);
or U14165 (N_14165,N_10880,N_11923);
or U14166 (N_14166,N_11183,N_10533);
nor U14167 (N_14167,N_11198,N_11715);
nand U14168 (N_14168,N_11307,N_9777);
nor U14169 (N_14169,N_10370,N_9753);
nor U14170 (N_14170,N_9596,N_9887);
or U14171 (N_14171,N_11073,N_11213);
nor U14172 (N_14172,N_11453,N_10213);
or U14173 (N_14173,N_10526,N_10993);
and U14174 (N_14174,N_10877,N_9636);
or U14175 (N_14175,N_9367,N_10836);
or U14176 (N_14176,N_9330,N_11409);
nand U14177 (N_14177,N_11984,N_9299);
nand U14178 (N_14178,N_10009,N_9671);
nor U14179 (N_14179,N_10477,N_9780);
xor U14180 (N_14180,N_11656,N_9708);
or U14181 (N_14181,N_10304,N_9835);
or U14182 (N_14182,N_10763,N_9105);
or U14183 (N_14183,N_11319,N_11488);
or U14184 (N_14184,N_10009,N_9055);
xor U14185 (N_14185,N_10047,N_9206);
nand U14186 (N_14186,N_9098,N_9946);
nand U14187 (N_14187,N_10600,N_11090);
nor U14188 (N_14188,N_9529,N_11193);
nor U14189 (N_14189,N_10122,N_11085);
and U14190 (N_14190,N_9832,N_10981);
nor U14191 (N_14191,N_10872,N_9305);
nor U14192 (N_14192,N_9295,N_10541);
and U14193 (N_14193,N_9519,N_10111);
or U14194 (N_14194,N_10620,N_11068);
nand U14195 (N_14195,N_9672,N_11829);
nor U14196 (N_14196,N_10864,N_9161);
nor U14197 (N_14197,N_10404,N_11794);
nor U14198 (N_14198,N_11399,N_9400);
nand U14199 (N_14199,N_11174,N_9806);
nand U14200 (N_14200,N_10474,N_10056);
nor U14201 (N_14201,N_11724,N_10647);
and U14202 (N_14202,N_11914,N_10809);
and U14203 (N_14203,N_9711,N_11046);
or U14204 (N_14204,N_10696,N_11680);
and U14205 (N_14205,N_11720,N_11264);
and U14206 (N_14206,N_10866,N_10628);
and U14207 (N_14207,N_10921,N_11080);
nor U14208 (N_14208,N_10619,N_9000);
nand U14209 (N_14209,N_11786,N_11873);
nor U14210 (N_14210,N_10420,N_10320);
nand U14211 (N_14211,N_9689,N_9430);
nand U14212 (N_14212,N_9008,N_11723);
nor U14213 (N_14213,N_11910,N_11131);
or U14214 (N_14214,N_11884,N_10753);
nor U14215 (N_14215,N_10248,N_11138);
nand U14216 (N_14216,N_9091,N_10019);
and U14217 (N_14217,N_10076,N_9468);
nand U14218 (N_14218,N_10245,N_9956);
nor U14219 (N_14219,N_9297,N_11597);
nor U14220 (N_14220,N_11637,N_9887);
nand U14221 (N_14221,N_9329,N_11290);
nor U14222 (N_14222,N_9464,N_11880);
nand U14223 (N_14223,N_9147,N_11352);
nand U14224 (N_14224,N_11184,N_9687);
or U14225 (N_14225,N_10493,N_10319);
nor U14226 (N_14226,N_10285,N_11234);
nor U14227 (N_14227,N_10879,N_11003);
nand U14228 (N_14228,N_9097,N_9056);
and U14229 (N_14229,N_11608,N_11281);
nand U14230 (N_14230,N_9241,N_9473);
or U14231 (N_14231,N_11875,N_10993);
and U14232 (N_14232,N_11807,N_9497);
and U14233 (N_14233,N_9324,N_9939);
or U14234 (N_14234,N_11414,N_10318);
nor U14235 (N_14235,N_11100,N_11229);
nor U14236 (N_14236,N_11719,N_11828);
or U14237 (N_14237,N_10902,N_10176);
nor U14238 (N_14238,N_10680,N_10245);
and U14239 (N_14239,N_11631,N_11430);
and U14240 (N_14240,N_10785,N_10232);
and U14241 (N_14241,N_9946,N_10935);
or U14242 (N_14242,N_10492,N_10440);
nor U14243 (N_14243,N_10999,N_9744);
and U14244 (N_14244,N_10978,N_10095);
and U14245 (N_14245,N_11430,N_11147);
or U14246 (N_14246,N_11831,N_9153);
nor U14247 (N_14247,N_11480,N_11318);
nand U14248 (N_14248,N_9002,N_9859);
or U14249 (N_14249,N_9480,N_10467);
nand U14250 (N_14250,N_9467,N_10214);
or U14251 (N_14251,N_9417,N_11686);
and U14252 (N_14252,N_9646,N_10508);
and U14253 (N_14253,N_9138,N_11000);
nor U14254 (N_14254,N_11997,N_9140);
nand U14255 (N_14255,N_9775,N_9156);
or U14256 (N_14256,N_9723,N_11996);
or U14257 (N_14257,N_11479,N_11823);
or U14258 (N_14258,N_11477,N_11052);
or U14259 (N_14259,N_10539,N_11686);
and U14260 (N_14260,N_10548,N_10464);
nand U14261 (N_14261,N_9940,N_10629);
nand U14262 (N_14262,N_11223,N_9644);
and U14263 (N_14263,N_11741,N_9232);
nand U14264 (N_14264,N_9107,N_9934);
or U14265 (N_14265,N_9279,N_11792);
and U14266 (N_14266,N_11990,N_10598);
nor U14267 (N_14267,N_11574,N_9154);
nor U14268 (N_14268,N_9312,N_11162);
and U14269 (N_14269,N_11761,N_9820);
nor U14270 (N_14270,N_10265,N_10550);
nand U14271 (N_14271,N_9483,N_10877);
xor U14272 (N_14272,N_9127,N_10162);
or U14273 (N_14273,N_10478,N_9488);
and U14274 (N_14274,N_10570,N_11981);
nand U14275 (N_14275,N_11501,N_11985);
nor U14276 (N_14276,N_11838,N_10828);
nand U14277 (N_14277,N_10750,N_10373);
nor U14278 (N_14278,N_9456,N_10040);
or U14279 (N_14279,N_11411,N_9810);
nor U14280 (N_14280,N_9479,N_9194);
nor U14281 (N_14281,N_10896,N_10701);
nor U14282 (N_14282,N_11905,N_10886);
nand U14283 (N_14283,N_9056,N_10302);
nand U14284 (N_14284,N_10581,N_10281);
nor U14285 (N_14285,N_9341,N_9657);
and U14286 (N_14286,N_11761,N_9192);
nand U14287 (N_14287,N_9858,N_9668);
or U14288 (N_14288,N_11902,N_9457);
nand U14289 (N_14289,N_11885,N_10345);
nand U14290 (N_14290,N_10935,N_11229);
or U14291 (N_14291,N_9569,N_9474);
and U14292 (N_14292,N_10294,N_11820);
nor U14293 (N_14293,N_11058,N_10842);
or U14294 (N_14294,N_10438,N_10333);
and U14295 (N_14295,N_11737,N_10602);
or U14296 (N_14296,N_10420,N_10888);
and U14297 (N_14297,N_9151,N_11602);
or U14298 (N_14298,N_10081,N_9929);
nand U14299 (N_14299,N_9880,N_9217);
or U14300 (N_14300,N_11055,N_11117);
nand U14301 (N_14301,N_11725,N_10314);
or U14302 (N_14302,N_11357,N_11659);
and U14303 (N_14303,N_10130,N_9873);
nor U14304 (N_14304,N_11663,N_10940);
or U14305 (N_14305,N_10523,N_10625);
nand U14306 (N_14306,N_9380,N_9640);
or U14307 (N_14307,N_11962,N_10216);
nand U14308 (N_14308,N_10458,N_10033);
nand U14309 (N_14309,N_11171,N_10153);
nand U14310 (N_14310,N_11965,N_10715);
and U14311 (N_14311,N_10661,N_9337);
or U14312 (N_14312,N_10783,N_9413);
or U14313 (N_14313,N_11761,N_9774);
nor U14314 (N_14314,N_9540,N_11552);
or U14315 (N_14315,N_9217,N_11411);
nand U14316 (N_14316,N_11110,N_10532);
nand U14317 (N_14317,N_11733,N_11085);
nand U14318 (N_14318,N_11218,N_11215);
or U14319 (N_14319,N_11325,N_10595);
or U14320 (N_14320,N_11592,N_10049);
or U14321 (N_14321,N_10431,N_9107);
or U14322 (N_14322,N_9051,N_11802);
nor U14323 (N_14323,N_11271,N_9539);
and U14324 (N_14324,N_11971,N_11910);
nand U14325 (N_14325,N_11854,N_10659);
nor U14326 (N_14326,N_10984,N_11637);
nand U14327 (N_14327,N_10966,N_11016);
or U14328 (N_14328,N_10895,N_9086);
and U14329 (N_14329,N_11964,N_10917);
and U14330 (N_14330,N_10573,N_9846);
or U14331 (N_14331,N_11624,N_11253);
or U14332 (N_14332,N_11880,N_11777);
and U14333 (N_14333,N_10593,N_9652);
nor U14334 (N_14334,N_10446,N_11394);
xor U14335 (N_14335,N_10752,N_10799);
xnor U14336 (N_14336,N_9381,N_10108);
and U14337 (N_14337,N_11773,N_9706);
and U14338 (N_14338,N_9557,N_11924);
and U14339 (N_14339,N_11556,N_9554);
or U14340 (N_14340,N_11866,N_11577);
and U14341 (N_14341,N_10695,N_11757);
nand U14342 (N_14342,N_11628,N_10151);
and U14343 (N_14343,N_10103,N_9373);
or U14344 (N_14344,N_11702,N_9740);
or U14345 (N_14345,N_9545,N_10475);
or U14346 (N_14346,N_9935,N_9667);
or U14347 (N_14347,N_11960,N_11677);
nor U14348 (N_14348,N_11574,N_10512);
and U14349 (N_14349,N_9152,N_11057);
nand U14350 (N_14350,N_10655,N_10950);
and U14351 (N_14351,N_11413,N_10671);
and U14352 (N_14352,N_9199,N_10724);
xnor U14353 (N_14353,N_10586,N_10303);
or U14354 (N_14354,N_9726,N_10123);
and U14355 (N_14355,N_9976,N_10687);
or U14356 (N_14356,N_9618,N_10016);
nand U14357 (N_14357,N_9996,N_11645);
nand U14358 (N_14358,N_10481,N_10190);
or U14359 (N_14359,N_10337,N_10997);
or U14360 (N_14360,N_11249,N_9343);
or U14361 (N_14361,N_9262,N_9208);
or U14362 (N_14362,N_9633,N_11534);
and U14363 (N_14363,N_9870,N_11083);
and U14364 (N_14364,N_11712,N_10679);
nor U14365 (N_14365,N_11192,N_9279);
and U14366 (N_14366,N_11821,N_10564);
nand U14367 (N_14367,N_9806,N_9210);
nand U14368 (N_14368,N_11960,N_9250);
or U14369 (N_14369,N_11867,N_9478);
and U14370 (N_14370,N_11631,N_10178);
nor U14371 (N_14371,N_9771,N_10276);
nor U14372 (N_14372,N_11918,N_9790);
nor U14373 (N_14373,N_9850,N_11865);
or U14374 (N_14374,N_10467,N_11807);
nor U14375 (N_14375,N_11326,N_10232);
or U14376 (N_14376,N_11888,N_11659);
nor U14377 (N_14377,N_9377,N_9739);
or U14378 (N_14378,N_9788,N_10308);
nand U14379 (N_14379,N_10008,N_10201);
nand U14380 (N_14380,N_10043,N_10972);
nand U14381 (N_14381,N_11414,N_10583);
and U14382 (N_14382,N_11931,N_10746);
or U14383 (N_14383,N_11604,N_11771);
nor U14384 (N_14384,N_9100,N_10579);
nor U14385 (N_14385,N_10885,N_11741);
and U14386 (N_14386,N_11462,N_11606);
and U14387 (N_14387,N_11400,N_9279);
and U14388 (N_14388,N_11089,N_10629);
or U14389 (N_14389,N_10933,N_10792);
and U14390 (N_14390,N_10660,N_11893);
and U14391 (N_14391,N_11138,N_11432);
or U14392 (N_14392,N_9521,N_10120);
nor U14393 (N_14393,N_11319,N_10971);
nand U14394 (N_14394,N_10552,N_9555);
nor U14395 (N_14395,N_11251,N_11709);
nor U14396 (N_14396,N_9037,N_9520);
nand U14397 (N_14397,N_9718,N_11824);
or U14398 (N_14398,N_11944,N_10787);
nor U14399 (N_14399,N_9242,N_10643);
nor U14400 (N_14400,N_10973,N_9490);
and U14401 (N_14401,N_9137,N_9667);
xnor U14402 (N_14402,N_11229,N_9709);
and U14403 (N_14403,N_11156,N_10307);
nor U14404 (N_14404,N_10613,N_9272);
or U14405 (N_14405,N_11086,N_10313);
and U14406 (N_14406,N_11730,N_9970);
or U14407 (N_14407,N_10577,N_9279);
or U14408 (N_14408,N_9598,N_11505);
nor U14409 (N_14409,N_10245,N_11880);
nor U14410 (N_14410,N_10950,N_9628);
nand U14411 (N_14411,N_11426,N_10083);
nand U14412 (N_14412,N_11928,N_9287);
nand U14413 (N_14413,N_9933,N_10880);
nand U14414 (N_14414,N_10930,N_9803);
nand U14415 (N_14415,N_11638,N_9859);
and U14416 (N_14416,N_11056,N_11042);
or U14417 (N_14417,N_9271,N_9488);
or U14418 (N_14418,N_10994,N_11158);
and U14419 (N_14419,N_9580,N_11364);
nor U14420 (N_14420,N_11346,N_10197);
nand U14421 (N_14421,N_9328,N_10502);
and U14422 (N_14422,N_10595,N_9695);
and U14423 (N_14423,N_9953,N_11098);
nand U14424 (N_14424,N_10809,N_9170);
and U14425 (N_14425,N_11981,N_10245);
nor U14426 (N_14426,N_9460,N_11594);
nand U14427 (N_14427,N_9927,N_9267);
nor U14428 (N_14428,N_10813,N_11499);
and U14429 (N_14429,N_9620,N_9964);
or U14430 (N_14430,N_10342,N_10978);
nor U14431 (N_14431,N_9911,N_9003);
nand U14432 (N_14432,N_10762,N_11906);
or U14433 (N_14433,N_9796,N_11488);
and U14434 (N_14434,N_11793,N_10984);
nand U14435 (N_14435,N_11228,N_10858);
nand U14436 (N_14436,N_11450,N_10219);
and U14437 (N_14437,N_9976,N_10644);
xor U14438 (N_14438,N_10564,N_10573);
nand U14439 (N_14439,N_10444,N_10722);
nand U14440 (N_14440,N_10113,N_10203);
nand U14441 (N_14441,N_9905,N_11001);
nand U14442 (N_14442,N_9937,N_10907);
nor U14443 (N_14443,N_9915,N_11912);
and U14444 (N_14444,N_10486,N_11274);
nand U14445 (N_14445,N_10338,N_11313);
nor U14446 (N_14446,N_11272,N_10597);
nand U14447 (N_14447,N_10167,N_10743);
or U14448 (N_14448,N_9336,N_10210);
or U14449 (N_14449,N_11129,N_10304);
nor U14450 (N_14450,N_11594,N_10181);
or U14451 (N_14451,N_11507,N_10131);
nand U14452 (N_14452,N_9642,N_9134);
nor U14453 (N_14453,N_11922,N_10128);
or U14454 (N_14454,N_11684,N_10705);
nor U14455 (N_14455,N_11328,N_11579);
nor U14456 (N_14456,N_9720,N_9370);
or U14457 (N_14457,N_10803,N_10332);
nand U14458 (N_14458,N_11240,N_9087);
and U14459 (N_14459,N_10048,N_10731);
or U14460 (N_14460,N_10589,N_11351);
and U14461 (N_14461,N_11005,N_10662);
nand U14462 (N_14462,N_10593,N_11448);
and U14463 (N_14463,N_10796,N_11109);
or U14464 (N_14464,N_9005,N_11588);
nand U14465 (N_14465,N_10126,N_11825);
and U14466 (N_14466,N_11476,N_9362);
xnor U14467 (N_14467,N_11042,N_9560);
and U14468 (N_14468,N_11972,N_11180);
or U14469 (N_14469,N_10240,N_10817);
and U14470 (N_14470,N_10832,N_11817);
and U14471 (N_14471,N_10497,N_9515);
and U14472 (N_14472,N_11482,N_10369);
or U14473 (N_14473,N_10245,N_10623);
nor U14474 (N_14474,N_11145,N_11143);
nand U14475 (N_14475,N_9676,N_9830);
nor U14476 (N_14476,N_11660,N_9381);
nor U14477 (N_14477,N_10094,N_11969);
nor U14478 (N_14478,N_9129,N_11876);
nor U14479 (N_14479,N_11310,N_11898);
or U14480 (N_14480,N_11070,N_11115);
or U14481 (N_14481,N_11157,N_9548);
nand U14482 (N_14482,N_10602,N_9981);
nand U14483 (N_14483,N_11121,N_10567);
nand U14484 (N_14484,N_11414,N_11976);
nor U14485 (N_14485,N_11779,N_11950);
nor U14486 (N_14486,N_10310,N_10821);
or U14487 (N_14487,N_11294,N_9842);
nand U14488 (N_14488,N_10717,N_10042);
nand U14489 (N_14489,N_10444,N_9455);
nand U14490 (N_14490,N_10536,N_11753);
or U14491 (N_14491,N_10051,N_9497);
or U14492 (N_14492,N_9106,N_9526);
nand U14493 (N_14493,N_11247,N_9805);
and U14494 (N_14494,N_9513,N_11621);
nor U14495 (N_14495,N_11992,N_10026);
or U14496 (N_14496,N_9266,N_9746);
and U14497 (N_14497,N_11340,N_10197);
nand U14498 (N_14498,N_10871,N_11479);
nand U14499 (N_14499,N_10326,N_10947);
nand U14500 (N_14500,N_10526,N_11224);
nor U14501 (N_14501,N_11602,N_9133);
nand U14502 (N_14502,N_10891,N_9514);
nand U14503 (N_14503,N_11104,N_10426);
nor U14504 (N_14504,N_9299,N_9863);
or U14505 (N_14505,N_11396,N_11062);
and U14506 (N_14506,N_10146,N_9984);
or U14507 (N_14507,N_9529,N_9248);
nand U14508 (N_14508,N_9703,N_10777);
or U14509 (N_14509,N_11733,N_11002);
nand U14510 (N_14510,N_9175,N_10374);
nand U14511 (N_14511,N_11705,N_10566);
or U14512 (N_14512,N_9439,N_9286);
nand U14513 (N_14513,N_9097,N_11194);
nor U14514 (N_14514,N_10377,N_11137);
or U14515 (N_14515,N_9685,N_11828);
nor U14516 (N_14516,N_9574,N_11741);
or U14517 (N_14517,N_11625,N_11088);
nor U14518 (N_14518,N_10103,N_10058);
or U14519 (N_14519,N_10690,N_9356);
nor U14520 (N_14520,N_11074,N_11346);
and U14521 (N_14521,N_11794,N_11810);
nor U14522 (N_14522,N_10811,N_10143);
nor U14523 (N_14523,N_10751,N_10218);
and U14524 (N_14524,N_11319,N_11952);
and U14525 (N_14525,N_9761,N_10658);
or U14526 (N_14526,N_10400,N_9265);
or U14527 (N_14527,N_10417,N_10070);
xnor U14528 (N_14528,N_10686,N_9442);
nor U14529 (N_14529,N_10105,N_9512);
or U14530 (N_14530,N_10025,N_11168);
nand U14531 (N_14531,N_9898,N_10668);
and U14532 (N_14532,N_11811,N_9819);
or U14533 (N_14533,N_10639,N_11140);
and U14534 (N_14534,N_11772,N_9315);
and U14535 (N_14535,N_10733,N_11399);
nor U14536 (N_14536,N_11056,N_9360);
nand U14537 (N_14537,N_10557,N_11967);
nor U14538 (N_14538,N_10618,N_9994);
or U14539 (N_14539,N_10032,N_11042);
nor U14540 (N_14540,N_10397,N_9403);
and U14541 (N_14541,N_9263,N_10941);
nand U14542 (N_14542,N_11085,N_10899);
nor U14543 (N_14543,N_9315,N_10861);
or U14544 (N_14544,N_11498,N_9445);
or U14545 (N_14545,N_11443,N_9699);
nand U14546 (N_14546,N_9856,N_9157);
nor U14547 (N_14547,N_11140,N_10315);
and U14548 (N_14548,N_9146,N_11987);
nor U14549 (N_14549,N_11199,N_10938);
nand U14550 (N_14550,N_11368,N_9393);
or U14551 (N_14551,N_9723,N_11980);
nor U14552 (N_14552,N_11218,N_10667);
nor U14553 (N_14553,N_10576,N_11435);
nand U14554 (N_14554,N_10038,N_10768);
or U14555 (N_14555,N_9379,N_11294);
nand U14556 (N_14556,N_10117,N_11200);
and U14557 (N_14557,N_9515,N_11749);
nor U14558 (N_14558,N_9639,N_11656);
nand U14559 (N_14559,N_9610,N_11858);
and U14560 (N_14560,N_10782,N_9684);
and U14561 (N_14561,N_11321,N_9641);
and U14562 (N_14562,N_11325,N_10517);
nor U14563 (N_14563,N_10564,N_10507);
or U14564 (N_14564,N_11476,N_10022);
nand U14565 (N_14565,N_10905,N_9293);
xor U14566 (N_14566,N_9585,N_9682);
nor U14567 (N_14567,N_9349,N_11901);
and U14568 (N_14568,N_9870,N_11159);
and U14569 (N_14569,N_10659,N_10231);
or U14570 (N_14570,N_9735,N_11516);
nand U14571 (N_14571,N_11497,N_9835);
nor U14572 (N_14572,N_9529,N_11380);
nand U14573 (N_14573,N_9324,N_10881);
or U14574 (N_14574,N_10649,N_10994);
nor U14575 (N_14575,N_9975,N_10599);
or U14576 (N_14576,N_10284,N_10756);
and U14577 (N_14577,N_9955,N_9554);
or U14578 (N_14578,N_11206,N_9964);
nor U14579 (N_14579,N_9930,N_10245);
nor U14580 (N_14580,N_11954,N_11337);
and U14581 (N_14581,N_10769,N_11265);
nor U14582 (N_14582,N_11097,N_10819);
nand U14583 (N_14583,N_9637,N_10747);
and U14584 (N_14584,N_11717,N_9401);
nor U14585 (N_14585,N_11656,N_9080);
nor U14586 (N_14586,N_10143,N_11352);
and U14587 (N_14587,N_9494,N_11818);
and U14588 (N_14588,N_11960,N_9673);
or U14589 (N_14589,N_11516,N_10587);
and U14590 (N_14590,N_11779,N_9221);
and U14591 (N_14591,N_10691,N_10331);
or U14592 (N_14592,N_10005,N_10293);
nand U14593 (N_14593,N_11706,N_10757);
or U14594 (N_14594,N_9071,N_11197);
nand U14595 (N_14595,N_11556,N_9623);
and U14596 (N_14596,N_9609,N_9850);
nand U14597 (N_14597,N_11659,N_9069);
or U14598 (N_14598,N_11037,N_10643);
and U14599 (N_14599,N_9368,N_10810);
xnor U14600 (N_14600,N_11953,N_10892);
or U14601 (N_14601,N_9005,N_11988);
or U14602 (N_14602,N_9127,N_10861);
and U14603 (N_14603,N_11315,N_9167);
or U14604 (N_14604,N_10803,N_11482);
nand U14605 (N_14605,N_10459,N_9508);
nor U14606 (N_14606,N_10719,N_9914);
or U14607 (N_14607,N_10557,N_10617);
nor U14608 (N_14608,N_9917,N_10502);
or U14609 (N_14609,N_11770,N_9416);
and U14610 (N_14610,N_10541,N_10100);
and U14611 (N_14611,N_11752,N_11995);
nor U14612 (N_14612,N_10647,N_11998);
nor U14613 (N_14613,N_9741,N_9232);
and U14614 (N_14614,N_9206,N_9328);
nor U14615 (N_14615,N_9868,N_10734);
and U14616 (N_14616,N_9182,N_10377);
nand U14617 (N_14617,N_10838,N_10627);
or U14618 (N_14618,N_11318,N_9365);
and U14619 (N_14619,N_9164,N_9823);
nor U14620 (N_14620,N_10513,N_9693);
and U14621 (N_14621,N_11496,N_10343);
nor U14622 (N_14622,N_9580,N_9405);
or U14623 (N_14623,N_11798,N_10211);
nor U14624 (N_14624,N_10571,N_11715);
nand U14625 (N_14625,N_11582,N_10772);
or U14626 (N_14626,N_10011,N_9703);
and U14627 (N_14627,N_9166,N_9479);
and U14628 (N_14628,N_11045,N_9195);
or U14629 (N_14629,N_11620,N_10344);
nor U14630 (N_14630,N_10250,N_11642);
nor U14631 (N_14631,N_9936,N_9876);
nor U14632 (N_14632,N_9949,N_11165);
and U14633 (N_14633,N_11594,N_10688);
nor U14634 (N_14634,N_11320,N_11088);
or U14635 (N_14635,N_10943,N_9699);
or U14636 (N_14636,N_10325,N_9522);
and U14637 (N_14637,N_11405,N_10578);
and U14638 (N_14638,N_10163,N_11828);
nor U14639 (N_14639,N_10084,N_11789);
and U14640 (N_14640,N_11199,N_10014);
or U14641 (N_14641,N_11601,N_10008);
xnor U14642 (N_14642,N_11958,N_11884);
and U14643 (N_14643,N_9414,N_9196);
and U14644 (N_14644,N_10386,N_10531);
nand U14645 (N_14645,N_11182,N_11291);
or U14646 (N_14646,N_10507,N_9293);
nor U14647 (N_14647,N_9105,N_10038);
and U14648 (N_14648,N_11421,N_11206);
nand U14649 (N_14649,N_10326,N_11174);
nand U14650 (N_14650,N_11593,N_10878);
and U14651 (N_14651,N_9712,N_10099);
or U14652 (N_14652,N_9955,N_10106);
and U14653 (N_14653,N_10412,N_11579);
or U14654 (N_14654,N_11492,N_10831);
and U14655 (N_14655,N_11853,N_9490);
and U14656 (N_14656,N_10026,N_9249);
nand U14657 (N_14657,N_10997,N_9970);
and U14658 (N_14658,N_10600,N_9217);
nand U14659 (N_14659,N_10376,N_10971);
nor U14660 (N_14660,N_10592,N_11987);
nor U14661 (N_14661,N_11713,N_9530);
or U14662 (N_14662,N_10272,N_9831);
nor U14663 (N_14663,N_10520,N_9032);
nand U14664 (N_14664,N_10551,N_11274);
nand U14665 (N_14665,N_10390,N_11171);
nand U14666 (N_14666,N_11480,N_10105);
or U14667 (N_14667,N_9809,N_10897);
or U14668 (N_14668,N_11959,N_11221);
nand U14669 (N_14669,N_11701,N_11175);
and U14670 (N_14670,N_10523,N_11410);
and U14671 (N_14671,N_9839,N_9663);
or U14672 (N_14672,N_10246,N_11732);
nor U14673 (N_14673,N_10290,N_9143);
nor U14674 (N_14674,N_9440,N_9876);
nor U14675 (N_14675,N_11044,N_11599);
or U14676 (N_14676,N_10242,N_9184);
and U14677 (N_14677,N_10928,N_9054);
and U14678 (N_14678,N_9449,N_11686);
and U14679 (N_14679,N_11755,N_10423);
nor U14680 (N_14680,N_11472,N_11833);
nor U14681 (N_14681,N_11917,N_10443);
or U14682 (N_14682,N_9333,N_11649);
and U14683 (N_14683,N_11649,N_9289);
nand U14684 (N_14684,N_10884,N_10747);
or U14685 (N_14685,N_10421,N_11511);
nand U14686 (N_14686,N_9986,N_9247);
or U14687 (N_14687,N_9917,N_10815);
and U14688 (N_14688,N_9257,N_10624);
nor U14689 (N_14689,N_10064,N_9177);
or U14690 (N_14690,N_10451,N_11820);
or U14691 (N_14691,N_9622,N_10344);
and U14692 (N_14692,N_11540,N_9502);
nor U14693 (N_14693,N_9260,N_9350);
or U14694 (N_14694,N_10273,N_11767);
nor U14695 (N_14695,N_9556,N_11037);
and U14696 (N_14696,N_9653,N_9100);
nand U14697 (N_14697,N_10203,N_11801);
or U14698 (N_14698,N_10340,N_11834);
or U14699 (N_14699,N_11378,N_11623);
nand U14700 (N_14700,N_11451,N_9223);
and U14701 (N_14701,N_10981,N_10086);
or U14702 (N_14702,N_11324,N_10609);
and U14703 (N_14703,N_11447,N_11590);
nand U14704 (N_14704,N_11800,N_10847);
nor U14705 (N_14705,N_10832,N_11512);
nand U14706 (N_14706,N_10946,N_11039);
and U14707 (N_14707,N_10563,N_9747);
nor U14708 (N_14708,N_9116,N_10415);
nor U14709 (N_14709,N_10396,N_11163);
nor U14710 (N_14710,N_10725,N_11900);
nor U14711 (N_14711,N_9195,N_10191);
or U14712 (N_14712,N_11392,N_10151);
nand U14713 (N_14713,N_10079,N_11660);
nand U14714 (N_14714,N_10132,N_11802);
nor U14715 (N_14715,N_10471,N_10558);
or U14716 (N_14716,N_9961,N_9291);
or U14717 (N_14717,N_9181,N_9119);
and U14718 (N_14718,N_11741,N_9279);
nor U14719 (N_14719,N_11718,N_9011);
nand U14720 (N_14720,N_10907,N_11810);
and U14721 (N_14721,N_9431,N_11009);
nand U14722 (N_14722,N_11150,N_9109);
nor U14723 (N_14723,N_10426,N_10637);
nor U14724 (N_14724,N_9854,N_9473);
or U14725 (N_14725,N_11153,N_11544);
nor U14726 (N_14726,N_10752,N_11989);
nor U14727 (N_14727,N_9168,N_9515);
and U14728 (N_14728,N_10764,N_9587);
nor U14729 (N_14729,N_9086,N_11218);
and U14730 (N_14730,N_11541,N_10074);
or U14731 (N_14731,N_9568,N_10749);
and U14732 (N_14732,N_9676,N_9085);
and U14733 (N_14733,N_10854,N_11655);
or U14734 (N_14734,N_10577,N_11544);
xnor U14735 (N_14735,N_9097,N_10024);
or U14736 (N_14736,N_10979,N_10708);
xnor U14737 (N_14737,N_11536,N_11339);
nor U14738 (N_14738,N_10370,N_10302);
nand U14739 (N_14739,N_11837,N_11766);
nand U14740 (N_14740,N_11477,N_11169);
and U14741 (N_14741,N_9428,N_11632);
or U14742 (N_14742,N_9092,N_9260);
and U14743 (N_14743,N_11306,N_10332);
nor U14744 (N_14744,N_10050,N_11770);
and U14745 (N_14745,N_10001,N_11790);
or U14746 (N_14746,N_11925,N_10183);
or U14747 (N_14747,N_9660,N_11668);
and U14748 (N_14748,N_10399,N_10238);
nor U14749 (N_14749,N_10141,N_11114);
or U14750 (N_14750,N_11500,N_9679);
and U14751 (N_14751,N_10241,N_9502);
or U14752 (N_14752,N_9692,N_10205);
or U14753 (N_14753,N_9422,N_10867);
or U14754 (N_14754,N_9833,N_11780);
nor U14755 (N_14755,N_10384,N_9409);
nor U14756 (N_14756,N_9446,N_11037);
nand U14757 (N_14757,N_9288,N_10093);
nor U14758 (N_14758,N_11088,N_10474);
and U14759 (N_14759,N_11380,N_9552);
or U14760 (N_14760,N_10189,N_9090);
nor U14761 (N_14761,N_11382,N_10604);
or U14762 (N_14762,N_11328,N_9242);
nor U14763 (N_14763,N_11513,N_9014);
and U14764 (N_14764,N_9355,N_11299);
and U14765 (N_14765,N_11990,N_11304);
nor U14766 (N_14766,N_11710,N_10376);
nand U14767 (N_14767,N_9784,N_9829);
and U14768 (N_14768,N_9043,N_9292);
and U14769 (N_14769,N_11486,N_9314);
or U14770 (N_14770,N_10789,N_11682);
nor U14771 (N_14771,N_11250,N_9861);
nand U14772 (N_14772,N_11770,N_10098);
nor U14773 (N_14773,N_10698,N_9019);
and U14774 (N_14774,N_11694,N_9094);
nand U14775 (N_14775,N_11002,N_10740);
nor U14776 (N_14776,N_11516,N_9338);
nor U14777 (N_14777,N_11699,N_10957);
or U14778 (N_14778,N_11316,N_10710);
nor U14779 (N_14779,N_10862,N_11495);
nor U14780 (N_14780,N_9175,N_10142);
nor U14781 (N_14781,N_11577,N_9739);
nand U14782 (N_14782,N_9435,N_9129);
nand U14783 (N_14783,N_9392,N_9048);
and U14784 (N_14784,N_11525,N_11586);
nor U14785 (N_14785,N_10732,N_11194);
and U14786 (N_14786,N_10997,N_11678);
nand U14787 (N_14787,N_10793,N_9994);
nor U14788 (N_14788,N_11803,N_10458);
nor U14789 (N_14789,N_9309,N_9570);
and U14790 (N_14790,N_11148,N_10723);
nor U14791 (N_14791,N_11780,N_9640);
or U14792 (N_14792,N_10179,N_11588);
or U14793 (N_14793,N_11661,N_10224);
nor U14794 (N_14794,N_9497,N_10059);
or U14795 (N_14795,N_11858,N_10312);
and U14796 (N_14796,N_11164,N_11982);
and U14797 (N_14797,N_9517,N_11152);
nor U14798 (N_14798,N_10562,N_11010);
and U14799 (N_14799,N_9424,N_10434);
nand U14800 (N_14800,N_11325,N_11351);
nor U14801 (N_14801,N_11387,N_9201);
nand U14802 (N_14802,N_10786,N_10669);
and U14803 (N_14803,N_11690,N_9112);
nand U14804 (N_14804,N_10329,N_9337);
or U14805 (N_14805,N_11554,N_11738);
nand U14806 (N_14806,N_9905,N_10544);
and U14807 (N_14807,N_10337,N_10134);
or U14808 (N_14808,N_11076,N_9603);
and U14809 (N_14809,N_11798,N_11088);
nand U14810 (N_14810,N_11862,N_10511);
and U14811 (N_14811,N_10055,N_10971);
or U14812 (N_14812,N_9782,N_11706);
nand U14813 (N_14813,N_10816,N_11986);
nor U14814 (N_14814,N_11868,N_9420);
nor U14815 (N_14815,N_10344,N_10793);
or U14816 (N_14816,N_11229,N_9375);
nor U14817 (N_14817,N_11660,N_11457);
nor U14818 (N_14818,N_9448,N_10125);
or U14819 (N_14819,N_9841,N_9281);
and U14820 (N_14820,N_9089,N_10741);
and U14821 (N_14821,N_11806,N_11318);
or U14822 (N_14822,N_9302,N_10037);
nand U14823 (N_14823,N_10964,N_10552);
nor U14824 (N_14824,N_11005,N_11967);
or U14825 (N_14825,N_11485,N_11993);
nor U14826 (N_14826,N_10675,N_10544);
nand U14827 (N_14827,N_11567,N_10886);
or U14828 (N_14828,N_11771,N_9643);
nor U14829 (N_14829,N_11043,N_10447);
and U14830 (N_14830,N_9822,N_11943);
or U14831 (N_14831,N_9091,N_9727);
nand U14832 (N_14832,N_10361,N_9508);
or U14833 (N_14833,N_10128,N_9264);
and U14834 (N_14834,N_10917,N_9587);
nand U14835 (N_14835,N_10966,N_9010);
or U14836 (N_14836,N_11216,N_9328);
or U14837 (N_14837,N_11324,N_10975);
or U14838 (N_14838,N_11129,N_11937);
nor U14839 (N_14839,N_11290,N_10171);
nor U14840 (N_14840,N_11422,N_10244);
nor U14841 (N_14841,N_10309,N_9140);
nor U14842 (N_14842,N_11579,N_10746);
nor U14843 (N_14843,N_9350,N_11717);
nor U14844 (N_14844,N_10906,N_11718);
nand U14845 (N_14845,N_11446,N_10633);
or U14846 (N_14846,N_11933,N_9965);
nor U14847 (N_14847,N_10538,N_11041);
and U14848 (N_14848,N_9014,N_11329);
nand U14849 (N_14849,N_11787,N_10119);
or U14850 (N_14850,N_10434,N_11350);
and U14851 (N_14851,N_10366,N_11003);
or U14852 (N_14852,N_10798,N_9038);
nor U14853 (N_14853,N_10053,N_11256);
or U14854 (N_14854,N_11968,N_11031);
and U14855 (N_14855,N_10748,N_10336);
nand U14856 (N_14856,N_10531,N_11085);
or U14857 (N_14857,N_9105,N_9161);
nor U14858 (N_14858,N_10928,N_10813);
xor U14859 (N_14859,N_9927,N_10790);
and U14860 (N_14860,N_9887,N_9903);
nand U14861 (N_14861,N_10193,N_11693);
nand U14862 (N_14862,N_11705,N_9090);
nor U14863 (N_14863,N_9693,N_10877);
nor U14864 (N_14864,N_11313,N_9576);
nand U14865 (N_14865,N_11555,N_11460);
or U14866 (N_14866,N_9157,N_10246);
nand U14867 (N_14867,N_10216,N_9564);
or U14868 (N_14868,N_10603,N_11110);
nor U14869 (N_14869,N_9221,N_9714);
or U14870 (N_14870,N_9947,N_9354);
or U14871 (N_14871,N_11938,N_9799);
nand U14872 (N_14872,N_10168,N_10775);
or U14873 (N_14873,N_9559,N_11871);
nand U14874 (N_14874,N_10008,N_11856);
nor U14875 (N_14875,N_11187,N_10629);
or U14876 (N_14876,N_9488,N_9112);
or U14877 (N_14877,N_10931,N_9569);
nor U14878 (N_14878,N_11249,N_10916);
nand U14879 (N_14879,N_10632,N_11620);
or U14880 (N_14880,N_10296,N_10067);
and U14881 (N_14881,N_10421,N_9265);
xor U14882 (N_14882,N_10476,N_11858);
nand U14883 (N_14883,N_9339,N_11898);
nand U14884 (N_14884,N_11713,N_11332);
and U14885 (N_14885,N_10866,N_10648);
nand U14886 (N_14886,N_11063,N_11460);
nand U14887 (N_14887,N_9150,N_10001);
nand U14888 (N_14888,N_11901,N_10500);
nor U14889 (N_14889,N_9864,N_9805);
nor U14890 (N_14890,N_9488,N_10665);
xor U14891 (N_14891,N_10689,N_9477);
or U14892 (N_14892,N_11234,N_10137);
and U14893 (N_14893,N_9682,N_11425);
nor U14894 (N_14894,N_10056,N_9643);
nor U14895 (N_14895,N_10862,N_9938);
nor U14896 (N_14896,N_9266,N_11848);
and U14897 (N_14897,N_11046,N_9194);
nand U14898 (N_14898,N_10936,N_11452);
nor U14899 (N_14899,N_11134,N_11686);
nand U14900 (N_14900,N_9071,N_11006);
or U14901 (N_14901,N_11537,N_10156);
nand U14902 (N_14902,N_10395,N_11300);
nor U14903 (N_14903,N_10276,N_11368);
nor U14904 (N_14904,N_9307,N_11573);
and U14905 (N_14905,N_9994,N_10149);
nand U14906 (N_14906,N_10578,N_9939);
or U14907 (N_14907,N_10305,N_9327);
and U14908 (N_14908,N_10837,N_9625);
nor U14909 (N_14909,N_9538,N_9318);
or U14910 (N_14910,N_9710,N_9139);
or U14911 (N_14911,N_10668,N_9635);
and U14912 (N_14912,N_9903,N_10925);
or U14913 (N_14913,N_10311,N_9431);
and U14914 (N_14914,N_9434,N_11470);
nor U14915 (N_14915,N_9669,N_11756);
and U14916 (N_14916,N_11206,N_11481);
and U14917 (N_14917,N_10815,N_10599);
nor U14918 (N_14918,N_10135,N_10219);
and U14919 (N_14919,N_10052,N_11445);
nand U14920 (N_14920,N_9180,N_10507);
nor U14921 (N_14921,N_10628,N_10178);
nor U14922 (N_14922,N_11118,N_10100);
nand U14923 (N_14923,N_9870,N_9531);
nor U14924 (N_14924,N_10840,N_11489);
or U14925 (N_14925,N_9304,N_10612);
nand U14926 (N_14926,N_9013,N_10285);
nand U14927 (N_14927,N_10483,N_10228);
nor U14928 (N_14928,N_9079,N_11110);
nand U14929 (N_14929,N_10239,N_11221);
nand U14930 (N_14930,N_11314,N_9076);
nand U14931 (N_14931,N_11046,N_10034);
nand U14932 (N_14932,N_10321,N_9667);
nor U14933 (N_14933,N_9202,N_10094);
nand U14934 (N_14934,N_9931,N_9895);
or U14935 (N_14935,N_11000,N_10340);
nand U14936 (N_14936,N_10851,N_9159);
nor U14937 (N_14937,N_10677,N_10856);
or U14938 (N_14938,N_11149,N_9127);
nor U14939 (N_14939,N_11860,N_11469);
and U14940 (N_14940,N_11780,N_9045);
and U14941 (N_14941,N_11602,N_11888);
nor U14942 (N_14942,N_11661,N_9682);
nor U14943 (N_14943,N_10429,N_11069);
and U14944 (N_14944,N_10117,N_10904);
or U14945 (N_14945,N_11974,N_11273);
nand U14946 (N_14946,N_11597,N_9317);
nand U14947 (N_14947,N_9101,N_10545);
nand U14948 (N_14948,N_9676,N_9189);
nor U14949 (N_14949,N_10089,N_11181);
or U14950 (N_14950,N_10347,N_9942);
nor U14951 (N_14951,N_10893,N_10301);
nor U14952 (N_14952,N_9574,N_10246);
or U14953 (N_14953,N_11076,N_10114);
and U14954 (N_14954,N_9314,N_10763);
nor U14955 (N_14955,N_11261,N_9656);
and U14956 (N_14956,N_9519,N_11189);
and U14957 (N_14957,N_9181,N_10406);
nand U14958 (N_14958,N_10862,N_10841);
and U14959 (N_14959,N_11343,N_10580);
nor U14960 (N_14960,N_11944,N_10532);
nor U14961 (N_14961,N_11930,N_10483);
and U14962 (N_14962,N_10595,N_11685);
nor U14963 (N_14963,N_9585,N_9855);
nand U14964 (N_14964,N_9899,N_11705);
or U14965 (N_14965,N_9548,N_9719);
nand U14966 (N_14966,N_9064,N_10838);
nand U14967 (N_14967,N_11436,N_10452);
nand U14968 (N_14968,N_10872,N_9930);
and U14969 (N_14969,N_11535,N_9921);
nor U14970 (N_14970,N_9876,N_10643);
or U14971 (N_14971,N_10615,N_9290);
and U14972 (N_14972,N_11982,N_10089);
and U14973 (N_14973,N_9694,N_10056);
and U14974 (N_14974,N_11988,N_10821);
nor U14975 (N_14975,N_10005,N_10306);
nor U14976 (N_14976,N_9332,N_10846);
or U14977 (N_14977,N_11090,N_11821);
or U14978 (N_14978,N_9415,N_9516);
nand U14979 (N_14979,N_10693,N_9585);
nor U14980 (N_14980,N_11519,N_10815);
nor U14981 (N_14981,N_9927,N_10990);
nor U14982 (N_14982,N_9014,N_9940);
and U14983 (N_14983,N_10436,N_9597);
or U14984 (N_14984,N_10920,N_10159);
nand U14985 (N_14985,N_11429,N_11007);
nor U14986 (N_14986,N_10059,N_10836);
nor U14987 (N_14987,N_11740,N_11363);
nor U14988 (N_14988,N_11853,N_11118);
nand U14989 (N_14989,N_11804,N_11377);
nand U14990 (N_14990,N_11660,N_10476);
nand U14991 (N_14991,N_9058,N_11234);
or U14992 (N_14992,N_10879,N_9086);
nand U14993 (N_14993,N_10024,N_10054);
nand U14994 (N_14994,N_10261,N_10882);
and U14995 (N_14995,N_10727,N_10406);
and U14996 (N_14996,N_11180,N_9392);
nand U14997 (N_14997,N_10893,N_11421);
and U14998 (N_14998,N_9899,N_10861);
nand U14999 (N_14999,N_10136,N_10018);
and UO_0 (O_0,N_14546,N_13440);
nand UO_1 (O_1,N_14126,N_12512);
nand UO_2 (O_2,N_12123,N_13920);
nor UO_3 (O_3,N_14912,N_12817);
nor UO_4 (O_4,N_14004,N_14099);
and UO_5 (O_5,N_13221,N_12815);
nor UO_6 (O_6,N_13529,N_14684);
or UO_7 (O_7,N_12059,N_12052);
nand UO_8 (O_8,N_12149,N_14272);
nor UO_9 (O_9,N_13864,N_12113);
or UO_10 (O_10,N_14111,N_14839);
nor UO_11 (O_11,N_14669,N_13714);
nor UO_12 (O_12,N_14398,N_14021);
and UO_13 (O_13,N_12619,N_14778);
and UO_14 (O_14,N_14532,N_13322);
and UO_15 (O_15,N_12582,N_12254);
or UO_16 (O_16,N_12450,N_13708);
or UO_17 (O_17,N_14377,N_14068);
nor UO_18 (O_18,N_12686,N_13715);
or UO_19 (O_19,N_12027,N_14062);
and UO_20 (O_20,N_14415,N_14446);
or UO_21 (O_21,N_12926,N_13147);
nor UO_22 (O_22,N_13995,N_13590);
nor UO_23 (O_23,N_12977,N_14540);
or UO_24 (O_24,N_13980,N_14615);
nand UO_25 (O_25,N_13117,N_12061);
and UO_26 (O_26,N_12289,N_12091);
nand UO_27 (O_27,N_14657,N_13088);
nor UO_28 (O_28,N_13061,N_12145);
nand UO_29 (O_29,N_13780,N_14789);
nor UO_30 (O_30,N_12367,N_12531);
nand UO_31 (O_31,N_12335,N_12894);
nor UO_32 (O_32,N_12180,N_13261);
and UO_33 (O_33,N_12471,N_12981);
or UO_34 (O_34,N_14599,N_14944);
nor UO_35 (O_35,N_13155,N_14592);
and UO_36 (O_36,N_13439,N_13934);
nor UO_37 (O_37,N_13614,N_12403);
or UO_38 (O_38,N_13139,N_14334);
nand UO_39 (O_39,N_13523,N_13024);
or UO_40 (O_40,N_14772,N_14116);
nor UO_41 (O_41,N_12908,N_12915);
nand UO_42 (O_42,N_12417,N_13230);
and UO_43 (O_43,N_12567,N_12905);
or UO_44 (O_44,N_14551,N_13095);
nand UO_45 (O_45,N_14775,N_14664);
nand UO_46 (O_46,N_14416,N_13876);
or UO_47 (O_47,N_12914,N_12881);
xor UO_48 (O_48,N_13459,N_14182);
nand UO_49 (O_49,N_12116,N_14779);
and UO_50 (O_50,N_12553,N_13537);
nor UO_51 (O_51,N_14635,N_14786);
and UO_52 (O_52,N_12080,N_14145);
nor UO_53 (O_53,N_14567,N_13329);
nor UO_54 (O_54,N_13145,N_12115);
and UO_55 (O_55,N_14503,N_12545);
or UO_56 (O_56,N_12279,N_12215);
and UO_57 (O_57,N_13732,N_13807);
nor UO_58 (O_58,N_13822,N_13427);
nor UO_59 (O_59,N_14086,N_13492);
nand UO_60 (O_60,N_12954,N_13607);
or UO_61 (O_61,N_14696,N_13481);
or UO_62 (O_62,N_14400,N_14777);
and UO_63 (O_63,N_12301,N_12277);
nor UO_64 (O_64,N_13343,N_12259);
nand UO_65 (O_65,N_12987,N_13847);
and UO_66 (O_66,N_13670,N_13078);
and UO_67 (O_67,N_14131,N_12672);
or UO_68 (O_68,N_12462,N_14000);
nor UO_69 (O_69,N_13806,N_14541);
or UO_70 (O_70,N_14699,N_13267);
nor UO_71 (O_71,N_12399,N_13579);
nor UO_72 (O_72,N_12962,N_14835);
nor UO_73 (O_73,N_12224,N_12135);
or UO_74 (O_74,N_12305,N_13393);
and UO_75 (O_75,N_12771,N_14476);
and UO_76 (O_76,N_12509,N_14629);
nor UO_77 (O_77,N_14878,N_13905);
or UO_78 (O_78,N_13130,N_14217);
or UO_79 (O_79,N_14469,N_12387);
nand UO_80 (O_80,N_14405,N_13777);
or UO_81 (O_81,N_14199,N_14349);
nand UO_82 (O_82,N_12868,N_13841);
and UO_83 (O_83,N_12420,N_14729);
nor UO_84 (O_84,N_13981,N_12453);
nor UO_85 (O_85,N_13101,N_14440);
or UO_86 (O_86,N_13052,N_13422);
nor UO_87 (O_87,N_13639,N_13031);
nand UO_88 (O_88,N_12381,N_12089);
nor UO_89 (O_89,N_13128,N_13034);
or UO_90 (O_90,N_14456,N_14876);
nor UO_91 (O_91,N_14641,N_13414);
or UO_92 (O_92,N_14151,N_13576);
nor UO_93 (O_93,N_13925,N_12950);
nand UO_94 (O_94,N_13328,N_14992);
or UO_95 (O_95,N_13265,N_12683);
or UO_96 (O_96,N_13235,N_14155);
and UO_97 (O_97,N_14363,N_12064);
nor UO_98 (O_98,N_14686,N_13884);
nor UO_99 (O_99,N_12704,N_13007);
or UO_100 (O_100,N_13069,N_13136);
or UO_101 (O_101,N_14981,N_13470);
or UO_102 (O_102,N_14003,N_14052);
nand UO_103 (O_103,N_12718,N_13955);
nor UO_104 (O_104,N_12848,N_13929);
or UO_105 (O_105,N_12142,N_12269);
or UO_106 (O_106,N_12320,N_13794);
nand UO_107 (O_107,N_12092,N_13245);
and UO_108 (O_108,N_14542,N_14110);
or UO_109 (O_109,N_13317,N_12897);
nand UO_110 (O_110,N_12228,N_12895);
nand UO_111 (O_111,N_12657,N_13342);
nand UO_112 (O_112,N_14601,N_13240);
or UO_113 (O_113,N_13933,N_13747);
nand UO_114 (O_114,N_12552,N_13928);
and UO_115 (O_115,N_12724,N_13562);
or UO_116 (O_116,N_12068,N_13950);
and UO_117 (O_117,N_12504,N_12985);
nor UO_118 (O_118,N_13721,N_13669);
and UO_119 (O_119,N_12513,N_13829);
and UO_120 (O_120,N_13972,N_13844);
nor UO_121 (O_121,N_14931,N_12484);
or UO_122 (O_122,N_12921,N_13943);
or UO_123 (O_123,N_13295,N_14848);
and UO_124 (O_124,N_13802,N_12096);
and UO_125 (O_125,N_13045,N_14809);
and UO_126 (O_126,N_14119,N_13213);
and UO_127 (O_127,N_12974,N_12392);
xor UO_128 (O_128,N_12422,N_14130);
and UO_129 (O_129,N_12725,N_12163);
or UO_130 (O_130,N_14431,N_14773);
or UO_131 (O_131,N_13953,N_14932);
or UO_132 (O_132,N_12465,N_13179);
nand UO_133 (O_133,N_14974,N_14327);
and UO_134 (O_134,N_12882,N_14160);
or UO_135 (O_135,N_12585,N_14082);
nand UO_136 (O_136,N_14675,N_14575);
and UO_137 (O_137,N_13615,N_13472);
or UO_138 (O_138,N_12010,N_14127);
and UO_139 (O_139,N_14547,N_13381);
nand UO_140 (O_140,N_14331,N_14113);
and UO_141 (O_141,N_14568,N_12664);
or UO_142 (O_142,N_14638,N_12046);
nand UO_143 (O_143,N_13200,N_12258);
nor UO_144 (O_144,N_13426,N_12999);
or UO_145 (O_145,N_14488,N_14459);
or UO_146 (O_146,N_12548,N_13525);
nor UO_147 (O_147,N_13908,N_14027);
nor UO_148 (O_148,N_13572,N_13020);
nor UO_149 (O_149,N_13759,N_12282);
and UO_150 (O_150,N_14692,N_12410);
or UO_151 (O_151,N_14015,N_14801);
and UO_152 (O_152,N_12171,N_14994);
nand UO_153 (O_153,N_14755,N_12408);
and UO_154 (O_154,N_12888,N_12896);
nand UO_155 (O_155,N_12839,N_12671);
and UO_156 (O_156,N_13868,N_12376);
and UO_157 (O_157,N_14760,N_13554);
nor UO_158 (O_158,N_13025,N_13313);
and UO_159 (O_159,N_12373,N_13538);
nand UO_160 (O_160,N_14572,N_13109);
and UO_161 (O_161,N_14057,N_14128);
nor UO_162 (O_162,N_13216,N_14862);
nor UO_163 (O_163,N_14263,N_13199);
nand UO_164 (O_164,N_13452,N_14103);
nor UO_165 (O_165,N_13819,N_13156);
nand UO_166 (O_166,N_12869,N_13580);
xor UO_167 (O_167,N_14163,N_13917);
nor UO_168 (O_168,N_14593,N_13341);
or UO_169 (O_169,N_14079,N_14354);
or UO_170 (O_170,N_12304,N_14608);
or UO_171 (O_171,N_13438,N_13236);
and UO_172 (O_172,N_12872,N_14428);
or UO_173 (O_173,N_14129,N_14124);
nor UO_174 (O_174,N_13373,N_14562);
nand UO_175 (O_175,N_12007,N_12943);
and UO_176 (O_176,N_12294,N_14971);
nand UO_177 (O_177,N_14856,N_13993);
nor UO_178 (O_178,N_12721,N_14041);
nor UO_179 (O_179,N_13134,N_13997);
nand UO_180 (O_180,N_13894,N_12267);
nor UO_181 (O_181,N_12098,N_13648);
and UO_182 (O_182,N_14759,N_12040);
nand UO_183 (O_183,N_13845,N_12645);
and UO_184 (O_184,N_14208,N_13234);
and UO_185 (O_185,N_12673,N_12391);
or UO_186 (O_186,N_12577,N_13241);
and UO_187 (O_187,N_12332,N_12611);
nand UO_188 (O_188,N_14998,N_13163);
or UO_189 (O_189,N_14123,N_12492);
and UO_190 (O_190,N_14868,N_12878);
and UO_191 (O_191,N_14770,N_12668);
and UO_192 (O_192,N_12958,N_14838);
nand UO_193 (O_193,N_13203,N_12866);
nor UO_194 (O_194,N_14081,N_13107);
nand UO_195 (O_195,N_14241,N_14105);
nor UO_196 (O_196,N_13799,N_12523);
and UO_197 (O_197,N_12374,N_14624);
and UO_198 (O_198,N_13703,N_12571);
and UO_199 (O_199,N_14067,N_13561);
or UO_200 (O_200,N_13314,N_13897);
or UO_201 (O_201,N_14576,N_12598);
or UO_202 (O_202,N_13263,N_12011);
nand UO_203 (O_203,N_13931,N_13971);
nand UO_204 (O_204,N_13044,N_12530);
nor UO_205 (O_205,N_12246,N_12883);
nor UO_206 (O_206,N_13181,N_12951);
and UO_207 (O_207,N_13753,N_14274);
and UO_208 (O_208,N_14765,N_12240);
and UO_209 (O_209,N_13290,N_13645);
and UO_210 (O_210,N_14697,N_12325);
or UO_211 (O_211,N_13969,N_12913);
and UO_212 (O_212,N_14399,N_14788);
and UO_213 (O_213,N_13640,N_14803);
or UO_214 (O_214,N_13012,N_12341);
nor UO_215 (O_215,N_14997,N_14351);
nand UO_216 (O_216,N_13258,N_12775);
nand UO_217 (O_217,N_12185,N_14648);
nor UO_218 (O_218,N_13110,N_12931);
nor UO_219 (O_219,N_13658,N_12752);
nand UO_220 (O_220,N_13996,N_12786);
nand UO_221 (O_221,N_12653,N_14884);
or UO_222 (O_222,N_14022,N_12284);
nand UO_223 (O_223,N_13783,N_14678);
or UO_224 (O_224,N_12085,N_14613);
nor UO_225 (O_225,N_13371,N_13690);
or UO_226 (O_226,N_14513,N_13064);
nor UO_227 (O_227,N_14187,N_13578);
and UO_228 (O_228,N_13403,N_13999);
nor UO_229 (O_229,N_12095,N_14925);
nand UO_230 (O_230,N_14284,N_12753);
nor UO_231 (O_231,N_13900,N_13906);
nand UO_232 (O_232,N_13520,N_12211);
or UO_233 (O_233,N_14036,N_12906);
nor UO_234 (O_234,N_14625,N_12699);
or UO_235 (O_235,N_14580,N_13142);
and UO_236 (O_236,N_14520,N_13453);
or UO_237 (O_237,N_13158,N_14637);
nand UO_238 (O_238,N_14013,N_14652);
and UO_239 (O_239,N_14911,N_13549);
nor UO_240 (O_240,N_12864,N_12566);
nand UO_241 (O_241,N_13089,N_12329);
nor UO_242 (O_242,N_12589,N_12125);
nand UO_243 (O_243,N_12776,N_13530);
or UO_244 (O_244,N_14813,N_12172);
nand UO_245 (O_245,N_12922,N_12073);
or UO_246 (O_246,N_13559,N_14883);
or UO_247 (O_247,N_13622,N_12500);
nor UO_248 (O_248,N_14268,N_12911);
nor UO_249 (O_249,N_12559,N_13512);
nor UO_250 (O_250,N_12290,N_14336);
nor UO_251 (O_251,N_14502,N_12798);
or UO_252 (O_252,N_13375,N_13923);
or UO_253 (O_253,N_12162,N_14597);
or UO_254 (O_254,N_12646,N_12744);
nor UO_255 (O_255,N_14453,N_12519);
nand UO_256 (O_256,N_14619,N_12885);
and UO_257 (O_257,N_14261,N_12077);
nand UO_258 (O_258,N_13967,N_13456);
or UO_259 (O_259,N_12472,N_14162);
nand UO_260 (O_260,N_13506,N_12261);
or UO_261 (O_261,N_13081,N_12438);
nand UO_262 (O_262,N_12680,N_13701);
nand UO_263 (O_263,N_13698,N_14161);
and UO_264 (O_264,N_14106,N_13601);
nor UO_265 (O_265,N_14357,N_14942);
or UO_266 (O_266,N_12837,N_14618);
xor UO_267 (O_267,N_14722,N_13469);
nand UO_268 (O_268,N_13152,N_12930);
or UO_269 (O_269,N_12265,N_12386);
nor UO_270 (O_270,N_12106,N_14726);
and UO_271 (O_271,N_12139,N_13226);
nor UO_272 (O_272,N_13168,N_13075);
or UO_273 (O_273,N_12212,N_12936);
nand UO_274 (O_274,N_13968,N_13678);
and UO_275 (O_275,N_14632,N_12967);
nand UO_276 (O_276,N_13097,N_12644);
nand UO_277 (O_277,N_14903,N_13617);
nand UO_278 (O_278,N_12017,N_14253);
nor UO_279 (O_279,N_12038,N_12594);
nor UO_280 (O_280,N_12409,N_12133);
nor UO_281 (O_281,N_12419,N_14249);
nor UO_282 (O_282,N_12433,N_12856);
or UO_283 (O_283,N_14531,N_12416);
nand UO_284 (O_284,N_14982,N_12747);
nor UO_285 (O_285,N_12855,N_12124);
and UO_286 (O_286,N_12250,N_12623);
nand UO_287 (O_287,N_14812,N_14096);
nand UO_288 (O_288,N_14907,N_14634);
and UO_289 (O_289,N_14859,N_13539);
nand UO_290 (O_290,N_12576,N_14100);
nand UO_291 (O_291,N_13090,N_14698);
and UO_292 (O_292,N_12076,N_12933);
nand UO_293 (O_293,N_14824,N_12498);
xnor UO_294 (O_294,N_12187,N_13555);
nand UO_295 (O_295,N_13803,N_12807);
nand UO_296 (O_296,N_14558,N_13387);
or UO_297 (O_297,N_13789,N_14149);
and UO_298 (O_298,N_13165,N_12455);
nor UO_299 (O_299,N_13630,N_12873);
or UO_300 (O_300,N_13938,N_13415);
and UO_301 (O_301,N_14554,N_14227);
nor UO_302 (O_302,N_12270,N_12961);
nor UO_303 (O_303,N_14511,N_13146);
or UO_304 (O_304,N_14138,N_13668);
nand UO_305 (O_305,N_12437,N_14417);
nor UO_306 (O_306,N_14960,N_13948);
xor UO_307 (O_307,N_14864,N_13390);
nand UO_308 (O_308,N_13962,N_14730);
and UO_309 (O_309,N_12009,N_14250);
nor UO_310 (O_310,N_14175,N_14251);
nand UO_311 (O_311,N_14737,N_13065);
nand UO_312 (O_312,N_12018,N_14359);
nor UO_313 (O_313,N_13086,N_12494);
nand UO_314 (O_314,N_14781,N_14260);
or UO_315 (O_315,N_14462,N_14202);
and UO_316 (O_316,N_13551,N_13141);
nand UO_317 (O_317,N_12247,N_12797);
and UO_318 (O_318,N_13793,N_12750);
nor UO_319 (O_319,N_14389,N_13495);
nand UO_320 (O_320,N_13533,N_12924);
or UO_321 (O_321,N_13030,N_14654);
or UO_322 (O_322,N_12278,N_13010);
or UO_323 (O_323,N_13547,N_14934);
nand UO_324 (O_324,N_13503,N_12062);
or UO_325 (O_325,N_12637,N_12748);
nor UO_326 (O_326,N_13818,N_12917);
and UO_327 (O_327,N_12841,N_14526);
and UO_328 (O_328,N_14661,N_12996);
nand UO_329 (O_329,N_14201,N_12385);
nor UO_330 (O_330,N_12971,N_14660);
and UO_331 (O_331,N_12165,N_13305);
nor UO_332 (O_332,N_14205,N_13935);
nand UO_333 (O_333,N_12430,N_12119);
nor UO_334 (O_334,N_13911,N_14559);
and UO_335 (O_335,N_12079,N_14953);
or UO_336 (O_336,N_13292,N_13727);
nand UO_337 (O_337,N_14853,N_14278);
and UO_338 (O_338,N_13631,N_12317);
and UO_339 (O_339,N_12501,N_14134);
xor UO_340 (O_340,N_12635,N_12375);
or UO_341 (O_341,N_12111,N_12469);
nand UO_342 (O_342,N_12157,N_13488);
and UO_343 (O_343,N_13374,N_12238);
nand UO_344 (O_344,N_13942,N_14317);
and UO_345 (O_345,N_14054,N_14071);
nand UO_346 (O_346,N_13445,N_14655);
nor UO_347 (O_347,N_12783,N_14011);
nand UO_348 (O_348,N_13652,N_14627);
or UO_349 (O_349,N_14478,N_13356);
and UO_350 (O_350,N_12712,N_14053);
nor UO_351 (O_351,N_13792,N_12078);
or UO_352 (O_352,N_14505,N_13796);
nand UO_353 (O_353,N_13050,N_12833);
nor UO_354 (O_354,N_13604,N_12760);
or UO_355 (O_355,N_12461,N_13872);
nor UO_356 (O_356,N_14107,N_13382);
nor UO_357 (O_357,N_14688,N_12218);
and UO_358 (O_358,N_13327,N_12800);
nand UO_359 (O_359,N_13707,N_14936);
or UO_360 (O_360,N_14154,N_13309);
and UO_361 (O_361,N_12412,N_14297);
and UO_362 (O_362,N_13149,N_12937);
or UO_363 (O_363,N_14744,N_14140);
or UO_364 (O_364,N_12207,N_12540);
or UO_365 (O_365,N_14065,N_12655);
nand UO_366 (O_366,N_12031,N_14653);
nor UO_367 (O_367,N_12847,N_13204);
or UO_368 (O_368,N_12466,N_14690);
and UO_369 (O_369,N_12845,N_12630);
and UO_370 (O_370,N_12380,N_14266);
and UO_371 (O_371,N_13471,N_12260);
or UO_372 (O_372,N_12057,N_13702);
nor UO_373 (O_373,N_14470,N_13037);
and UO_374 (O_374,N_14097,N_12217);
nand UO_375 (O_375,N_14851,N_12182);
xor UO_376 (O_376,N_12107,N_12805);
or UO_377 (O_377,N_13157,N_13264);
or UO_378 (O_378,N_14303,N_13974);
nor UO_379 (O_379,N_13205,N_14311);
or UO_380 (O_380,N_13180,N_12255);
or UO_381 (O_381,N_12489,N_14525);
and UO_382 (O_382,N_14479,N_12121);
or UO_383 (O_383,N_13713,N_13366);
and UO_384 (O_384,N_13804,N_14247);
nand UO_385 (O_385,N_12322,N_12205);
nor UO_386 (O_386,N_14668,N_14296);
nand UO_387 (O_387,N_14704,N_14508);
and UO_388 (O_388,N_14957,N_12607);
nand UO_389 (O_389,N_13891,N_13865);
nand UO_390 (O_390,N_14939,N_12534);
nand UO_391 (O_391,N_12615,N_13451);
nand UO_392 (O_392,N_14800,N_13635);
nand UO_393 (O_393,N_14677,N_13323);
and UO_394 (O_394,N_14120,N_12909);
and UO_395 (O_395,N_12362,N_12081);
and UO_396 (O_396,N_12904,N_13407);
nand UO_397 (O_397,N_14849,N_12901);
nand UO_398 (O_398,N_12342,N_14092);
nor UO_399 (O_399,N_13666,N_14854);
or UO_400 (O_400,N_12648,N_13377);
and UO_401 (O_401,N_12138,N_13653);
or UO_402 (O_402,N_13540,N_12732);
and UO_403 (O_403,N_13123,N_12499);
and UO_404 (O_404,N_13102,N_13486);
nor UO_405 (O_405,N_12424,N_12717);
or UO_406 (O_406,N_13354,N_12075);
nand UO_407 (O_407,N_12525,N_12431);
nand UO_408 (O_408,N_14477,N_13368);
and UO_409 (O_409,N_12487,N_12407);
and UO_410 (O_410,N_13386,N_14611);
nand UO_411 (O_411,N_14017,N_13741);
nor UO_412 (O_412,N_13770,N_14472);
nand UO_413 (O_413,N_12352,N_14340);
or UO_414 (O_414,N_12330,N_13124);
nor UO_415 (O_415,N_13692,N_14796);
and UO_416 (O_416,N_14834,N_14132);
nand UO_417 (O_417,N_12094,N_14191);
nand UO_418 (O_418,N_12857,N_13224);
and UO_419 (O_419,N_12563,N_13397);
nor UO_420 (O_420,N_13823,N_14924);
nor UO_421 (O_421,N_13154,N_12168);
and UO_422 (O_422,N_13567,N_13705);
or UO_423 (O_423,N_12573,N_14607);
and UO_424 (O_424,N_12599,N_12204);
and UO_425 (O_425,N_12758,N_12702);
or UO_426 (O_426,N_14346,N_12264);
nor UO_427 (O_427,N_14913,N_14406);
nand UO_428 (O_428,N_12398,N_14527);
or UO_429 (O_429,N_12141,N_13005);
nand UO_430 (O_430,N_12378,N_14147);
nor UO_431 (O_431,N_14108,N_12879);
nand UO_432 (O_432,N_13877,N_13300);
nor UO_433 (O_433,N_13642,N_13306);
or UO_434 (O_434,N_12912,N_12656);
or UO_435 (O_435,N_13003,N_14783);
and UO_436 (O_436,N_13231,N_14970);
nand UO_437 (O_437,N_12001,N_14229);
nor UO_438 (O_438,N_12314,N_13207);
nand UO_439 (O_439,N_13766,N_13710);
nor UO_440 (O_440,N_12521,N_14948);
or UO_441 (O_441,N_13310,N_12876);
and UO_442 (O_442,N_14586,N_14837);
or UO_443 (O_443,N_12877,N_13115);
and UO_444 (O_444,N_14705,N_13083);
nand UO_445 (O_445,N_14656,N_12236);
nor UO_446 (O_446,N_12597,N_14798);
nor UO_447 (O_447,N_12813,N_13956);
and UO_448 (O_448,N_13514,N_12287);
nand UO_449 (O_449,N_14221,N_14679);
xnor UO_450 (O_450,N_13270,N_13720);
nand UO_451 (O_451,N_13276,N_14432);
nor UO_452 (O_452,N_12891,N_12790);
nand UO_453 (O_453,N_14609,N_13712);
and UO_454 (O_454,N_13001,N_14651);
or UO_455 (O_455,N_13667,N_14522);
nand UO_456 (O_456,N_12252,N_14626);
nor UO_457 (O_457,N_13965,N_13162);
and UO_458 (O_458,N_13885,N_12740);
or UO_459 (O_459,N_13913,N_12044);
nor UO_460 (O_460,N_13277,N_14345);
nor UO_461 (O_461,N_12442,N_13746);
or UO_462 (O_462,N_13662,N_13062);
or UO_463 (O_463,N_12271,N_14945);
or UO_464 (O_464,N_13238,N_14235);
or UO_465 (O_465,N_14538,N_12249);
or UO_466 (O_466,N_14200,N_14159);
nand UO_467 (O_467,N_13160,N_14647);
or UO_468 (O_468,N_13623,N_13961);
nand UO_469 (O_469,N_14891,N_12476);
nor UO_470 (O_470,N_13518,N_14226);
and UO_471 (O_471,N_14139,N_12041);
nor UO_472 (O_472,N_14921,N_12899);
xor UO_473 (O_473,N_12160,N_14169);
nor UO_474 (O_474,N_13596,N_14392);
nor UO_475 (O_475,N_14174,N_14136);
nor UO_476 (O_476,N_14860,N_13210);
nand UO_477 (O_477,N_12199,N_14330);
nor UO_478 (O_478,N_12678,N_12436);
or UO_479 (O_479,N_14791,N_13524);
nor UO_480 (O_480,N_14858,N_12852);
and UO_481 (O_481,N_14371,N_12628);
nor UO_482 (O_482,N_13326,N_12892);
nor UO_483 (O_483,N_12156,N_12929);
or UO_484 (O_484,N_12789,N_14673);
and UO_485 (O_485,N_14564,N_14257);
and UO_486 (O_486,N_14587,N_12475);
nand UO_487 (O_487,N_12243,N_14588);
and UO_488 (O_488,N_12023,N_12263);
or UO_489 (O_489,N_14375,N_13545);
and UO_490 (O_490,N_14448,N_13244);
nand UO_491 (O_491,N_12539,N_13289);
and UO_492 (O_492,N_12507,N_14797);
nand UO_493 (O_493,N_13603,N_14402);
or UO_494 (O_494,N_13125,N_13417);
or UO_495 (O_495,N_13412,N_14179);
and UO_496 (O_496,N_12975,N_14886);
nand UO_497 (O_497,N_13291,N_13535);
nand UO_498 (O_498,N_14749,N_12794);
nand UO_499 (O_499,N_12291,N_13063);
and UO_500 (O_500,N_13716,N_14270);
and UO_501 (O_501,N_12136,N_12510);
nand UO_502 (O_502,N_13634,N_14395);
nor UO_503 (O_503,N_12629,N_13552);
nor UO_504 (O_504,N_14189,N_13042);
and UO_505 (O_505,N_12793,N_14276);
or UO_506 (O_506,N_14324,N_13443);
nor UO_507 (O_507,N_14764,N_13032);
and UO_508 (O_508,N_14560,N_13744);
nor UO_509 (O_509,N_12354,N_13564);
nor UO_510 (O_510,N_14421,N_13599);
nand UO_511 (O_511,N_13223,N_14289);
or UO_512 (O_512,N_12257,N_12982);
and UO_513 (O_513,N_14636,N_12870);
nor UO_514 (O_514,N_13915,N_13939);
nand UO_515 (O_515,N_13480,N_14033);
or UO_516 (O_516,N_14940,N_12143);
or UO_517 (O_517,N_14602,N_14198);
nor UO_518 (O_518,N_13421,N_12175);
nor UO_519 (O_519,N_12522,N_12546);
or UO_520 (O_520,N_12483,N_13786);
nor UO_521 (O_521,N_14776,N_14935);
nand UO_522 (O_522,N_13378,N_13098);
and UO_523 (O_523,N_12272,N_13360);
and UO_524 (O_524,N_13970,N_14418);
and UO_525 (O_525,N_14080,N_14492);
nor UO_526 (O_526,N_12886,N_13093);
nand UO_527 (O_527,N_13167,N_13482);
and UO_528 (O_528,N_14927,N_14329);
and UO_529 (O_529,N_14785,N_14628);
or UO_530 (O_530,N_12543,N_14711);
or UO_531 (O_531,N_12323,N_12208);
nand UO_532 (O_532,N_12346,N_13857);
and UO_533 (O_533,N_14180,N_13056);
or UO_534 (O_534,N_12741,N_14964);
and UO_535 (O_535,N_14712,N_14847);
nor UO_536 (O_536,N_13748,N_12490);
and UO_537 (O_537,N_12679,N_12588);
and UO_538 (O_538,N_13779,N_13571);
and UO_539 (O_539,N_13233,N_14237);
xnor UO_540 (O_540,N_14058,N_12229);
nand UO_541 (O_541,N_12714,N_14279);
nor UO_542 (O_542,N_14183,N_14390);
nand UO_543 (O_543,N_14646,N_12302);
and UO_544 (O_544,N_13418,N_12659);
nand UO_545 (O_545,N_14826,N_14211);
nor UO_546 (O_546,N_12233,N_12348);
or UO_547 (O_547,N_12210,N_12293);
nor UO_548 (O_548,N_13504,N_12670);
and UO_549 (O_549,N_12043,N_14093);
nor UO_550 (O_550,N_14366,N_14309);
nand UO_551 (O_551,N_14283,N_13333);
nor UO_552 (O_552,N_13304,N_14423);
and UO_553 (O_553,N_12202,N_14984);
and UO_554 (O_554,N_13113,N_13269);
and UO_555 (O_555,N_14739,N_13080);
nor UO_556 (O_556,N_13194,N_14995);
or UO_557 (O_557,N_12343,N_12998);
nor UO_558 (O_558,N_12390,N_13404);
nand UO_559 (O_559,N_14828,N_12144);
and UO_560 (O_560,N_13553,N_14926);
nor UO_561 (O_561,N_14214,N_13271);
or UO_562 (O_562,N_12890,N_13764);
or UO_563 (O_563,N_12112,N_12150);
nand UO_564 (O_564,N_13455,N_14269);
nor UO_565 (O_565,N_13605,N_14143);
or UO_566 (O_566,N_12900,N_14874);
nand UO_567 (O_567,N_12826,N_14193);
xnor UO_568 (O_568,N_14090,N_12618);
or UO_569 (O_569,N_13719,N_12344);
nor UO_570 (O_570,N_14915,N_13542);
nand UO_571 (O_571,N_13135,N_12292);
nand UO_572 (O_572,N_12485,N_14954);
and UO_573 (O_573,N_13851,N_12429);
nor UO_574 (O_574,N_13602,N_13801);
and UO_575 (O_575,N_14682,N_12624);
and UO_576 (O_576,N_13916,N_13259);
and UO_577 (O_577,N_12966,N_14715);
or UO_578 (O_578,N_13380,N_13890);
nand UO_579 (O_579,N_14246,N_13337);
or UO_580 (O_580,N_13391,N_12197);
or UO_581 (O_581,N_13986,N_13644);
or UO_582 (O_582,N_14481,N_14869);
or UO_583 (O_583,N_14952,N_14005);
nand UO_584 (O_584,N_13958,N_14614);
and UO_585 (O_585,N_13026,N_14441);
nor UO_586 (O_586,N_13858,N_13650);
nand UO_587 (O_587,N_13307,N_13137);
nor UO_588 (O_588,N_13060,N_13202);
and UO_589 (O_589,N_13629,N_14890);
and UO_590 (O_590,N_12316,N_12058);
or UO_591 (O_591,N_14742,N_14548);
nand UO_592 (O_592,N_14146,N_14294);
nor UO_593 (O_593,N_12858,N_13619);
or UO_594 (O_594,N_14795,N_12331);
and UO_595 (O_595,N_14967,N_13071);
and UO_596 (O_596,N_12581,N_14732);
nand UO_597 (O_597,N_14996,N_13573);
or UO_598 (O_598,N_12336,N_14181);
xnor UO_599 (O_599,N_14333,N_12764);
or UO_600 (O_600,N_14494,N_13787);
and UO_601 (O_601,N_12012,N_14896);
nor UO_602 (O_602,N_14676,N_12251);
and UO_603 (O_603,N_12762,N_13575);
nand UO_604 (O_604,N_14823,N_12654);
nor UO_605 (O_605,N_12321,N_13039);
xnor UO_606 (O_606,N_13379,N_12434);
or UO_607 (O_607,N_12902,N_12675);
nor UO_608 (O_608,N_13724,N_14016);
or UO_609 (O_609,N_12942,N_13840);
nor UO_610 (O_610,N_14028,N_13177);
or UO_611 (O_611,N_14857,N_13187);
and UO_612 (O_612,N_14137,N_14443);
and UO_613 (O_613,N_13301,N_14745);
or UO_614 (O_614,N_14288,N_14521);
nand UO_615 (O_615,N_13718,N_12830);
nand UO_616 (O_616,N_12393,N_13355);
or UO_617 (O_617,N_12308,N_13489);
or UO_618 (O_618,N_12154,N_14735);
and UO_619 (O_619,N_14691,N_12127);
nand UO_620 (O_620,N_12583,N_14285);
and UO_621 (O_621,N_12164,N_13978);
nor UO_622 (O_622,N_14552,N_12757);
and UO_623 (O_623,N_13106,N_12622);
nand UO_624 (O_624,N_13870,N_12312);
xnor UO_625 (O_625,N_13830,N_14379);
nor UO_626 (O_626,N_13987,N_13336);
and UO_627 (O_627,N_12910,N_12486);
or UO_628 (O_628,N_14060,N_13035);
and UO_629 (O_629,N_13116,N_14401);
nor UO_630 (O_630,N_14064,N_12777);
nand UO_631 (O_631,N_12169,N_14056);
and UO_632 (O_632,N_13148,N_14396);
nand UO_633 (O_633,N_13508,N_12458);
nor UO_634 (O_634,N_14579,N_14708);
nor UO_635 (O_635,N_12578,N_13896);
nand UO_636 (O_636,N_12448,N_14464);
nor UO_637 (O_637,N_12158,N_14748);
nor UO_638 (O_638,N_13612,N_14885);
or UO_639 (O_639,N_12413,N_13433);
and UO_640 (O_640,N_14014,N_12722);
nor UO_641 (O_641,N_13346,N_14897);
nor UO_642 (O_642,N_13153,N_14372);
nand UO_643 (O_643,N_12025,N_13038);
nor UO_644 (O_644,N_12935,N_14165);
nand UO_645 (O_645,N_13460,N_13437);
or UO_646 (O_646,N_14498,N_14434);
nor UO_647 (O_647,N_13941,N_13677);
nor UO_648 (O_648,N_12749,N_12418);
and UO_649 (O_649,N_14212,N_12428);
or UO_650 (O_650,N_12549,N_14943);
or UO_651 (O_651,N_12884,N_12666);
nor UO_652 (O_652,N_13006,N_12460);
nand UO_653 (O_653,N_13468,N_13027);
nand UO_654 (O_654,N_13082,N_12503);
nand UO_655 (O_655,N_12518,N_14902);
nor UO_656 (O_656,N_13242,N_13952);
nand UO_657 (O_657,N_14037,N_14482);
xnor UO_658 (O_658,N_14724,N_14436);
nor UO_659 (O_659,N_12824,N_14102);
nand UO_660 (O_660,N_12533,N_13275);
nor UO_661 (O_661,N_13402,N_12328);
nor UO_662 (O_662,N_12652,N_13922);
nand UO_663 (O_663,N_14196,N_14667);
xor UO_664 (O_664,N_14225,N_13247);
and UO_665 (O_665,N_13511,N_13009);
nor UO_666 (O_666,N_12862,N_13268);
nor UO_667 (O_667,N_14176,N_13798);
or UO_668 (O_668,N_12440,N_13757);
and UO_669 (O_669,N_13926,N_14458);
nor UO_670 (O_670,N_12568,N_12692);
nor UO_671 (O_671,N_13362,N_12688);
or UO_672 (O_672,N_14710,N_14447);
and UO_673 (O_673,N_12880,N_14243);
xor UO_674 (O_674,N_12083,N_12372);
nand UO_675 (O_675,N_12767,N_13811);
and UO_676 (O_676,N_12808,N_14497);
and UO_677 (O_677,N_12432,N_13608);
nor UO_678 (O_678,N_13094,N_13531);
xnor UO_679 (O_679,N_12853,N_13394);
and UO_680 (O_680,N_12600,N_13143);
nand UO_681 (O_681,N_13253,N_13861);
nand UO_682 (O_682,N_13696,N_14843);
nand UO_683 (O_683,N_14524,N_14955);
or UO_684 (O_684,N_12021,N_13385);
nand UO_685 (O_685,N_14215,N_14008);
nor UO_686 (O_686,N_13334,N_12941);
nand UO_687 (O_687,N_14507,N_13127);
nor UO_688 (O_688,N_12071,N_14277);
and UO_689 (O_689,N_12634,N_12716);
nor UO_690 (O_690,N_12370,N_13454);
nor UO_691 (O_691,N_12361,N_12988);
or UO_692 (O_692,N_13945,N_14962);
or UO_693 (O_693,N_14846,N_12013);
and UO_694 (O_694,N_12221,N_13944);
nand UO_695 (O_695,N_13855,N_12700);
nand UO_696 (O_696,N_13367,N_13189);
and UO_697 (O_697,N_12351,N_14714);
and UO_698 (O_698,N_12050,N_12557);
nand UO_699 (O_699,N_14117,N_12445);
and UO_700 (O_700,N_14338,N_12687);
and UO_701 (O_701,N_14585,N_13767);
nor UO_702 (O_702,N_13076,N_13600);
nand UO_703 (O_703,N_14245,N_14035);
or UO_704 (O_704,N_14973,N_14254);
and UO_705 (O_705,N_14666,N_14665);
or UO_706 (O_706,N_12049,N_13467);
and UO_707 (O_707,N_14516,N_12726);
and UO_708 (O_708,N_13474,N_12035);
or UO_709 (O_709,N_12606,N_13348);
or UO_710 (O_710,N_14917,N_12402);
nand UO_711 (O_711,N_12658,N_14411);
nor UO_712 (O_712,N_12636,N_14049);
nor UO_713 (O_713,N_14424,N_14487);
nand UO_714 (O_714,N_12065,N_13016);
or UO_715 (O_715,N_12153,N_12339);
and UO_716 (O_716,N_12918,N_12167);
or UO_717 (O_717,N_14233,N_14403);
or UO_718 (O_718,N_13464,N_13641);
or UO_719 (O_719,N_13758,N_12691);
nor UO_720 (O_720,N_13998,N_12209);
nand UO_721 (O_721,N_12151,N_12861);
nor UO_722 (O_722,N_13023,N_14792);
or UO_723 (O_723,N_13633,N_13850);
and UO_724 (O_724,N_13015,N_14717);
nor UO_725 (O_725,N_14950,N_14353);
and UO_726 (O_726,N_14444,N_12591);
nor UO_727 (O_727,N_14118,N_13358);
and UO_728 (O_728,N_14206,N_12268);
or UO_729 (O_729,N_14658,N_12569);
or UO_730 (O_730,N_12161,N_12821);
or UO_731 (O_731,N_13598,N_12306);
nor UO_732 (O_732,N_12838,N_12253);
nor UO_733 (O_733,N_14388,N_14582);
and UO_734 (O_734,N_13797,N_13004);
nor UO_735 (O_735,N_12796,N_12364);
nor UO_736 (O_736,N_12174,N_12464);
nand UO_737 (O_737,N_12190,N_12016);
nor UO_738 (O_738,N_13190,N_14133);
nor UO_739 (O_739,N_14550,N_14304);
nor UO_740 (O_740,N_12196,N_14671);
and UO_741 (O_741,N_12538,N_12481);
nand UO_742 (O_742,N_12574,N_14975);
and UO_743 (O_743,N_14573,N_13957);
nand UO_744 (O_744,N_12621,N_12754);
nand UO_745 (O_745,N_13577,N_14050);
nand UO_746 (O_746,N_12235,N_13879);
nand UO_747 (O_747,N_12047,N_12613);
nor UO_748 (O_748,N_12769,N_12667);
and UO_749 (O_749,N_12008,N_13663);
nor UO_750 (O_750,N_12032,N_14055);
nor UO_751 (O_751,N_13331,N_12761);
and UO_752 (O_752,N_13425,N_12295);
and UO_753 (O_753,N_12608,N_14310);
nand UO_754 (O_754,N_12105,N_14293);
nand UO_755 (O_755,N_12927,N_14299);
or UO_756 (O_756,N_14763,N_13195);
nand UO_757 (O_757,N_12551,N_14020);
or UO_758 (O_758,N_13584,N_14980);
nor UO_759 (O_759,N_12356,N_12811);
nand UO_760 (O_760,N_12787,N_14898);
nand UO_761 (O_761,N_12441,N_14549);
nand UO_762 (O_762,N_13172,N_14281);
nand UO_763 (O_763,N_13100,N_12780);
and UO_764 (O_764,N_14620,N_14413);
or UO_765 (O_765,N_14387,N_12685);
nand UO_766 (O_766,N_13975,N_13827);
nand UO_767 (O_767,N_13297,N_12556);
and UO_768 (O_768,N_14539,N_13737);
and UO_769 (O_769,N_12447,N_14471);
and UO_770 (O_770,N_13126,N_13930);
and UO_771 (O_771,N_14889,N_14639);
or UO_772 (O_772,N_14817,N_13087);
or UO_773 (O_773,N_12439,N_14892);
nor UO_774 (O_774,N_13303,N_12003);
nand UO_775 (O_775,N_13735,N_14951);
and UO_776 (O_776,N_13751,N_14435);
nand UO_777 (O_777,N_13656,N_14881);
and UO_778 (O_778,N_13351,N_12480);
nand UO_779 (O_779,N_12358,N_14818);
and UO_780 (O_780,N_14298,N_12334);
or UO_781 (O_781,N_12694,N_12427);
nand UO_782 (O_782,N_13182,N_12479);
nand UO_783 (O_783,N_12756,N_13388);
nor UO_784 (O_784,N_12575,N_13501);
xor UO_785 (O_785,N_12707,N_13606);
or UO_786 (O_786,N_12920,N_13543);
nand UO_787 (O_787,N_14807,N_13339);
nor UO_788 (O_788,N_14426,N_12829);
nand UO_789 (O_789,N_13228,N_14976);
nor UO_790 (O_790,N_13686,N_14318);
and UO_791 (O_791,N_14204,N_14001);
nand UO_792 (O_792,N_14171,N_14946);
or UO_793 (O_793,N_13624,N_14073);
or UO_794 (O_794,N_13054,N_14873);
nor UO_795 (O_795,N_12147,N_13733);
and UO_796 (O_796,N_13161,N_14177);
or UO_797 (O_797,N_14098,N_13406);
or UO_798 (O_798,N_13260,N_14612);
nand UO_799 (O_799,N_13497,N_13740);
nand UO_800 (O_800,N_13046,N_14820);
nor UO_801 (O_801,N_12166,N_13196);
and UO_802 (O_802,N_13742,N_13790);
nor UO_803 (O_803,N_12082,N_13493);
nand UO_804 (O_804,N_12946,N_14007);
nand UO_805 (O_805,N_14213,N_13218);
nor UO_806 (O_806,N_12188,N_13266);
and UO_807 (O_807,N_12256,N_14043);
nand UO_808 (O_808,N_13914,N_13416);
nor UO_809 (O_809,N_14302,N_13131);
or UO_810 (O_810,N_12980,N_12728);
and UO_811 (O_811,N_13325,N_14929);
nand UO_812 (O_812,N_13462,N_12632);
and UO_813 (O_813,N_12763,N_13029);
and UO_814 (O_814,N_14344,N_12024);
nand UO_815 (O_815,N_12554,N_14600);
nand UO_816 (O_816,N_14530,N_13835);
or UO_817 (O_817,N_12176,N_14074);
nor UO_818 (O_818,N_14173,N_13949);
nand UO_819 (O_819,N_13112,N_13685);
nand UO_820 (O_820,N_12626,N_12338);
nor UO_821 (O_821,N_13515,N_12661);
and UO_822 (O_822,N_13984,N_14410);
nand UO_823 (O_823,N_12110,N_13647);
or UO_824 (O_824,N_12069,N_13183);
and UO_825 (O_825,N_13709,N_12126);
and UO_826 (O_826,N_12495,N_14156);
and UO_827 (O_827,N_14234,N_13866);
nor UO_828 (O_828,N_12701,N_12297);
nor UO_829 (O_829,N_13768,N_14218);
or UO_830 (O_830,N_14821,N_14244);
nor UO_831 (O_831,N_12311,N_14326);
and UO_832 (O_832,N_13487,N_14910);
or UO_833 (O_833,N_12170,N_14920);
or UO_834 (O_834,N_14042,N_14914);
or UO_835 (O_835,N_14461,N_12693);
or UO_836 (O_836,N_13215,N_13679);
or UO_837 (O_837,N_13655,N_12463);
nand UO_838 (O_838,N_14373,N_14622);
or UO_839 (O_839,N_13616,N_12345);
nand UO_840 (O_840,N_13294,N_14535);
nor UO_841 (O_841,N_14077,N_12191);
nor UO_842 (O_842,N_12042,N_14977);
nand UO_843 (O_843,N_12274,N_14219);
and UO_844 (O_844,N_12401,N_14966);
or UO_845 (O_845,N_14166,N_12642);
and UO_846 (O_846,N_12803,N_13420);
nor UO_847 (O_847,N_14325,N_12843);
and UO_848 (O_848,N_12515,N_14031);
or UO_849 (O_849,N_14561,N_14590);
or UO_850 (O_850,N_14850,N_13833);
nor UO_851 (O_851,N_14186,N_14808);
nand UO_852 (O_852,N_13220,N_13546);
or UO_853 (O_853,N_13700,N_12784);
nand UO_854 (O_854,N_13296,N_13805);
nor UO_855 (O_855,N_12313,N_14793);
or UO_856 (O_856,N_14815,N_14831);
and UO_857 (O_857,N_13816,N_14991);
nand UO_858 (O_858,N_14906,N_14830);
nand UO_859 (O_859,N_12713,N_13585);
nor UO_860 (O_860,N_12394,N_14574);
nor UO_861 (O_861,N_12604,N_12067);
or UO_862 (O_862,N_14841,N_12214);
nand UO_863 (O_863,N_12425,N_12184);
nor UO_864 (O_864,N_13138,N_14152);
and UO_865 (O_865,N_12834,N_12063);
nand UO_866 (O_866,N_14419,N_12863);
nor UO_867 (O_867,N_12772,N_14501);
nor UO_868 (O_868,N_12871,N_12120);
nand UO_869 (O_869,N_13383,N_14475);
or UO_870 (O_870,N_12867,N_14364);
nor UO_871 (O_871,N_14670,N_13907);
nand UO_872 (O_872,N_14335,N_12132);
and UO_873 (O_873,N_13762,N_14623);
or UO_874 (O_874,N_12703,N_13252);
nor UO_875 (O_875,N_14231,N_12949);
nor UO_876 (O_876,N_12972,N_14937);
nor UO_877 (O_877,N_14190,N_14583);
nor UO_878 (O_878,N_13222,N_12854);
or UO_879 (O_879,N_13413,N_13809);
nand UO_880 (O_880,N_12751,N_12755);
nor UO_881 (O_881,N_13649,N_14790);
and UO_882 (O_882,N_13442,N_13370);
and UO_883 (O_883,N_12266,N_13119);
or UO_884 (O_884,N_13824,N_13171);
nor UO_885 (O_885,N_14457,N_14369);
nor UO_886 (O_886,N_13919,N_13832);
nor UO_887 (O_887,N_13729,N_13283);
nor UO_888 (O_888,N_12651,N_13484);
nand UO_889 (O_889,N_13435,N_14365);
nor UO_890 (O_890,N_13785,N_12831);
and UO_891 (O_891,N_13910,N_14640);
or UO_892 (O_892,N_14880,N_14752);
xor UO_893 (O_893,N_12333,N_13396);
nor UO_894 (O_894,N_14566,N_12641);
nor UO_895 (O_895,N_14537,N_14061);
and UO_896 (O_896,N_12446,N_12201);
nor UO_897 (O_897,N_14286,N_12030);
nor UO_898 (O_898,N_14347,N_12819);
nand UO_899 (O_899,N_12874,N_14445);
or UO_900 (O_900,N_12477,N_14762);
and UO_901 (O_901,N_13284,N_12231);
nand UO_902 (O_902,N_14861,N_13664);
and UO_903 (O_903,N_13212,N_12932);
nor UO_904 (O_904,N_12706,N_13800);
nand UO_905 (O_905,N_14070,N_14633);
or UO_906 (O_906,N_14731,N_13496);
nor UO_907 (O_907,N_13772,N_12225);
or UO_908 (O_908,N_13457,N_12122);
nor UO_909 (O_909,N_14355,N_14046);
nor UO_910 (O_910,N_14414,N_14972);
and UO_911 (O_911,N_14723,N_12697);
nor UO_912 (O_912,N_13660,N_13320);
nor UO_913 (O_913,N_12388,N_14222);
xnor UO_914 (O_914,N_12404,N_12603);
nand UO_915 (O_915,N_13409,N_13017);
and UO_916 (O_916,N_14978,N_13408);
or UO_917 (O_917,N_12005,N_14700);
and UO_918 (O_918,N_12482,N_13722);
nor UO_919 (O_919,N_13754,N_12823);
nand UO_920 (O_920,N_13548,N_14184);
or UO_921 (O_921,N_14076,N_12779);
and UO_922 (O_922,N_12070,N_14969);
nor UO_923 (O_923,N_13775,N_13760);
or UO_924 (O_924,N_12226,N_14144);
and UO_925 (O_925,N_12101,N_13058);
nor UO_926 (O_926,N_14040,N_13681);
nand UO_927 (O_927,N_12088,N_14584);
and UO_928 (O_928,N_13675,N_14743);
or UO_929 (O_929,N_14545,N_13966);
and UO_930 (O_930,N_13319,N_12595);
or UO_931 (O_931,N_14832,N_13755);
nand UO_932 (O_932,N_13286,N_13140);
or UO_933 (O_933,N_12529,N_13924);
nand UO_934 (O_934,N_14733,N_13643);
and UO_935 (O_935,N_14543,N_12411);
nand UO_936 (O_936,N_12955,N_13033);
xor UO_937 (O_937,N_13051,N_14756);
nor UO_938 (O_938,N_14767,N_14157);
or UO_939 (O_939,N_14468,N_13256);
nor UO_940 (O_940,N_12689,N_13475);
and UO_941 (O_941,N_12849,N_13449);
nand UO_942 (O_942,N_12708,N_14774);
nand UO_943 (O_943,N_13049,N_12006);
and UO_944 (O_944,N_14404,N_13502);
nor UO_945 (O_945,N_12198,N_12109);
and UO_946 (O_946,N_13494,N_14827);
and UO_947 (O_947,N_12093,N_14986);
nand UO_948 (O_948,N_13281,N_13363);
or UO_949 (O_949,N_13085,N_13621);
or UO_950 (O_950,N_14569,N_12889);
and UO_951 (O_951,N_14556,N_13316);
and UO_952 (O_952,N_13178,N_14879);
or UO_953 (O_953,N_14577,N_12785);
nand UO_954 (O_954,N_13736,N_14514);
or UO_955 (O_955,N_13960,N_13516);
or UO_956 (O_956,N_14300,N_14305);
nor UO_957 (O_957,N_12371,N_14771);
nand UO_958 (O_958,N_12759,N_12239);
or UO_959 (O_959,N_14875,N_12818);
nand UO_960 (O_960,N_14384,N_13726);
nor UO_961 (O_961,N_13887,N_14989);
and UO_962 (O_962,N_12850,N_13927);
and UO_963 (O_963,N_12451,N_14923);
nand UO_964 (O_964,N_14063,N_13784);
and UO_965 (O_965,N_12952,N_14239);
and UO_966 (O_966,N_13174,N_14207);
and UO_967 (O_967,N_13092,N_13883);
nor UO_968 (O_968,N_13932,N_14442);
nand UO_969 (O_969,N_13769,N_14242);
or UO_970 (O_970,N_14158,N_13862);
nor UO_971 (O_971,N_13903,N_12986);
or UO_972 (O_972,N_12804,N_13878);
nor UO_973 (O_973,N_12053,N_13350);
and UO_974 (O_974,N_13990,N_14034);
or UO_975 (O_975,N_14570,N_13699);
and UO_976 (O_976,N_13432,N_13627);
nor UO_977 (O_977,N_13510,N_13659);
and UO_978 (O_978,N_14988,N_13781);
and UO_979 (O_979,N_13973,N_13447);
nand UO_980 (O_980,N_14987,N_13311);
or UO_981 (O_981,N_13353,N_14918);
and UO_982 (O_982,N_12097,N_13626);
and UO_983 (O_983,N_13372,N_14529);
and UO_984 (O_984,N_12488,N_14010);
or UO_985 (O_985,N_13401,N_14866);
nand UO_986 (O_986,N_12028,N_13246);
nand UO_987 (O_987,N_13689,N_12572);
nand UO_988 (O_988,N_12596,N_13361);
or UO_989 (O_989,N_14610,N_14167);
or UO_990 (O_990,N_14115,N_12505);
or UO_991 (O_991,N_14045,N_12791);
and UO_992 (O_992,N_13282,N_12532);
and UO_993 (O_993,N_13047,N_14192);
or UO_994 (O_994,N_12514,N_14203);
or UO_995 (O_995,N_13749,N_13569);
or UO_996 (O_996,N_14909,N_12310);
nand UO_997 (O_997,N_14378,N_12561);
or UO_998 (O_998,N_13651,N_12137);
and UO_999 (O_999,N_12426,N_14339);
and UO_1000 (O_1000,N_12283,N_13983);
nand UO_1001 (O_1001,N_13239,N_14709);
or UO_1002 (O_1002,N_13463,N_13834);
and UO_1003 (O_1003,N_13411,N_13490);
nand UO_1004 (O_1004,N_14716,N_14919);
and UO_1005 (O_1005,N_14500,N_12558);
and UO_1006 (O_1006,N_13262,N_12526);
or UO_1007 (O_1007,N_14019,N_14504);
nand UO_1008 (O_1008,N_13392,N_14397);
or UO_1009 (O_1009,N_13410,N_13232);
nor UO_1010 (O_1010,N_14947,N_14643);
or UO_1011 (O_1011,N_14510,N_12177);
and UO_1012 (O_1012,N_13485,N_14706);
or UO_1013 (O_1013,N_13022,N_13068);
and UO_1014 (O_1014,N_13133,N_13114);
and UO_1015 (O_1015,N_12774,N_12383);
nand UO_1016 (O_1016,N_14352,N_12363);
or UO_1017 (O_1017,N_14240,N_12565);
nand UO_1018 (O_1018,N_12978,N_13197);
and UO_1019 (O_1019,N_13873,N_13465);
nor UO_1020 (O_1020,N_14747,N_12234);
nor UO_1021 (O_1021,N_14591,N_12802);
or UO_1022 (O_1022,N_13077,N_12570);
nor UO_1023 (O_1023,N_14044,N_14301);
or UO_1024 (O_1024,N_13441,N_12467);
or UO_1025 (O_1025,N_13173,N_13237);
nor UO_1026 (O_1026,N_12809,N_12959);
and UO_1027 (O_1027,N_13184,N_13904);
or UO_1028 (O_1028,N_14452,N_13977);
nor UO_1029 (O_1029,N_14408,N_13066);
nor UO_1030 (O_1030,N_14141,N_12155);
or UO_1031 (O_1031,N_14707,N_13321);
xnor UO_1032 (O_1032,N_12973,N_12074);
and UO_1033 (O_1033,N_14422,N_12842);
and UO_1034 (O_1034,N_14322,N_12938);
and UO_1035 (O_1035,N_12192,N_12640);
and UO_1036 (O_1036,N_14727,N_12262);
and UO_1037 (O_1037,N_12421,N_12580);
and UO_1038 (O_1038,N_12195,N_14220);
and UO_1039 (O_1039,N_13901,N_14985);
and UO_1040 (O_1040,N_13763,N_13795);
and UO_1041 (O_1041,N_12669,N_13691);
or UO_1042 (O_1042,N_12537,N_12288);
nor UO_1043 (O_1043,N_14517,N_13521);
nor UO_1044 (O_1044,N_12562,N_13889);
or UO_1045 (O_1045,N_14455,N_14308);
nor UO_1046 (O_1046,N_12925,N_13302);
and UO_1047 (O_1047,N_12340,N_13191);
and UO_1048 (O_1048,N_13638,N_12382);
nor UO_1049 (O_1049,N_12099,N_13192);
nand UO_1050 (O_1050,N_14905,N_12609);
nand UO_1051 (O_1051,N_12090,N_13359);
nand UO_1052 (O_1052,N_13728,N_12733);
nor UO_1053 (O_1053,N_14663,N_13812);
xor UO_1054 (O_1054,N_12919,N_13863);
or UO_1055 (O_1055,N_12130,N_14750);
nand UO_1056 (O_1056,N_13478,N_14490);
or UO_1057 (O_1057,N_13837,N_13188);
nor UO_1058 (O_1058,N_14870,N_14433);
or UO_1059 (O_1059,N_14533,N_12840);
or UO_1060 (O_1060,N_12719,N_14386);
nor UO_1061 (O_1061,N_12893,N_12720);
nand UO_1062 (O_1062,N_14258,N_13164);
nand UO_1063 (O_1063,N_14644,N_13959);
or UO_1064 (O_1064,N_13665,N_13436);
nor UO_1065 (O_1065,N_14259,N_13505);
or UO_1066 (O_1066,N_12051,N_13208);
nand UO_1067 (O_1067,N_12612,N_14348);
nor UO_1068 (O_1068,N_13991,N_14210);
nor UO_1069 (O_1069,N_12152,N_13671);
and UO_1070 (O_1070,N_14893,N_13122);
and UO_1071 (O_1071,N_14307,N_12377);
nor UO_1072 (O_1072,N_13661,N_14804);
or UO_1073 (O_1073,N_14780,N_12535);
or UO_1074 (O_1074,N_14557,N_14840);
and UO_1075 (O_1075,N_12643,N_12633);
and UO_1076 (O_1076,N_13723,N_14095);
nor UO_1077 (O_1077,N_12550,N_13597);
xnor UO_1078 (O_1078,N_12508,N_12506);
nor UO_1079 (O_1079,N_14719,N_13684);
and UO_1080 (O_1080,N_12743,N_13843);
and UO_1081 (O_1081,N_14829,N_13821);
nand UO_1082 (O_1082,N_13859,N_13429);
nand UO_1083 (O_1083,N_12536,N_12690);
or UO_1084 (O_1084,N_12734,N_12347);
and UO_1085 (O_1085,N_13674,N_13588);
nand UO_1086 (O_1086,N_14787,N_14553);
nand UO_1087 (O_1087,N_14993,N_13018);
or UO_1088 (O_1088,N_12617,N_14672);
nand UO_1089 (O_1089,N_12592,N_13185);
and UO_1090 (O_1090,N_12990,N_12528);
nand UO_1091 (O_1091,N_12502,N_12953);
nand UO_1092 (O_1092,N_12812,N_13450);
nor UO_1093 (O_1093,N_14084,N_13299);
and UO_1094 (O_1094,N_13565,N_13013);
nor UO_1095 (O_1095,N_14275,N_14265);
or UO_1096 (O_1096,N_12281,N_13424);
nand UO_1097 (O_1097,N_12456,N_12186);
nor UO_1098 (O_1098,N_12060,N_12349);
nor UO_1099 (O_1099,N_14718,N_13695);
nor UO_1100 (O_1100,N_12898,N_12048);
nand UO_1101 (O_1101,N_13053,N_13111);
nor UO_1102 (O_1102,N_12614,N_14938);
or UO_1103 (O_1103,N_12836,N_14224);
and UO_1104 (O_1104,N_12660,N_13186);
or UO_1105 (O_1105,N_12627,N_14509);
nor UO_1106 (O_1106,N_14928,N_12736);
xor UO_1107 (O_1107,N_12544,N_13854);
nand UO_1108 (O_1108,N_12396,N_13592);
and UO_1109 (O_1109,N_12245,N_13198);
or UO_1110 (O_1110,N_12944,N_13750);
nand UO_1111 (O_1111,N_13057,N_13344);
or UO_1112 (O_1112,N_14882,N_14342);
nand UO_1113 (O_1113,N_13704,N_13620);
and UO_1114 (O_1114,N_13808,N_13509);
nand UO_1115 (O_1115,N_12605,N_13654);
nor UO_1116 (O_1116,N_12739,N_13637);
nand UO_1117 (O_1117,N_12232,N_12887);
and UO_1118 (O_1118,N_13581,N_14088);
nand UO_1119 (O_1119,N_12542,N_14754);
and UO_1120 (O_1120,N_14295,N_14571);
or UO_1121 (O_1121,N_14358,N_13214);
nor UO_1122 (O_1122,N_13219,N_12036);
nand UO_1123 (O_1123,N_14871,N_13055);
nor UO_1124 (O_1124,N_13682,N_14506);
nand UO_1125 (O_1125,N_12916,N_12103);
and UO_1126 (O_1126,N_12631,N_13398);
and UO_1127 (O_1127,N_12825,N_12319);
nand UO_1128 (O_1128,N_13849,N_14877);
or UO_1129 (O_1129,N_12275,N_13227);
nor UO_1130 (O_1130,N_14029,N_12369);
or UO_1131 (O_1131,N_14361,N_14589);
nand UO_1132 (O_1132,N_12730,N_13888);
nand UO_1133 (O_1133,N_12859,N_13711);
or UO_1134 (O_1134,N_14512,N_14519);
nand UO_1135 (O_1135,N_14292,N_12117);
or UO_1136 (O_1136,N_13251,N_14153);
nor UO_1137 (O_1137,N_13255,N_14930);
and UO_1138 (O_1138,N_13519,N_14681);
nand UO_1139 (O_1139,N_12992,N_14328);
nor UO_1140 (O_1140,N_14075,N_13528);
and UO_1141 (O_1141,N_14023,N_14842);
xnor UO_1142 (O_1142,N_14894,N_12002);
and UO_1143 (O_1143,N_14374,N_14232);
nor UO_1144 (O_1144,N_12746,N_14425);
and UO_1145 (O_1145,N_13479,N_14197);
nor UO_1146 (O_1146,N_12280,N_14280);
and UO_1147 (O_1147,N_14844,N_13814);
or UO_1148 (O_1148,N_14262,N_12474);
and UO_1149 (O_1149,N_14290,N_14746);
nor UO_1150 (O_1150,N_13340,N_13739);
nor UO_1151 (O_1151,N_14381,N_13761);
nand UO_1152 (O_1152,N_13586,N_12695);
and UO_1153 (O_1153,N_12768,N_14941);
nand UO_1154 (O_1154,N_12327,N_14594);
and UO_1155 (O_1155,N_14649,N_12034);
or UO_1156 (O_1156,N_14694,N_14486);
nand UO_1157 (O_1157,N_14761,N_14702);
nand UO_1158 (O_1158,N_14794,N_12365);
nor UO_1159 (O_1159,N_13312,N_13048);
or UO_1160 (O_1160,N_13937,N_14499);
and UO_1161 (O_1161,N_13491,N_12939);
nand UO_1162 (O_1162,N_14267,N_14230);
nor UO_1163 (O_1163,N_12989,N_13028);
and UO_1164 (O_1164,N_14236,N_14662);
and UO_1165 (O_1165,N_12851,N_12193);
and UO_1166 (O_1166,N_14544,N_14383);
nor UO_1167 (O_1167,N_14382,N_14429);
nor UO_1168 (O_1168,N_13458,N_14078);
nor UO_1169 (O_1169,N_12541,N_14104);
nor UO_1170 (O_1170,N_14799,N_12956);
or UO_1171 (O_1171,N_13982,N_12286);
or UO_1172 (O_1172,N_13170,N_14493);
nor UO_1173 (O_1173,N_13683,N_13352);
nand UO_1174 (O_1174,N_14563,N_13257);
nor UO_1175 (O_1175,N_12491,N_13132);
or UO_1176 (O_1176,N_14385,N_13752);
and UO_1177 (O_1177,N_13688,N_14757);
or UO_1178 (O_1178,N_13169,N_12178);
nor UO_1179 (O_1179,N_13206,N_12957);
nor UO_1180 (O_1180,N_14865,N_14687);
or UO_1181 (O_1181,N_12735,N_12248);
xor UO_1182 (O_1182,N_12242,N_12128);
and UO_1183 (O_1183,N_14047,N_14631);
and UO_1184 (O_1184,N_14438,N_13193);
nand UO_1185 (O_1185,N_14087,N_12835);
nor UO_1186 (O_1186,N_12397,N_14713);
or UO_1187 (O_1187,N_12773,N_12860);
or UO_1188 (O_1188,N_12315,N_13376);
or UO_1189 (O_1189,N_13384,N_14194);
xnor UO_1190 (O_1190,N_12584,N_12696);
and UO_1191 (O_1191,N_13499,N_13150);
nor UO_1192 (O_1192,N_14836,N_12729);
and UO_1193 (O_1193,N_14685,N_14802);
nor UO_1194 (O_1194,N_14172,N_12148);
nor UO_1195 (O_1195,N_14901,N_14738);
nor UO_1196 (O_1196,N_13108,N_13293);
nand UO_1197 (O_1197,N_14863,N_14474);
and UO_1198 (O_1198,N_13365,N_13298);
or UO_1199 (O_1199,N_12663,N_13249);
and UO_1200 (O_1200,N_13278,N_12799);
nand UO_1201 (O_1201,N_12298,N_12241);
nand UO_1202 (O_1202,N_13104,N_13332);
nor UO_1203 (O_1203,N_12194,N_12159);
or UO_1204 (O_1204,N_14463,N_13159);
nor UO_1205 (O_1205,N_12995,N_14728);
nand UO_1206 (O_1206,N_14581,N_13217);
or UO_1207 (O_1207,N_14248,N_12709);
and UO_1208 (O_1208,N_14072,N_14523);
nor UO_1209 (O_1209,N_14032,N_13364);
or UO_1210 (O_1210,N_13825,N_13568);
nand UO_1211 (O_1211,N_12414,N_12022);
nor UO_1212 (O_1212,N_13610,N_14908);
or UO_1213 (O_1213,N_12055,N_14195);
nor UO_1214 (O_1214,N_12200,N_14038);
nor UO_1215 (O_1215,N_12948,N_12206);
nor UO_1216 (O_1216,N_12649,N_13544);
or UO_1217 (O_1217,N_13773,N_13330);
and UO_1218 (O_1218,N_13285,N_13582);
nor UO_1219 (O_1219,N_12907,N_12355);
and UO_1220 (O_1220,N_12086,N_12555);
and UO_1221 (O_1221,N_13613,N_13036);
nand UO_1222 (O_1222,N_12677,N_13209);
nand UO_1223 (O_1223,N_13680,N_12244);
and UO_1224 (O_1224,N_13308,N_13706);
or UO_1225 (O_1225,N_12727,N_12979);
or UO_1226 (O_1226,N_12792,N_14282);
nor UO_1227 (O_1227,N_14185,N_12066);
and UO_1228 (O_1228,N_12827,N_13895);
nand UO_1229 (O_1229,N_14314,N_12602);
nand UO_1230 (O_1230,N_13166,N_12865);
and UO_1231 (O_1231,N_13144,N_14528);
nor UO_1232 (O_1232,N_12810,N_13853);
or UO_1233 (O_1233,N_12524,N_14112);
and UO_1234 (O_1234,N_13517,N_12087);
and UO_1235 (O_1235,N_13096,N_13676);
nand UO_1236 (O_1236,N_14164,N_13151);
and UO_1237 (O_1237,N_13079,N_14370);
nor UO_1238 (O_1238,N_12705,N_12681);
nor UO_1239 (O_1239,N_14701,N_13881);
nor UO_1240 (O_1240,N_13395,N_12104);
nand UO_1241 (O_1241,N_14693,N_14256);
nor UO_1242 (O_1242,N_12738,N_13287);
or UO_1243 (O_1243,N_12639,N_13583);
or UO_1244 (O_1244,N_12353,N_12875);
nand UO_1245 (O_1245,N_14895,N_13274);
or UO_1246 (O_1246,N_12056,N_14811);
nor UO_1247 (O_1247,N_13557,N_14819);
or UO_1248 (O_1248,N_13625,N_12216);
and UO_1249 (O_1249,N_12903,N_12940);
or UO_1250 (O_1250,N_14209,N_14150);
nor UO_1251 (O_1251,N_14595,N_12102);
and UO_1252 (O_1252,N_14825,N_13399);
nor UO_1253 (O_1253,N_13014,N_12219);
nand UO_1254 (O_1254,N_14450,N_13498);
nand UO_1255 (O_1255,N_13839,N_14025);
or UO_1256 (O_1256,N_13315,N_14473);
or UO_1257 (O_1257,N_14142,N_13473);
nor UO_1258 (O_1258,N_12527,N_12822);
nor UO_1259 (O_1259,N_14887,N_13423);
or UO_1260 (O_1260,N_12814,N_12665);
and UO_1261 (O_1261,N_13243,N_12698);
nor UO_1262 (O_1262,N_12309,N_13657);
or UO_1263 (O_1263,N_14223,N_13541);
and UO_1264 (O_1264,N_12766,N_13335);
or UO_1265 (O_1265,N_12276,N_14555);
and UO_1266 (O_1266,N_14703,N_13918);
or UO_1267 (O_1267,N_13587,N_14725);
and UO_1268 (O_1268,N_13476,N_13810);
nand UO_1269 (O_1269,N_14271,N_14467);
nand UO_1270 (O_1270,N_13070,N_13357);
nand UO_1271 (O_1271,N_14323,N_14051);
and UO_1272 (O_1272,N_13964,N_13534);
nor UO_1273 (O_1273,N_14736,N_13869);
nor UO_1274 (O_1274,N_14491,N_14009);
nand UO_1275 (O_1275,N_14451,N_12934);
or UO_1276 (O_1276,N_13225,N_12285);
nor UO_1277 (O_1277,N_13782,N_13947);
nor UO_1278 (O_1278,N_13570,N_12468);
nor UO_1279 (O_1279,N_13002,N_13738);
nor UO_1280 (O_1280,N_13563,N_14956);
and UO_1281 (O_1281,N_12173,N_14026);
nand UO_1282 (O_1282,N_12223,N_12493);
nor UO_1283 (O_1283,N_13011,N_14321);
and UO_1284 (O_1284,N_12620,N_14949);
nand UO_1285 (O_1285,N_13431,N_13522);
nand UO_1286 (O_1286,N_13400,N_13507);
nand UO_1287 (O_1287,N_13040,N_13813);
nor UO_1288 (O_1288,N_13778,N_13008);
nand UO_1289 (O_1289,N_14255,N_13526);
and UO_1290 (O_1290,N_12520,N_12443);
nor UO_1291 (O_1291,N_13902,N_14782);
and UO_1292 (O_1292,N_14753,N_12765);
nand UO_1293 (O_1293,N_13513,N_13084);
nor UO_1294 (O_1294,N_13734,N_13105);
nor UO_1295 (O_1295,N_12029,N_14319);
and UO_1296 (O_1296,N_14059,N_12179);
nand UO_1297 (O_1297,N_13593,N_12435);
nor UO_1298 (O_1298,N_14598,N_13730);
nor UO_1299 (O_1299,N_12806,N_13693);
and UO_1300 (O_1300,N_13566,N_14606);
or UO_1301 (O_1301,N_13788,N_12560);
nor UO_1302 (O_1302,N_12045,N_12478);
nor UO_1303 (O_1303,N_12994,N_14367);
nand UO_1304 (O_1304,N_12203,N_14999);
or UO_1305 (O_1305,N_13338,N_12579);
and UO_1306 (O_1306,N_13019,N_14979);
and UO_1307 (O_1307,N_14605,N_14806);
nand UO_1308 (O_1308,N_13279,N_13856);
or UO_1309 (O_1309,N_14689,N_12928);
or UO_1310 (O_1310,N_13550,N_12945);
nand UO_1311 (O_1311,N_14168,N_14316);
and UO_1312 (O_1312,N_14933,N_13791);
nand UO_1313 (O_1313,N_13909,N_12832);
nand UO_1314 (O_1314,N_13461,N_14394);
nor UO_1315 (O_1315,N_14465,N_12406);
and UO_1316 (O_1316,N_13954,N_12715);
nor UO_1317 (O_1317,N_14855,N_13349);
nand UO_1318 (O_1318,N_14900,N_12997);
nand UO_1319 (O_1319,N_13756,N_14888);
nor UO_1320 (O_1320,N_14617,N_13560);
xor UO_1321 (O_1321,N_12054,N_12983);
or UO_1322 (O_1322,N_13898,N_13073);
nor UO_1323 (O_1323,N_12183,N_13103);
nor UO_1324 (O_1324,N_12300,N_12004);
or UO_1325 (O_1325,N_14483,N_13532);
or UO_1326 (O_1326,N_13921,N_13820);
nand UO_1327 (O_1327,N_13672,N_14252);
nand UO_1328 (O_1328,N_12711,N_13636);
and UO_1329 (O_1329,N_13500,N_13880);
or UO_1330 (O_1330,N_14002,N_14485);
xor UO_1331 (O_1331,N_14805,N_12146);
or UO_1332 (O_1332,N_12395,N_14313);
nand UO_1333 (O_1333,N_14515,N_13860);
or UO_1334 (O_1334,N_14343,N_13446);
or UO_1335 (O_1335,N_14006,N_12601);
and UO_1336 (O_1336,N_12511,N_13875);
nand UO_1337 (O_1337,N_14645,N_14489);
or UO_1338 (O_1338,N_12517,N_14135);
or UO_1339 (O_1339,N_14534,N_12100);
or UO_1340 (O_1340,N_14822,N_13611);
nor UO_1341 (O_1341,N_13574,N_14784);
nand UO_1342 (O_1342,N_13405,N_14264);
or UO_1343 (O_1343,N_14216,N_12026);
nand UO_1344 (O_1344,N_13946,N_12360);
nand UO_1345 (O_1345,N_13434,N_13595);
nor UO_1346 (O_1346,N_14460,N_13121);
nor UO_1347 (O_1347,N_12114,N_14961);
or UO_1348 (O_1348,N_13288,N_14965);
nor UO_1349 (O_1349,N_13771,N_13369);
and UO_1350 (O_1350,N_14273,N_12449);
or UO_1351 (O_1351,N_14768,N_13646);
nor UO_1352 (O_1352,N_12444,N_12710);
and UO_1353 (O_1353,N_12745,N_12731);
xor UO_1354 (O_1354,N_14958,N_13389);
nand UO_1355 (O_1355,N_14659,N_12662);
or UO_1356 (O_1356,N_13992,N_13871);
nand UO_1357 (O_1357,N_12222,N_13817);
or UO_1358 (O_1358,N_14420,N_14362);
nand UO_1359 (O_1359,N_14091,N_12547);
nor UO_1360 (O_1360,N_14454,N_14766);
and UO_1361 (O_1361,N_12000,N_13979);
nand UO_1362 (O_1362,N_12781,N_13176);
nor UO_1363 (O_1363,N_13867,N_14852);
and UO_1364 (O_1364,N_14963,N_12923);
nor UO_1365 (O_1365,N_14430,N_14959);
nor UO_1366 (O_1366,N_12963,N_12019);
nor UO_1367 (O_1367,N_12650,N_12991);
and UO_1368 (O_1368,N_12337,N_13988);
xor UO_1369 (O_1369,N_12368,N_14872);
or UO_1370 (O_1370,N_13743,N_13687);
nor UO_1371 (O_1371,N_12303,N_14148);
nand UO_1372 (O_1372,N_14332,N_12415);
nand UO_1373 (O_1373,N_13074,N_13886);
nor UO_1374 (O_1374,N_14066,N_13838);
or UO_1375 (O_1375,N_14916,N_12072);
or UO_1376 (O_1376,N_14291,N_14674);
nand UO_1377 (O_1377,N_13118,N_14393);
nand UO_1378 (O_1378,N_13072,N_14069);
nor UO_1379 (O_1379,N_14740,N_13280);
nand UO_1380 (O_1380,N_14565,N_13254);
nand UO_1381 (O_1381,N_13848,N_12846);
or UO_1382 (O_1382,N_14466,N_14721);
nand UO_1383 (O_1383,N_14125,N_14312);
nor UO_1384 (O_1384,N_14320,N_12452);
and UO_1385 (O_1385,N_14603,N_12033);
nor UO_1386 (O_1386,N_12379,N_12586);
or UO_1387 (O_1387,N_12801,N_14306);
and UO_1388 (O_1388,N_12015,N_13936);
nand UO_1389 (O_1389,N_13989,N_12084);
and UO_1390 (O_1390,N_12593,N_14409);
or UO_1391 (O_1391,N_12788,N_14109);
and UO_1392 (O_1392,N_12496,N_12984);
nand UO_1393 (O_1393,N_13430,N_13963);
and UO_1394 (O_1394,N_13536,N_12969);
nor UO_1395 (O_1395,N_12118,N_14228);
or UO_1396 (O_1396,N_13725,N_13828);
or UO_1397 (O_1397,N_13912,N_13324);
nand UO_1398 (O_1398,N_14368,N_13272);
and UO_1399 (O_1399,N_12610,N_12976);
nor UO_1400 (O_1400,N_14039,N_13893);
nand UO_1401 (O_1401,N_14018,N_12816);
or UO_1402 (O_1402,N_13618,N_14899);
nor UO_1403 (O_1403,N_13717,N_12237);
or UO_1404 (O_1404,N_13589,N_14983);
nor UO_1405 (O_1405,N_12227,N_13609);
and UO_1406 (O_1406,N_14427,N_12140);
or UO_1407 (O_1407,N_12129,N_12405);
or UO_1408 (O_1408,N_12134,N_12296);
xor UO_1409 (O_1409,N_12820,N_14814);
nor UO_1410 (O_1410,N_14596,N_14616);
or UO_1411 (O_1411,N_12795,N_12366);
nor UO_1412 (O_1412,N_14867,N_13558);
nand UO_1413 (O_1413,N_12037,N_14380);
nor UO_1414 (O_1414,N_14922,N_14407);
and UO_1415 (O_1415,N_13021,N_14094);
and UO_1416 (O_1416,N_14741,N_12616);
and UO_1417 (O_1417,N_12400,N_14437);
nor UO_1418 (O_1418,N_12459,N_13347);
nor UO_1419 (O_1419,N_12638,N_12020);
or UO_1420 (O_1420,N_13874,N_13774);
and UO_1421 (O_1421,N_13250,N_13985);
nand UO_1422 (O_1422,N_13229,N_14048);
or UO_1423 (O_1423,N_14758,N_13831);
and UO_1424 (O_1424,N_13099,N_13041);
nor UO_1425 (O_1425,N_14680,N_14816);
and UO_1426 (O_1426,N_12318,N_14170);
nand UO_1427 (O_1427,N_12782,N_13211);
nor UO_1428 (O_1428,N_14480,N_12564);
and UO_1429 (O_1429,N_12964,N_12684);
nor UO_1430 (O_1430,N_13976,N_12307);
or UO_1431 (O_1431,N_14188,N_12181);
nand UO_1432 (O_1432,N_12516,N_12039);
nand UO_1433 (O_1433,N_14536,N_13842);
nand UO_1434 (O_1434,N_12960,N_13899);
nand UO_1435 (O_1435,N_12674,N_13175);
or UO_1436 (O_1436,N_12326,N_14114);
nand UO_1437 (O_1437,N_14734,N_13776);
and UO_1438 (O_1438,N_12389,N_14030);
nor UO_1439 (O_1439,N_14089,N_14845);
nand UO_1440 (O_1440,N_14720,N_13273);
and UO_1441 (O_1441,N_14101,N_13951);
nor UO_1442 (O_1442,N_12454,N_13129);
nor UO_1443 (O_1443,N_14833,N_13745);
nor UO_1444 (O_1444,N_14356,N_14122);
and UO_1445 (O_1445,N_13765,N_12968);
or UO_1446 (O_1446,N_12844,N_12473);
nand UO_1447 (O_1447,N_13419,N_14810);
nor UO_1448 (O_1448,N_12189,N_14337);
nor UO_1449 (O_1449,N_14904,N_12590);
xnor UO_1450 (O_1450,N_13556,N_14350);
and UO_1451 (O_1451,N_12947,N_13731);
or UO_1452 (O_1452,N_14360,N_14650);
nand UO_1453 (O_1453,N_14024,N_14376);
or UO_1454 (O_1454,N_13815,N_12213);
nand UO_1455 (O_1455,N_14968,N_12770);
nor UO_1456 (O_1456,N_12470,N_14121);
nor UO_1457 (O_1457,N_13477,N_12970);
and UO_1458 (O_1458,N_13591,N_13846);
nand UO_1459 (O_1459,N_14683,N_14495);
or UO_1460 (O_1460,N_12220,N_12676);
nor UO_1461 (O_1461,N_13428,N_12742);
nor UO_1462 (O_1462,N_14341,N_13527);
nand UO_1463 (O_1463,N_14012,N_12108);
xnor UO_1464 (O_1464,N_12273,N_14642);
nand UO_1465 (O_1465,N_12682,N_13444);
nand UO_1466 (O_1466,N_12014,N_14238);
nand UO_1467 (O_1467,N_13091,N_14085);
nor UO_1468 (O_1468,N_12359,N_14496);
nand UO_1469 (O_1469,N_14621,N_12423);
or UO_1470 (O_1470,N_13248,N_13120);
or UO_1471 (O_1471,N_13632,N_12131);
and UO_1472 (O_1472,N_13594,N_13673);
nand UO_1473 (O_1473,N_14287,N_13466);
nor UO_1474 (O_1474,N_13628,N_14178);
nand UO_1475 (O_1475,N_14391,N_13852);
or UO_1476 (O_1476,N_13836,N_13940);
and UO_1477 (O_1477,N_12230,N_14578);
or UO_1478 (O_1478,N_13994,N_13000);
or UO_1479 (O_1479,N_12299,N_13483);
and UO_1480 (O_1480,N_12497,N_12647);
or UO_1481 (O_1481,N_14439,N_14412);
nor UO_1482 (O_1482,N_12993,N_12723);
nand UO_1483 (O_1483,N_12324,N_14604);
nor UO_1484 (O_1484,N_14769,N_13882);
or UO_1485 (O_1485,N_14315,N_13345);
nor UO_1486 (O_1486,N_13067,N_12737);
or UO_1487 (O_1487,N_12384,N_13694);
nand UO_1488 (O_1488,N_14518,N_13448);
or UO_1489 (O_1489,N_12350,N_13826);
nor UO_1490 (O_1490,N_12965,N_13059);
nand UO_1491 (O_1491,N_13043,N_13318);
nor UO_1492 (O_1492,N_13892,N_13697);
nor UO_1493 (O_1493,N_12457,N_12587);
nand UO_1494 (O_1494,N_13201,N_14695);
nand UO_1495 (O_1495,N_14990,N_12828);
nand UO_1496 (O_1496,N_14449,N_14630);
and UO_1497 (O_1497,N_14484,N_12778);
and UO_1498 (O_1498,N_14751,N_14083);
and UO_1499 (O_1499,N_12625,N_12357);
nor UO_1500 (O_1500,N_12238,N_14868);
nor UO_1501 (O_1501,N_14484,N_14253);
nand UO_1502 (O_1502,N_12816,N_13212);
or UO_1503 (O_1503,N_13349,N_14431);
or UO_1504 (O_1504,N_13910,N_13050);
xnor UO_1505 (O_1505,N_13829,N_13671);
and UO_1506 (O_1506,N_14391,N_14619);
or UO_1507 (O_1507,N_13034,N_13829);
nor UO_1508 (O_1508,N_13411,N_12820);
and UO_1509 (O_1509,N_12728,N_14623);
nor UO_1510 (O_1510,N_13988,N_12456);
or UO_1511 (O_1511,N_13982,N_12432);
nor UO_1512 (O_1512,N_14300,N_13069);
nor UO_1513 (O_1513,N_13351,N_12117);
xor UO_1514 (O_1514,N_12343,N_12110);
nand UO_1515 (O_1515,N_13401,N_13623);
nand UO_1516 (O_1516,N_14437,N_12125);
or UO_1517 (O_1517,N_12043,N_14688);
or UO_1518 (O_1518,N_13117,N_14348);
nor UO_1519 (O_1519,N_14701,N_13046);
nand UO_1520 (O_1520,N_14800,N_14748);
or UO_1521 (O_1521,N_14032,N_12508);
nor UO_1522 (O_1522,N_12345,N_14791);
and UO_1523 (O_1523,N_13079,N_13838);
and UO_1524 (O_1524,N_14060,N_12456);
nand UO_1525 (O_1525,N_14712,N_14355);
nand UO_1526 (O_1526,N_14726,N_12310);
nand UO_1527 (O_1527,N_13185,N_14217);
or UO_1528 (O_1528,N_14610,N_14806);
and UO_1529 (O_1529,N_14635,N_14079);
nand UO_1530 (O_1530,N_13279,N_13645);
nor UO_1531 (O_1531,N_14248,N_14158);
and UO_1532 (O_1532,N_13531,N_13941);
nand UO_1533 (O_1533,N_14310,N_14440);
and UO_1534 (O_1534,N_13950,N_14559);
nor UO_1535 (O_1535,N_12958,N_13866);
nor UO_1536 (O_1536,N_12174,N_13174);
nand UO_1537 (O_1537,N_13657,N_14785);
and UO_1538 (O_1538,N_14640,N_13536);
and UO_1539 (O_1539,N_13837,N_14360);
nand UO_1540 (O_1540,N_13888,N_14754);
nor UO_1541 (O_1541,N_13549,N_14859);
nand UO_1542 (O_1542,N_13972,N_13184);
and UO_1543 (O_1543,N_12400,N_12012);
nor UO_1544 (O_1544,N_12721,N_14733);
nand UO_1545 (O_1545,N_12367,N_12284);
or UO_1546 (O_1546,N_12727,N_12289);
nor UO_1547 (O_1547,N_13540,N_12658);
or UO_1548 (O_1548,N_13350,N_14177);
xnor UO_1549 (O_1549,N_12292,N_14855);
and UO_1550 (O_1550,N_14439,N_13837);
and UO_1551 (O_1551,N_14145,N_13617);
nor UO_1552 (O_1552,N_13207,N_13524);
nand UO_1553 (O_1553,N_14078,N_13756);
or UO_1554 (O_1554,N_12158,N_13688);
nand UO_1555 (O_1555,N_14403,N_12510);
or UO_1556 (O_1556,N_13213,N_14471);
and UO_1557 (O_1557,N_14592,N_13602);
or UO_1558 (O_1558,N_12308,N_13784);
and UO_1559 (O_1559,N_13332,N_14512);
nand UO_1560 (O_1560,N_13887,N_13652);
or UO_1561 (O_1561,N_13766,N_14689);
or UO_1562 (O_1562,N_12982,N_13811);
and UO_1563 (O_1563,N_12849,N_12010);
nand UO_1564 (O_1564,N_12037,N_12879);
nor UO_1565 (O_1565,N_14347,N_14283);
nand UO_1566 (O_1566,N_13943,N_13114);
and UO_1567 (O_1567,N_12811,N_14907);
nor UO_1568 (O_1568,N_14375,N_12171);
nor UO_1569 (O_1569,N_13692,N_12080);
nor UO_1570 (O_1570,N_14375,N_12225);
and UO_1571 (O_1571,N_14533,N_12035);
or UO_1572 (O_1572,N_14637,N_12303);
and UO_1573 (O_1573,N_12052,N_12152);
nor UO_1574 (O_1574,N_14943,N_12649);
or UO_1575 (O_1575,N_14795,N_12138);
nand UO_1576 (O_1576,N_13331,N_14021);
xor UO_1577 (O_1577,N_13657,N_14015);
nand UO_1578 (O_1578,N_13304,N_14687);
nor UO_1579 (O_1579,N_13380,N_14612);
nor UO_1580 (O_1580,N_13778,N_14230);
nand UO_1581 (O_1581,N_13695,N_14024);
nor UO_1582 (O_1582,N_13390,N_14201);
or UO_1583 (O_1583,N_13902,N_14567);
nand UO_1584 (O_1584,N_14474,N_12949);
xor UO_1585 (O_1585,N_12015,N_12947);
nand UO_1586 (O_1586,N_14266,N_13942);
or UO_1587 (O_1587,N_12731,N_14294);
nor UO_1588 (O_1588,N_12117,N_12801);
or UO_1589 (O_1589,N_12975,N_12012);
or UO_1590 (O_1590,N_12969,N_12610);
nor UO_1591 (O_1591,N_13868,N_14615);
and UO_1592 (O_1592,N_12996,N_12168);
and UO_1593 (O_1593,N_12106,N_13316);
or UO_1594 (O_1594,N_12615,N_13096);
or UO_1595 (O_1595,N_14038,N_12256);
and UO_1596 (O_1596,N_14383,N_13485);
and UO_1597 (O_1597,N_14292,N_13378);
nor UO_1598 (O_1598,N_12145,N_13915);
nor UO_1599 (O_1599,N_14535,N_13215);
and UO_1600 (O_1600,N_13758,N_12810);
nor UO_1601 (O_1601,N_12631,N_13112);
and UO_1602 (O_1602,N_12803,N_14924);
nor UO_1603 (O_1603,N_14266,N_14006);
and UO_1604 (O_1604,N_13068,N_14512);
nor UO_1605 (O_1605,N_12899,N_13712);
and UO_1606 (O_1606,N_12375,N_12571);
nand UO_1607 (O_1607,N_14327,N_14423);
and UO_1608 (O_1608,N_14634,N_14002);
and UO_1609 (O_1609,N_12831,N_14488);
nand UO_1610 (O_1610,N_13788,N_12247);
or UO_1611 (O_1611,N_14329,N_12072);
nand UO_1612 (O_1612,N_14316,N_14270);
or UO_1613 (O_1613,N_14038,N_13434);
or UO_1614 (O_1614,N_14196,N_12063);
or UO_1615 (O_1615,N_13842,N_12874);
or UO_1616 (O_1616,N_14358,N_13604);
and UO_1617 (O_1617,N_12750,N_14426);
or UO_1618 (O_1618,N_14290,N_12213);
nor UO_1619 (O_1619,N_13979,N_13479);
and UO_1620 (O_1620,N_12585,N_14347);
and UO_1621 (O_1621,N_14999,N_14568);
and UO_1622 (O_1622,N_12045,N_13601);
or UO_1623 (O_1623,N_12037,N_13745);
and UO_1624 (O_1624,N_12149,N_12493);
and UO_1625 (O_1625,N_14756,N_12874);
nor UO_1626 (O_1626,N_13887,N_13202);
nor UO_1627 (O_1627,N_14524,N_12757);
nand UO_1628 (O_1628,N_12346,N_14152);
nand UO_1629 (O_1629,N_14156,N_12080);
and UO_1630 (O_1630,N_14264,N_13467);
and UO_1631 (O_1631,N_14442,N_12280);
and UO_1632 (O_1632,N_13617,N_14590);
and UO_1633 (O_1633,N_14296,N_14469);
nand UO_1634 (O_1634,N_14127,N_13397);
nor UO_1635 (O_1635,N_14137,N_14782);
and UO_1636 (O_1636,N_13116,N_12907);
nor UO_1637 (O_1637,N_12687,N_14015);
nand UO_1638 (O_1638,N_13917,N_14329);
and UO_1639 (O_1639,N_12401,N_14272);
nor UO_1640 (O_1640,N_13778,N_12630);
nor UO_1641 (O_1641,N_14081,N_14591);
nand UO_1642 (O_1642,N_14496,N_14230);
or UO_1643 (O_1643,N_13455,N_12924);
and UO_1644 (O_1644,N_13435,N_14734);
nor UO_1645 (O_1645,N_13721,N_12114);
or UO_1646 (O_1646,N_14100,N_12074);
nor UO_1647 (O_1647,N_12939,N_12311);
nand UO_1648 (O_1648,N_13272,N_13845);
nand UO_1649 (O_1649,N_14175,N_12504);
and UO_1650 (O_1650,N_14153,N_14642);
and UO_1651 (O_1651,N_13758,N_13125);
nor UO_1652 (O_1652,N_14063,N_14122);
nor UO_1653 (O_1653,N_13514,N_12814);
or UO_1654 (O_1654,N_13039,N_13381);
and UO_1655 (O_1655,N_13973,N_14278);
or UO_1656 (O_1656,N_13304,N_13936);
nor UO_1657 (O_1657,N_12600,N_13552);
xor UO_1658 (O_1658,N_14386,N_14086);
or UO_1659 (O_1659,N_12950,N_12686);
and UO_1660 (O_1660,N_14420,N_12459);
nor UO_1661 (O_1661,N_12199,N_13410);
and UO_1662 (O_1662,N_13962,N_13715);
and UO_1663 (O_1663,N_14921,N_14211);
or UO_1664 (O_1664,N_14145,N_13634);
and UO_1665 (O_1665,N_13773,N_14432);
nand UO_1666 (O_1666,N_12296,N_14488);
or UO_1667 (O_1667,N_12903,N_13246);
nand UO_1668 (O_1668,N_12717,N_13578);
and UO_1669 (O_1669,N_14752,N_14067);
nor UO_1670 (O_1670,N_14196,N_12462);
and UO_1671 (O_1671,N_14826,N_14218);
xor UO_1672 (O_1672,N_14299,N_13279);
or UO_1673 (O_1673,N_13684,N_14053);
and UO_1674 (O_1674,N_12164,N_14573);
or UO_1675 (O_1675,N_13757,N_12941);
or UO_1676 (O_1676,N_14254,N_12275);
nand UO_1677 (O_1677,N_12620,N_12140);
or UO_1678 (O_1678,N_14837,N_14651);
nand UO_1679 (O_1679,N_12273,N_12875);
or UO_1680 (O_1680,N_12107,N_12221);
or UO_1681 (O_1681,N_14862,N_14590);
and UO_1682 (O_1682,N_14279,N_12910);
or UO_1683 (O_1683,N_14950,N_13415);
and UO_1684 (O_1684,N_13199,N_12080);
or UO_1685 (O_1685,N_14170,N_12747);
and UO_1686 (O_1686,N_14322,N_13785);
nor UO_1687 (O_1687,N_12714,N_13634);
or UO_1688 (O_1688,N_12489,N_13783);
and UO_1689 (O_1689,N_14563,N_12390);
nor UO_1690 (O_1690,N_14376,N_12655);
nand UO_1691 (O_1691,N_14695,N_12814);
nand UO_1692 (O_1692,N_12463,N_13951);
nand UO_1693 (O_1693,N_14690,N_13860);
xor UO_1694 (O_1694,N_12439,N_13786);
or UO_1695 (O_1695,N_13588,N_12563);
or UO_1696 (O_1696,N_12169,N_14592);
nor UO_1697 (O_1697,N_13855,N_14707);
and UO_1698 (O_1698,N_13921,N_13280);
nor UO_1699 (O_1699,N_12333,N_13215);
and UO_1700 (O_1700,N_14513,N_13157);
nor UO_1701 (O_1701,N_14142,N_13325);
or UO_1702 (O_1702,N_13592,N_13376);
and UO_1703 (O_1703,N_12131,N_14618);
or UO_1704 (O_1704,N_12057,N_13819);
nor UO_1705 (O_1705,N_12562,N_13473);
or UO_1706 (O_1706,N_13811,N_14306);
nand UO_1707 (O_1707,N_14213,N_13596);
nor UO_1708 (O_1708,N_13981,N_14453);
nand UO_1709 (O_1709,N_13612,N_12501);
nand UO_1710 (O_1710,N_14818,N_14837);
and UO_1711 (O_1711,N_12307,N_12092);
and UO_1712 (O_1712,N_14797,N_14315);
nand UO_1713 (O_1713,N_13785,N_14479);
nor UO_1714 (O_1714,N_13767,N_14096);
nor UO_1715 (O_1715,N_14814,N_13174);
and UO_1716 (O_1716,N_12641,N_13072);
nor UO_1717 (O_1717,N_12910,N_14724);
or UO_1718 (O_1718,N_13436,N_14961);
and UO_1719 (O_1719,N_13044,N_14485);
nor UO_1720 (O_1720,N_12462,N_12306);
and UO_1721 (O_1721,N_13648,N_14499);
nor UO_1722 (O_1722,N_13752,N_14780);
nor UO_1723 (O_1723,N_14257,N_12783);
nor UO_1724 (O_1724,N_14541,N_14954);
nor UO_1725 (O_1725,N_14319,N_14872);
nand UO_1726 (O_1726,N_12736,N_13231);
and UO_1727 (O_1727,N_12876,N_14940);
nor UO_1728 (O_1728,N_14356,N_14664);
nand UO_1729 (O_1729,N_12062,N_14650);
and UO_1730 (O_1730,N_12004,N_13563);
nand UO_1731 (O_1731,N_13221,N_12428);
nor UO_1732 (O_1732,N_13312,N_12909);
nor UO_1733 (O_1733,N_14279,N_14316);
and UO_1734 (O_1734,N_14671,N_12017);
and UO_1735 (O_1735,N_12533,N_12385);
nand UO_1736 (O_1736,N_14468,N_14785);
nand UO_1737 (O_1737,N_14912,N_13848);
or UO_1738 (O_1738,N_14436,N_12024);
and UO_1739 (O_1739,N_13726,N_14340);
nor UO_1740 (O_1740,N_12542,N_12705);
and UO_1741 (O_1741,N_13959,N_14124);
nor UO_1742 (O_1742,N_13478,N_13042);
nand UO_1743 (O_1743,N_14925,N_14721);
or UO_1744 (O_1744,N_12739,N_14231);
xnor UO_1745 (O_1745,N_12526,N_14614);
nor UO_1746 (O_1746,N_13492,N_12119);
xor UO_1747 (O_1747,N_13329,N_14427);
or UO_1748 (O_1748,N_13659,N_12941);
and UO_1749 (O_1749,N_13107,N_14692);
and UO_1750 (O_1750,N_14854,N_13715);
or UO_1751 (O_1751,N_12056,N_12939);
nor UO_1752 (O_1752,N_14022,N_13997);
nand UO_1753 (O_1753,N_14147,N_14838);
and UO_1754 (O_1754,N_14223,N_12196);
or UO_1755 (O_1755,N_14251,N_12780);
nor UO_1756 (O_1756,N_14192,N_14923);
or UO_1757 (O_1757,N_13012,N_12229);
nand UO_1758 (O_1758,N_12172,N_14619);
nor UO_1759 (O_1759,N_14257,N_13867);
or UO_1760 (O_1760,N_14476,N_14153);
and UO_1761 (O_1761,N_14752,N_14487);
nand UO_1762 (O_1762,N_12058,N_14284);
nor UO_1763 (O_1763,N_12664,N_13386);
and UO_1764 (O_1764,N_13534,N_12928);
and UO_1765 (O_1765,N_12942,N_13653);
xnor UO_1766 (O_1766,N_14228,N_14490);
and UO_1767 (O_1767,N_12646,N_13533);
nor UO_1768 (O_1768,N_14275,N_13949);
nand UO_1769 (O_1769,N_12512,N_12275);
nor UO_1770 (O_1770,N_12898,N_14686);
nor UO_1771 (O_1771,N_12000,N_12224);
or UO_1772 (O_1772,N_14113,N_12598);
nand UO_1773 (O_1773,N_13472,N_14117);
nor UO_1774 (O_1774,N_13453,N_12392);
or UO_1775 (O_1775,N_12409,N_12337);
nor UO_1776 (O_1776,N_13916,N_12774);
or UO_1777 (O_1777,N_13008,N_13079);
nor UO_1778 (O_1778,N_14024,N_14133);
nor UO_1779 (O_1779,N_13191,N_14168);
nand UO_1780 (O_1780,N_14936,N_12574);
and UO_1781 (O_1781,N_14564,N_12666);
nor UO_1782 (O_1782,N_14155,N_14460);
nand UO_1783 (O_1783,N_13402,N_13578);
nor UO_1784 (O_1784,N_12854,N_12461);
and UO_1785 (O_1785,N_12690,N_12140);
or UO_1786 (O_1786,N_13347,N_13164);
nor UO_1787 (O_1787,N_13404,N_12376);
and UO_1788 (O_1788,N_12300,N_14073);
nand UO_1789 (O_1789,N_13630,N_13749);
and UO_1790 (O_1790,N_14573,N_13482);
nor UO_1791 (O_1791,N_12432,N_12163);
and UO_1792 (O_1792,N_14849,N_12849);
nand UO_1793 (O_1793,N_14184,N_12350);
or UO_1794 (O_1794,N_14078,N_14580);
or UO_1795 (O_1795,N_12308,N_14486);
nand UO_1796 (O_1796,N_14013,N_12171);
or UO_1797 (O_1797,N_12642,N_14808);
nand UO_1798 (O_1798,N_14949,N_13123);
or UO_1799 (O_1799,N_14988,N_13629);
or UO_1800 (O_1800,N_14511,N_13136);
or UO_1801 (O_1801,N_13543,N_14092);
nor UO_1802 (O_1802,N_12901,N_13549);
nor UO_1803 (O_1803,N_12025,N_14513);
and UO_1804 (O_1804,N_12438,N_13883);
and UO_1805 (O_1805,N_12243,N_12922);
or UO_1806 (O_1806,N_12266,N_14027);
nor UO_1807 (O_1807,N_13292,N_12868);
or UO_1808 (O_1808,N_13263,N_13617);
nor UO_1809 (O_1809,N_14054,N_13829);
nand UO_1810 (O_1810,N_12701,N_14400);
or UO_1811 (O_1811,N_14256,N_14093);
nand UO_1812 (O_1812,N_14445,N_13733);
nor UO_1813 (O_1813,N_13632,N_14194);
and UO_1814 (O_1814,N_14520,N_12467);
nand UO_1815 (O_1815,N_14171,N_13690);
or UO_1816 (O_1816,N_12914,N_12503);
nor UO_1817 (O_1817,N_14982,N_14202);
nor UO_1818 (O_1818,N_12741,N_13641);
or UO_1819 (O_1819,N_12364,N_12311);
or UO_1820 (O_1820,N_14843,N_13315);
nand UO_1821 (O_1821,N_13472,N_14488);
or UO_1822 (O_1822,N_14509,N_13104);
nor UO_1823 (O_1823,N_12670,N_14481);
or UO_1824 (O_1824,N_13049,N_12902);
or UO_1825 (O_1825,N_13773,N_13263);
and UO_1826 (O_1826,N_14693,N_13994);
or UO_1827 (O_1827,N_12408,N_13065);
and UO_1828 (O_1828,N_13868,N_13376);
and UO_1829 (O_1829,N_14253,N_14048);
nor UO_1830 (O_1830,N_14008,N_14566);
nor UO_1831 (O_1831,N_12735,N_13031);
nand UO_1832 (O_1832,N_14665,N_14470);
or UO_1833 (O_1833,N_13145,N_12884);
nand UO_1834 (O_1834,N_13370,N_12536);
or UO_1835 (O_1835,N_12339,N_14729);
nand UO_1836 (O_1836,N_13855,N_13049);
or UO_1837 (O_1837,N_12051,N_12670);
nand UO_1838 (O_1838,N_12712,N_13693);
and UO_1839 (O_1839,N_13927,N_13820);
and UO_1840 (O_1840,N_12678,N_14485);
or UO_1841 (O_1841,N_12571,N_14039);
or UO_1842 (O_1842,N_14450,N_14396);
nand UO_1843 (O_1843,N_14925,N_13686);
nor UO_1844 (O_1844,N_12160,N_13705);
nand UO_1845 (O_1845,N_12785,N_13424);
and UO_1846 (O_1846,N_13529,N_13825);
nor UO_1847 (O_1847,N_12232,N_12364);
or UO_1848 (O_1848,N_13910,N_12783);
and UO_1849 (O_1849,N_12944,N_13686);
or UO_1850 (O_1850,N_12111,N_12434);
and UO_1851 (O_1851,N_13328,N_13578);
nand UO_1852 (O_1852,N_13994,N_13936);
and UO_1853 (O_1853,N_12457,N_12610);
or UO_1854 (O_1854,N_13804,N_12049);
nor UO_1855 (O_1855,N_14472,N_12573);
nand UO_1856 (O_1856,N_14674,N_13610);
nand UO_1857 (O_1857,N_12888,N_12762);
nor UO_1858 (O_1858,N_13746,N_12124);
nor UO_1859 (O_1859,N_12145,N_12609);
and UO_1860 (O_1860,N_14270,N_12579);
nand UO_1861 (O_1861,N_12073,N_13863);
and UO_1862 (O_1862,N_13469,N_14725);
nor UO_1863 (O_1863,N_14025,N_14965);
nand UO_1864 (O_1864,N_13856,N_12455);
nand UO_1865 (O_1865,N_12416,N_13191);
nand UO_1866 (O_1866,N_14936,N_12370);
nor UO_1867 (O_1867,N_14093,N_14929);
nand UO_1868 (O_1868,N_14211,N_14351);
and UO_1869 (O_1869,N_14226,N_13102);
nand UO_1870 (O_1870,N_13739,N_12551);
or UO_1871 (O_1871,N_14526,N_12499);
or UO_1872 (O_1872,N_12054,N_14837);
nand UO_1873 (O_1873,N_12927,N_12005);
or UO_1874 (O_1874,N_13658,N_14675);
and UO_1875 (O_1875,N_14234,N_13252);
or UO_1876 (O_1876,N_14536,N_13568);
and UO_1877 (O_1877,N_13291,N_12195);
nor UO_1878 (O_1878,N_12061,N_13699);
or UO_1879 (O_1879,N_12972,N_13902);
and UO_1880 (O_1880,N_14512,N_13064);
nand UO_1881 (O_1881,N_12012,N_12303);
or UO_1882 (O_1882,N_14449,N_13178);
nand UO_1883 (O_1883,N_14971,N_13768);
nor UO_1884 (O_1884,N_14204,N_14391);
and UO_1885 (O_1885,N_12189,N_12869);
nor UO_1886 (O_1886,N_14757,N_12900);
nand UO_1887 (O_1887,N_14730,N_12676);
nor UO_1888 (O_1888,N_13175,N_13279);
nand UO_1889 (O_1889,N_12370,N_12951);
or UO_1890 (O_1890,N_12425,N_13422);
nand UO_1891 (O_1891,N_14863,N_12798);
or UO_1892 (O_1892,N_14765,N_12282);
and UO_1893 (O_1893,N_12742,N_12792);
nor UO_1894 (O_1894,N_12263,N_13196);
nand UO_1895 (O_1895,N_12387,N_12126);
nor UO_1896 (O_1896,N_14675,N_12466);
nor UO_1897 (O_1897,N_13016,N_12944);
nor UO_1898 (O_1898,N_14814,N_12818);
nor UO_1899 (O_1899,N_14955,N_12423);
nand UO_1900 (O_1900,N_13212,N_13337);
nor UO_1901 (O_1901,N_12006,N_13422);
nand UO_1902 (O_1902,N_12436,N_12724);
nand UO_1903 (O_1903,N_13607,N_12457);
and UO_1904 (O_1904,N_14377,N_13975);
nor UO_1905 (O_1905,N_14895,N_12352);
and UO_1906 (O_1906,N_12432,N_13564);
nand UO_1907 (O_1907,N_13393,N_13844);
or UO_1908 (O_1908,N_14879,N_13791);
nor UO_1909 (O_1909,N_13317,N_13594);
nor UO_1910 (O_1910,N_12544,N_14434);
or UO_1911 (O_1911,N_14394,N_12766);
nand UO_1912 (O_1912,N_12823,N_12846);
or UO_1913 (O_1913,N_13465,N_12801);
and UO_1914 (O_1914,N_12469,N_14817);
or UO_1915 (O_1915,N_13891,N_14559);
or UO_1916 (O_1916,N_12323,N_12693);
and UO_1917 (O_1917,N_14560,N_13309);
or UO_1918 (O_1918,N_12091,N_12304);
nor UO_1919 (O_1919,N_12942,N_12971);
and UO_1920 (O_1920,N_12973,N_13236);
nand UO_1921 (O_1921,N_13501,N_12545);
and UO_1922 (O_1922,N_12771,N_13388);
nand UO_1923 (O_1923,N_13714,N_13832);
nor UO_1924 (O_1924,N_14145,N_14929);
and UO_1925 (O_1925,N_14859,N_14992);
nand UO_1926 (O_1926,N_13556,N_13725);
nor UO_1927 (O_1927,N_14991,N_13443);
or UO_1928 (O_1928,N_13574,N_14125);
nand UO_1929 (O_1929,N_13969,N_13148);
or UO_1930 (O_1930,N_12887,N_14448);
and UO_1931 (O_1931,N_14915,N_12807);
or UO_1932 (O_1932,N_12218,N_13274);
nand UO_1933 (O_1933,N_13995,N_12217);
nor UO_1934 (O_1934,N_13305,N_14419);
nor UO_1935 (O_1935,N_12062,N_12663);
nor UO_1936 (O_1936,N_13471,N_14141);
nand UO_1937 (O_1937,N_13488,N_14272);
or UO_1938 (O_1938,N_12375,N_12367);
and UO_1939 (O_1939,N_13944,N_13555);
nor UO_1940 (O_1940,N_12483,N_14827);
and UO_1941 (O_1941,N_14623,N_14613);
nand UO_1942 (O_1942,N_14054,N_13622);
and UO_1943 (O_1943,N_12967,N_14867);
or UO_1944 (O_1944,N_14380,N_14583);
nor UO_1945 (O_1945,N_12548,N_12563);
or UO_1946 (O_1946,N_13174,N_14889);
and UO_1947 (O_1947,N_12619,N_14262);
and UO_1948 (O_1948,N_14501,N_14996);
or UO_1949 (O_1949,N_12986,N_13886);
and UO_1950 (O_1950,N_14188,N_12698);
and UO_1951 (O_1951,N_14698,N_12477);
nand UO_1952 (O_1952,N_14585,N_13620);
and UO_1953 (O_1953,N_13085,N_13134);
nor UO_1954 (O_1954,N_14727,N_14578);
nand UO_1955 (O_1955,N_12845,N_13547);
and UO_1956 (O_1956,N_13737,N_13693);
or UO_1957 (O_1957,N_14903,N_14160);
or UO_1958 (O_1958,N_12390,N_13586);
or UO_1959 (O_1959,N_14795,N_12958);
or UO_1960 (O_1960,N_14735,N_13419);
or UO_1961 (O_1961,N_13492,N_14070);
and UO_1962 (O_1962,N_13951,N_13616);
nand UO_1963 (O_1963,N_12917,N_13665);
nand UO_1964 (O_1964,N_12689,N_14785);
nand UO_1965 (O_1965,N_13728,N_14269);
nor UO_1966 (O_1966,N_12498,N_14622);
and UO_1967 (O_1967,N_13003,N_13100);
and UO_1968 (O_1968,N_12712,N_13024);
or UO_1969 (O_1969,N_13362,N_14791);
and UO_1970 (O_1970,N_13496,N_13526);
nor UO_1971 (O_1971,N_12946,N_12408);
and UO_1972 (O_1972,N_13246,N_13377);
and UO_1973 (O_1973,N_14967,N_13990);
and UO_1974 (O_1974,N_13921,N_13220);
nand UO_1975 (O_1975,N_12812,N_14096);
or UO_1976 (O_1976,N_13873,N_12610);
nor UO_1977 (O_1977,N_12741,N_13721);
nand UO_1978 (O_1978,N_12830,N_12488);
nand UO_1979 (O_1979,N_12501,N_12119);
or UO_1980 (O_1980,N_13342,N_12020);
or UO_1981 (O_1981,N_13265,N_12679);
nand UO_1982 (O_1982,N_14252,N_14409);
and UO_1983 (O_1983,N_12650,N_13099);
and UO_1984 (O_1984,N_12250,N_12219);
nor UO_1985 (O_1985,N_13683,N_14710);
nand UO_1986 (O_1986,N_14484,N_12800);
nand UO_1987 (O_1987,N_14337,N_14161);
nor UO_1988 (O_1988,N_14164,N_13017);
or UO_1989 (O_1989,N_14005,N_13161);
nand UO_1990 (O_1990,N_12273,N_13313);
nand UO_1991 (O_1991,N_14394,N_12293);
and UO_1992 (O_1992,N_12111,N_13613);
nand UO_1993 (O_1993,N_12761,N_12808);
nor UO_1994 (O_1994,N_13765,N_13289);
xor UO_1995 (O_1995,N_14028,N_12007);
nand UO_1996 (O_1996,N_13744,N_12513);
and UO_1997 (O_1997,N_14733,N_12248);
and UO_1998 (O_1998,N_12737,N_12647);
and UO_1999 (O_1999,N_14890,N_12731);
endmodule