module basic_500_3000_500_6_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_341,In_245);
nor U1 (N_1,In_150,In_56);
and U2 (N_2,In_71,In_432);
xnor U3 (N_3,In_73,In_433);
nand U4 (N_4,In_440,In_463);
nor U5 (N_5,In_237,In_193);
nand U6 (N_6,In_422,In_89);
and U7 (N_7,In_457,In_207);
and U8 (N_8,In_498,In_389);
xor U9 (N_9,In_59,In_31);
and U10 (N_10,In_214,In_372);
and U11 (N_11,In_343,In_0);
and U12 (N_12,In_19,In_197);
or U13 (N_13,In_24,In_32);
nor U14 (N_14,In_52,In_88);
xor U15 (N_15,In_278,In_83);
and U16 (N_16,In_431,In_441);
nor U17 (N_17,In_240,In_228);
nand U18 (N_18,In_231,In_98);
nand U19 (N_19,In_413,In_455);
nand U20 (N_20,In_232,In_419);
nand U21 (N_21,In_315,In_253);
nor U22 (N_22,In_279,In_406);
xnor U23 (N_23,In_70,In_388);
nand U24 (N_24,In_85,In_143);
xor U25 (N_25,In_472,In_181);
or U26 (N_26,In_484,In_421);
nand U27 (N_27,In_66,In_105);
xnor U28 (N_28,In_20,In_302);
and U29 (N_29,In_120,In_111);
or U30 (N_30,In_121,In_179);
nand U31 (N_31,In_86,In_337);
nor U32 (N_32,In_74,In_368);
or U33 (N_33,In_470,In_411);
nor U34 (N_34,In_362,In_53);
nor U35 (N_35,In_13,In_471);
or U36 (N_36,In_108,In_359);
nor U37 (N_37,In_296,In_187);
and U38 (N_38,In_447,In_162);
xor U39 (N_39,In_233,In_6);
xnor U40 (N_40,In_48,In_129);
or U41 (N_41,In_499,In_361);
or U42 (N_42,In_346,In_356);
or U43 (N_43,In_387,In_271);
or U44 (N_44,In_424,In_306);
xor U45 (N_45,In_436,In_177);
xnor U46 (N_46,In_286,In_115);
nor U47 (N_47,In_252,In_178);
or U48 (N_48,In_327,In_109);
or U49 (N_49,In_60,In_138);
nand U50 (N_50,In_204,In_225);
and U51 (N_51,In_423,In_324);
xnor U52 (N_52,In_259,In_325);
nand U53 (N_53,In_23,In_191);
and U54 (N_54,In_209,In_134);
or U55 (N_55,In_65,In_301);
or U56 (N_56,In_78,In_404);
nor U57 (N_57,In_84,In_442);
or U58 (N_58,In_276,In_412);
nor U59 (N_59,In_418,In_45);
nand U60 (N_60,In_62,In_349);
and U61 (N_61,In_320,In_336);
nor U62 (N_62,In_246,In_257);
or U63 (N_63,In_54,In_303);
or U64 (N_64,In_307,In_364);
xnor U65 (N_65,In_168,In_132);
nand U66 (N_66,In_77,In_353);
nor U67 (N_67,In_100,In_399);
and U68 (N_68,In_415,In_216);
or U69 (N_69,In_288,In_348);
xor U70 (N_70,In_36,In_358);
nor U71 (N_71,In_392,In_158);
or U72 (N_72,In_99,In_127);
xor U73 (N_73,In_313,In_354);
and U74 (N_74,In_213,In_194);
and U75 (N_75,In_163,In_277);
xor U76 (N_76,In_68,In_117);
or U77 (N_77,In_275,In_160);
and U78 (N_78,In_322,In_211);
or U79 (N_79,In_481,In_185);
nand U80 (N_80,In_227,In_161);
and U81 (N_81,In_333,In_487);
and U82 (N_82,In_192,In_310);
nor U83 (N_83,In_55,In_126);
nand U84 (N_84,In_450,In_130);
xor U85 (N_85,In_5,In_135);
or U86 (N_86,In_328,In_61);
nand U87 (N_87,In_355,In_8);
or U88 (N_88,In_287,In_189);
or U89 (N_89,In_492,In_294);
nand U90 (N_90,In_262,In_391);
xor U91 (N_91,In_87,In_308);
or U92 (N_92,In_34,In_144);
xor U93 (N_93,In_403,In_488);
nor U94 (N_94,In_1,In_344);
xnor U95 (N_95,In_370,In_67);
and U96 (N_96,In_254,In_201);
nor U97 (N_97,In_205,In_206);
nor U98 (N_98,In_235,In_125);
or U99 (N_99,In_184,In_37);
or U100 (N_100,In_223,In_311);
and U101 (N_101,In_9,In_429);
or U102 (N_102,In_167,In_405);
and U103 (N_103,In_29,In_285);
nor U104 (N_104,In_342,In_293);
or U105 (N_105,In_480,In_122);
or U106 (N_106,In_208,In_81);
nor U107 (N_107,In_321,In_238);
nor U108 (N_108,In_467,In_452);
nor U109 (N_109,In_203,In_281);
or U110 (N_110,In_451,In_393);
nand U111 (N_111,In_35,In_239);
nand U112 (N_112,In_420,In_292);
nor U113 (N_113,In_448,In_381);
xor U114 (N_114,In_289,In_114);
nand U115 (N_115,In_494,In_458);
and U116 (N_116,In_386,In_106);
xor U117 (N_117,In_124,In_260);
xnor U118 (N_118,In_475,In_80);
nand U119 (N_119,In_16,In_15);
or U120 (N_120,In_107,In_305);
nor U121 (N_121,In_384,In_30);
and U122 (N_122,In_402,In_473);
nor U123 (N_123,In_247,In_335);
and U124 (N_124,In_215,In_338);
xor U125 (N_125,In_397,In_493);
nor U126 (N_126,In_266,In_425);
nand U127 (N_127,In_261,In_490);
xnor U128 (N_128,In_92,In_497);
or U129 (N_129,In_176,In_434);
xor U130 (N_130,In_159,In_196);
or U131 (N_131,In_438,In_17);
nor U132 (N_132,In_445,In_334);
nor U133 (N_133,In_118,In_50);
nand U134 (N_134,In_186,In_79);
and U135 (N_135,In_446,In_299);
xnor U136 (N_136,In_329,In_477);
xor U137 (N_137,In_116,In_38);
and U138 (N_138,In_456,In_256);
nand U139 (N_139,In_142,In_241);
xor U140 (N_140,In_222,In_251);
xnor U141 (N_141,In_464,In_273);
or U142 (N_142,In_283,In_270);
and U143 (N_143,In_435,In_146);
nand U144 (N_144,In_172,In_268);
or U145 (N_145,In_495,In_409);
xnor U146 (N_146,In_263,In_466);
and U147 (N_147,In_380,In_82);
nor U148 (N_148,In_11,In_234);
xor U149 (N_149,In_290,In_382);
nor U150 (N_150,In_377,In_258);
or U151 (N_151,In_376,In_443);
nor U152 (N_152,In_465,In_141);
nor U153 (N_153,In_375,In_102);
or U154 (N_154,In_7,In_408);
nor U155 (N_155,In_264,In_154);
and U156 (N_156,In_230,In_332);
or U157 (N_157,In_58,In_345);
nand U158 (N_158,In_212,In_42);
nand U159 (N_159,In_317,In_486);
or U160 (N_160,In_295,In_280);
or U161 (N_161,In_414,In_309);
nor U162 (N_162,In_369,In_416);
and U163 (N_163,In_323,In_491);
nand U164 (N_164,In_427,In_255);
xnor U165 (N_165,In_198,In_319);
xnor U166 (N_166,In_69,In_33);
xnor U167 (N_167,In_43,In_22);
nand U168 (N_168,In_395,In_312);
and U169 (N_169,In_156,In_357);
xnor U170 (N_170,In_26,In_27);
xor U171 (N_171,In_390,In_454);
nor U172 (N_172,In_166,In_482);
nor U173 (N_173,In_367,In_4);
nor U174 (N_174,In_284,In_76);
or U175 (N_175,In_373,In_94);
or U176 (N_176,In_152,In_366);
or U177 (N_177,In_330,In_331);
nor U178 (N_178,In_226,In_3);
and U179 (N_179,In_479,In_244);
nor U180 (N_180,In_63,In_183);
nor U181 (N_181,In_151,In_25);
nand U182 (N_182,In_385,In_137);
and U183 (N_183,In_47,In_170);
or U184 (N_184,In_430,In_378);
or U185 (N_185,In_426,In_272);
nand U186 (N_186,In_282,In_363);
xor U187 (N_187,In_39,In_379);
and U188 (N_188,In_173,In_171);
nor U189 (N_189,In_97,In_371);
and U190 (N_190,In_136,In_483);
nand U191 (N_191,In_10,In_417);
xnor U192 (N_192,In_439,In_360);
nor U193 (N_193,In_91,In_453);
nand U194 (N_194,In_220,In_123);
and U195 (N_195,In_219,In_224);
and U196 (N_196,In_218,In_131);
xnor U197 (N_197,In_14,In_51);
nor U198 (N_198,In_95,In_155);
nand U199 (N_199,In_304,In_41);
nor U200 (N_200,In_374,In_140);
nor U201 (N_201,In_103,In_242);
or U202 (N_202,In_119,In_221);
xor U203 (N_203,In_110,In_474);
nor U204 (N_204,In_326,In_298);
xor U205 (N_205,In_229,In_188);
and U206 (N_206,In_274,In_316);
nor U207 (N_207,In_265,In_396);
xor U208 (N_208,In_460,In_180);
or U209 (N_209,In_93,In_57);
nand U210 (N_210,In_407,In_365);
and U211 (N_211,In_478,In_28);
and U212 (N_212,In_496,In_400);
nand U213 (N_213,In_190,In_40);
nor U214 (N_214,In_199,In_145);
and U215 (N_215,In_462,In_394);
xnor U216 (N_216,In_291,In_164);
and U217 (N_217,In_182,In_398);
nand U218 (N_218,In_174,In_18);
nor U219 (N_219,In_459,In_485);
nand U220 (N_220,In_72,In_49);
nand U221 (N_221,In_243,In_21);
nand U222 (N_222,In_449,In_437);
xnor U223 (N_223,In_200,In_269);
and U224 (N_224,In_350,In_428);
xor U225 (N_225,In_153,In_64);
xnor U226 (N_226,In_157,In_113);
nor U227 (N_227,In_12,In_250);
nand U228 (N_228,In_2,In_401);
nand U229 (N_229,In_169,In_351);
nand U230 (N_230,In_44,In_46);
nor U231 (N_231,In_210,In_468);
or U232 (N_232,In_314,In_175);
xnor U233 (N_233,In_489,In_469);
or U234 (N_234,In_128,In_410);
nor U235 (N_235,In_217,In_195);
nor U236 (N_236,In_202,In_75);
and U237 (N_237,In_347,In_340);
nor U238 (N_238,In_339,In_318);
nor U239 (N_239,In_444,In_96);
nor U240 (N_240,In_149,In_476);
and U241 (N_241,In_101,In_165);
xor U242 (N_242,In_249,In_248);
nor U243 (N_243,In_383,In_112);
nor U244 (N_244,In_267,In_461);
xnor U245 (N_245,In_148,In_90);
xnor U246 (N_246,In_352,In_300);
nor U247 (N_247,In_104,In_133);
and U248 (N_248,In_297,In_139);
and U249 (N_249,In_147,In_236);
and U250 (N_250,In_91,In_387);
xor U251 (N_251,In_104,In_74);
xor U252 (N_252,In_114,In_70);
nor U253 (N_253,In_46,In_427);
and U254 (N_254,In_457,In_201);
nor U255 (N_255,In_224,In_498);
nand U256 (N_256,In_10,In_220);
nand U257 (N_257,In_183,In_112);
nor U258 (N_258,In_266,In_485);
xor U259 (N_259,In_349,In_175);
and U260 (N_260,In_277,In_288);
or U261 (N_261,In_424,In_328);
or U262 (N_262,In_109,In_375);
nor U263 (N_263,In_491,In_80);
nand U264 (N_264,In_52,In_335);
nand U265 (N_265,In_402,In_224);
nor U266 (N_266,In_47,In_24);
nor U267 (N_267,In_55,In_89);
nor U268 (N_268,In_347,In_213);
and U269 (N_269,In_387,In_359);
nor U270 (N_270,In_51,In_333);
or U271 (N_271,In_135,In_158);
nor U272 (N_272,In_92,In_45);
or U273 (N_273,In_325,In_295);
and U274 (N_274,In_264,In_267);
or U275 (N_275,In_37,In_124);
xor U276 (N_276,In_18,In_351);
nor U277 (N_277,In_309,In_389);
or U278 (N_278,In_496,In_346);
or U279 (N_279,In_346,In_200);
xnor U280 (N_280,In_489,In_123);
or U281 (N_281,In_196,In_164);
and U282 (N_282,In_55,In_95);
xor U283 (N_283,In_404,In_472);
nand U284 (N_284,In_273,In_92);
and U285 (N_285,In_15,In_152);
nand U286 (N_286,In_7,In_278);
or U287 (N_287,In_157,In_331);
nand U288 (N_288,In_66,In_470);
nor U289 (N_289,In_115,In_419);
nor U290 (N_290,In_414,In_322);
xor U291 (N_291,In_279,In_2);
xor U292 (N_292,In_470,In_455);
or U293 (N_293,In_272,In_231);
nor U294 (N_294,In_428,In_279);
xor U295 (N_295,In_34,In_200);
and U296 (N_296,In_165,In_308);
and U297 (N_297,In_169,In_196);
xnor U298 (N_298,In_86,In_241);
xnor U299 (N_299,In_326,In_220);
or U300 (N_300,In_36,In_369);
xnor U301 (N_301,In_450,In_4);
nand U302 (N_302,In_149,In_469);
xnor U303 (N_303,In_33,In_372);
nor U304 (N_304,In_17,In_268);
and U305 (N_305,In_23,In_414);
nor U306 (N_306,In_213,In_61);
nor U307 (N_307,In_216,In_277);
or U308 (N_308,In_192,In_357);
or U309 (N_309,In_242,In_234);
xnor U310 (N_310,In_468,In_388);
and U311 (N_311,In_204,In_130);
or U312 (N_312,In_419,In_108);
and U313 (N_313,In_72,In_147);
or U314 (N_314,In_278,In_343);
xor U315 (N_315,In_1,In_339);
and U316 (N_316,In_389,In_419);
nand U317 (N_317,In_392,In_479);
or U318 (N_318,In_481,In_215);
or U319 (N_319,In_208,In_397);
or U320 (N_320,In_491,In_84);
or U321 (N_321,In_394,In_47);
nand U322 (N_322,In_196,In_489);
nor U323 (N_323,In_148,In_435);
xnor U324 (N_324,In_373,In_367);
nand U325 (N_325,In_3,In_436);
or U326 (N_326,In_211,In_361);
and U327 (N_327,In_145,In_68);
nand U328 (N_328,In_191,In_256);
or U329 (N_329,In_335,In_391);
nor U330 (N_330,In_88,In_15);
xor U331 (N_331,In_59,In_277);
nor U332 (N_332,In_328,In_400);
xnor U333 (N_333,In_300,In_82);
nor U334 (N_334,In_402,In_85);
and U335 (N_335,In_421,In_206);
nor U336 (N_336,In_2,In_39);
or U337 (N_337,In_161,In_311);
and U338 (N_338,In_286,In_331);
nor U339 (N_339,In_467,In_84);
nand U340 (N_340,In_24,In_388);
xnor U341 (N_341,In_480,In_412);
and U342 (N_342,In_72,In_132);
and U343 (N_343,In_398,In_222);
and U344 (N_344,In_360,In_293);
xor U345 (N_345,In_145,In_438);
and U346 (N_346,In_406,In_44);
nor U347 (N_347,In_106,In_185);
nor U348 (N_348,In_308,In_397);
xnor U349 (N_349,In_150,In_212);
nand U350 (N_350,In_209,In_269);
nand U351 (N_351,In_21,In_165);
nor U352 (N_352,In_458,In_188);
nor U353 (N_353,In_324,In_458);
and U354 (N_354,In_348,In_425);
xor U355 (N_355,In_148,In_352);
nand U356 (N_356,In_440,In_183);
and U357 (N_357,In_353,In_429);
nand U358 (N_358,In_494,In_368);
xnor U359 (N_359,In_494,In_312);
xor U360 (N_360,In_24,In_471);
nand U361 (N_361,In_408,In_323);
or U362 (N_362,In_43,In_292);
nor U363 (N_363,In_313,In_197);
or U364 (N_364,In_37,In_49);
or U365 (N_365,In_20,In_157);
nor U366 (N_366,In_495,In_437);
nand U367 (N_367,In_465,In_340);
nand U368 (N_368,In_144,In_229);
nor U369 (N_369,In_99,In_75);
nor U370 (N_370,In_122,In_328);
nor U371 (N_371,In_351,In_477);
or U372 (N_372,In_324,In_464);
nand U373 (N_373,In_219,In_345);
nand U374 (N_374,In_82,In_416);
xor U375 (N_375,In_273,In_442);
or U376 (N_376,In_459,In_188);
and U377 (N_377,In_386,In_33);
and U378 (N_378,In_324,In_181);
and U379 (N_379,In_127,In_314);
or U380 (N_380,In_3,In_103);
nand U381 (N_381,In_40,In_174);
nor U382 (N_382,In_410,In_164);
or U383 (N_383,In_192,In_466);
nor U384 (N_384,In_349,In_75);
or U385 (N_385,In_391,In_229);
nor U386 (N_386,In_148,In_344);
and U387 (N_387,In_281,In_308);
or U388 (N_388,In_180,In_129);
nor U389 (N_389,In_138,In_374);
and U390 (N_390,In_360,In_254);
nor U391 (N_391,In_101,In_315);
and U392 (N_392,In_171,In_162);
or U393 (N_393,In_372,In_24);
or U394 (N_394,In_408,In_406);
or U395 (N_395,In_54,In_27);
nor U396 (N_396,In_286,In_465);
and U397 (N_397,In_73,In_134);
nand U398 (N_398,In_212,In_443);
xor U399 (N_399,In_405,In_366);
nand U400 (N_400,In_348,In_328);
or U401 (N_401,In_436,In_360);
nor U402 (N_402,In_219,In_307);
and U403 (N_403,In_349,In_393);
or U404 (N_404,In_279,In_184);
nor U405 (N_405,In_326,In_104);
xnor U406 (N_406,In_318,In_206);
nor U407 (N_407,In_456,In_453);
xnor U408 (N_408,In_24,In_145);
or U409 (N_409,In_62,In_209);
and U410 (N_410,In_456,In_475);
nand U411 (N_411,In_449,In_348);
or U412 (N_412,In_20,In_177);
or U413 (N_413,In_3,In_324);
and U414 (N_414,In_386,In_274);
xnor U415 (N_415,In_296,In_290);
nand U416 (N_416,In_115,In_57);
nor U417 (N_417,In_151,In_254);
xor U418 (N_418,In_476,In_265);
and U419 (N_419,In_221,In_443);
nor U420 (N_420,In_148,In_12);
xnor U421 (N_421,In_114,In_238);
nand U422 (N_422,In_359,In_307);
nor U423 (N_423,In_61,In_282);
xnor U424 (N_424,In_147,In_56);
xnor U425 (N_425,In_86,In_327);
and U426 (N_426,In_308,In_326);
nor U427 (N_427,In_139,In_318);
nand U428 (N_428,In_485,In_150);
nand U429 (N_429,In_402,In_345);
or U430 (N_430,In_244,In_68);
and U431 (N_431,In_153,In_192);
nand U432 (N_432,In_338,In_86);
xor U433 (N_433,In_472,In_119);
nor U434 (N_434,In_57,In_455);
and U435 (N_435,In_464,In_240);
or U436 (N_436,In_216,In_96);
nor U437 (N_437,In_381,In_254);
or U438 (N_438,In_128,In_341);
nand U439 (N_439,In_178,In_355);
xnor U440 (N_440,In_470,In_164);
nor U441 (N_441,In_472,In_7);
nor U442 (N_442,In_136,In_111);
nand U443 (N_443,In_204,In_106);
nand U444 (N_444,In_37,In_98);
xnor U445 (N_445,In_436,In_248);
and U446 (N_446,In_474,In_371);
and U447 (N_447,In_215,In_357);
xor U448 (N_448,In_37,In_489);
and U449 (N_449,In_496,In_238);
or U450 (N_450,In_318,In_313);
nand U451 (N_451,In_297,In_160);
nor U452 (N_452,In_57,In_165);
nor U453 (N_453,In_405,In_157);
nand U454 (N_454,In_95,In_377);
or U455 (N_455,In_130,In_12);
xor U456 (N_456,In_372,In_46);
xnor U457 (N_457,In_144,In_90);
xnor U458 (N_458,In_11,In_463);
nor U459 (N_459,In_208,In_185);
nor U460 (N_460,In_106,In_376);
nor U461 (N_461,In_167,In_375);
nor U462 (N_462,In_246,In_412);
nand U463 (N_463,In_31,In_195);
and U464 (N_464,In_458,In_401);
nand U465 (N_465,In_301,In_36);
nor U466 (N_466,In_290,In_9);
nand U467 (N_467,In_168,In_163);
nand U468 (N_468,In_136,In_4);
nor U469 (N_469,In_161,In_381);
or U470 (N_470,In_135,In_70);
and U471 (N_471,In_277,In_251);
xor U472 (N_472,In_441,In_217);
xnor U473 (N_473,In_51,In_25);
or U474 (N_474,In_345,In_115);
xnor U475 (N_475,In_305,In_48);
nor U476 (N_476,In_364,In_411);
or U477 (N_477,In_90,In_193);
nand U478 (N_478,In_240,In_138);
and U479 (N_479,In_365,In_234);
and U480 (N_480,In_200,In_169);
and U481 (N_481,In_388,In_333);
or U482 (N_482,In_488,In_301);
and U483 (N_483,In_487,In_120);
or U484 (N_484,In_408,In_55);
or U485 (N_485,In_28,In_30);
xnor U486 (N_486,In_132,In_135);
nand U487 (N_487,In_327,In_275);
nand U488 (N_488,In_356,In_338);
or U489 (N_489,In_331,In_402);
xnor U490 (N_490,In_142,In_437);
nor U491 (N_491,In_144,In_63);
and U492 (N_492,In_181,In_339);
and U493 (N_493,In_332,In_294);
xor U494 (N_494,In_130,In_437);
and U495 (N_495,In_399,In_123);
nor U496 (N_496,In_246,In_344);
xor U497 (N_497,In_492,In_379);
and U498 (N_498,In_401,In_209);
nand U499 (N_499,In_414,In_428);
or U500 (N_500,N_174,N_265);
nor U501 (N_501,N_210,N_492);
xnor U502 (N_502,N_273,N_457);
xor U503 (N_503,N_333,N_236);
nor U504 (N_504,N_446,N_369);
nand U505 (N_505,N_226,N_381);
xnor U506 (N_506,N_376,N_338);
nand U507 (N_507,N_342,N_349);
and U508 (N_508,N_81,N_461);
nor U509 (N_509,N_148,N_26);
or U510 (N_510,N_485,N_10);
xnor U511 (N_511,N_326,N_147);
or U512 (N_512,N_256,N_29);
and U513 (N_513,N_77,N_254);
xor U514 (N_514,N_483,N_490);
nor U515 (N_515,N_292,N_208);
nand U516 (N_516,N_137,N_387);
or U517 (N_517,N_94,N_334);
nand U518 (N_518,N_180,N_74);
and U519 (N_519,N_318,N_97);
nor U520 (N_520,N_340,N_34);
or U521 (N_521,N_282,N_451);
and U522 (N_522,N_319,N_305);
nand U523 (N_523,N_38,N_179);
or U524 (N_524,N_206,N_9);
or U525 (N_525,N_441,N_279);
nand U526 (N_526,N_310,N_371);
xor U527 (N_527,N_455,N_23);
or U528 (N_528,N_31,N_330);
nand U529 (N_529,N_413,N_225);
nor U530 (N_530,N_303,N_395);
nand U531 (N_531,N_471,N_11);
or U532 (N_532,N_307,N_216);
and U533 (N_533,N_96,N_86);
and U534 (N_534,N_90,N_76);
or U535 (N_535,N_394,N_211);
nor U536 (N_536,N_24,N_411);
and U537 (N_537,N_419,N_377);
xnor U538 (N_538,N_190,N_87);
and U539 (N_539,N_8,N_274);
nand U540 (N_540,N_129,N_169);
nor U541 (N_541,N_57,N_170);
or U542 (N_542,N_146,N_250);
nand U543 (N_543,N_162,N_16);
nand U544 (N_544,N_198,N_214);
or U545 (N_545,N_314,N_270);
and U546 (N_546,N_391,N_52);
or U547 (N_547,N_407,N_161);
and U548 (N_548,N_325,N_175);
and U549 (N_549,N_486,N_475);
xor U550 (N_550,N_405,N_164);
xor U551 (N_551,N_271,N_150);
nand U552 (N_552,N_71,N_215);
nand U553 (N_553,N_103,N_228);
nor U554 (N_554,N_131,N_470);
and U555 (N_555,N_439,N_158);
or U556 (N_556,N_312,N_429);
nand U557 (N_557,N_375,N_499);
xor U558 (N_558,N_384,N_6);
nor U559 (N_559,N_324,N_130);
xor U560 (N_560,N_336,N_35);
or U561 (N_561,N_496,N_67);
nor U562 (N_562,N_427,N_328);
nand U563 (N_563,N_252,N_347);
and U564 (N_564,N_68,N_444);
xor U565 (N_565,N_266,N_400);
nor U566 (N_566,N_308,N_493);
and U567 (N_567,N_187,N_61);
xor U568 (N_568,N_197,N_237);
xor U569 (N_569,N_351,N_346);
and U570 (N_570,N_465,N_431);
and U571 (N_571,N_232,N_79);
and U572 (N_572,N_433,N_401);
or U573 (N_573,N_443,N_293);
or U574 (N_574,N_116,N_337);
nand U575 (N_575,N_422,N_370);
xnor U576 (N_576,N_18,N_277);
nor U577 (N_577,N_269,N_434);
or U578 (N_578,N_218,N_188);
and U579 (N_579,N_481,N_70);
or U580 (N_580,N_123,N_363);
nor U581 (N_581,N_472,N_396);
xnor U582 (N_582,N_262,N_53);
or U583 (N_583,N_5,N_278);
nand U584 (N_584,N_113,N_44);
nor U585 (N_585,N_88,N_452);
nand U586 (N_586,N_403,N_260);
nand U587 (N_587,N_288,N_112);
xor U588 (N_588,N_120,N_241);
nand U589 (N_589,N_295,N_219);
nor U590 (N_590,N_311,N_320);
or U591 (N_591,N_152,N_244);
xor U592 (N_592,N_366,N_181);
nand U593 (N_593,N_64,N_383);
xor U594 (N_594,N_408,N_117);
xor U595 (N_595,N_423,N_454);
nor U596 (N_596,N_440,N_447);
and U597 (N_597,N_193,N_171);
or U598 (N_598,N_176,N_357);
nor U599 (N_599,N_378,N_107);
and U600 (N_600,N_235,N_41);
or U601 (N_601,N_425,N_209);
nand U602 (N_602,N_258,N_109);
nor U603 (N_603,N_283,N_361);
nand U604 (N_604,N_92,N_362);
nor U605 (N_605,N_259,N_478);
xnor U606 (N_606,N_205,N_255);
or U607 (N_607,N_54,N_48);
and U608 (N_608,N_168,N_105);
xnor U609 (N_609,N_257,N_416);
nor U610 (N_610,N_343,N_459);
nor U611 (N_611,N_217,N_195);
or U612 (N_612,N_263,N_368);
xor U613 (N_613,N_484,N_463);
nand U614 (N_614,N_315,N_138);
xor U615 (N_615,N_331,N_382);
xnor U616 (N_616,N_15,N_58);
or U617 (N_617,N_335,N_156);
xor U618 (N_618,N_294,N_108);
or U619 (N_619,N_221,N_245);
nand U620 (N_620,N_313,N_22);
and U621 (N_621,N_379,N_157);
and U622 (N_622,N_133,N_173);
nor U623 (N_623,N_40,N_359);
nor U624 (N_624,N_442,N_497);
nor U625 (N_625,N_80,N_111);
or U626 (N_626,N_115,N_280);
nand U627 (N_627,N_223,N_2);
and U628 (N_628,N_17,N_240);
nor U629 (N_629,N_358,N_426);
nand U630 (N_630,N_234,N_281);
xnor U631 (N_631,N_19,N_230);
xnor U632 (N_632,N_365,N_207);
or U633 (N_633,N_364,N_389);
and U634 (N_634,N_125,N_399);
or U635 (N_635,N_183,N_202);
nand U636 (N_636,N_247,N_144);
xor U637 (N_637,N_185,N_409);
nor U638 (N_638,N_388,N_78);
and U639 (N_639,N_178,N_200);
and U640 (N_640,N_300,N_151);
xor U641 (N_641,N_153,N_448);
xor U642 (N_642,N_229,N_332);
nand U643 (N_643,N_126,N_233);
or U644 (N_644,N_321,N_12);
and U645 (N_645,N_69,N_121);
nor U646 (N_646,N_424,N_415);
and U647 (N_647,N_37,N_380);
xor U648 (N_648,N_341,N_291);
and U649 (N_649,N_32,N_449);
nor U650 (N_650,N_199,N_201);
nor U651 (N_651,N_458,N_194);
xnor U652 (N_652,N_373,N_102);
nand U653 (N_653,N_212,N_385);
nand U654 (N_654,N_345,N_43);
and U655 (N_655,N_420,N_249);
nand U656 (N_656,N_127,N_353);
xor U657 (N_657,N_1,N_428);
or U658 (N_658,N_239,N_297);
or U659 (N_659,N_139,N_56);
xor U660 (N_660,N_322,N_272);
or U661 (N_661,N_390,N_268);
nand U662 (N_662,N_432,N_104);
nor U663 (N_663,N_404,N_356);
or U664 (N_664,N_145,N_75);
nand U665 (N_665,N_99,N_154);
and U666 (N_666,N_482,N_309);
nor U667 (N_667,N_298,N_39);
nor U668 (N_668,N_45,N_89);
nand U669 (N_669,N_82,N_73);
and U670 (N_670,N_438,N_242);
nand U671 (N_671,N_72,N_196);
or U672 (N_672,N_479,N_20);
or U673 (N_673,N_55,N_473);
or U674 (N_674,N_430,N_50);
xnor U675 (N_675,N_317,N_128);
xnor U676 (N_676,N_30,N_119);
xor U677 (N_677,N_98,N_464);
or U678 (N_678,N_192,N_495);
nand U679 (N_679,N_344,N_453);
nor U680 (N_680,N_163,N_60);
xor U681 (N_681,N_167,N_489);
xor U682 (N_682,N_110,N_287);
and U683 (N_683,N_142,N_477);
or U684 (N_684,N_460,N_227);
nor U685 (N_685,N_327,N_172);
and U686 (N_686,N_246,N_402);
or U687 (N_687,N_21,N_159);
or U688 (N_688,N_392,N_350);
nor U689 (N_689,N_231,N_301);
or U690 (N_690,N_186,N_323);
or U691 (N_691,N_397,N_49);
nor U692 (N_692,N_118,N_290);
and U693 (N_693,N_304,N_238);
xor U694 (N_694,N_42,N_136);
nand U695 (N_695,N_275,N_220);
or U696 (N_696,N_95,N_435);
nor U697 (N_697,N_184,N_135);
and U698 (N_698,N_134,N_84);
xor U699 (N_699,N_398,N_65);
xnor U700 (N_700,N_316,N_46);
and U701 (N_701,N_498,N_354);
xnor U702 (N_702,N_355,N_412);
xnor U703 (N_703,N_348,N_329);
xor U704 (N_704,N_421,N_306);
nand U705 (N_705,N_469,N_253);
nor U706 (N_706,N_166,N_367);
or U707 (N_707,N_47,N_468);
nor U708 (N_708,N_160,N_488);
nand U709 (N_709,N_393,N_480);
nor U710 (N_710,N_189,N_91);
nor U711 (N_711,N_261,N_66);
nand U712 (N_712,N_467,N_149);
nor U713 (N_713,N_28,N_182);
nand U714 (N_714,N_14,N_296);
and U715 (N_715,N_124,N_466);
xnor U716 (N_716,N_487,N_62);
nand U717 (N_717,N_33,N_25);
xor U718 (N_718,N_248,N_456);
or U719 (N_719,N_93,N_251);
and U720 (N_720,N_36,N_289);
xnor U721 (N_721,N_286,N_132);
nand U722 (N_722,N_222,N_4);
xor U723 (N_723,N_386,N_491);
nand U724 (N_724,N_140,N_285);
xor U725 (N_725,N_3,N_51);
or U726 (N_726,N_59,N_445);
nand U727 (N_727,N_203,N_191);
nor U728 (N_728,N_114,N_418);
nand U729 (N_729,N_437,N_374);
nor U730 (N_730,N_141,N_284);
nor U731 (N_731,N_436,N_165);
nor U732 (N_732,N_410,N_267);
nor U733 (N_733,N_0,N_462);
nand U734 (N_734,N_352,N_264);
nand U735 (N_735,N_100,N_414);
and U736 (N_736,N_339,N_276);
and U737 (N_737,N_302,N_177);
and U738 (N_738,N_450,N_406);
xnor U739 (N_739,N_299,N_27);
nor U740 (N_740,N_63,N_85);
nor U741 (N_741,N_360,N_417);
or U742 (N_742,N_243,N_122);
nor U743 (N_743,N_476,N_106);
nand U744 (N_744,N_143,N_224);
nor U745 (N_745,N_13,N_7);
and U746 (N_746,N_474,N_372);
and U747 (N_747,N_213,N_101);
or U748 (N_748,N_204,N_83);
or U749 (N_749,N_494,N_155);
nand U750 (N_750,N_218,N_301);
nor U751 (N_751,N_338,N_399);
nor U752 (N_752,N_340,N_497);
nand U753 (N_753,N_193,N_432);
xnor U754 (N_754,N_460,N_492);
xor U755 (N_755,N_401,N_414);
nand U756 (N_756,N_34,N_252);
or U757 (N_757,N_440,N_104);
xnor U758 (N_758,N_253,N_235);
nand U759 (N_759,N_148,N_314);
xnor U760 (N_760,N_491,N_59);
xnor U761 (N_761,N_332,N_16);
nor U762 (N_762,N_488,N_276);
nor U763 (N_763,N_341,N_249);
xor U764 (N_764,N_190,N_337);
and U765 (N_765,N_473,N_345);
nand U766 (N_766,N_43,N_454);
nand U767 (N_767,N_391,N_492);
or U768 (N_768,N_496,N_310);
and U769 (N_769,N_375,N_217);
xor U770 (N_770,N_305,N_310);
xnor U771 (N_771,N_363,N_347);
or U772 (N_772,N_18,N_90);
nor U773 (N_773,N_395,N_45);
xnor U774 (N_774,N_83,N_461);
or U775 (N_775,N_420,N_225);
or U776 (N_776,N_235,N_46);
xnor U777 (N_777,N_145,N_22);
or U778 (N_778,N_95,N_387);
nor U779 (N_779,N_6,N_9);
nand U780 (N_780,N_315,N_158);
and U781 (N_781,N_232,N_53);
nand U782 (N_782,N_50,N_452);
xnor U783 (N_783,N_346,N_94);
and U784 (N_784,N_220,N_309);
nand U785 (N_785,N_451,N_46);
nor U786 (N_786,N_451,N_56);
xor U787 (N_787,N_279,N_130);
xor U788 (N_788,N_216,N_386);
xor U789 (N_789,N_58,N_463);
and U790 (N_790,N_363,N_78);
nand U791 (N_791,N_306,N_458);
nand U792 (N_792,N_374,N_184);
or U793 (N_793,N_2,N_60);
xor U794 (N_794,N_221,N_400);
nand U795 (N_795,N_298,N_484);
nand U796 (N_796,N_324,N_360);
and U797 (N_797,N_358,N_8);
and U798 (N_798,N_217,N_220);
xor U799 (N_799,N_150,N_490);
xor U800 (N_800,N_278,N_149);
nand U801 (N_801,N_91,N_161);
nand U802 (N_802,N_264,N_143);
nor U803 (N_803,N_499,N_135);
nand U804 (N_804,N_329,N_346);
or U805 (N_805,N_148,N_333);
nand U806 (N_806,N_325,N_193);
or U807 (N_807,N_433,N_89);
nor U808 (N_808,N_295,N_226);
or U809 (N_809,N_255,N_212);
nand U810 (N_810,N_62,N_437);
and U811 (N_811,N_81,N_477);
nor U812 (N_812,N_120,N_157);
nor U813 (N_813,N_494,N_49);
and U814 (N_814,N_172,N_270);
and U815 (N_815,N_153,N_10);
xnor U816 (N_816,N_476,N_220);
or U817 (N_817,N_48,N_431);
nor U818 (N_818,N_199,N_15);
and U819 (N_819,N_361,N_380);
nand U820 (N_820,N_318,N_314);
nor U821 (N_821,N_410,N_26);
or U822 (N_822,N_169,N_430);
or U823 (N_823,N_315,N_178);
nor U824 (N_824,N_400,N_251);
and U825 (N_825,N_353,N_256);
nand U826 (N_826,N_263,N_255);
nand U827 (N_827,N_497,N_315);
or U828 (N_828,N_75,N_119);
nor U829 (N_829,N_328,N_241);
nand U830 (N_830,N_128,N_444);
or U831 (N_831,N_488,N_203);
and U832 (N_832,N_32,N_345);
and U833 (N_833,N_272,N_447);
nor U834 (N_834,N_140,N_474);
and U835 (N_835,N_210,N_105);
nand U836 (N_836,N_412,N_263);
nand U837 (N_837,N_124,N_191);
and U838 (N_838,N_258,N_36);
xnor U839 (N_839,N_30,N_3);
nand U840 (N_840,N_406,N_441);
and U841 (N_841,N_273,N_94);
and U842 (N_842,N_183,N_459);
or U843 (N_843,N_347,N_190);
or U844 (N_844,N_265,N_339);
nor U845 (N_845,N_323,N_69);
nand U846 (N_846,N_390,N_163);
xor U847 (N_847,N_392,N_98);
nor U848 (N_848,N_3,N_404);
and U849 (N_849,N_313,N_197);
nor U850 (N_850,N_354,N_266);
nand U851 (N_851,N_96,N_104);
xnor U852 (N_852,N_366,N_425);
nand U853 (N_853,N_271,N_456);
and U854 (N_854,N_268,N_12);
nor U855 (N_855,N_93,N_434);
xor U856 (N_856,N_353,N_345);
or U857 (N_857,N_349,N_272);
nand U858 (N_858,N_227,N_252);
or U859 (N_859,N_198,N_431);
xnor U860 (N_860,N_163,N_197);
and U861 (N_861,N_204,N_139);
nor U862 (N_862,N_40,N_60);
and U863 (N_863,N_168,N_346);
or U864 (N_864,N_313,N_52);
xnor U865 (N_865,N_362,N_344);
xnor U866 (N_866,N_429,N_146);
nor U867 (N_867,N_280,N_323);
and U868 (N_868,N_481,N_170);
or U869 (N_869,N_119,N_296);
and U870 (N_870,N_256,N_487);
nand U871 (N_871,N_453,N_409);
or U872 (N_872,N_36,N_17);
xnor U873 (N_873,N_108,N_57);
and U874 (N_874,N_304,N_432);
and U875 (N_875,N_382,N_456);
and U876 (N_876,N_37,N_402);
or U877 (N_877,N_420,N_65);
and U878 (N_878,N_427,N_296);
nor U879 (N_879,N_307,N_403);
or U880 (N_880,N_73,N_491);
xor U881 (N_881,N_346,N_462);
nor U882 (N_882,N_12,N_498);
xor U883 (N_883,N_228,N_274);
or U884 (N_884,N_55,N_200);
nand U885 (N_885,N_73,N_464);
or U886 (N_886,N_158,N_374);
and U887 (N_887,N_442,N_411);
nor U888 (N_888,N_222,N_458);
and U889 (N_889,N_263,N_266);
nor U890 (N_890,N_212,N_486);
nand U891 (N_891,N_178,N_44);
or U892 (N_892,N_375,N_238);
and U893 (N_893,N_495,N_190);
nand U894 (N_894,N_105,N_465);
xnor U895 (N_895,N_275,N_164);
xor U896 (N_896,N_285,N_221);
nand U897 (N_897,N_240,N_470);
xnor U898 (N_898,N_18,N_269);
and U899 (N_899,N_56,N_485);
nor U900 (N_900,N_408,N_329);
nand U901 (N_901,N_416,N_342);
xnor U902 (N_902,N_294,N_321);
or U903 (N_903,N_368,N_458);
nor U904 (N_904,N_115,N_402);
nand U905 (N_905,N_111,N_380);
or U906 (N_906,N_39,N_236);
nand U907 (N_907,N_126,N_360);
nand U908 (N_908,N_279,N_168);
and U909 (N_909,N_498,N_182);
nand U910 (N_910,N_314,N_170);
and U911 (N_911,N_56,N_105);
nor U912 (N_912,N_464,N_140);
or U913 (N_913,N_213,N_170);
nand U914 (N_914,N_337,N_158);
or U915 (N_915,N_195,N_495);
xor U916 (N_916,N_433,N_458);
nand U917 (N_917,N_399,N_73);
nand U918 (N_918,N_467,N_167);
and U919 (N_919,N_103,N_363);
xor U920 (N_920,N_5,N_197);
xor U921 (N_921,N_352,N_13);
nand U922 (N_922,N_431,N_381);
nand U923 (N_923,N_167,N_119);
xnor U924 (N_924,N_31,N_104);
and U925 (N_925,N_120,N_383);
and U926 (N_926,N_91,N_179);
or U927 (N_927,N_130,N_379);
nand U928 (N_928,N_132,N_428);
xnor U929 (N_929,N_401,N_447);
nor U930 (N_930,N_201,N_148);
nand U931 (N_931,N_173,N_67);
xor U932 (N_932,N_455,N_348);
and U933 (N_933,N_141,N_295);
nand U934 (N_934,N_478,N_43);
or U935 (N_935,N_496,N_364);
nand U936 (N_936,N_241,N_429);
nor U937 (N_937,N_490,N_144);
and U938 (N_938,N_442,N_445);
or U939 (N_939,N_423,N_358);
xor U940 (N_940,N_148,N_354);
nor U941 (N_941,N_312,N_435);
nor U942 (N_942,N_92,N_169);
or U943 (N_943,N_402,N_96);
xnor U944 (N_944,N_467,N_225);
nor U945 (N_945,N_56,N_67);
nand U946 (N_946,N_208,N_347);
nand U947 (N_947,N_154,N_137);
nand U948 (N_948,N_466,N_229);
nor U949 (N_949,N_170,N_464);
xnor U950 (N_950,N_96,N_12);
or U951 (N_951,N_99,N_398);
xnor U952 (N_952,N_280,N_380);
xor U953 (N_953,N_212,N_473);
or U954 (N_954,N_263,N_437);
xor U955 (N_955,N_366,N_73);
and U956 (N_956,N_4,N_34);
nor U957 (N_957,N_251,N_133);
or U958 (N_958,N_32,N_28);
and U959 (N_959,N_362,N_499);
xnor U960 (N_960,N_171,N_4);
and U961 (N_961,N_497,N_260);
nand U962 (N_962,N_161,N_210);
nand U963 (N_963,N_60,N_103);
xor U964 (N_964,N_183,N_190);
nor U965 (N_965,N_37,N_443);
nand U966 (N_966,N_315,N_486);
or U967 (N_967,N_222,N_413);
or U968 (N_968,N_321,N_393);
or U969 (N_969,N_297,N_351);
xor U970 (N_970,N_200,N_230);
and U971 (N_971,N_436,N_179);
nor U972 (N_972,N_345,N_84);
or U973 (N_973,N_353,N_312);
or U974 (N_974,N_52,N_338);
xnor U975 (N_975,N_284,N_222);
xnor U976 (N_976,N_37,N_170);
xnor U977 (N_977,N_240,N_310);
nor U978 (N_978,N_393,N_198);
or U979 (N_979,N_267,N_484);
or U980 (N_980,N_54,N_320);
nor U981 (N_981,N_17,N_182);
xnor U982 (N_982,N_258,N_473);
xnor U983 (N_983,N_309,N_424);
xor U984 (N_984,N_332,N_463);
nor U985 (N_985,N_164,N_132);
nor U986 (N_986,N_403,N_189);
and U987 (N_987,N_403,N_380);
nand U988 (N_988,N_160,N_78);
xnor U989 (N_989,N_332,N_150);
and U990 (N_990,N_160,N_135);
or U991 (N_991,N_437,N_396);
and U992 (N_992,N_446,N_83);
nor U993 (N_993,N_47,N_462);
nor U994 (N_994,N_261,N_423);
nand U995 (N_995,N_64,N_127);
nor U996 (N_996,N_337,N_137);
and U997 (N_997,N_290,N_36);
nand U998 (N_998,N_277,N_244);
and U999 (N_999,N_213,N_58);
xnor U1000 (N_1000,N_668,N_857);
xnor U1001 (N_1001,N_625,N_880);
nor U1002 (N_1002,N_643,N_995);
xor U1003 (N_1003,N_715,N_652);
xor U1004 (N_1004,N_861,N_934);
nor U1005 (N_1005,N_859,N_766);
nand U1006 (N_1006,N_521,N_554);
nand U1007 (N_1007,N_568,N_669);
or U1008 (N_1008,N_624,N_633);
nor U1009 (N_1009,N_908,N_732);
or U1010 (N_1010,N_751,N_680);
nand U1011 (N_1011,N_875,N_822);
xor U1012 (N_1012,N_761,N_639);
and U1013 (N_1013,N_737,N_983);
nand U1014 (N_1014,N_963,N_872);
and U1015 (N_1015,N_551,N_864);
nand U1016 (N_1016,N_539,N_956);
and U1017 (N_1017,N_515,N_973);
nor U1018 (N_1018,N_637,N_506);
nor U1019 (N_1019,N_722,N_758);
or U1020 (N_1020,N_712,N_999);
nor U1021 (N_1021,N_505,N_666);
nor U1022 (N_1022,N_776,N_667);
or U1023 (N_1023,N_977,N_882);
nor U1024 (N_1024,N_940,N_721);
or U1025 (N_1025,N_501,N_985);
nor U1026 (N_1026,N_904,N_553);
nor U1027 (N_1027,N_965,N_949);
nand U1028 (N_1028,N_524,N_964);
or U1029 (N_1029,N_707,N_797);
nand U1030 (N_1030,N_723,N_510);
nor U1031 (N_1031,N_783,N_961);
or U1032 (N_1032,N_803,N_762);
nor U1033 (N_1033,N_610,N_815);
nor U1034 (N_1034,N_926,N_763);
xor U1035 (N_1035,N_583,N_552);
or U1036 (N_1036,N_688,N_805);
and U1037 (N_1037,N_559,N_991);
xor U1038 (N_1038,N_795,N_578);
or U1039 (N_1039,N_976,N_544);
nand U1040 (N_1040,N_513,N_874);
and U1041 (N_1041,N_546,N_791);
and U1042 (N_1042,N_945,N_811);
or U1043 (N_1043,N_603,N_519);
and U1044 (N_1044,N_567,N_591);
nand U1045 (N_1045,N_614,N_627);
nor U1046 (N_1046,N_767,N_612);
or U1047 (N_1047,N_787,N_598);
nor U1048 (N_1048,N_745,N_818);
xnor U1049 (N_1049,N_773,N_717);
xnor U1050 (N_1050,N_938,N_593);
nand U1051 (N_1051,N_935,N_529);
nand U1052 (N_1052,N_611,N_532);
or U1053 (N_1053,N_768,N_570);
nand U1054 (N_1054,N_565,N_631);
nor U1055 (N_1055,N_786,N_996);
nor U1056 (N_1056,N_670,N_747);
and U1057 (N_1057,N_760,N_871);
nor U1058 (N_1058,N_947,N_974);
nand U1059 (N_1059,N_993,N_933);
nand U1060 (N_1060,N_847,N_750);
and U1061 (N_1061,N_527,N_500);
or U1062 (N_1062,N_809,N_700);
xnor U1063 (N_1063,N_780,N_792);
or U1064 (N_1064,N_957,N_915);
nand U1065 (N_1065,N_692,N_769);
nor U1066 (N_1066,N_869,N_579);
nor U1067 (N_1067,N_699,N_672);
nor U1068 (N_1068,N_924,N_946);
nor U1069 (N_1069,N_619,N_648);
xor U1070 (N_1070,N_753,N_657);
nand U1071 (N_1071,N_581,N_748);
xor U1072 (N_1072,N_560,N_897);
nor U1073 (N_1073,N_623,N_903);
or U1074 (N_1074,N_647,N_588);
nor U1075 (N_1075,N_816,N_833);
and U1076 (N_1076,N_960,N_734);
or U1077 (N_1077,N_548,N_609);
nor U1078 (N_1078,N_731,N_728);
nand U1079 (N_1079,N_689,N_621);
or U1080 (N_1080,N_817,N_952);
xor U1081 (N_1081,N_577,N_914);
xnor U1082 (N_1082,N_726,N_879);
xnor U1083 (N_1083,N_858,N_981);
and U1084 (N_1084,N_895,N_909);
or U1085 (N_1085,N_646,N_517);
or U1086 (N_1086,N_906,N_573);
and U1087 (N_1087,N_622,N_912);
xor U1088 (N_1088,N_542,N_899);
and U1089 (N_1089,N_825,N_704);
nand U1090 (N_1090,N_739,N_572);
nand U1091 (N_1091,N_971,N_536);
xnor U1092 (N_1092,N_642,N_812);
and U1093 (N_1093,N_932,N_777);
or U1094 (N_1094,N_804,N_574);
nand U1095 (N_1095,N_867,N_713);
or U1096 (N_1096,N_820,N_606);
and U1097 (N_1097,N_929,N_526);
nor U1098 (N_1098,N_679,N_853);
nor U1099 (N_1099,N_562,N_590);
nand U1100 (N_1100,N_547,N_535);
nand U1101 (N_1101,N_978,N_881);
or U1102 (N_1102,N_873,N_520);
xnor U1103 (N_1103,N_785,N_814);
or U1104 (N_1104,N_665,N_675);
nor U1105 (N_1105,N_921,N_752);
and U1106 (N_1106,N_595,N_866);
xnor U1107 (N_1107,N_617,N_892);
and U1108 (N_1108,N_564,N_923);
xnor U1109 (N_1109,N_930,N_555);
nand U1110 (N_1110,N_703,N_658);
and U1111 (N_1111,N_898,N_917);
nand U1112 (N_1112,N_741,N_759);
nor U1113 (N_1113,N_522,N_905);
and U1114 (N_1114,N_835,N_528);
and U1115 (N_1115,N_708,N_735);
nor U1116 (N_1116,N_994,N_685);
and U1117 (N_1117,N_860,N_876);
xor U1118 (N_1118,N_798,N_813);
nor U1119 (N_1119,N_629,N_808);
and U1120 (N_1120,N_509,N_620);
and U1121 (N_1121,N_770,N_671);
nor U1122 (N_1122,N_788,N_877);
nand U1123 (N_1123,N_523,N_702);
xnor U1124 (N_1124,N_807,N_677);
xor U1125 (N_1125,N_749,N_635);
nor U1126 (N_1126,N_508,N_782);
nor U1127 (N_1127,N_587,N_774);
nor U1128 (N_1128,N_634,N_885);
xnor U1129 (N_1129,N_594,N_569);
nand U1130 (N_1130,N_775,N_684);
nand U1131 (N_1131,N_829,N_796);
nand U1132 (N_1132,N_800,N_602);
nand U1133 (N_1133,N_931,N_799);
xor U1134 (N_1134,N_705,N_980);
nor U1135 (N_1135,N_695,N_984);
xor U1136 (N_1136,N_706,N_831);
nand U1137 (N_1137,N_756,N_742);
and U1138 (N_1138,N_846,N_533);
and U1139 (N_1139,N_663,N_597);
or U1140 (N_1140,N_541,N_969);
xnor U1141 (N_1141,N_887,N_902);
nand U1142 (N_1142,N_661,N_640);
nand U1143 (N_1143,N_806,N_607);
nand U1144 (N_1144,N_870,N_514);
nor U1145 (N_1145,N_557,N_918);
xnor U1146 (N_1146,N_836,N_709);
or U1147 (N_1147,N_538,N_950);
xnor U1148 (N_1148,N_693,N_919);
nor U1149 (N_1149,N_589,N_615);
and U1150 (N_1150,N_990,N_710);
or U1151 (N_1151,N_504,N_848);
nor U1152 (N_1152,N_948,N_525);
nor U1153 (N_1153,N_596,N_678);
nand U1154 (N_1154,N_600,N_936);
xnor U1155 (N_1155,N_608,N_937);
xor U1156 (N_1156,N_862,N_841);
nor U1157 (N_1157,N_613,N_585);
xor U1158 (N_1158,N_545,N_540);
nand U1159 (N_1159,N_698,N_828);
xor U1160 (N_1160,N_802,N_910);
and U1161 (N_1161,N_823,N_718);
and U1162 (N_1162,N_660,N_863);
and U1163 (N_1163,N_743,N_824);
and U1164 (N_1164,N_778,N_771);
nand U1165 (N_1165,N_674,N_503);
nand U1166 (N_1166,N_911,N_730);
nor U1167 (N_1167,N_781,N_975);
and U1168 (N_1168,N_832,N_972);
nand U1169 (N_1169,N_865,N_507);
nand U1170 (N_1170,N_764,N_638);
nand U1171 (N_1171,N_605,N_694);
xnor U1172 (N_1172,N_959,N_890);
or U1173 (N_1173,N_714,N_900);
xnor U1174 (N_1174,N_821,N_951);
nand U1175 (N_1175,N_687,N_746);
nor U1176 (N_1176,N_650,N_954);
and U1177 (N_1177,N_645,N_883);
nand U1178 (N_1178,N_916,N_896);
nor U1179 (N_1179,N_691,N_592);
nor U1180 (N_1180,N_894,N_556);
nand U1181 (N_1181,N_928,N_837);
nand U1182 (N_1182,N_989,N_654);
xor U1183 (N_1183,N_659,N_582);
and U1184 (N_1184,N_801,N_537);
xor U1185 (N_1185,N_966,N_901);
nand U1186 (N_1186,N_849,N_922);
xor U1187 (N_1187,N_843,N_913);
and U1188 (N_1188,N_686,N_601);
nor U1189 (N_1189,N_757,N_834);
nand U1190 (N_1190,N_852,N_632);
xor U1191 (N_1191,N_744,N_868);
nand U1192 (N_1192,N_839,N_530);
and U1193 (N_1193,N_676,N_827);
and U1194 (N_1194,N_793,N_855);
nand U1195 (N_1195,N_907,N_844);
or U1196 (N_1196,N_673,N_939);
xnor U1197 (N_1197,N_740,N_580);
and U1198 (N_1198,N_719,N_518);
nand U1199 (N_1199,N_830,N_958);
or U1200 (N_1200,N_779,N_772);
nand U1201 (N_1201,N_696,N_571);
or U1202 (N_1202,N_878,N_851);
xnor U1203 (N_1203,N_644,N_549);
and U1204 (N_1204,N_738,N_511);
nor U1205 (N_1205,N_998,N_641);
xnor U1206 (N_1206,N_943,N_986);
xnor U1207 (N_1207,N_531,N_988);
or U1208 (N_1208,N_604,N_558);
nor U1209 (N_1209,N_736,N_599);
nor U1210 (N_1210,N_810,N_955);
and U1211 (N_1211,N_941,N_826);
nand U1212 (N_1212,N_664,N_701);
nor U1213 (N_1213,N_886,N_789);
nand U1214 (N_1214,N_856,N_566);
nand U1215 (N_1215,N_725,N_819);
and U1216 (N_1216,N_845,N_794);
and U1217 (N_1217,N_655,N_720);
nor U1218 (N_1218,N_724,N_512);
xor U1219 (N_1219,N_784,N_618);
or U1220 (N_1220,N_682,N_891);
nand U1221 (N_1221,N_683,N_982);
and U1222 (N_1222,N_711,N_649);
xnor U1223 (N_1223,N_962,N_561);
nand U1224 (N_1224,N_888,N_628);
xnor U1225 (N_1225,N_651,N_729);
nor U1226 (N_1226,N_942,N_626);
xnor U1227 (N_1227,N_681,N_979);
nor U1228 (N_1228,N_754,N_584);
nor U1229 (N_1229,N_987,N_889);
nand U1230 (N_1230,N_884,N_576);
or U1231 (N_1231,N_690,N_838);
nand U1232 (N_1232,N_944,N_765);
nor U1233 (N_1233,N_697,N_970);
xor U1234 (N_1234,N_534,N_997);
xor U1235 (N_1235,N_850,N_840);
nand U1236 (N_1236,N_755,N_586);
nand U1237 (N_1237,N_854,N_543);
and U1238 (N_1238,N_516,N_636);
nor U1239 (N_1239,N_630,N_563);
nand U1240 (N_1240,N_927,N_992);
nor U1241 (N_1241,N_716,N_653);
xnor U1242 (N_1242,N_893,N_656);
and U1243 (N_1243,N_616,N_925);
xor U1244 (N_1244,N_953,N_575);
or U1245 (N_1245,N_968,N_733);
nor U1246 (N_1246,N_967,N_727);
nand U1247 (N_1247,N_662,N_790);
and U1248 (N_1248,N_502,N_842);
and U1249 (N_1249,N_550,N_920);
or U1250 (N_1250,N_682,N_674);
or U1251 (N_1251,N_639,N_621);
nor U1252 (N_1252,N_933,N_578);
or U1253 (N_1253,N_652,N_552);
and U1254 (N_1254,N_704,N_539);
xnor U1255 (N_1255,N_662,N_795);
nand U1256 (N_1256,N_639,N_869);
xnor U1257 (N_1257,N_740,N_564);
nor U1258 (N_1258,N_541,N_576);
xor U1259 (N_1259,N_541,N_772);
nand U1260 (N_1260,N_735,N_531);
nand U1261 (N_1261,N_904,N_549);
nand U1262 (N_1262,N_898,N_859);
nand U1263 (N_1263,N_828,N_540);
nor U1264 (N_1264,N_875,N_952);
nor U1265 (N_1265,N_892,N_721);
xnor U1266 (N_1266,N_597,N_683);
nor U1267 (N_1267,N_828,N_666);
and U1268 (N_1268,N_805,N_691);
nor U1269 (N_1269,N_696,N_546);
and U1270 (N_1270,N_760,N_999);
or U1271 (N_1271,N_991,N_935);
xor U1272 (N_1272,N_733,N_673);
xor U1273 (N_1273,N_851,N_751);
xor U1274 (N_1274,N_598,N_518);
and U1275 (N_1275,N_500,N_760);
or U1276 (N_1276,N_831,N_862);
xnor U1277 (N_1277,N_762,N_593);
xor U1278 (N_1278,N_519,N_676);
nand U1279 (N_1279,N_657,N_668);
nand U1280 (N_1280,N_856,N_907);
and U1281 (N_1281,N_570,N_556);
or U1282 (N_1282,N_882,N_577);
xor U1283 (N_1283,N_819,N_945);
nand U1284 (N_1284,N_990,N_676);
nor U1285 (N_1285,N_950,N_792);
xor U1286 (N_1286,N_705,N_593);
xnor U1287 (N_1287,N_620,N_991);
xnor U1288 (N_1288,N_789,N_607);
or U1289 (N_1289,N_733,N_634);
and U1290 (N_1290,N_818,N_750);
nand U1291 (N_1291,N_886,N_876);
or U1292 (N_1292,N_904,N_893);
xor U1293 (N_1293,N_850,N_816);
xor U1294 (N_1294,N_606,N_912);
nor U1295 (N_1295,N_764,N_538);
or U1296 (N_1296,N_798,N_551);
xor U1297 (N_1297,N_626,N_885);
nor U1298 (N_1298,N_946,N_527);
nor U1299 (N_1299,N_646,N_698);
nor U1300 (N_1300,N_943,N_717);
or U1301 (N_1301,N_616,N_624);
nand U1302 (N_1302,N_785,N_624);
or U1303 (N_1303,N_618,N_880);
xnor U1304 (N_1304,N_695,N_909);
nand U1305 (N_1305,N_780,N_890);
nor U1306 (N_1306,N_869,N_647);
xor U1307 (N_1307,N_629,N_855);
or U1308 (N_1308,N_643,N_910);
nor U1309 (N_1309,N_709,N_726);
nand U1310 (N_1310,N_958,N_926);
nand U1311 (N_1311,N_686,N_872);
nand U1312 (N_1312,N_618,N_764);
or U1313 (N_1313,N_928,N_617);
nand U1314 (N_1314,N_975,N_575);
and U1315 (N_1315,N_676,N_603);
nor U1316 (N_1316,N_513,N_843);
nor U1317 (N_1317,N_619,N_514);
and U1318 (N_1318,N_766,N_823);
xnor U1319 (N_1319,N_595,N_810);
nor U1320 (N_1320,N_604,N_742);
or U1321 (N_1321,N_722,N_518);
nor U1322 (N_1322,N_821,N_524);
and U1323 (N_1323,N_712,N_920);
xnor U1324 (N_1324,N_744,N_957);
nor U1325 (N_1325,N_631,N_907);
or U1326 (N_1326,N_529,N_713);
nor U1327 (N_1327,N_567,N_794);
and U1328 (N_1328,N_572,N_875);
xnor U1329 (N_1329,N_513,N_927);
or U1330 (N_1330,N_836,N_529);
xor U1331 (N_1331,N_669,N_851);
xor U1332 (N_1332,N_803,N_511);
nor U1333 (N_1333,N_519,N_691);
or U1334 (N_1334,N_548,N_592);
nand U1335 (N_1335,N_884,N_504);
xnor U1336 (N_1336,N_889,N_999);
and U1337 (N_1337,N_740,N_920);
nor U1338 (N_1338,N_733,N_686);
and U1339 (N_1339,N_995,N_785);
nor U1340 (N_1340,N_750,N_799);
xor U1341 (N_1341,N_723,N_558);
nand U1342 (N_1342,N_696,N_848);
and U1343 (N_1343,N_981,N_861);
or U1344 (N_1344,N_940,N_502);
xnor U1345 (N_1345,N_804,N_769);
and U1346 (N_1346,N_680,N_896);
nand U1347 (N_1347,N_779,N_599);
xnor U1348 (N_1348,N_619,N_546);
or U1349 (N_1349,N_549,N_794);
and U1350 (N_1350,N_648,N_988);
nand U1351 (N_1351,N_798,N_760);
nand U1352 (N_1352,N_890,N_569);
or U1353 (N_1353,N_906,N_804);
and U1354 (N_1354,N_602,N_603);
nand U1355 (N_1355,N_997,N_757);
nand U1356 (N_1356,N_767,N_820);
or U1357 (N_1357,N_761,N_891);
and U1358 (N_1358,N_750,N_704);
xor U1359 (N_1359,N_918,N_780);
nor U1360 (N_1360,N_800,N_517);
nand U1361 (N_1361,N_872,N_924);
or U1362 (N_1362,N_692,N_884);
nor U1363 (N_1363,N_659,N_899);
or U1364 (N_1364,N_909,N_997);
and U1365 (N_1365,N_845,N_738);
or U1366 (N_1366,N_737,N_734);
xor U1367 (N_1367,N_700,N_899);
nand U1368 (N_1368,N_866,N_845);
and U1369 (N_1369,N_736,N_605);
or U1370 (N_1370,N_782,N_701);
nand U1371 (N_1371,N_932,N_521);
xor U1372 (N_1372,N_721,N_784);
or U1373 (N_1373,N_601,N_643);
nor U1374 (N_1374,N_826,N_871);
or U1375 (N_1375,N_586,N_886);
nor U1376 (N_1376,N_775,N_686);
nor U1377 (N_1377,N_576,N_944);
and U1378 (N_1378,N_827,N_744);
or U1379 (N_1379,N_569,N_593);
or U1380 (N_1380,N_740,N_602);
nand U1381 (N_1381,N_727,N_985);
and U1382 (N_1382,N_645,N_698);
nor U1383 (N_1383,N_586,N_539);
nand U1384 (N_1384,N_608,N_713);
nand U1385 (N_1385,N_796,N_743);
nor U1386 (N_1386,N_550,N_744);
nand U1387 (N_1387,N_882,N_746);
nor U1388 (N_1388,N_793,N_542);
nor U1389 (N_1389,N_985,N_986);
nor U1390 (N_1390,N_908,N_789);
and U1391 (N_1391,N_853,N_894);
nor U1392 (N_1392,N_624,N_552);
and U1393 (N_1393,N_916,N_962);
nor U1394 (N_1394,N_957,N_952);
nor U1395 (N_1395,N_717,N_723);
or U1396 (N_1396,N_830,N_998);
xnor U1397 (N_1397,N_857,N_916);
or U1398 (N_1398,N_588,N_661);
nand U1399 (N_1399,N_841,N_653);
or U1400 (N_1400,N_609,N_567);
nand U1401 (N_1401,N_833,N_893);
nor U1402 (N_1402,N_981,N_562);
nand U1403 (N_1403,N_673,N_959);
nand U1404 (N_1404,N_955,N_870);
xor U1405 (N_1405,N_587,N_728);
and U1406 (N_1406,N_830,N_963);
nor U1407 (N_1407,N_725,N_985);
xnor U1408 (N_1408,N_632,N_729);
xnor U1409 (N_1409,N_581,N_784);
xnor U1410 (N_1410,N_636,N_776);
or U1411 (N_1411,N_912,N_567);
and U1412 (N_1412,N_680,N_809);
or U1413 (N_1413,N_654,N_641);
nand U1414 (N_1414,N_650,N_927);
nand U1415 (N_1415,N_503,N_875);
nand U1416 (N_1416,N_685,N_953);
and U1417 (N_1417,N_699,N_670);
or U1418 (N_1418,N_564,N_665);
xnor U1419 (N_1419,N_730,N_891);
xor U1420 (N_1420,N_521,N_600);
and U1421 (N_1421,N_839,N_866);
nand U1422 (N_1422,N_712,N_559);
xnor U1423 (N_1423,N_989,N_813);
xor U1424 (N_1424,N_844,N_737);
or U1425 (N_1425,N_640,N_826);
nor U1426 (N_1426,N_754,N_685);
nand U1427 (N_1427,N_625,N_729);
or U1428 (N_1428,N_900,N_794);
nand U1429 (N_1429,N_996,N_676);
nor U1430 (N_1430,N_735,N_576);
xnor U1431 (N_1431,N_777,N_902);
and U1432 (N_1432,N_697,N_854);
and U1433 (N_1433,N_929,N_530);
and U1434 (N_1434,N_744,N_848);
nand U1435 (N_1435,N_764,N_619);
nand U1436 (N_1436,N_655,N_565);
and U1437 (N_1437,N_780,N_810);
and U1438 (N_1438,N_953,N_771);
nand U1439 (N_1439,N_826,N_720);
nand U1440 (N_1440,N_625,N_602);
and U1441 (N_1441,N_799,N_629);
nor U1442 (N_1442,N_850,N_717);
or U1443 (N_1443,N_645,N_639);
and U1444 (N_1444,N_701,N_968);
xnor U1445 (N_1445,N_723,N_851);
and U1446 (N_1446,N_648,N_609);
or U1447 (N_1447,N_975,N_908);
xor U1448 (N_1448,N_607,N_954);
or U1449 (N_1449,N_871,N_856);
and U1450 (N_1450,N_644,N_581);
or U1451 (N_1451,N_845,N_581);
and U1452 (N_1452,N_970,N_838);
and U1453 (N_1453,N_706,N_597);
xnor U1454 (N_1454,N_774,N_662);
nand U1455 (N_1455,N_873,N_986);
nor U1456 (N_1456,N_599,N_692);
or U1457 (N_1457,N_819,N_993);
and U1458 (N_1458,N_541,N_737);
xor U1459 (N_1459,N_800,N_705);
or U1460 (N_1460,N_743,N_546);
nand U1461 (N_1461,N_984,N_567);
and U1462 (N_1462,N_609,N_809);
xor U1463 (N_1463,N_791,N_966);
xor U1464 (N_1464,N_675,N_803);
and U1465 (N_1465,N_795,N_732);
nand U1466 (N_1466,N_710,N_500);
nand U1467 (N_1467,N_737,N_701);
nor U1468 (N_1468,N_662,N_793);
nor U1469 (N_1469,N_918,N_715);
nand U1470 (N_1470,N_938,N_880);
and U1471 (N_1471,N_703,N_928);
and U1472 (N_1472,N_733,N_660);
nor U1473 (N_1473,N_517,N_806);
xor U1474 (N_1474,N_566,N_894);
and U1475 (N_1475,N_926,N_753);
nor U1476 (N_1476,N_913,N_980);
xor U1477 (N_1477,N_895,N_960);
or U1478 (N_1478,N_580,N_565);
nor U1479 (N_1479,N_813,N_740);
nor U1480 (N_1480,N_798,N_660);
nor U1481 (N_1481,N_740,N_609);
nand U1482 (N_1482,N_863,N_847);
nand U1483 (N_1483,N_604,N_994);
or U1484 (N_1484,N_961,N_865);
nand U1485 (N_1485,N_806,N_546);
nand U1486 (N_1486,N_817,N_847);
and U1487 (N_1487,N_940,N_501);
and U1488 (N_1488,N_979,N_618);
nor U1489 (N_1489,N_920,N_590);
and U1490 (N_1490,N_509,N_604);
nor U1491 (N_1491,N_920,N_900);
nand U1492 (N_1492,N_556,N_751);
or U1493 (N_1493,N_703,N_619);
or U1494 (N_1494,N_546,N_652);
nor U1495 (N_1495,N_783,N_941);
and U1496 (N_1496,N_707,N_660);
and U1497 (N_1497,N_736,N_904);
or U1498 (N_1498,N_794,N_832);
nor U1499 (N_1499,N_973,N_661);
xor U1500 (N_1500,N_1337,N_1100);
nand U1501 (N_1501,N_1368,N_1469);
nor U1502 (N_1502,N_1470,N_1431);
nand U1503 (N_1503,N_1082,N_1244);
xor U1504 (N_1504,N_1018,N_1375);
nor U1505 (N_1505,N_1365,N_1027);
nand U1506 (N_1506,N_1467,N_1250);
nor U1507 (N_1507,N_1045,N_1150);
xor U1508 (N_1508,N_1141,N_1424);
nand U1509 (N_1509,N_1489,N_1090);
nor U1510 (N_1510,N_1483,N_1355);
nand U1511 (N_1511,N_1227,N_1190);
and U1512 (N_1512,N_1006,N_1019);
nand U1513 (N_1513,N_1387,N_1130);
or U1514 (N_1514,N_1005,N_1218);
nor U1515 (N_1515,N_1322,N_1290);
xor U1516 (N_1516,N_1443,N_1129);
or U1517 (N_1517,N_1468,N_1243);
or U1518 (N_1518,N_1157,N_1374);
nor U1519 (N_1519,N_1184,N_1125);
or U1520 (N_1520,N_1025,N_1034);
or U1521 (N_1521,N_1095,N_1418);
and U1522 (N_1522,N_1167,N_1340);
and U1523 (N_1523,N_1474,N_1354);
nand U1524 (N_1524,N_1203,N_1239);
or U1525 (N_1525,N_1384,N_1316);
xor U1526 (N_1526,N_1358,N_1098);
nand U1527 (N_1527,N_1292,N_1388);
xnor U1528 (N_1528,N_1484,N_1212);
nor U1529 (N_1529,N_1260,N_1194);
and U1530 (N_1530,N_1080,N_1459);
xnor U1531 (N_1531,N_1229,N_1170);
and U1532 (N_1532,N_1366,N_1158);
nand U1533 (N_1533,N_1155,N_1007);
nor U1534 (N_1534,N_1056,N_1140);
and U1535 (N_1535,N_1023,N_1178);
nand U1536 (N_1536,N_1187,N_1196);
nor U1537 (N_1537,N_1348,N_1153);
or U1538 (N_1538,N_1179,N_1268);
or U1539 (N_1539,N_1057,N_1495);
or U1540 (N_1540,N_1273,N_1144);
nand U1541 (N_1541,N_1121,N_1165);
xor U1542 (N_1542,N_1498,N_1116);
nor U1543 (N_1543,N_1325,N_1482);
nand U1544 (N_1544,N_1436,N_1142);
xnor U1545 (N_1545,N_1181,N_1208);
nand U1546 (N_1546,N_1259,N_1289);
and U1547 (N_1547,N_1377,N_1298);
nand U1548 (N_1548,N_1312,N_1457);
xor U1549 (N_1549,N_1438,N_1075);
or U1550 (N_1550,N_1405,N_1283);
and U1551 (N_1551,N_1039,N_1177);
nand U1552 (N_1552,N_1462,N_1256);
nand U1553 (N_1553,N_1126,N_1058);
and U1554 (N_1554,N_1303,N_1067);
nand U1555 (N_1555,N_1323,N_1456);
xor U1556 (N_1556,N_1373,N_1055);
nor U1557 (N_1557,N_1171,N_1064);
xnor U1558 (N_1558,N_1106,N_1411);
or U1559 (N_1559,N_1347,N_1416);
nand U1560 (N_1560,N_1395,N_1291);
and U1561 (N_1561,N_1162,N_1475);
xnor U1562 (N_1562,N_1240,N_1371);
xor U1563 (N_1563,N_1216,N_1101);
nor U1564 (N_1564,N_1205,N_1231);
nand U1565 (N_1565,N_1399,N_1321);
or U1566 (N_1566,N_1254,N_1186);
and U1567 (N_1567,N_1004,N_1147);
nor U1568 (N_1568,N_1015,N_1441);
nand U1569 (N_1569,N_1339,N_1285);
nand U1570 (N_1570,N_1085,N_1050);
nand U1571 (N_1571,N_1040,N_1401);
nand U1572 (N_1572,N_1282,N_1145);
xor U1573 (N_1573,N_1136,N_1473);
and U1574 (N_1574,N_1253,N_1191);
or U1575 (N_1575,N_1343,N_1406);
or U1576 (N_1576,N_1234,N_1241);
xor U1577 (N_1577,N_1331,N_1204);
nor U1578 (N_1578,N_1275,N_1166);
nor U1579 (N_1579,N_1264,N_1262);
xnor U1580 (N_1580,N_1396,N_1041);
nor U1581 (N_1581,N_1326,N_1103);
xnor U1582 (N_1582,N_1003,N_1120);
nor U1583 (N_1583,N_1242,N_1011);
xnor U1584 (N_1584,N_1478,N_1486);
and U1585 (N_1585,N_1028,N_1219);
and U1586 (N_1586,N_1132,N_1112);
nor U1587 (N_1587,N_1369,N_1074);
nor U1588 (N_1588,N_1367,N_1161);
nor U1589 (N_1589,N_1214,N_1012);
nand U1590 (N_1590,N_1393,N_1414);
xnor U1591 (N_1591,N_1193,N_1213);
nand U1592 (N_1592,N_1359,N_1247);
nor U1593 (N_1593,N_1288,N_1420);
and U1594 (N_1594,N_1432,N_1378);
nand U1595 (N_1595,N_1134,N_1296);
or U1596 (N_1596,N_1311,N_1345);
nand U1597 (N_1597,N_1448,N_1445);
or U1598 (N_1598,N_1118,N_1385);
or U1599 (N_1599,N_1381,N_1328);
xor U1600 (N_1600,N_1046,N_1222);
or U1601 (N_1601,N_1463,N_1391);
or U1602 (N_1602,N_1175,N_1002);
xnor U1603 (N_1603,N_1089,N_1376);
nand U1604 (N_1604,N_1033,N_1008);
nor U1605 (N_1605,N_1038,N_1278);
nand U1606 (N_1606,N_1454,N_1070);
or U1607 (N_1607,N_1138,N_1274);
and U1608 (N_1608,N_1245,N_1319);
nand U1609 (N_1609,N_1295,N_1429);
or U1610 (N_1610,N_1284,N_1320);
and U1611 (N_1611,N_1096,N_1048);
nand U1612 (N_1612,N_1077,N_1010);
nand U1613 (N_1613,N_1447,N_1065);
or U1614 (N_1614,N_1020,N_1297);
nand U1615 (N_1615,N_1412,N_1269);
nand U1616 (N_1616,N_1476,N_1225);
xnor U1617 (N_1617,N_1172,N_1160);
nand U1618 (N_1618,N_1341,N_1188);
and U1619 (N_1619,N_1499,N_1472);
or U1620 (N_1620,N_1014,N_1332);
or U1621 (N_1621,N_1455,N_1465);
and U1622 (N_1622,N_1163,N_1249);
nand U1623 (N_1623,N_1361,N_1380);
nand U1624 (N_1624,N_1437,N_1049);
nor U1625 (N_1625,N_1054,N_1016);
nand U1626 (N_1626,N_1185,N_1183);
and U1627 (N_1627,N_1081,N_1021);
or U1628 (N_1628,N_1350,N_1494);
nor U1629 (N_1629,N_1117,N_1353);
nor U1630 (N_1630,N_1428,N_1092);
or U1631 (N_1631,N_1257,N_1449);
nand U1632 (N_1632,N_1107,N_1270);
nand U1633 (N_1633,N_1230,N_1265);
xor U1634 (N_1634,N_1304,N_1061);
xor U1635 (N_1635,N_1079,N_1306);
xor U1636 (N_1636,N_1037,N_1444);
and U1637 (N_1637,N_1279,N_1154);
nor U1638 (N_1638,N_1430,N_1488);
xnor U1639 (N_1639,N_1029,N_1001);
or U1640 (N_1640,N_1330,N_1176);
nand U1641 (N_1641,N_1422,N_1071);
nand U1642 (N_1642,N_1315,N_1093);
xnor U1643 (N_1643,N_1143,N_1417);
or U1644 (N_1644,N_1392,N_1210);
and U1645 (N_1645,N_1228,N_1127);
nand U1646 (N_1646,N_1199,N_1419);
or U1647 (N_1647,N_1258,N_1173);
and U1648 (N_1648,N_1281,N_1440);
nor U1649 (N_1649,N_1073,N_1099);
or U1650 (N_1650,N_1485,N_1197);
xor U1651 (N_1651,N_1232,N_1174);
nor U1652 (N_1652,N_1314,N_1156);
or U1653 (N_1653,N_1386,N_1083);
xnor U1654 (N_1654,N_1479,N_1063);
nand U1655 (N_1655,N_1481,N_1492);
nand U1656 (N_1656,N_1301,N_1336);
nor U1657 (N_1657,N_1047,N_1464);
nor U1658 (N_1658,N_1017,N_1195);
or U1659 (N_1659,N_1403,N_1491);
xor U1660 (N_1660,N_1097,N_1349);
and U1661 (N_1661,N_1035,N_1105);
xnor U1662 (N_1662,N_1490,N_1206);
nand U1663 (N_1663,N_1372,N_1182);
nand U1664 (N_1664,N_1069,N_1094);
nand U1665 (N_1665,N_1442,N_1110);
or U1666 (N_1666,N_1276,N_1066);
nor U1667 (N_1667,N_1223,N_1072);
or U1668 (N_1668,N_1453,N_1329);
and U1669 (N_1669,N_1450,N_1458);
nand U1670 (N_1670,N_1271,N_1200);
nand U1671 (N_1671,N_1159,N_1334);
nor U1672 (N_1672,N_1086,N_1043);
or U1673 (N_1673,N_1272,N_1266);
nor U1674 (N_1674,N_1133,N_1032);
nor U1675 (N_1675,N_1169,N_1333);
nor U1676 (N_1676,N_1201,N_1124);
and U1677 (N_1677,N_1435,N_1324);
nand U1678 (N_1678,N_1139,N_1287);
xnor U1679 (N_1679,N_1137,N_1310);
nand U1680 (N_1680,N_1415,N_1477);
and U1681 (N_1681,N_1233,N_1076);
xor U1682 (N_1682,N_1398,N_1180);
nand U1683 (N_1683,N_1421,N_1426);
or U1684 (N_1684,N_1427,N_1211);
nor U1685 (N_1685,N_1389,N_1168);
xnor U1686 (N_1686,N_1044,N_1031);
xor U1687 (N_1687,N_1215,N_1087);
xnor U1688 (N_1688,N_1446,N_1255);
and U1689 (N_1689,N_1237,N_1383);
nor U1690 (N_1690,N_1496,N_1313);
and U1691 (N_1691,N_1026,N_1164);
or U1692 (N_1692,N_1379,N_1471);
nor U1693 (N_1693,N_1293,N_1198);
or U1694 (N_1694,N_1246,N_1400);
nand U1695 (N_1695,N_1084,N_1305);
xnor U1696 (N_1696,N_1407,N_1277);
nand U1697 (N_1697,N_1115,N_1413);
xor U1698 (N_1698,N_1238,N_1308);
nand U1699 (N_1699,N_1036,N_1261);
or U1700 (N_1700,N_1434,N_1360);
and U1701 (N_1701,N_1362,N_1327);
and U1702 (N_1702,N_1480,N_1235);
xnor U1703 (N_1703,N_1409,N_1226);
and U1704 (N_1704,N_1382,N_1122);
and U1705 (N_1705,N_1135,N_1408);
xor U1706 (N_1706,N_1338,N_1356);
or U1707 (N_1707,N_1013,N_1466);
nor U1708 (N_1708,N_1299,N_1113);
xnor U1709 (N_1709,N_1030,N_1433);
or U1710 (N_1710,N_1451,N_1335);
and U1711 (N_1711,N_1280,N_1059);
and U1712 (N_1712,N_1051,N_1423);
nor U1713 (N_1713,N_1146,N_1397);
xor U1714 (N_1714,N_1425,N_1220);
nor U1715 (N_1715,N_1221,N_1439);
nor U1716 (N_1716,N_1152,N_1307);
nand U1717 (N_1717,N_1052,N_1394);
and U1718 (N_1718,N_1461,N_1248);
xor U1719 (N_1719,N_1410,N_1024);
nand U1720 (N_1720,N_1128,N_1346);
and U1721 (N_1721,N_1300,N_1318);
and U1722 (N_1722,N_1286,N_1487);
and U1723 (N_1723,N_1119,N_1102);
nand U1724 (N_1724,N_1104,N_1009);
or U1725 (N_1725,N_1342,N_1352);
or U1726 (N_1726,N_1060,N_1357);
and U1727 (N_1727,N_1209,N_1317);
and U1728 (N_1728,N_1108,N_1251);
or U1729 (N_1729,N_1114,N_1404);
nand U1730 (N_1730,N_1363,N_1402);
nor U1731 (N_1731,N_1263,N_1148);
or U1732 (N_1732,N_1460,N_1042);
or U1733 (N_1733,N_1022,N_1302);
xnor U1734 (N_1734,N_1000,N_1364);
or U1735 (N_1735,N_1351,N_1390);
xnor U1736 (N_1736,N_1217,N_1053);
nand U1737 (N_1737,N_1309,N_1344);
nor U1738 (N_1738,N_1151,N_1109);
xor U1739 (N_1739,N_1236,N_1189);
nor U1740 (N_1740,N_1224,N_1062);
nor U1741 (N_1741,N_1078,N_1497);
or U1742 (N_1742,N_1149,N_1294);
nor U1743 (N_1743,N_1370,N_1192);
xor U1744 (N_1744,N_1202,N_1493);
and U1745 (N_1745,N_1091,N_1111);
nor U1746 (N_1746,N_1267,N_1131);
xor U1747 (N_1747,N_1068,N_1207);
and U1748 (N_1748,N_1088,N_1252);
and U1749 (N_1749,N_1123,N_1452);
xnor U1750 (N_1750,N_1244,N_1302);
and U1751 (N_1751,N_1311,N_1388);
xor U1752 (N_1752,N_1101,N_1218);
or U1753 (N_1753,N_1162,N_1033);
xnor U1754 (N_1754,N_1352,N_1459);
xor U1755 (N_1755,N_1329,N_1013);
nand U1756 (N_1756,N_1375,N_1218);
xor U1757 (N_1757,N_1124,N_1394);
nor U1758 (N_1758,N_1151,N_1464);
and U1759 (N_1759,N_1175,N_1023);
nor U1760 (N_1760,N_1284,N_1179);
or U1761 (N_1761,N_1224,N_1034);
or U1762 (N_1762,N_1355,N_1403);
nand U1763 (N_1763,N_1451,N_1336);
and U1764 (N_1764,N_1061,N_1194);
or U1765 (N_1765,N_1150,N_1139);
xnor U1766 (N_1766,N_1088,N_1115);
nor U1767 (N_1767,N_1477,N_1021);
and U1768 (N_1768,N_1254,N_1275);
nor U1769 (N_1769,N_1070,N_1208);
xor U1770 (N_1770,N_1073,N_1070);
nand U1771 (N_1771,N_1297,N_1082);
nand U1772 (N_1772,N_1105,N_1450);
nand U1773 (N_1773,N_1310,N_1436);
nor U1774 (N_1774,N_1274,N_1162);
nor U1775 (N_1775,N_1382,N_1470);
or U1776 (N_1776,N_1410,N_1327);
nor U1777 (N_1777,N_1183,N_1103);
nand U1778 (N_1778,N_1050,N_1364);
or U1779 (N_1779,N_1478,N_1219);
xor U1780 (N_1780,N_1115,N_1449);
nand U1781 (N_1781,N_1481,N_1465);
nor U1782 (N_1782,N_1499,N_1446);
nor U1783 (N_1783,N_1366,N_1033);
nor U1784 (N_1784,N_1168,N_1184);
or U1785 (N_1785,N_1223,N_1287);
or U1786 (N_1786,N_1347,N_1091);
nand U1787 (N_1787,N_1401,N_1247);
nor U1788 (N_1788,N_1417,N_1142);
or U1789 (N_1789,N_1070,N_1447);
or U1790 (N_1790,N_1381,N_1002);
nor U1791 (N_1791,N_1341,N_1273);
and U1792 (N_1792,N_1462,N_1463);
nor U1793 (N_1793,N_1467,N_1348);
xor U1794 (N_1794,N_1079,N_1488);
and U1795 (N_1795,N_1403,N_1142);
and U1796 (N_1796,N_1067,N_1259);
xor U1797 (N_1797,N_1220,N_1454);
nand U1798 (N_1798,N_1206,N_1191);
and U1799 (N_1799,N_1251,N_1218);
or U1800 (N_1800,N_1196,N_1173);
nor U1801 (N_1801,N_1068,N_1105);
and U1802 (N_1802,N_1023,N_1087);
nand U1803 (N_1803,N_1311,N_1163);
nand U1804 (N_1804,N_1141,N_1302);
or U1805 (N_1805,N_1497,N_1432);
nand U1806 (N_1806,N_1393,N_1195);
or U1807 (N_1807,N_1065,N_1482);
nor U1808 (N_1808,N_1244,N_1153);
nor U1809 (N_1809,N_1386,N_1176);
and U1810 (N_1810,N_1138,N_1397);
nor U1811 (N_1811,N_1049,N_1326);
xor U1812 (N_1812,N_1272,N_1019);
nand U1813 (N_1813,N_1316,N_1453);
and U1814 (N_1814,N_1282,N_1239);
nor U1815 (N_1815,N_1396,N_1482);
nand U1816 (N_1816,N_1087,N_1005);
or U1817 (N_1817,N_1217,N_1497);
or U1818 (N_1818,N_1379,N_1438);
xnor U1819 (N_1819,N_1357,N_1417);
or U1820 (N_1820,N_1381,N_1450);
xnor U1821 (N_1821,N_1268,N_1005);
nand U1822 (N_1822,N_1033,N_1242);
and U1823 (N_1823,N_1182,N_1132);
xor U1824 (N_1824,N_1121,N_1014);
nor U1825 (N_1825,N_1412,N_1072);
nor U1826 (N_1826,N_1199,N_1406);
xor U1827 (N_1827,N_1124,N_1172);
nand U1828 (N_1828,N_1223,N_1181);
or U1829 (N_1829,N_1452,N_1110);
xor U1830 (N_1830,N_1366,N_1314);
nor U1831 (N_1831,N_1044,N_1264);
nand U1832 (N_1832,N_1252,N_1087);
nand U1833 (N_1833,N_1059,N_1494);
nor U1834 (N_1834,N_1388,N_1108);
nand U1835 (N_1835,N_1153,N_1453);
and U1836 (N_1836,N_1395,N_1245);
nor U1837 (N_1837,N_1100,N_1074);
and U1838 (N_1838,N_1409,N_1269);
xnor U1839 (N_1839,N_1175,N_1051);
xor U1840 (N_1840,N_1201,N_1249);
nor U1841 (N_1841,N_1066,N_1097);
nor U1842 (N_1842,N_1476,N_1475);
or U1843 (N_1843,N_1321,N_1256);
nor U1844 (N_1844,N_1454,N_1377);
xor U1845 (N_1845,N_1178,N_1370);
or U1846 (N_1846,N_1255,N_1095);
xnor U1847 (N_1847,N_1316,N_1181);
xnor U1848 (N_1848,N_1470,N_1156);
or U1849 (N_1849,N_1403,N_1139);
nor U1850 (N_1850,N_1464,N_1401);
or U1851 (N_1851,N_1176,N_1021);
or U1852 (N_1852,N_1279,N_1157);
nor U1853 (N_1853,N_1333,N_1053);
nand U1854 (N_1854,N_1192,N_1057);
and U1855 (N_1855,N_1318,N_1158);
xor U1856 (N_1856,N_1356,N_1459);
nand U1857 (N_1857,N_1078,N_1286);
and U1858 (N_1858,N_1183,N_1105);
nor U1859 (N_1859,N_1030,N_1128);
nor U1860 (N_1860,N_1175,N_1254);
nand U1861 (N_1861,N_1392,N_1240);
nand U1862 (N_1862,N_1495,N_1377);
nor U1863 (N_1863,N_1089,N_1476);
nand U1864 (N_1864,N_1350,N_1488);
xnor U1865 (N_1865,N_1367,N_1238);
and U1866 (N_1866,N_1151,N_1167);
nor U1867 (N_1867,N_1129,N_1054);
nor U1868 (N_1868,N_1018,N_1456);
xnor U1869 (N_1869,N_1391,N_1430);
nor U1870 (N_1870,N_1091,N_1360);
nand U1871 (N_1871,N_1178,N_1441);
and U1872 (N_1872,N_1445,N_1442);
nand U1873 (N_1873,N_1365,N_1458);
nand U1874 (N_1874,N_1339,N_1114);
xnor U1875 (N_1875,N_1090,N_1491);
xor U1876 (N_1876,N_1457,N_1299);
or U1877 (N_1877,N_1472,N_1245);
nand U1878 (N_1878,N_1236,N_1011);
or U1879 (N_1879,N_1156,N_1162);
nor U1880 (N_1880,N_1142,N_1375);
or U1881 (N_1881,N_1155,N_1148);
and U1882 (N_1882,N_1234,N_1289);
or U1883 (N_1883,N_1340,N_1281);
or U1884 (N_1884,N_1197,N_1310);
and U1885 (N_1885,N_1104,N_1141);
xor U1886 (N_1886,N_1140,N_1365);
nor U1887 (N_1887,N_1274,N_1037);
nor U1888 (N_1888,N_1063,N_1420);
xnor U1889 (N_1889,N_1166,N_1032);
nand U1890 (N_1890,N_1144,N_1293);
or U1891 (N_1891,N_1216,N_1058);
and U1892 (N_1892,N_1309,N_1080);
or U1893 (N_1893,N_1293,N_1265);
nor U1894 (N_1894,N_1480,N_1108);
nor U1895 (N_1895,N_1428,N_1354);
nand U1896 (N_1896,N_1119,N_1279);
nor U1897 (N_1897,N_1183,N_1445);
and U1898 (N_1898,N_1371,N_1487);
nor U1899 (N_1899,N_1456,N_1270);
nor U1900 (N_1900,N_1360,N_1151);
nand U1901 (N_1901,N_1031,N_1258);
xnor U1902 (N_1902,N_1446,N_1398);
xor U1903 (N_1903,N_1366,N_1168);
xor U1904 (N_1904,N_1493,N_1381);
and U1905 (N_1905,N_1074,N_1253);
nand U1906 (N_1906,N_1029,N_1063);
nor U1907 (N_1907,N_1380,N_1046);
xnor U1908 (N_1908,N_1239,N_1026);
or U1909 (N_1909,N_1274,N_1337);
xor U1910 (N_1910,N_1367,N_1133);
nand U1911 (N_1911,N_1129,N_1275);
xor U1912 (N_1912,N_1466,N_1080);
nor U1913 (N_1913,N_1397,N_1216);
or U1914 (N_1914,N_1225,N_1204);
or U1915 (N_1915,N_1483,N_1028);
nor U1916 (N_1916,N_1144,N_1161);
nand U1917 (N_1917,N_1410,N_1413);
nor U1918 (N_1918,N_1044,N_1423);
or U1919 (N_1919,N_1027,N_1258);
xnor U1920 (N_1920,N_1241,N_1300);
nor U1921 (N_1921,N_1318,N_1223);
nor U1922 (N_1922,N_1251,N_1107);
nand U1923 (N_1923,N_1440,N_1082);
nand U1924 (N_1924,N_1439,N_1240);
nand U1925 (N_1925,N_1490,N_1128);
xor U1926 (N_1926,N_1298,N_1495);
nor U1927 (N_1927,N_1188,N_1436);
nor U1928 (N_1928,N_1089,N_1107);
or U1929 (N_1929,N_1330,N_1035);
or U1930 (N_1930,N_1499,N_1017);
xor U1931 (N_1931,N_1180,N_1490);
xor U1932 (N_1932,N_1484,N_1186);
nor U1933 (N_1933,N_1152,N_1457);
nor U1934 (N_1934,N_1286,N_1111);
nand U1935 (N_1935,N_1095,N_1126);
or U1936 (N_1936,N_1137,N_1258);
nor U1937 (N_1937,N_1314,N_1200);
nor U1938 (N_1938,N_1418,N_1437);
and U1939 (N_1939,N_1273,N_1010);
or U1940 (N_1940,N_1245,N_1042);
nor U1941 (N_1941,N_1323,N_1130);
and U1942 (N_1942,N_1409,N_1116);
xor U1943 (N_1943,N_1218,N_1449);
xor U1944 (N_1944,N_1259,N_1471);
nor U1945 (N_1945,N_1158,N_1087);
xnor U1946 (N_1946,N_1367,N_1469);
or U1947 (N_1947,N_1365,N_1003);
or U1948 (N_1948,N_1229,N_1013);
nand U1949 (N_1949,N_1029,N_1474);
nor U1950 (N_1950,N_1085,N_1489);
nand U1951 (N_1951,N_1438,N_1483);
or U1952 (N_1952,N_1308,N_1045);
and U1953 (N_1953,N_1050,N_1463);
and U1954 (N_1954,N_1372,N_1364);
or U1955 (N_1955,N_1053,N_1029);
nor U1956 (N_1956,N_1338,N_1329);
or U1957 (N_1957,N_1178,N_1460);
nand U1958 (N_1958,N_1180,N_1265);
and U1959 (N_1959,N_1075,N_1173);
nor U1960 (N_1960,N_1306,N_1185);
or U1961 (N_1961,N_1002,N_1406);
nand U1962 (N_1962,N_1468,N_1134);
xor U1963 (N_1963,N_1370,N_1174);
and U1964 (N_1964,N_1231,N_1066);
nand U1965 (N_1965,N_1117,N_1177);
nor U1966 (N_1966,N_1051,N_1140);
nand U1967 (N_1967,N_1175,N_1490);
nand U1968 (N_1968,N_1266,N_1119);
and U1969 (N_1969,N_1140,N_1091);
xor U1970 (N_1970,N_1004,N_1462);
xnor U1971 (N_1971,N_1017,N_1401);
nor U1972 (N_1972,N_1315,N_1495);
nand U1973 (N_1973,N_1378,N_1394);
and U1974 (N_1974,N_1042,N_1128);
nand U1975 (N_1975,N_1287,N_1171);
or U1976 (N_1976,N_1293,N_1024);
nor U1977 (N_1977,N_1399,N_1496);
nor U1978 (N_1978,N_1010,N_1137);
xnor U1979 (N_1979,N_1142,N_1042);
nand U1980 (N_1980,N_1387,N_1154);
xnor U1981 (N_1981,N_1447,N_1298);
nand U1982 (N_1982,N_1426,N_1027);
xor U1983 (N_1983,N_1279,N_1264);
or U1984 (N_1984,N_1400,N_1323);
xnor U1985 (N_1985,N_1322,N_1261);
or U1986 (N_1986,N_1288,N_1485);
or U1987 (N_1987,N_1245,N_1442);
xnor U1988 (N_1988,N_1134,N_1172);
xor U1989 (N_1989,N_1012,N_1055);
and U1990 (N_1990,N_1261,N_1020);
nand U1991 (N_1991,N_1024,N_1465);
xor U1992 (N_1992,N_1229,N_1327);
xor U1993 (N_1993,N_1351,N_1342);
nor U1994 (N_1994,N_1164,N_1422);
nor U1995 (N_1995,N_1201,N_1028);
and U1996 (N_1996,N_1315,N_1472);
and U1997 (N_1997,N_1490,N_1119);
or U1998 (N_1998,N_1051,N_1395);
nand U1999 (N_1999,N_1321,N_1013);
nor U2000 (N_2000,N_1901,N_1509);
nor U2001 (N_2001,N_1757,N_1745);
nor U2002 (N_2002,N_1650,N_1906);
nor U2003 (N_2003,N_1779,N_1782);
xor U2004 (N_2004,N_1784,N_1935);
nand U2005 (N_2005,N_1515,N_1795);
or U2006 (N_2006,N_1950,N_1880);
or U2007 (N_2007,N_1549,N_1584);
and U2008 (N_2008,N_1920,N_1553);
xnor U2009 (N_2009,N_1653,N_1883);
or U2010 (N_2010,N_1774,N_1873);
and U2011 (N_2011,N_1634,N_1556);
and U2012 (N_2012,N_1933,N_1843);
or U2013 (N_2013,N_1851,N_1909);
nand U2014 (N_2014,N_1945,N_1504);
nor U2015 (N_2015,N_1559,N_1862);
nor U2016 (N_2016,N_1815,N_1731);
xnor U2017 (N_2017,N_1594,N_1661);
nand U2018 (N_2018,N_1550,N_1937);
or U2019 (N_2019,N_1834,N_1613);
and U2020 (N_2020,N_1656,N_1925);
nand U2021 (N_2021,N_1989,N_1615);
xnor U2022 (N_2022,N_1742,N_1887);
and U2023 (N_2023,N_1930,N_1671);
nor U2024 (N_2024,N_1564,N_1810);
and U2025 (N_2025,N_1966,N_1589);
and U2026 (N_2026,N_1639,N_1970);
nor U2027 (N_2027,N_1555,N_1766);
xnor U2028 (N_2028,N_1809,N_1974);
nor U2029 (N_2029,N_1725,N_1599);
nand U2030 (N_2030,N_1947,N_1957);
or U2031 (N_2031,N_1645,N_1793);
nand U2032 (N_2032,N_1619,N_1510);
and U2033 (N_2033,N_1832,N_1863);
or U2034 (N_2034,N_1526,N_1631);
or U2035 (N_2035,N_1718,N_1750);
or U2036 (N_2036,N_1899,N_1850);
or U2037 (N_2037,N_1708,N_1743);
nor U2038 (N_2038,N_1758,N_1733);
and U2039 (N_2039,N_1605,N_1734);
nand U2040 (N_2040,N_1719,N_1787);
or U2041 (N_2041,N_1765,N_1700);
or U2042 (N_2042,N_1581,N_1866);
or U2043 (N_2043,N_1643,N_1754);
or U2044 (N_2044,N_1764,N_1525);
xor U2045 (N_2045,N_1516,N_1833);
nand U2046 (N_2046,N_1622,N_1612);
nor U2047 (N_2047,N_1629,N_1987);
nand U2048 (N_2048,N_1500,N_1885);
and U2049 (N_2049,N_1805,N_1895);
nand U2050 (N_2050,N_1724,N_1768);
or U2051 (N_2051,N_1951,N_1968);
nand U2052 (N_2052,N_1735,N_1667);
and U2053 (N_2053,N_1858,N_1871);
nor U2054 (N_2054,N_1691,N_1928);
xor U2055 (N_2055,N_1820,N_1938);
or U2056 (N_2056,N_1771,N_1641);
and U2057 (N_2057,N_1630,N_1702);
and U2058 (N_2058,N_1682,N_1929);
nand U2059 (N_2059,N_1620,N_1535);
nand U2060 (N_2060,N_1816,N_1633);
and U2061 (N_2061,N_1759,N_1867);
and U2062 (N_2062,N_1696,N_1777);
or U2063 (N_2063,N_1818,N_1824);
and U2064 (N_2064,N_1943,N_1614);
nor U2065 (N_2065,N_1528,N_1911);
xor U2066 (N_2066,N_1756,N_1994);
nand U2067 (N_2067,N_1587,N_1904);
nor U2068 (N_2068,N_1872,N_1940);
or U2069 (N_2069,N_1915,N_1761);
nor U2070 (N_2070,N_1907,N_1664);
xor U2071 (N_2071,N_1882,N_1511);
nor U2072 (N_2072,N_1790,N_1651);
nand U2073 (N_2073,N_1604,N_1997);
and U2074 (N_2074,N_1644,N_1905);
and U2075 (N_2075,N_1737,N_1886);
and U2076 (N_2076,N_1804,N_1699);
nor U2077 (N_2077,N_1532,N_1729);
nand U2078 (N_2078,N_1964,N_1654);
or U2079 (N_2079,N_1678,N_1590);
and U2080 (N_2080,N_1632,N_1919);
nand U2081 (N_2081,N_1783,N_1813);
xor U2082 (N_2082,N_1593,N_1694);
nand U2083 (N_2083,N_1686,N_1990);
nor U2084 (N_2084,N_1865,N_1753);
nand U2085 (N_2085,N_1709,N_1983);
and U2086 (N_2086,N_1772,N_1857);
nor U2087 (N_2087,N_1922,N_1638);
or U2088 (N_2088,N_1931,N_1652);
or U2089 (N_2089,N_1798,N_1781);
nand U2090 (N_2090,N_1898,N_1831);
xnor U2091 (N_2091,N_1946,N_1854);
nor U2092 (N_2092,N_1996,N_1568);
and U2093 (N_2093,N_1675,N_1927);
nor U2094 (N_2094,N_1827,N_1881);
or U2095 (N_2095,N_1954,N_1910);
or U2096 (N_2096,N_1517,N_1514);
xnor U2097 (N_2097,N_1681,N_1884);
nor U2098 (N_2098,N_1748,N_1977);
nand U2099 (N_2099,N_1845,N_1864);
or U2100 (N_2100,N_1621,N_1665);
nor U2101 (N_2101,N_1539,N_1890);
xnor U2102 (N_2102,N_1600,N_1860);
nand U2103 (N_2103,N_1602,N_1981);
nand U2104 (N_2104,N_1672,N_1698);
xnor U2105 (N_2105,N_1939,N_1684);
or U2106 (N_2106,N_1730,N_1623);
nand U2107 (N_2107,N_1531,N_1912);
and U2108 (N_2108,N_1926,N_1579);
or U2109 (N_2109,N_1591,N_1685);
xor U2110 (N_2110,N_1707,N_1806);
xnor U2111 (N_2111,N_1746,N_1932);
xnor U2112 (N_2112,N_1585,N_1849);
or U2113 (N_2113,N_1507,N_1807);
or U2114 (N_2114,N_1952,N_1786);
nand U2115 (N_2115,N_1519,N_1846);
and U2116 (N_2116,N_1868,N_1993);
nor U2117 (N_2117,N_1659,N_1780);
nand U2118 (N_2118,N_1878,N_1658);
or U2119 (N_2119,N_1776,N_1738);
xor U2120 (N_2120,N_1529,N_1712);
nand U2121 (N_2121,N_1836,N_1670);
nor U2122 (N_2122,N_1575,N_1603);
and U2123 (N_2123,N_1875,N_1829);
nor U2124 (N_2124,N_1856,N_1635);
nor U2125 (N_2125,N_1923,N_1891);
nor U2126 (N_2126,N_1897,N_1545);
or U2127 (N_2127,N_1900,N_1979);
or U2128 (N_2128,N_1588,N_1869);
nand U2129 (N_2129,N_1705,N_1811);
nand U2130 (N_2130,N_1668,N_1908);
xor U2131 (N_2131,N_1788,N_1578);
and U2132 (N_2132,N_1543,N_1547);
and U2133 (N_2133,N_1755,N_1502);
nand U2134 (N_2134,N_1794,N_1689);
and U2135 (N_2135,N_1592,N_1551);
xor U2136 (N_2136,N_1506,N_1797);
or U2137 (N_2137,N_1582,N_1893);
nand U2138 (N_2138,N_1640,N_1527);
nor U2139 (N_2139,N_1695,N_1728);
nand U2140 (N_2140,N_1544,N_1717);
xnor U2141 (N_2141,N_1595,N_1518);
nand U2142 (N_2142,N_1844,N_1914);
and U2143 (N_2143,N_1978,N_1601);
and U2144 (N_2144,N_1999,N_1889);
and U2145 (N_2145,N_1980,N_1649);
xor U2146 (N_2146,N_1982,N_1789);
nand U2147 (N_2147,N_1840,N_1962);
xnor U2148 (N_2148,N_1655,N_1870);
nand U2149 (N_2149,N_1975,N_1775);
or U2150 (N_2150,N_1720,N_1577);
and U2151 (N_2151,N_1835,N_1533);
or U2152 (N_2152,N_1558,N_1741);
nor U2153 (N_2153,N_1625,N_1596);
or U2154 (N_2154,N_1610,N_1913);
and U2155 (N_2155,N_1740,N_1540);
or U2156 (N_2156,N_1956,N_1902);
xnor U2157 (N_2157,N_1744,N_1648);
nand U2158 (N_2158,N_1713,N_1965);
or U2159 (N_2159,N_1791,N_1916);
xor U2160 (N_2160,N_1837,N_1876);
or U2161 (N_2161,N_1680,N_1942);
or U2162 (N_2162,N_1611,N_1732);
or U2163 (N_2163,N_1606,N_1716);
and U2164 (N_2164,N_1972,N_1542);
nor U2165 (N_2165,N_1953,N_1995);
nand U2166 (N_2166,N_1683,N_1936);
or U2167 (N_2167,N_1848,N_1616);
nand U2168 (N_2168,N_1874,N_1752);
nor U2169 (N_2169,N_1536,N_1823);
nor U2170 (N_2170,N_1546,N_1751);
or U2171 (N_2171,N_1958,N_1574);
nor U2172 (N_2172,N_1608,N_1971);
nor U2173 (N_2173,N_1800,N_1598);
xnor U2174 (N_2174,N_1674,N_1676);
or U2175 (N_2175,N_1687,N_1839);
xnor U2176 (N_2176,N_1853,N_1892);
and U2177 (N_2177,N_1692,N_1513);
or U2178 (N_2178,N_1657,N_1855);
xor U2179 (N_2179,N_1830,N_1524);
nand U2180 (N_2180,N_1802,N_1739);
nor U2181 (N_2181,N_1917,N_1646);
and U2182 (N_2182,N_1666,N_1573);
or U2183 (N_2183,N_1773,N_1859);
and U2184 (N_2184,N_1530,N_1814);
nand U2185 (N_2185,N_1697,N_1714);
and U2186 (N_2186,N_1557,N_1618);
xor U2187 (N_2187,N_1715,N_1921);
nand U2188 (N_2188,N_1988,N_1736);
or U2189 (N_2189,N_1896,N_1537);
nand U2190 (N_2190,N_1948,N_1501);
nand U2191 (N_2191,N_1503,N_1726);
nand U2192 (N_2192,N_1960,N_1894);
nand U2193 (N_2193,N_1763,N_1969);
or U2194 (N_2194,N_1944,N_1941);
xnor U2195 (N_2195,N_1986,N_1548);
xnor U2196 (N_2196,N_1647,N_1505);
or U2197 (N_2197,N_1583,N_1808);
and U2198 (N_2198,N_1523,N_1770);
xnor U2199 (N_2199,N_1747,N_1961);
and U2200 (N_2200,N_1821,N_1992);
xnor U2201 (N_2201,N_1976,N_1955);
xor U2202 (N_2202,N_1826,N_1597);
xnor U2203 (N_2203,N_1949,N_1673);
nor U2204 (N_2204,N_1801,N_1803);
or U2205 (N_2205,N_1792,N_1903);
and U2206 (N_2206,N_1521,N_1998);
and U2207 (N_2207,N_1567,N_1552);
or U2208 (N_2208,N_1677,N_1819);
nor U2209 (N_2209,N_1569,N_1723);
or U2210 (N_2210,N_1825,N_1522);
or U2211 (N_2211,N_1959,N_1534);
nand U2212 (N_2212,N_1565,N_1704);
and U2213 (N_2213,N_1560,N_1609);
nand U2214 (N_2214,N_1984,N_1693);
xor U2215 (N_2215,N_1626,N_1679);
xor U2216 (N_2216,N_1512,N_1538);
or U2217 (N_2217,N_1877,N_1918);
or U2218 (N_2218,N_1607,N_1688);
nand U2219 (N_2219,N_1690,N_1711);
and U2220 (N_2220,N_1760,N_1571);
xor U2221 (N_2221,N_1520,N_1554);
and U2222 (N_2222,N_1828,N_1508);
or U2223 (N_2223,N_1624,N_1662);
xnor U2224 (N_2224,N_1572,N_1817);
xor U2225 (N_2225,N_1785,N_1637);
or U2226 (N_2226,N_1934,N_1778);
nor U2227 (N_2227,N_1838,N_1586);
nand U2228 (N_2228,N_1636,N_1985);
nand U2229 (N_2229,N_1566,N_1842);
nand U2230 (N_2230,N_1628,N_1796);
or U2231 (N_2231,N_1991,N_1563);
and U2232 (N_2232,N_1924,N_1973);
nor U2233 (N_2233,N_1879,N_1642);
nand U2234 (N_2234,N_1710,N_1722);
or U2235 (N_2235,N_1703,N_1852);
xor U2236 (N_2236,N_1799,N_1861);
nor U2237 (N_2237,N_1561,N_1822);
xnor U2238 (N_2238,N_1769,N_1888);
and U2239 (N_2239,N_1762,N_1660);
xor U2240 (N_2240,N_1580,N_1727);
xnor U2241 (N_2241,N_1570,N_1812);
nor U2242 (N_2242,N_1576,N_1767);
nand U2243 (N_2243,N_1663,N_1627);
or U2244 (N_2244,N_1749,N_1967);
nand U2245 (N_2245,N_1562,N_1721);
and U2246 (N_2246,N_1701,N_1541);
or U2247 (N_2247,N_1963,N_1706);
and U2248 (N_2248,N_1847,N_1669);
nand U2249 (N_2249,N_1617,N_1841);
and U2250 (N_2250,N_1784,N_1597);
xor U2251 (N_2251,N_1822,N_1865);
or U2252 (N_2252,N_1958,N_1768);
nor U2253 (N_2253,N_1728,N_1820);
or U2254 (N_2254,N_1923,N_1547);
nand U2255 (N_2255,N_1818,N_1614);
nor U2256 (N_2256,N_1591,N_1567);
or U2257 (N_2257,N_1843,N_1955);
xor U2258 (N_2258,N_1824,N_1784);
nand U2259 (N_2259,N_1929,N_1563);
xnor U2260 (N_2260,N_1811,N_1986);
or U2261 (N_2261,N_1984,N_1844);
xor U2262 (N_2262,N_1935,N_1982);
nand U2263 (N_2263,N_1815,N_1559);
or U2264 (N_2264,N_1886,N_1740);
xor U2265 (N_2265,N_1954,N_1561);
and U2266 (N_2266,N_1676,N_1502);
nor U2267 (N_2267,N_1558,N_1776);
xor U2268 (N_2268,N_1566,N_1533);
xor U2269 (N_2269,N_1827,N_1897);
nand U2270 (N_2270,N_1885,N_1507);
and U2271 (N_2271,N_1720,N_1671);
nor U2272 (N_2272,N_1827,N_1739);
nand U2273 (N_2273,N_1828,N_1819);
or U2274 (N_2274,N_1970,N_1825);
and U2275 (N_2275,N_1544,N_1966);
nor U2276 (N_2276,N_1898,N_1560);
and U2277 (N_2277,N_1724,N_1568);
and U2278 (N_2278,N_1985,N_1676);
and U2279 (N_2279,N_1985,N_1887);
nor U2280 (N_2280,N_1937,N_1619);
nand U2281 (N_2281,N_1625,N_1932);
nand U2282 (N_2282,N_1930,N_1749);
nor U2283 (N_2283,N_1678,N_1600);
or U2284 (N_2284,N_1634,N_1683);
nor U2285 (N_2285,N_1702,N_1752);
and U2286 (N_2286,N_1821,N_1974);
xnor U2287 (N_2287,N_1819,N_1525);
nand U2288 (N_2288,N_1957,N_1659);
nand U2289 (N_2289,N_1973,N_1728);
xnor U2290 (N_2290,N_1766,N_1654);
xor U2291 (N_2291,N_1837,N_1580);
xnor U2292 (N_2292,N_1680,N_1827);
and U2293 (N_2293,N_1779,N_1929);
nor U2294 (N_2294,N_1733,N_1532);
nand U2295 (N_2295,N_1774,N_1976);
and U2296 (N_2296,N_1501,N_1516);
and U2297 (N_2297,N_1732,N_1782);
and U2298 (N_2298,N_1969,N_1533);
xnor U2299 (N_2299,N_1746,N_1597);
nand U2300 (N_2300,N_1733,N_1933);
and U2301 (N_2301,N_1708,N_1875);
nor U2302 (N_2302,N_1554,N_1874);
and U2303 (N_2303,N_1864,N_1893);
or U2304 (N_2304,N_1726,N_1642);
xnor U2305 (N_2305,N_1784,N_1945);
or U2306 (N_2306,N_1858,N_1774);
and U2307 (N_2307,N_1774,N_1798);
xnor U2308 (N_2308,N_1800,N_1820);
nor U2309 (N_2309,N_1923,N_1924);
nand U2310 (N_2310,N_1517,N_1995);
nor U2311 (N_2311,N_1703,N_1984);
nand U2312 (N_2312,N_1939,N_1875);
nand U2313 (N_2313,N_1694,N_1677);
xor U2314 (N_2314,N_1916,N_1781);
or U2315 (N_2315,N_1901,N_1694);
and U2316 (N_2316,N_1583,N_1658);
nand U2317 (N_2317,N_1687,N_1525);
xor U2318 (N_2318,N_1621,N_1842);
nor U2319 (N_2319,N_1758,N_1649);
and U2320 (N_2320,N_1898,N_1587);
and U2321 (N_2321,N_1743,N_1798);
or U2322 (N_2322,N_1739,N_1616);
and U2323 (N_2323,N_1739,N_1883);
nand U2324 (N_2324,N_1774,N_1796);
nor U2325 (N_2325,N_1680,N_1582);
nor U2326 (N_2326,N_1662,N_1804);
and U2327 (N_2327,N_1825,N_1719);
xnor U2328 (N_2328,N_1703,N_1908);
and U2329 (N_2329,N_1641,N_1984);
nand U2330 (N_2330,N_1678,N_1927);
nand U2331 (N_2331,N_1950,N_1586);
nor U2332 (N_2332,N_1736,N_1846);
xor U2333 (N_2333,N_1526,N_1562);
or U2334 (N_2334,N_1720,N_1979);
nor U2335 (N_2335,N_1953,N_1753);
xnor U2336 (N_2336,N_1523,N_1657);
nor U2337 (N_2337,N_1758,N_1635);
or U2338 (N_2338,N_1849,N_1550);
xor U2339 (N_2339,N_1889,N_1874);
nand U2340 (N_2340,N_1776,N_1686);
nand U2341 (N_2341,N_1644,N_1864);
nor U2342 (N_2342,N_1716,N_1551);
xor U2343 (N_2343,N_1702,N_1871);
nor U2344 (N_2344,N_1757,N_1641);
xnor U2345 (N_2345,N_1785,N_1952);
or U2346 (N_2346,N_1963,N_1903);
and U2347 (N_2347,N_1804,N_1745);
or U2348 (N_2348,N_1945,N_1771);
nor U2349 (N_2349,N_1591,N_1959);
or U2350 (N_2350,N_1804,N_1586);
nand U2351 (N_2351,N_1928,N_1925);
nand U2352 (N_2352,N_1792,N_1693);
nor U2353 (N_2353,N_1990,N_1923);
nor U2354 (N_2354,N_1786,N_1798);
nand U2355 (N_2355,N_1609,N_1632);
xor U2356 (N_2356,N_1672,N_1797);
nor U2357 (N_2357,N_1518,N_1893);
and U2358 (N_2358,N_1946,N_1721);
xor U2359 (N_2359,N_1952,N_1560);
xor U2360 (N_2360,N_1521,N_1557);
or U2361 (N_2361,N_1550,N_1985);
xnor U2362 (N_2362,N_1607,N_1535);
and U2363 (N_2363,N_1501,N_1947);
xnor U2364 (N_2364,N_1878,N_1758);
or U2365 (N_2365,N_1705,N_1555);
nand U2366 (N_2366,N_1511,N_1524);
and U2367 (N_2367,N_1680,N_1707);
nand U2368 (N_2368,N_1571,N_1713);
and U2369 (N_2369,N_1893,N_1736);
nand U2370 (N_2370,N_1830,N_1746);
or U2371 (N_2371,N_1527,N_1578);
nand U2372 (N_2372,N_1756,N_1667);
or U2373 (N_2373,N_1974,N_1816);
xor U2374 (N_2374,N_1751,N_1585);
nor U2375 (N_2375,N_1831,N_1876);
and U2376 (N_2376,N_1546,N_1695);
nand U2377 (N_2377,N_1971,N_1973);
xor U2378 (N_2378,N_1999,N_1881);
and U2379 (N_2379,N_1664,N_1827);
or U2380 (N_2380,N_1859,N_1647);
xor U2381 (N_2381,N_1605,N_1772);
nand U2382 (N_2382,N_1713,N_1536);
or U2383 (N_2383,N_1760,N_1585);
or U2384 (N_2384,N_1806,N_1676);
nand U2385 (N_2385,N_1705,N_1899);
xor U2386 (N_2386,N_1584,N_1854);
nand U2387 (N_2387,N_1576,N_1812);
or U2388 (N_2388,N_1973,N_1780);
and U2389 (N_2389,N_1778,N_1928);
nor U2390 (N_2390,N_1911,N_1520);
and U2391 (N_2391,N_1889,N_1843);
xor U2392 (N_2392,N_1714,N_1826);
or U2393 (N_2393,N_1710,N_1943);
or U2394 (N_2394,N_1936,N_1741);
xnor U2395 (N_2395,N_1863,N_1573);
xnor U2396 (N_2396,N_1787,N_1714);
nor U2397 (N_2397,N_1943,N_1879);
and U2398 (N_2398,N_1930,N_1601);
nor U2399 (N_2399,N_1869,N_1920);
nand U2400 (N_2400,N_1563,N_1515);
nor U2401 (N_2401,N_1885,N_1601);
xor U2402 (N_2402,N_1603,N_1822);
or U2403 (N_2403,N_1777,N_1903);
or U2404 (N_2404,N_1648,N_1640);
xnor U2405 (N_2405,N_1516,N_1844);
nand U2406 (N_2406,N_1555,N_1631);
nor U2407 (N_2407,N_1981,N_1503);
nand U2408 (N_2408,N_1956,N_1605);
or U2409 (N_2409,N_1791,N_1810);
and U2410 (N_2410,N_1913,N_1704);
or U2411 (N_2411,N_1539,N_1565);
xnor U2412 (N_2412,N_1620,N_1617);
nand U2413 (N_2413,N_1841,N_1703);
xor U2414 (N_2414,N_1739,N_1902);
or U2415 (N_2415,N_1555,N_1825);
and U2416 (N_2416,N_1534,N_1737);
or U2417 (N_2417,N_1795,N_1592);
and U2418 (N_2418,N_1719,N_1502);
xor U2419 (N_2419,N_1939,N_1954);
and U2420 (N_2420,N_1540,N_1828);
nor U2421 (N_2421,N_1590,N_1601);
or U2422 (N_2422,N_1997,N_1852);
nor U2423 (N_2423,N_1517,N_1856);
xor U2424 (N_2424,N_1896,N_1760);
nor U2425 (N_2425,N_1539,N_1821);
or U2426 (N_2426,N_1661,N_1981);
xnor U2427 (N_2427,N_1509,N_1677);
nor U2428 (N_2428,N_1873,N_1582);
nand U2429 (N_2429,N_1891,N_1740);
nor U2430 (N_2430,N_1916,N_1590);
and U2431 (N_2431,N_1815,N_1646);
and U2432 (N_2432,N_1574,N_1702);
nand U2433 (N_2433,N_1953,N_1768);
nand U2434 (N_2434,N_1691,N_1696);
or U2435 (N_2435,N_1818,N_1952);
or U2436 (N_2436,N_1945,N_1988);
xnor U2437 (N_2437,N_1824,N_1610);
and U2438 (N_2438,N_1505,N_1893);
nand U2439 (N_2439,N_1877,N_1978);
nand U2440 (N_2440,N_1773,N_1874);
nor U2441 (N_2441,N_1562,N_1529);
nand U2442 (N_2442,N_1801,N_1554);
xnor U2443 (N_2443,N_1690,N_1856);
nand U2444 (N_2444,N_1918,N_1773);
and U2445 (N_2445,N_1843,N_1828);
nor U2446 (N_2446,N_1876,N_1616);
and U2447 (N_2447,N_1771,N_1973);
nor U2448 (N_2448,N_1545,N_1872);
nand U2449 (N_2449,N_1741,N_1891);
nor U2450 (N_2450,N_1689,N_1532);
nor U2451 (N_2451,N_1826,N_1679);
or U2452 (N_2452,N_1706,N_1780);
nand U2453 (N_2453,N_1526,N_1872);
nor U2454 (N_2454,N_1713,N_1800);
and U2455 (N_2455,N_1783,N_1552);
xnor U2456 (N_2456,N_1947,N_1517);
or U2457 (N_2457,N_1986,N_1962);
xnor U2458 (N_2458,N_1945,N_1605);
and U2459 (N_2459,N_1554,N_1728);
nor U2460 (N_2460,N_1894,N_1971);
and U2461 (N_2461,N_1719,N_1782);
or U2462 (N_2462,N_1506,N_1901);
xor U2463 (N_2463,N_1506,N_1969);
xor U2464 (N_2464,N_1958,N_1728);
xor U2465 (N_2465,N_1688,N_1875);
xnor U2466 (N_2466,N_1962,N_1901);
xor U2467 (N_2467,N_1672,N_1796);
xor U2468 (N_2468,N_1692,N_1655);
nand U2469 (N_2469,N_1731,N_1523);
and U2470 (N_2470,N_1654,N_1524);
xnor U2471 (N_2471,N_1583,N_1750);
nand U2472 (N_2472,N_1837,N_1892);
or U2473 (N_2473,N_1838,N_1568);
xor U2474 (N_2474,N_1668,N_1886);
and U2475 (N_2475,N_1819,N_1714);
and U2476 (N_2476,N_1516,N_1694);
and U2477 (N_2477,N_1563,N_1832);
nand U2478 (N_2478,N_1645,N_1815);
xnor U2479 (N_2479,N_1838,N_1726);
or U2480 (N_2480,N_1844,N_1556);
or U2481 (N_2481,N_1598,N_1803);
or U2482 (N_2482,N_1673,N_1957);
nor U2483 (N_2483,N_1708,N_1703);
or U2484 (N_2484,N_1750,N_1917);
nand U2485 (N_2485,N_1692,N_1662);
nor U2486 (N_2486,N_1762,N_1940);
nor U2487 (N_2487,N_1897,N_1569);
nor U2488 (N_2488,N_1849,N_1789);
xnor U2489 (N_2489,N_1722,N_1753);
nand U2490 (N_2490,N_1707,N_1934);
or U2491 (N_2491,N_1952,N_1599);
nand U2492 (N_2492,N_1863,N_1697);
or U2493 (N_2493,N_1933,N_1849);
or U2494 (N_2494,N_1508,N_1623);
and U2495 (N_2495,N_1958,N_1571);
or U2496 (N_2496,N_1525,N_1912);
nor U2497 (N_2497,N_1725,N_1517);
and U2498 (N_2498,N_1864,N_1747);
nand U2499 (N_2499,N_1587,N_1919);
and U2500 (N_2500,N_2102,N_2066);
nand U2501 (N_2501,N_2442,N_2385);
nand U2502 (N_2502,N_2423,N_2071);
xor U2503 (N_2503,N_2336,N_2193);
xor U2504 (N_2504,N_2450,N_2279);
xor U2505 (N_2505,N_2120,N_2402);
nand U2506 (N_2506,N_2098,N_2386);
nor U2507 (N_2507,N_2333,N_2277);
xnor U2508 (N_2508,N_2150,N_2311);
nor U2509 (N_2509,N_2398,N_2353);
xor U2510 (N_2510,N_2130,N_2367);
and U2511 (N_2511,N_2181,N_2217);
nand U2512 (N_2512,N_2406,N_2087);
and U2513 (N_2513,N_2004,N_2001);
or U2514 (N_2514,N_2077,N_2223);
and U2515 (N_2515,N_2021,N_2464);
or U2516 (N_2516,N_2170,N_2415);
or U2517 (N_2517,N_2421,N_2005);
nor U2518 (N_2518,N_2092,N_2349);
and U2519 (N_2519,N_2467,N_2069);
and U2520 (N_2520,N_2422,N_2202);
and U2521 (N_2521,N_2324,N_2251);
nor U2522 (N_2522,N_2381,N_2143);
nor U2523 (N_2523,N_2297,N_2178);
xor U2524 (N_2524,N_2265,N_2055);
and U2525 (N_2525,N_2335,N_2195);
xnor U2526 (N_2526,N_2475,N_2135);
and U2527 (N_2527,N_2225,N_2300);
or U2528 (N_2528,N_2028,N_2363);
or U2529 (N_2529,N_2167,N_2462);
nor U2530 (N_2530,N_2303,N_2444);
nor U2531 (N_2531,N_2240,N_2292);
nor U2532 (N_2532,N_2085,N_2219);
and U2533 (N_2533,N_2316,N_2089);
xor U2534 (N_2534,N_2378,N_2308);
or U2535 (N_2535,N_2076,N_2272);
xor U2536 (N_2536,N_2156,N_2228);
nand U2537 (N_2537,N_2137,N_2203);
nand U2538 (N_2538,N_2013,N_2037);
and U2539 (N_2539,N_2326,N_2086);
or U2540 (N_2540,N_2112,N_2245);
or U2541 (N_2541,N_2115,N_2371);
nor U2542 (N_2542,N_2059,N_2169);
nor U2543 (N_2543,N_2382,N_2270);
xor U2544 (N_2544,N_2068,N_2343);
nor U2545 (N_2545,N_2006,N_2206);
or U2546 (N_2546,N_2124,N_2480);
xor U2547 (N_2547,N_2332,N_2249);
or U2548 (N_2548,N_2489,N_2294);
nor U2549 (N_2549,N_2080,N_2290);
and U2550 (N_2550,N_2458,N_2027);
nand U2551 (N_2551,N_2397,N_2466);
nor U2552 (N_2552,N_2067,N_2024);
nor U2553 (N_2553,N_2084,N_2015);
xor U2554 (N_2554,N_2045,N_2168);
nand U2555 (N_2555,N_2498,N_2393);
nand U2556 (N_2556,N_2446,N_2131);
xor U2557 (N_2557,N_2012,N_2351);
and U2558 (N_2558,N_2109,N_2495);
nand U2559 (N_2559,N_2305,N_2185);
and U2560 (N_2560,N_2145,N_2481);
nand U2561 (N_2561,N_2419,N_2197);
or U2562 (N_2562,N_2493,N_2039);
nor U2563 (N_2563,N_2038,N_2320);
nor U2564 (N_2564,N_2123,N_2389);
and U2565 (N_2565,N_2042,N_2162);
nand U2566 (N_2566,N_2079,N_2409);
nand U2567 (N_2567,N_2288,N_2044);
and U2568 (N_2568,N_2205,N_2065);
xnor U2569 (N_2569,N_2016,N_2091);
xnor U2570 (N_2570,N_2298,N_2163);
nor U2571 (N_2571,N_2494,N_2025);
or U2572 (N_2572,N_2113,N_2058);
nand U2573 (N_2573,N_2242,N_2449);
and U2574 (N_2574,N_2034,N_2201);
or U2575 (N_2575,N_2139,N_2325);
nand U2576 (N_2576,N_2400,N_2022);
or U2577 (N_2577,N_2267,N_2438);
nor U2578 (N_2578,N_2281,N_2032);
nand U2579 (N_2579,N_2246,N_2072);
xor U2580 (N_2580,N_2470,N_2296);
or U2581 (N_2581,N_2008,N_2054);
nor U2582 (N_2582,N_2261,N_2010);
and U2583 (N_2583,N_2282,N_2184);
nand U2584 (N_2584,N_2314,N_2429);
or U2585 (N_2585,N_2097,N_2134);
xnor U2586 (N_2586,N_2274,N_2317);
and U2587 (N_2587,N_2117,N_2018);
nor U2588 (N_2588,N_2148,N_2153);
xor U2589 (N_2589,N_2142,N_2176);
xnor U2590 (N_2590,N_2183,N_2486);
nor U2591 (N_2591,N_2035,N_2328);
or U2592 (N_2592,N_2252,N_2331);
nor U2593 (N_2593,N_2499,N_2154);
nor U2594 (N_2594,N_2126,N_2323);
nand U2595 (N_2595,N_2443,N_2469);
nor U2596 (N_2596,N_2330,N_2302);
nor U2597 (N_2597,N_2241,N_2362);
xnor U2598 (N_2598,N_2374,N_2285);
or U2599 (N_2599,N_2144,N_2430);
nand U2600 (N_2600,N_2243,N_2310);
nor U2601 (N_2601,N_2436,N_2239);
nand U2602 (N_2602,N_2479,N_2408);
or U2603 (N_2603,N_2482,N_2187);
and U2604 (N_2604,N_2266,N_2114);
or U2605 (N_2605,N_2488,N_2361);
nor U2606 (N_2606,N_2158,N_2365);
or U2607 (N_2607,N_2405,N_2198);
nand U2608 (N_2608,N_2452,N_2108);
or U2609 (N_2609,N_2368,N_2439);
and U2610 (N_2610,N_2020,N_2254);
xnor U2611 (N_2611,N_2295,N_2062);
nand U2612 (N_2612,N_2453,N_2061);
or U2613 (N_2613,N_2403,N_2064);
nand U2614 (N_2614,N_2356,N_2411);
nand U2615 (N_2615,N_2358,N_2096);
nand U2616 (N_2616,N_2428,N_2172);
nand U2617 (N_2617,N_2136,N_2485);
nand U2618 (N_2618,N_2433,N_2159);
xnor U2619 (N_2619,N_2461,N_2132);
nand U2620 (N_2620,N_2370,N_2026);
nor U2621 (N_2621,N_2211,N_2291);
and U2622 (N_2622,N_2401,N_2111);
xor U2623 (N_2623,N_2214,N_2196);
nor U2624 (N_2624,N_2399,N_2250);
nor U2625 (N_2625,N_2372,N_2074);
and U2626 (N_2626,N_2152,N_2334);
or U2627 (N_2627,N_2000,N_2396);
and U2628 (N_2628,N_2116,N_2424);
or U2629 (N_2629,N_2346,N_2051);
or U2630 (N_2630,N_2057,N_2341);
and U2631 (N_2631,N_2427,N_2283);
nor U2632 (N_2632,N_2221,N_2070);
or U2633 (N_2633,N_2262,N_2047);
and U2634 (N_2634,N_2041,N_2431);
and U2635 (N_2635,N_2484,N_2344);
or U2636 (N_2636,N_2379,N_2440);
nand U2637 (N_2637,N_2191,N_2149);
or U2638 (N_2638,N_2229,N_2208);
or U2639 (N_2639,N_2235,N_2233);
or U2640 (N_2640,N_2164,N_2471);
xnor U2641 (N_2641,N_2321,N_2147);
nand U2642 (N_2642,N_2391,N_2293);
xor U2643 (N_2643,N_2210,N_2383);
nand U2644 (N_2644,N_2204,N_2448);
nor U2645 (N_2645,N_2138,N_2434);
or U2646 (N_2646,N_2190,N_2040);
and U2647 (N_2647,N_2073,N_2258);
and U2648 (N_2648,N_2118,N_2175);
xnor U2649 (N_2649,N_2390,N_2269);
nand U2650 (N_2650,N_2141,N_2151);
or U2651 (N_2651,N_2425,N_2460);
and U2652 (N_2652,N_2451,N_2490);
or U2653 (N_2653,N_2327,N_2188);
and U2654 (N_2654,N_2271,N_2412);
xor U2655 (N_2655,N_2286,N_2180);
nand U2656 (N_2656,N_2338,N_2209);
xor U2657 (N_2657,N_2220,N_2093);
and U2658 (N_2658,N_2146,N_2119);
nor U2659 (N_2659,N_2230,N_2056);
nor U2660 (N_2660,N_2031,N_2174);
nand U2661 (N_2661,N_2046,N_2043);
or U2662 (N_2662,N_2432,N_2359);
and U2663 (N_2663,N_2030,N_2459);
nand U2664 (N_2664,N_2416,N_2226);
nand U2665 (N_2665,N_2002,N_2478);
or U2666 (N_2666,N_2088,N_2369);
xor U2667 (N_2667,N_2420,N_2468);
and U2668 (N_2668,N_2352,N_2248);
and U2669 (N_2669,N_2003,N_2384);
or U2670 (N_2670,N_2099,N_2127);
and U2671 (N_2671,N_2105,N_2173);
xor U2672 (N_2672,N_2125,N_2380);
nand U2673 (N_2673,N_2456,N_2160);
xnor U2674 (N_2674,N_2418,N_2340);
and U2675 (N_2675,N_2081,N_2094);
or U2676 (N_2676,N_2048,N_2253);
and U2677 (N_2677,N_2011,N_2238);
nor U2678 (N_2678,N_2360,N_2445);
nand U2679 (N_2679,N_2216,N_2417);
and U2680 (N_2680,N_2414,N_2104);
xor U2681 (N_2681,N_2082,N_2435);
xor U2682 (N_2682,N_2273,N_2410);
xnor U2683 (N_2683,N_2301,N_2194);
xnor U2684 (N_2684,N_2244,N_2395);
xnor U2685 (N_2685,N_2213,N_2189);
and U2686 (N_2686,N_2007,N_2166);
or U2687 (N_2687,N_2036,N_2155);
nor U2688 (N_2688,N_2318,N_2312);
or U2689 (N_2689,N_2257,N_2052);
and U2690 (N_2690,N_2095,N_2437);
nor U2691 (N_2691,N_2276,N_2465);
or U2692 (N_2692,N_2483,N_2247);
and U2693 (N_2693,N_2263,N_2171);
or U2694 (N_2694,N_2284,N_2280);
xnor U2695 (N_2695,N_2121,N_2177);
nor U2696 (N_2696,N_2100,N_2497);
and U2697 (N_2697,N_2023,N_2345);
nor U2698 (N_2698,N_2377,N_2060);
and U2699 (N_2699,N_2492,N_2347);
or U2700 (N_2700,N_2049,N_2259);
xnor U2701 (N_2701,N_2256,N_2165);
or U2702 (N_2702,N_2207,N_2222);
xor U2703 (N_2703,N_2236,N_2426);
nor U2704 (N_2704,N_2237,N_2199);
or U2705 (N_2705,N_2014,N_2392);
nor U2706 (N_2706,N_2476,N_2388);
or U2707 (N_2707,N_2179,N_2491);
and U2708 (N_2708,N_2106,N_2348);
and U2709 (N_2709,N_2029,N_2234);
or U2710 (N_2710,N_2387,N_2107);
xnor U2711 (N_2711,N_2140,N_2350);
nand U2712 (N_2712,N_2161,N_2101);
nor U2713 (N_2713,N_2200,N_2224);
nand U2714 (N_2714,N_2315,N_2313);
xor U2715 (N_2715,N_2009,N_2231);
nor U2716 (N_2716,N_2355,N_2404);
and U2717 (N_2717,N_2376,N_2413);
or U2718 (N_2718,N_2110,N_2455);
or U2719 (N_2719,N_2053,N_2322);
xor U2720 (N_2720,N_2050,N_2182);
nor U2721 (N_2721,N_2186,N_2477);
xor U2722 (N_2722,N_2473,N_2337);
or U2723 (N_2723,N_2366,N_2255);
nor U2724 (N_2724,N_2487,N_2129);
or U2725 (N_2725,N_2472,N_2373);
xnor U2726 (N_2726,N_2090,N_2227);
nand U2727 (N_2727,N_2122,N_2463);
and U2728 (N_2728,N_2457,N_2304);
xor U2729 (N_2729,N_2063,N_2375);
xor U2730 (N_2730,N_2232,N_2278);
nand U2731 (N_2731,N_2128,N_2441);
xnor U2732 (N_2732,N_2289,N_2329);
xnor U2733 (N_2733,N_2342,N_2299);
xnor U2734 (N_2734,N_2017,N_2474);
nand U2735 (N_2735,N_2275,N_2496);
and U2736 (N_2736,N_2407,N_2078);
xor U2737 (N_2737,N_2103,N_2192);
and U2738 (N_2738,N_2075,N_2354);
nor U2739 (N_2739,N_2019,N_2157);
nor U2740 (N_2740,N_2319,N_2339);
nor U2741 (N_2741,N_2309,N_2447);
or U2742 (N_2742,N_2306,N_2357);
nor U2743 (N_2743,N_2287,N_2212);
or U2744 (N_2744,N_2364,N_2033);
or U2745 (N_2745,N_2083,N_2260);
and U2746 (N_2746,N_2218,N_2133);
and U2747 (N_2747,N_2454,N_2394);
or U2748 (N_2748,N_2264,N_2307);
xor U2749 (N_2749,N_2268,N_2215);
and U2750 (N_2750,N_2143,N_2053);
and U2751 (N_2751,N_2230,N_2209);
or U2752 (N_2752,N_2046,N_2445);
and U2753 (N_2753,N_2257,N_2025);
or U2754 (N_2754,N_2015,N_2017);
xnor U2755 (N_2755,N_2293,N_2446);
or U2756 (N_2756,N_2281,N_2408);
xnor U2757 (N_2757,N_2300,N_2195);
and U2758 (N_2758,N_2330,N_2109);
xnor U2759 (N_2759,N_2337,N_2263);
nor U2760 (N_2760,N_2485,N_2420);
or U2761 (N_2761,N_2371,N_2413);
and U2762 (N_2762,N_2405,N_2017);
nor U2763 (N_2763,N_2434,N_2314);
nand U2764 (N_2764,N_2176,N_2113);
nor U2765 (N_2765,N_2448,N_2285);
nor U2766 (N_2766,N_2376,N_2362);
or U2767 (N_2767,N_2352,N_2249);
and U2768 (N_2768,N_2398,N_2215);
xnor U2769 (N_2769,N_2219,N_2283);
xnor U2770 (N_2770,N_2148,N_2261);
and U2771 (N_2771,N_2381,N_2173);
nand U2772 (N_2772,N_2034,N_2033);
and U2773 (N_2773,N_2177,N_2451);
nor U2774 (N_2774,N_2451,N_2013);
and U2775 (N_2775,N_2096,N_2286);
or U2776 (N_2776,N_2337,N_2421);
or U2777 (N_2777,N_2376,N_2358);
nand U2778 (N_2778,N_2218,N_2251);
or U2779 (N_2779,N_2215,N_2064);
and U2780 (N_2780,N_2280,N_2345);
nand U2781 (N_2781,N_2422,N_2091);
or U2782 (N_2782,N_2481,N_2267);
or U2783 (N_2783,N_2393,N_2326);
and U2784 (N_2784,N_2477,N_2036);
or U2785 (N_2785,N_2123,N_2173);
nand U2786 (N_2786,N_2092,N_2262);
or U2787 (N_2787,N_2405,N_2117);
nand U2788 (N_2788,N_2051,N_2020);
or U2789 (N_2789,N_2362,N_2104);
and U2790 (N_2790,N_2279,N_2067);
and U2791 (N_2791,N_2134,N_2104);
nor U2792 (N_2792,N_2294,N_2344);
or U2793 (N_2793,N_2154,N_2032);
xnor U2794 (N_2794,N_2177,N_2384);
xnor U2795 (N_2795,N_2323,N_2022);
nand U2796 (N_2796,N_2093,N_2290);
and U2797 (N_2797,N_2179,N_2247);
or U2798 (N_2798,N_2352,N_2477);
xor U2799 (N_2799,N_2041,N_2090);
and U2800 (N_2800,N_2116,N_2033);
nand U2801 (N_2801,N_2468,N_2083);
nand U2802 (N_2802,N_2361,N_2065);
or U2803 (N_2803,N_2124,N_2173);
xnor U2804 (N_2804,N_2288,N_2100);
nand U2805 (N_2805,N_2195,N_2188);
nor U2806 (N_2806,N_2408,N_2192);
xnor U2807 (N_2807,N_2385,N_2286);
xor U2808 (N_2808,N_2171,N_2220);
nand U2809 (N_2809,N_2432,N_2257);
xor U2810 (N_2810,N_2385,N_2365);
xnor U2811 (N_2811,N_2405,N_2359);
nor U2812 (N_2812,N_2467,N_2432);
xnor U2813 (N_2813,N_2151,N_2022);
nand U2814 (N_2814,N_2107,N_2287);
and U2815 (N_2815,N_2021,N_2460);
nor U2816 (N_2816,N_2478,N_2057);
or U2817 (N_2817,N_2360,N_2082);
nand U2818 (N_2818,N_2428,N_2348);
or U2819 (N_2819,N_2221,N_2114);
xor U2820 (N_2820,N_2408,N_2092);
or U2821 (N_2821,N_2306,N_2212);
nand U2822 (N_2822,N_2354,N_2112);
or U2823 (N_2823,N_2150,N_2201);
nor U2824 (N_2824,N_2133,N_2157);
xor U2825 (N_2825,N_2347,N_2070);
nor U2826 (N_2826,N_2130,N_2356);
or U2827 (N_2827,N_2450,N_2146);
nand U2828 (N_2828,N_2460,N_2421);
xor U2829 (N_2829,N_2283,N_2151);
nor U2830 (N_2830,N_2103,N_2021);
xor U2831 (N_2831,N_2177,N_2333);
xnor U2832 (N_2832,N_2003,N_2125);
xor U2833 (N_2833,N_2268,N_2281);
xnor U2834 (N_2834,N_2446,N_2167);
or U2835 (N_2835,N_2322,N_2371);
nor U2836 (N_2836,N_2269,N_2412);
and U2837 (N_2837,N_2445,N_2126);
or U2838 (N_2838,N_2368,N_2326);
nand U2839 (N_2839,N_2035,N_2418);
nor U2840 (N_2840,N_2091,N_2272);
xor U2841 (N_2841,N_2175,N_2363);
nand U2842 (N_2842,N_2036,N_2323);
xnor U2843 (N_2843,N_2401,N_2252);
nor U2844 (N_2844,N_2216,N_2304);
nand U2845 (N_2845,N_2256,N_2393);
and U2846 (N_2846,N_2327,N_2152);
xnor U2847 (N_2847,N_2127,N_2398);
or U2848 (N_2848,N_2197,N_2183);
or U2849 (N_2849,N_2145,N_2224);
nand U2850 (N_2850,N_2052,N_2218);
nand U2851 (N_2851,N_2147,N_2262);
nor U2852 (N_2852,N_2269,N_2175);
nand U2853 (N_2853,N_2444,N_2209);
nand U2854 (N_2854,N_2416,N_2040);
and U2855 (N_2855,N_2042,N_2322);
nor U2856 (N_2856,N_2263,N_2155);
xnor U2857 (N_2857,N_2489,N_2110);
and U2858 (N_2858,N_2060,N_2246);
xor U2859 (N_2859,N_2283,N_2333);
nor U2860 (N_2860,N_2379,N_2195);
and U2861 (N_2861,N_2260,N_2101);
nand U2862 (N_2862,N_2431,N_2069);
nand U2863 (N_2863,N_2123,N_2444);
xor U2864 (N_2864,N_2214,N_2117);
nand U2865 (N_2865,N_2312,N_2325);
and U2866 (N_2866,N_2004,N_2483);
nor U2867 (N_2867,N_2337,N_2054);
nor U2868 (N_2868,N_2396,N_2227);
or U2869 (N_2869,N_2402,N_2260);
nand U2870 (N_2870,N_2173,N_2386);
or U2871 (N_2871,N_2464,N_2230);
and U2872 (N_2872,N_2041,N_2143);
xor U2873 (N_2873,N_2090,N_2016);
nor U2874 (N_2874,N_2406,N_2048);
and U2875 (N_2875,N_2021,N_2220);
and U2876 (N_2876,N_2307,N_2167);
nor U2877 (N_2877,N_2044,N_2358);
nand U2878 (N_2878,N_2105,N_2221);
xor U2879 (N_2879,N_2132,N_2010);
nand U2880 (N_2880,N_2380,N_2415);
or U2881 (N_2881,N_2298,N_2153);
or U2882 (N_2882,N_2442,N_2199);
nand U2883 (N_2883,N_2045,N_2287);
xor U2884 (N_2884,N_2382,N_2293);
and U2885 (N_2885,N_2367,N_2361);
and U2886 (N_2886,N_2145,N_2451);
or U2887 (N_2887,N_2331,N_2291);
nand U2888 (N_2888,N_2274,N_2233);
nand U2889 (N_2889,N_2166,N_2330);
nand U2890 (N_2890,N_2480,N_2365);
nor U2891 (N_2891,N_2441,N_2111);
xor U2892 (N_2892,N_2272,N_2124);
nor U2893 (N_2893,N_2249,N_2451);
and U2894 (N_2894,N_2368,N_2042);
nand U2895 (N_2895,N_2374,N_2068);
or U2896 (N_2896,N_2109,N_2010);
and U2897 (N_2897,N_2422,N_2426);
and U2898 (N_2898,N_2116,N_2287);
or U2899 (N_2899,N_2027,N_2359);
nand U2900 (N_2900,N_2044,N_2256);
nand U2901 (N_2901,N_2175,N_2278);
and U2902 (N_2902,N_2306,N_2165);
nand U2903 (N_2903,N_2050,N_2362);
xnor U2904 (N_2904,N_2260,N_2053);
or U2905 (N_2905,N_2324,N_2286);
and U2906 (N_2906,N_2013,N_2462);
and U2907 (N_2907,N_2079,N_2132);
nand U2908 (N_2908,N_2288,N_2140);
xnor U2909 (N_2909,N_2197,N_2427);
and U2910 (N_2910,N_2017,N_2448);
nand U2911 (N_2911,N_2367,N_2185);
nor U2912 (N_2912,N_2154,N_2242);
nor U2913 (N_2913,N_2030,N_2106);
and U2914 (N_2914,N_2284,N_2361);
and U2915 (N_2915,N_2448,N_2166);
xor U2916 (N_2916,N_2174,N_2400);
xor U2917 (N_2917,N_2152,N_2298);
nand U2918 (N_2918,N_2417,N_2383);
or U2919 (N_2919,N_2251,N_2449);
xnor U2920 (N_2920,N_2187,N_2443);
and U2921 (N_2921,N_2023,N_2067);
nor U2922 (N_2922,N_2113,N_2419);
nor U2923 (N_2923,N_2105,N_2096);
or U2924 (N_2924,N_2214,N_2399);
nand U2925 (N_2925,N_2003,N_2414);
xor U2926 (N_2926,N_2465,N_2135);
nor U2927 (N_2927,N_2378,N_2089);
and U2928 (N_2928,N_2288,N_2028);
or U2929 (N_2929,N_2033,N_2159);
xnor U2930 (N_2930,N_2248,N_2497);
and U2931 (N_2931,N_2153,N_2293);
nand U2932 (N_2932,N_2478,N_2347);
nand U2933 (N_2933,N_2467,N_2427);
nor U2934 (N_2934,N_2442,N_2037);
nor U2935 (N_2935,N_2015,N_2298);
xnor U2936 (N_2936,N_2388,N_2451);
nor U2937 (N_2937,N_2438,N_2323);
nor U2938 (N_2938,N_2315,N_2285);
and U2939 (N_2939,N_2240,N_2428);
or U2940 (N_2940,N_2210,N_2384);
and U2941 (N_2941,N_2114,N_2246);
xnor U2942 (N_2942,N_2266,N_2265);
and U2943 (N_2943,N_2208,N_2095);
nand U2944 (N_2944,N_2203,N_2067);
and U2945 (N_2945,N_2166,N_2493);
and U2946 (N_2946,N_2359,N_2444);
nand U2947 (N_2947,N_2336,N_2313);
nand U2948 (N_2948,N_2214,N_2365);
and U2949 (N_2949,N_2039,N_2221);
xnor U2950 (N_2950,N_2231,N_2487);
nand U2951 (N_2951,N_2090,N_2085);
and U2952 (N_2952,N_2280,N_2096);
xor U2953 (N_2953,N_2250,N_2085);
and U2954 (N_2954,N_2050,N_2177);
xnor U2955 (N_2955,N_2066,N_2069);
or U2956 (N_2956,N_2452,N_2059);
and U2957 (N_2957,N_2450,N_2120);
xor U2958 (N_2958,N_2470,N_2203);
nand U2959 (N_2959,N_2063,N_2110);
xor U2960 (N_2960,N_2012,N_2137);
and U2961 (N_2961,N_2395,N_2006);
or U2962 (N_2962,N_2323,N_2416);
xor U2963 (N_2963,N_2258,N_2400);
nand U2964 (N_2964,N_2106,N_2027);
or U2965 (N_2965,N_2262,N_2368);
or U2966 (N_2966,N_2413,N_2317);
nand U2967 (N_2967,N_2211,N_2112);
nand U2968 (N_2968,N_2100,N_2268);
or U2969 (N_2969,N_2161,N_2456);
nor U2970 (N_2970,N_2406,N_2449);
and U2971 (N_2971,N_2022,N_2415);
nand U2972 (N_2972,N_2133,N_2363);
or U2973 (N_2973,N_2033,N_2120);
and U2974 (N_2974,N_2281,N_2188);
nand U2975 (N_2975,N_2113,N_2064);
nor U2976 (N_2976,N_2190,N_2228);
and U2977 (N_2977,N_2263,N_2114);
nor U2978 (N_2978,N_2382,N_2474);
or U2979 (N_2979,N_2087,N_2333);
and U2980 (N_2980,N_2369,N_2383);
or U2981 (N_2981,N_2228,N_2108);
xnor U2982 (N_2982,N_2098,N_2418);
and U2983 (N_2983,N_2355,N_2331);
and U2984 (N_2984,N_2261,N_2358);
and U2985 (N_2985,N_2257,N_2022);
nand U2986 (N_2986,N_2325,N_2110);
and U2987 (N_2987,N_2470,N_2029);
xor U2988 (N_2988,N_2161,N_2487);
xnor U2989 (N_2989,N_2213,N_2185);
xnor U2990 (N_2990,N_2245,N_2106);
nand U2991 (N_2991,N_2189,N_2426);
nand U2992 (N_2992,N_2384,N_2201);
and U2993 (N_2993,N_2000,N_2429);
xor U2994 (N_2994,N_2227,N_2438);
nand U2995 (N_2995,N_2455,N_2334);
nand U2996 (N_2996,N_2433,N_2055);
nor U2997 (N_2997,N_2178,N_2186);
or U2998 (N_2998,N_2187,N_2196);
or U2999 (N_2999,N_2166,N_2459);
nor UO_0 (O_0,N_2613,N_2875);
nand UO_1 (O_1,N_2722,N_2746);
and UO_2 (O_2,N_2820,N_2514);
xnor UO_3 (O_3,N_2927,N_2633);
nand UO_4 (O_4,N_2830,N_2534);
xor UO_5 (O_5,N_2705,N_2603);
or UO_6 (O_6,N_2944,N_2846);
nand UO_7 (O_7,N_2965,N_2630);
nor UO_8 (O_8,N_2536,N_2931);
nand UO_9 (O_9,N_2509,N_2672);
nor UO_10 (O_10,N_2643,N_2858);
and UO_11 (O_11,N_2512,N_2808);
and UO_12 (O_12,N_2991,N_2584);
xnor UO_13 (O_13,N_2761,N_2979);
nand UO_14 (O_14,N_2850,N_2974);
nand UO_15 (O_15,N_2992,N_2550);
and UO_16 (O_16,N_2701,N_2551);
or UO_17 (O_17,N_2753,N_2657);
nand UO_18 (O_18,N_2933,N_2598);
or UO_19 (O_19,N_2513,N_2986);
or UO_20 (O_20,N_2975,N_2525);
and UO_21 (O_21,N_2520,N_2577);
nor UO_22 (O_22,N_2893,N_2531);
nand UO_23 (O_23,N_2956,N_2669);
nor UO_24 (O_24,N_2812,N_2922);
nand UO_25 (O_25,N_2844,N_2569);
nor UO_26 (O_26,N_2904,N_2727);
nand UO_27 (O_27,N_2608,N_2687);
or UO_28 (O_28,N_2511,N_2612);
and UO_29 (O_29,N_2868,N_2545);
and UO_30 (O_30,N_2754,N_2817);
or UO_31 (O_31,N_2610,N_2831);
or UO_32 (O_32,N_2563,N_2823);
nor UO_33 (O_33,N_2818,N_2535);
xnor UO_34 (O_34,N_2686,N_2937);
xor UO_35 (O_35,N_2959,N_2886);
or UO_36 (O_36,N_2955,N_2622);
xor UO_37 (O_37,N_2703,N_2556);
xnor UO_38 (O_38,N_2856,N_2683);
nand UO_39 (O_39,N_2571,N_2673);
xor UO_40 (O_40,N_2735,N_2611);
and UO_41 (O_41,N_2656,N_2601);
xor UO_42 (O_42,N_2607,N_2691);
and UO_43 (O_43,N_2859,N_2950);
nor UO_44 (O_44,N_2659,N_2902);
nor UO_45 (O_45,N_2614,N_2898);
and UO_46 (O_46,N_2695,N_2790);
xor UO_47 (O_47,N_2935,N_2967);
and UO_48 (O_48,N_2797,N_2606);
or UO_49 (O_49,N_2855,N_2892);
and UO_50 (O_50,N_2662,N_2777);
xnor UO_51 (O_51,N_2888,N_2515);
or UO_52 (O_52,N_2772,N_2674);
nand UO_53 (O_53,N_2504,N_2762);
nor UO_54 (O_54,N_2739,N_2936);
xor UO_55 (O_55,N_2838,N_2912);
and UO_56 (O_56,N_2816,N_2896);
nor UO_57 (O_57,N_2693,N_2899);
nor UO_58 (O_58,N_2985,N_2783);
and UO_59 (O_59,N_2594,N_2652);
nor UO_60 (O_60,N_2802,N_2923);
nor UO_61 (O_61,N_2828,N_2984);
nand UO_62 (O_62,N_2524,N_2887);
and UO_63 (O_63,N_2940,N_2963);
nand UO_64 (O_64,N_2579,N_2609);
nor UO_65 (O_65,N_2806,N_2720);
or UO_66 (O_66,N_2747,N_2730);
nor UO_67 (O_67,N_2913,N_2919);
nand UO_68 (O_68,N_2872,N_2781);
xor UO_69 (O_69,N_2682,N_2891);
or UO_70 (O_70,N_2676,N_2784);
xnor UO_71 (O_71,N_2758,N_2702);
xnor UO_72 (O_72,N_2755,N_2996);
xnor UO_73 (O_73,N_2995,N_2748);
nand UO_74 (O_74,N_2507,N_2900);
nand UO_75 (O_75,N_2798,N_2770);
or UO_76 (O_76,N_2629,N_2663);
nand UO_77 (O_77,N_2717,N_2616);
xnor UO_78 (O_78,N_2501,N_2533);
nor UO_79 (O_79,N_2759,N_2848);
or UO_80 (O_80,N_2764,N_2660);
or UO_81 (O_81,N_2597,N_2926);
xor UO_82 (O_82,N_2842,N_2775);
and UO_83 (O_83,N_2526,N_2993);
xnor UO_84 (O_84,N_2821,N_2977);
nand UO_85 (O_85,N_2617,N_2707);
nor UO_86 (O_86,N_2654,N_2723);
xor UO_87 (O_87,N_2810,N_2724);
nor UO_88 (O_88,N_2518,N_2671);
nand UO_89 (O_89,N_2521,N_2837);
nor UO_90 (O_90,N_2742,N_2824);
nand UO_91 (O_91,N_2508,N_2641);
xnor UO_92 (O_92,N_2636,N_2989);
or UO_93 (O_93,N_2756,N_2819);
and UO_94 (O_94,N_2541,N_2964);
nor UO_95 (O_95,N_2668,N_2881);
xnor UO_96 (O_96,N_2885,N_2568);
nand UO_97 (O_97,N_2953,N_2527);
and UO_98 (O_98,N_2882,N_2814);
nand UO_99 (O_99,N_2757,N_2949);
nor UO_100 (O_100,N_2832,N_2983);
xor UO_101 (O_101,N_2714,N_2646);
and UO_102 (O_102,N_2920,N_2916);
nor UO_103 (O_103,N_2538,N_2980);
xor UO_104 (O_104,N_2645,N_2736);
xnor UO_105 (O_105,N_2681,N_2679);
nand UO_106 (O_106,N_2751,N_2696);
or UO_107 (O_107,N_2807,N_2910);
xnor UO_108 (O_108,N_2860,N_2804);
nor UO_109 (O_109,N_2729,N_2811);
xor UO_110 (O_110,N_2778,N_2952);
nor UO_111 (O_111,N_2528,N_2960);
xor UO_112 (O_112,N_2620,N_2500);
nand UO_113 (O_113,N_2769,N_2625);
nor UO_114 (O_114,N_2690,N_2516);
nor UO_115 (O_115,N_2853,N_2795);
or UO_116 (O_116,N_2994,N_2851);
or UO_117 (O_117,N_2870,N_2743);
or UO_118 (O_118,N_2575,N_2698);
or UO_119 (O_119,N_2566,N_2911);
xor UO_120 (O_120,N_2634,N_2947);
nor UO_121 (O_121,N_2618,N_2697);
and UO_122 (O_122,N_2667,N_2574);
xnor UO_123 (O_123,N_2801,N_2962);
nor UO_124 (O_124,N_2879,N_2655);
xor UO_125 (O_125,N_2649,N_2680);
or UO_126 (O_126,N_2715,N_2780);
nand UO_127 (O_127,N_2591,N_2589);
or UO_128 (O_128,N_2675,N_2505);
xor UO_129 (O_129,N_2670,N_2908);
and UO_130 (O_130,N_2889,N_2685);
or UO_131 (O_131,N_2951,N_2564);
nand UO_132 (O_132,N_2523,N_2576);
xor UO_133 (O_133,N_2544,N_2878);
and UO_134 (O_134,N_2626,N_2578);
or UO_135 (O_135,N_2638,N_2585);
and UO_136 (O_136,N_2688,N_2517);
nor UO_137 (O_137,N_2903,N_2961);
nand UO_138 (O_138,N_2867,N_2813);
and UO_139 (O_139,N_2864,N_2588);
nand UO_140 (O_140,N_2726,N_2704);
and UO_141 (O_141,N_2941,N_2958);
xor UO_142 (O_142,N_2917,N_2829);
xor UO_143 (O_143,N_2948,N_2738);
nand UO_144 (O_144,N_2786,N_2570);
nand UO_145 (O_145,N_2918,N_2639);
or UO_146 (O_146,N_2623,N_2901);
nand UO_147 (O_147,N_2737,N_2689);
nand UO_148 (O_148,N_2631,N_2938);
or UO_149 (O_149,N_2815,N_2592);
nor UO_150 (O_150,N_2745,N_2794);
nor UO_151 (O_151,N_2734,N_2866);
or UO_152 (O_152,N_2627,N_2708);
nor UO_153 (O_153,N_2880,N_2973);
or UO_154 (O_154,N_2529,N_2954);
and UO_155 (O_155,N_2788,N_2785);
nand UO_156 (O_156,N_2637,N_2557);
xnor UO_157 (O_157,N_2642,N_2854);
and UO_158 (O_158,N_2718,N_2624);
nor UO_159 (O_159,N_2547,N_2539);
xor UO_160 (O_160,N_2978,N_2648);
or UO_161 (O_161,N_2749,N_2537);
and UO_162 (O_162,N_2763,N_2827);
or UO_163 (O_163,N_2914,N_2628);
xnor UO_164 (O_164,N_2530,N_2826);
or UO_165 (O_165,N_2694,N_2849);
and UO_166 (O_166,N_2664,N_2621);
and UO_167 (O_167,N_2750,N_2957);
and UO_168 (O_168,N_2877,N_2939);
xor UO_169 (O_169,N_2921,N_2839);
nor UO_170 (O_170,N_2873,N_2604);
xnor UO_171 (O_171,N_2555,N_2605);
xnor UO_172 (O_172,N_2852,N_2562);
xnor UO_173 (O_173,N_2776,N_2968);
nand UO_174 (O_174,N_2650,N_2857);
nor UO_175 (O_175,N_2560,N_2587);
nand UO_176 (O_176,N_2600,N_2658);
nor UO_177 (O_177,N_2861,N_2946);
xnor UO_178 (O_178,N_2590,N_2930);
or UO_179 (O_179,N_2895,N_2988);
nor UO_180 (O_180,N_2847,N_2710);
xor UO_181 (O_181,N_2665,N_2789);
and UO_182 (O_182,N_2945,N_2640);
xnor UO_183 (O_183,N_2833,N_2791);
nand UO_184 (O_184,N_2792,N_2596);
xnor UO_185 (O_185,N_2805,N_2987);
xnor UO_186 (O_186,N_2894,N_2803);
xnor UO_187 (O_187,N_2744,N_2874);
nor UO_188 (O_188,N_2540,N_2981);
nand UO_189 (O_189,N_2619,N_2969);
xnor UO_190 (O_190,N_2572,N_2719);
nor UO_191 (O_191,N_2583,N_2519);
or UO_192 (O_192,N_2580,N_2599);
or UO_193 (O_193,N_2506,N_2998);
xnor UO_194 (O_194,N_2976,N_2934);
xnor UO_195 (O_195,N_2595,N_2836);
and UO_196 (O_196,N_2542,N_2779);
or UO_197 (O_197,N_2943,N_2567);
and UO_198 (O_198,N_2799,N_2760);
or UO_199 (O_199,N_2647,N_2928);
and UO_200 (O_200,N_2543,N_2644);
or UO_201 (O_201,N_2796,N_2782);
or UO_202 (O_202,N_2653,N_2822);
or UO_203 (O_203,N_2552,N_2774);
and UO_204 (O_204,N_2752,N_2546);
and UO_205 (O_205,N_2932,N_2522);
nand UO_206 (O_206,N_2971,N_2766);
and UO_207 (O_207,N_2787,N_2999);
and UO_208 (O_208,N_2906,N_2997);
and UO_209 (O_209,N_2966,N_2559);
nor UO_210 (O_210,N_2711,N_2843);
and UO_211 (O_211,N_2532,N_2661);
xor UO_212 (O_212,N_2876,N_2884);
or UO_213 (O_213,N_2502,N_2713);
nor UO_214 (O_214,N_2586,N_2972);
nand UO_215 (O_215,N_2712,N_2602);
nor UO_216 (O_216,N_2863,N_2666);
and UO_217 (O_217,N_2554,N_2553);
xnor UO_218 (O_218,N_2871,N_2728);
nand UO_219 (O_219,N_2883,N_2925);
nor UO_220 (O_220,N_2862,N_2684);
nand UO_221 (O_221,N_2699,N_2593);
and UO_222 (O_222,N_2692,N_2582);
nand UO_223 (O_223,N_2840,N_2865);
and UO_224 (O_224,N_2725,N_2565);
or UO_225 (O_225,N_2733,N_2503);
xnor UO_226 (O_226,N_2869,N_2890);
or UO_227 (O_227,N_2773,N_2700);
nor UO_228 (O_228,N_2767,N_2732);
and UO_229 (O_229,N_2741,N_2793);
and UO_230 (O_230,N_2800,N_2731);
nand UO_231 (O_231,N_2970,N_2834);
nor UO_232 (O_232,N_2924,N_2632);
nor UO_233 (O_233,N_2573,N_2835);
nand UO_234 (O_234,N_2510,N_2548);
nor UO_235 (O_235,N_2740,N_2561);
or UO_236 (O_236,N_2716,N_2635);
or UO_237 (O_237,N_2845,N_2721);
xor UO_238 (O_238,N_2915,N_2765);
xnor UO_239 (O_239,N_2706,N_2982);
or UO_240 (O_240,N_2581,N_2677);
and UO_241 (O_241,N_2771,N_2841);
nor UO_242 (O_242,N_2651,N_2905);
nor UO_243 (O_243,N_2990,N_2942);
or UO_244 (O_244,N_2897,N_2549);
or UO_245 (O_245,N_2809,N_2907);
nand UO_246 (O_246,N_2768,N_2709);
and UO_247 (O_247,N_2678,N_2825);
or UO_248 (O_248,N_2929,N_2909);
nor UO_249 (O_249,N_2558,N_2615);
and UO_250 (O_250,N_2725,N_2623);
and UO_251 (O_251,N_2801,N_2671);
nor UO_252 (O_252,N_2739,N_2650);
xnor UO_253 (O_253,N_2937,N_2771);
nand UO_254 (O_254,N_2799,N_2642);
and UO_255 (O_255,N_2503,N_2585);
nor UO_256 (O_256,N_2557,N_2893);
or UO_257 (O_257,N_2532,N_2616);
nand UO_258 (O_258,N_2886,N_2832);
or UO_259 (O_259,N_2825,N_2603);
nor UO_260 (O_260,N_2880,N_2656);
nor UO_261 (O_261,N_2897,N_2961);
nand UO_262 (O_262,N_2627,N_2932);
and UO_263 (O_263,N_2759,N_2585);
and UO_264 (O_264,N_2577,N_2882);
nand UO_265 (O_265,N_2747,N_2845);
and UO_266 (O_266,N_2985,N_2631);
xor UO_267 (O_267,N_2705,N_2709);
or UO_268 (O_268,N_2805,N_2871);
and UO_269 (O_269,N_2896,N_2584);
nor UO_270 (O_270,N_2831,N_2609);
nor UO_271 (O_271,N_2696,N_2633);
and UO_272 (O_272,N_2706,N_2864);
nor UO_273 (O_273,N_2961,N_2587);
or UO_274 (O_274,N_2803,N_2771);
or UO_275 (O_275,N_2973,N_2991);
and UO_276 (O_276,N_2940,N_2690);
xnor UO_277 (O_277,N_2535,N_2750);
nand UO_278 (O_278,N_2978,N_2718);
nor UO_279 (O_279,N_2942,N_2558);
nor UO_280 (O_280,N_2745,N_2677);
or UO_281 (O_281,N_2623,N_2752);
nand UO_282 (O_282,N_2685,N_2598);
nand UO_283 (O_283,N_2778,N_2904);
nand UO_284 (O_284,N_2763,N_2549);
or UO_285 (O_285,N_2571,N_2815);
or UO_286 (O_286,N_2863,N_2758);
nor UO_287 (O_287,N_2852,N_2990);
nor UO_288 (O_288,N_2815,N_2752);
xnor UO_289 (O_289,N_2648,N_2806);
or UO_290 (O_290,N_2765,N_2867);
and UO_291 (O_291,N_2735,N_2861);
and UO_292 (O_292,N_2888,N_2878);
and UO_293 (O_293,N_2506,N_2693);
and UO_294 (O_294,N_2728,N_2655);
and UO_295 (O_295,N_2624,N_2852);
nand UO_296 (O_296,N_2643,N_2836);
nor UO_297 (O_297,N_2958,N_2886);
nand UO_298 (O_298,N_2733,N_2529);
or UO_299 (O_299,N_2768,N_2704);
nor UO_300 (O_300,N_2545,N_2636);
nand UO_301 (O_301,N_2809,N_2799);
nand UO_302 (O_302,N_2678,N_2888);
nor UO_303 (O_303,N_2640,N_2513);
xnor UO_304 (O_304,N_2640,N_2911);
nand UO_305 (O_305,N_2964,N_2985);
nor UO_306 (O_306,N_2799,N_2775);
and UO_307 (O_307,N_2590,N_2685);
nand UO_308 (O_308,N_2991,N_2668);
or UO_309 (O_309,N_2608,N_2927);
or UO_310 (O_310,N_2979,N_2509);
nand UO_311 (O_311,N_2650,N_2841);
nand UO_312 (O_312,N_2776,N_2641);
and UO_313 (O_313,N_2583,N_2717);
xnor UO_314 (O_314,N_2514,N_2811);
or UO_315 (O_315,N_2849,N_2573);
nor UO_316 (O_316,N_2817,N_2566);
xnor UO_317 (O_317,N_2833,N_2691);
nand UO_318 (O_318,N_2649,N_2851);
or UO_319 (O_319,N_2813,N_2788);
or UO_320 (O_320,N_2829,N_2976);
xnor UO_321 (O_321,N_2706,N_2541);
xnor UO_322 (O_322,N_2514,N_2805);
or UO_323 (O_323,N_2916,N_2793);
or UO_324 (O_324,N_2857,N_2945);
or UO_325 (O_325,N_2934,N_2706);
nand UO_326 (O_326,N_2526,N_2900);
nor UO_327 (O_327,N_2746,N_2943);
nand UO_328 (O_328,N_2781,N_2644);
or UO_329 (O_329,N_2869,N_2534);
nor UO_330 (O_330,N_2595,N_2664);
xor UO_331 (O_331,N_2665,N_2535);
or UO_332 (O_332,N_2855,N_2959);
or UO_333 (O_333,N_2855,N_2588);
or UO_334 (O_334,N_2595,N_2920);
nand UO_335 (O_335,N_2984,N_2500);
and UO_336 (O_336,N_2779,N_2776);
and UO_337 (O_337,N_2572,N_2542);
nand UO_338 (O_338,N_2704,N_2663);
or UO_339 (O_339,N_2776,N_2664);
nand UO_340 (O_340,N_2760,N_2751);
nand UO_341 (O_341,N_2807,N_2845);
nand UO_342 (O_342,N_2740,N_2812);
nor UO_343 (O_343,N_2841,N_2840);
xor UO_344 (O_344,N_2774,N_2780);
or UO_345 (O_345,N_2503,N_2630);
or UO_346 (O_346,N_2691,N_2567);
and UO_347 (O_347,N_2617,N_2953);
nor UO_348 (O_348,N_2676,N_2768);
nand UO_349 (O_349,N_2883,N_2545);
xor UO_350 (O_350,N_2594,N_2875);
or UO_351 (O_351,N_2561,N_2986);
or UO_352 (O_352,N_2643,N_2660);
xor UO_353 (O_353,N_2589,N_2617);
xor UO_354 (O_354,N_2668,N_2706);
nor UO_355 (O_355,N_2722,N_2701);
nand UO_356 (O_356,N_2616,N_2526);
xnor UO_357 (O_357,N_2590,N_2888);
nor UO_358 (O_358,N_2523,N_2532);
and UO_359 (O_359,N_2641,N_2764);
nor UO_360 (O_360,N_2583,N_2679);
nand UO_361 (O_361,N_2941,N_2662);
and UO_362 (O_362,N_2840,N_2769);
and UO_363 (O_363,N_2548,N_2650);
xor UO_364 (O_364,N_2581,N_2657);
or UO_365 (O_365,N_2905,N_2863);
or UO_366 (O_366,N_2709,N_2614);
and UO_367 (O_367,N_2593,N_2652);
nor UO_368 (O_368,N_2563,N_2613);
nand UO_369 (O_369,N_2653,N_2976);
nand UO_370 (O_370,N_2855,N_2634);
xor UO_371 (O_371,N_2719,N_2766);
nand UO_372 (O_372,N_2657,N_2505);
nor UO_373 (O_373,N_2965,N_2653);
and UO_374 (O_374,N_2908,N_2592);
nor UO_375 (O_375,N_2574,N_2613);
or UO_376 (O_376,N_2663,N_2734);
or UO_377 (O_377,N_2535,N_2852);
nor UO_378 (O_378,N_2985,N_2617);
and UO_379 (O_379,N_2825,N_2793);
and UO_380 (O_380,N_2903,N_2813);
or UO_381 (O_381,N_2883,N_2736);
or UO_382 (O_382,N_2709,N_2748);
nor UO_383 (O_383,N_2930,N_2951);
nand UO_384 (O_384,N_2919,N_2665);
nand UO_385 (O_385,N_2562,N_2699);
or UO_386 (O_386,N_2519,N_2935);
and UO_387 (O_387,N_2581,N_2501);
nor UO_388 (O_388,N_2512,N_2525);
and UO_389 (O_389,N_2934,N_2874);
and UO_390 (O_390,N_2647,N_2753);
xor UO_391 (O_391,N_2580,N_2617);
or UO_392 (O_392,N_2959,N_2962);
and UO_393 (O_393,N_2833,N_2819);
nor UO_394 (O_394,N_2656,N_2568);
xor UO_395 (O_395,N_2523,N_2700);
and UO_396 (O_396,N_2913,N_2773);
or UO_397 (O_397,N_2769,N_2511);
xor UO_398 (O_398,N_2691,N_2892);
nor UO_399 (O_399,N_2593,N_2795);
nor UO_400 (O_400,N_2766,N_2733);
xor UO_401 (O_401,N_2526,N_2767);
nor UO_402 (O_402,N_2706,N_2590);
nand UO_403 (O_403,N_2561,N_2581);
or UO_404 (O_404,N_2533,N_2863);
and UO_405 (O_405,N_2893,N_2877);
xor UO_406 (O_406,N_2818,N_2914);
nor UO_407 (O_407,N_2888,N_2989);
nor UO_408 (O_408,N_2689,N_2605);
nand UO_409 (O_409,N_2951,N_2633);
nand UO_410 (O_410,N_2924,N_2928);
nand UO_411 (O_411,N_2599,N_2754);
xnor UO_412 (O_412,N_2957,N_2834);
nand UO_413 (O_413,N_2723,N_2510);
nor UO_414 (O_414,N_2513,N_2616);
xnor UO_415 (O_415,N_2723,N_2846);
nand UO_416 (O_416,N_2875,N_2890);
nand UO_417 (O_417,N_2791,N_2983);
and UO_418 (O_418,N_2922,N_2515);
nor UO_419 (O_419,N_2979,N_2586);
and UO_420 (O_420,N_2563,N_2634);
nand UO_421 (O_421,N_2689,N_2980);
or UO_422 (O_422,N_2523,N_2508);
nand UO_423 (O_423,N_2743,N_2544);
xnor UO_424 (O_424,N_2622,N_2806);
and UO_425 (O_425,N_2943,N_2823);
or UO_426 (O_426,N_2523,N_2997);
nand UO_427 (O_427,N_2814,N_2852);
nand UO_428 (O_428,N_2574,N_2583);
and UO_429 (O_429,N_2573,N_2585);
or UO_430 (O_430,N_2806,N_2511);
nand UO_431 (O_431,N_2565,N_2586);
nand UO_432 (O_432,N_2987,N_2861);
nor UO_433 (O_433,N_2573,N_2867);
nor UO_434 (O_434,N_2501,N_2547);
nand UO_435 (O_435,N_2817,N_2725);
and UO_436 (O_436,N_2505,N_2937);
nand UO_437 (O_437,N_2637,N_2502);
nor UO_438 (O_438,N_2895,N_2740);
nor UO_439 (O_439,N_2763,N_2946);
or UO_440 (O_440,N_2887,N_2703);
nand UO_441 (O_441,N_2787,N_2767);
and UO_442 (O_442,N_2593,N_2980);
nor UO_443 (O_443,N_2807,N_2601);
and UO_444 (O_444,N_2508,N_2629);
or UO_445 (O_445,N_2897,N_2928);
nand UO_446 (O_446,N_2866,N_2802);
nand UO_447 (O_447,N_2629,N_2511);
xor UO_448 (O_448,N_2800,N_2545);
and UO_449 (O_449,N_2899,N_2696);
nor UO_450 (O_450,N_2850,N_2562);
xor UO_451 (O_451,N_2810,N_2848);
nand UO_452 (O_452,N_2603,N_2614);
and UO_453 (O_453,N_2637,N_2917);
or UO_454 (O_454,N_2974,N_2841);
nand UO_455 (O_455,N_2989,N_2981);
or UO_456 (O_456,N_2933,N_2537);
nand UO_457 (O_457,N_2688,N_2611);
nand UO_458 (O_458,N_2503,N_2706);
nor UO_459 (O_459,N_2774,N_2584);
nor UO_460 (O_460,N_2809,N_2539);
xnor UO_461 (O_461,N_2719,N_2951);
nand UO_462 (O_462,N_2615,N_2628);
or UO_463 (O_463,N_2526,N_2784);
nand UO_464 (O_464,N_2632,N_2939);
or UO_465 (O_465,N_2567,N_2769);
and UO_466 (O_466,N_2678,N_2512);
and UO_467 (O_467,N_2505,N_2599);
nor UO_468 (O_468,N_2955,N_2634);
and UO_469 (O_469,N_2755,N_2759);
nor UO_470 (O_470,N_2860,N_2886);
and UO_471 (O_471,N_2820,N_2714);
xnor UO_472 (O_472,N_2943,N_2691);
or UO_473 (O_473,N_2523,N_2769);
nor UO_474 (O_474,N_2795,N_2553);
or UO_475 (O_475,N_2889,N_2956);
xor UO_476 (O_476,N_2711,N_2695);
and UO_477 (O_477,N_2875,N_2553);
and UO_478 (O_478,N_2656,N_2715);
xnor UO_479 (O_479,N_2735,N_2654);
nand UO_480 (O_480,N_2722,N_2902);
or UO_481 (O_481,N_2999,N_2962);
xor UO_482 (O_482,N_2918,N_2608);
and UO_483 (O_483,N_2967,N_2636);
nand UO_484 (O_484,N_2922,N_2761);
xor UO_485 (O_485,N_2859,N_2915);
and UO_486 (O_486,N_2534,N_2511);
nor UO_487 (O_487,N_2529,N_2739);
xnor UO_488 (O_488,N_2763,N_2909);
or UO_489 (O_489,N_2576,N_2951);
or UO_490 (O_490,N_2659,N_2595);
xnor UO_491 (O_491,N_2711,N_2571);
or UO_492 (O_492,N_2792,N_2567);
nor UO_493 (O_493,N_2628,N_2886);
or UO_494 (O_494,N_2984,N_2583);
nor UO_495 (O_495,N_2832,N_2624);
nor UO_496 (O_496,N_2755,N_2530);
nand UO_497 (O_497,N_2921,N_2944);
xnor UO_498 (O_498,N_2687,N_2731);
nand UO_499 (O_499,N_2605,N_2546);
endmodule