module basic_2000_20000_2500_5_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1266,In_1771);
or U1 (N_1,In_1631,In_873);
and U2 (N_2,In_319,In_1196);
nor U3 (N_3,In_368,In_1650);
nand U4 (N_4,In_1788,In_340);
nand U5 (N_5,In_1523,In_1529);
or U6 (N_6,In_54,In_1011);
or U7 (N_7,In_1983,In_1894);
nand U8 (N_8,In_1378,In_554);
nand U9 (N_9,In_1883,In_1527);
nand U10 (N_10,In_432,In_1211);
and U11 (N_11,In_817,In_1720);
nand U12 (N_12,In_784,In_925);
nor U13 (N_13,In_737,In_1175);
nand U14 (N_14,In_1094,In_574);
or U15 (N_15,In_95,In_1706);
and U16 (N_16,In_1025,In_639);
nand U17 (N_17,In_646,In_1560);
and U18 (N_18,In_549,In_1925);
or U19 (N_19,In_662,In_1200);
and U20 (N_20,In_1626,In_1831);
nor U21 (N_21,In_423,In_1235);
and U22 (N_22,In_1362,In_722);
and U23 (N_23,In_1046,In_78);
and U24 (N_24,In_1402,In_427);
and U25 (N_25,In_1098,In_1822);
or U26 (N_26,In_1816,In_756);
nand U27 (N_27,In_422,In_1619);
nand U28 (N_28,In_292,In_1132);
and U29 (N_29,In_1153,In_1045);
nor U30 (N_30,In_1877,In_260);
nand U31 (N_31,In_295,In_1798);
nor U32 (N_32,In_1099,In_668);
nor U33 (N_33,In_39,In_1762);
nor U34 (N_34,In_1286,In_471);
nand U35 (N_35,In_989,In_55);
or U36 (N_36,In_526,In_715);
or U37 (N_37,In_1353,In_1616);
and U38 (N_38,In_46,In_410);
or U39 (N_39,In_1791,In_1693);
nor U40 (N_40,In_1172,In_919);
nand U41 (N_41,In_1360,In_659);
nand U42 (N_42,In_564,In_1775);
and U43 (N_43,In_28,In_491);
and U44 (N_44,In_1740,In_1916);
nand U45 (N_45,In_941,In_1888);
or U46 (N_46,In_1428,In_377);
nor U47 (N_47,In_1271,In_146);
nor U48 (N_48,In_591,In_839);
or U49 (N_49,In_1388,In_623);
nor U50 (N_50,In_515,In_987);
nor U51 (N_51,In_677,In_1371);
nand U52 (N_52,In_730,In_1670);
nand U53 (N_53,In_790,In_233);
or U54 (N_54,In_1760,In_495);
and U55 (N_55,In_1505,In_1151);
and U56 (N_56,In_1574,In_1569);
or U57 (N_57,In_198,In_996);
or U58 (N_58,In_1672,In_1677);
nor U59 (N_59,In_690,In_1189);
and U60 (N_60,In_80,In_1969);
nand U61 (N_61,In_56,In_398);
and U62 (N_62,In_1407,In_1023);
nor U63 (N_63,In_207,In_1159);
and U64 (N_64,In_434,In_889);
nand U65 (N_65,In_1448,In_986);
nand U66 (N_66,In_838,In_707);
and U67 (N_67,In_1756,In_1264);
nand U68 (N_68,In_540,In_1051);
or U69 (N_69,In_1870,In_345);
and U70 (N_70,In_940,In_261);
nor U71 (N_71,In_1814,In_878);
or U72 (N_72,In_264,In_1296);
and U73 (N_73,In_1783,In_1781);
nor U74 (N_74,In_1878,In_1803);
nand U75 (N_75,In_974,In_1735);
and U76 (N_76,In_252,In_185);
nand U77 (N_77,In_1795,In_809);
nor U78 (N_78,In_1589,In_1738);
nor U79 (N_79,In_590,In_792);
nand U80 (N_80,In_903,In_965);
and U81 (N_81,In_73,In_164);
and U82 (N_82,In_411,In_758);
nor U83 (N_83,In_812,In_1833);
nand U84 (N_84,In_1225,In_99);
nor U85 (N_85,In_1608,In_908);
nor U86 (N_86,In_875,In_40);
and U87 (N_87,In_76,In_301);
nor U88 (N_88,In_457,In_769);
nand U89 (N_89,In_430,In_504);
and U90 (N_90,In_1900,In_713);
or U91 (N_91,In_230,In_517);
and U92 (N_92,In_1800,In_1578);
and U93 (N_93,In_300,In_429);
nand U94 (N_94,In_244,In_1864);
and U95 (N_95,In_744,In_174);
nand U96 (N_96,In_886,In_1038);
or U97 (N_97,In_1852,In_1587);
and U98 (N_98,In_837,In_293);
or U99 (N_99,In_1949,In_197);
nand U100 (N_100,In_1862,In_213);
nand U101 (N_101,In_1824,In_716);
nand U102 (N_102,In_1807,In_961);
and U103 (N_103,In_81,In_1806);
xnor U104 (N_104,In_938,In_1968);
nor U105 (N_105,In_16,In_33);
and U106 (N_106,In_665,In_1328);
and U107 (N_107,In_1521,In_893);
nor U108 (N_108,In_1029,In_1964);
and U109 (N_109,In_957,In_1143);
nor U110 (N_110,In_1437,In_152);
and U111 (N_111,In_1996,In_1270);
or U112 (N_112,In_1936,In_426);
or U113 (N_113,In_832,In_1041);
and U114 (N_114,In_1630,In_881);
nand U115 (N_115,In_1239,In_802);
or U116 (N_116,In_787,In_982);
and U117 (N_117,In_414,In_236);
nor U118 (N_118,In_1674,In_1543);
nor U119 (N_119,In_1942,In_1333);
and U120 (N_120,In_1823,In_1145);
nor U121 (N_121,In_1203,In_329);
and U122 (N_122,In_587,In_543);
nand U123 (N_123,In_1343,In_1147);
nand U124 (N_124,In_1133,In_640);
and U125 (N_125,In_1963,In_1739);
nand U126 (N_126,In_1726,In_311);
and U127 (N_127,In_1403,In_1390);
nand U128 (N_128,In_914,In_1349);
or U129 (N_129,In_194,In_1982);
nand U130 (N_130,In_1861,In_406);
and U131 (N_131,In_1395,In_1931);
and U132 (N_132,In_5,In_303);
or U133 (N_133,In_1606,In_1231);
and U134 (N_134,In_1240,In_1979);
and U135 (N_135,In_419,In_454);
or U136 (N_136,In_1450,In_242);
nor U137 (N_137,In_496,In_992);
or U138 (N_138,In_958,In_1799);
or U139 (N_139,In_1742,In_420);
nor U140 (N_140,In_4,In_1267);
nor U141 (N_141,In_1697,In_1346);
nor U142 (N_142,In_1217,In_356);
nand U143 (N_143,In_1700,In_1042);
nand U144 (N_144,In_1792,In_1923);
or U145 (N_145,In_905,In_577);
nor U146 (N_146,In_202,In_281);
nor U147 (N_147,In_1386,In_1912);
or U148 (N_148,In_109,In_966);
nor U149 (N_149,In_970,In_1926);
or U150 (N_150,In_1306,In_972);
and U151 (N_151,In_1489,In_921);
nand U152 (N_152,In_1310,In_830);
xor U153 (N_153,In_1681,In_1398);
and U154 (N_154,In_1855,In_1929);
and U155 (N_155,In_1255,In_488);
nand U156 (N_156,In_1166,In_1503);
and U157 (N_157,In_876,In_1052);
or U158 (N_158,In_1617,In_527);
nand U159 (N_159,In_147,In_592);
nor U160 (N_160,In_387,In_1506);
or U161 (N_161,In_1120,In_1321);
nand U162 (N_162,In_1443,In_775);
nor U163 (N_163,In_1647,In_1854);
nand U164 (N_164,In_928,In_1640);
or U165 (N_165,In_1887,In_205);
nand U166 (N_166,In_456,In_685);
or U167 (N_167,In_1566,In_0);
or U168 (N_168,In_1810,In_1684);
nand U169 (N_169,In_476,In_1119);
nand U170 (N_170,In_1860,In_1063);
and U171 (N_171,In_1224,In_1076);
nand U172 (N_172,In_1898,In_20);
and U173 (N_173,In_1184,In_1113);
or U174 (N_174,In_859,In_150);
nor U175 (N_175,In_1307,In_177);
and U176 (N_176,In_1243,In_774);
nor U177 (N_177,In_666,In_7);
and U178 (N_178,In_1304,In_1478);
or U179 (N_179,In_1641,In_308);
and U180 (N_180,In_1208,In_1138);
nand U181 (N_181,In_1975,In_753);
or U182 (N_182,In_1100,In_1185);
nor U183 (N_183,In_887,In_1385);
and U184 (N_184,In_800,In_1117);
nand U185 (N_185,In_464,In_976);
nor U186 (N_186,In_489,In_34);
or U187 (N_187,In_1858,In_641);
nand U188 (N_188,In_117,In_1556);
or U189 (N_189,In_127,In_663);
and U190 (N_190,In_1469,In_1376);
and U191 (N_191,In_224,In_118);
nand U192 (N_192,In_1876,In_1055);
xnor U193 (N_193,In_1363,In_1223);
nand U194 (N_194,In_783,In_371);
or U195 (N_195,In_1186,In_386);
nand U196 (N_196,In_614,In_1790);
xnor U197 (N_197,In_952,In_1381);
or U198 (N_198,In_497,In_693);
nand U199 (N_199,In_253,In_733);
nand U200 (N_200,In_959,In_612);
nor U201 (N_201,In_1789,In_206);
or U202 (N_202,In_1519,In_669);
and U203 (N_203,In_1541,In_954);
nand U204 (N_204,In_739,In_296);
or U205 (N_205,In_1970,In_1733);
nor U206 (N_206,In_1897,In_1655);
nor U207 (N_207,In_1911,In_581);
and U208 (N_208,In_1188,In_788);
and U209 (N_209,In_1993,In_107);
nor U210 (N_210,In_535,In_53);
or U211 (N_211,In_232,In_359);
and U212 (N_212,In_1127,In_1199);
nor U213 (N_213,In_1167,In_1462);
nor U214 (N_214,In_776,In_872);
or U215 (N_215,In_1347,In_1471);
or U216 (N_216,In_1397,In_858);
and U217 (N_217,In_1338,In_828);
nand U218 (N_218,In_979,In_636);
and U219 (N_219,In_1744,In_948);
and U220 (N_220,In_1031,In_1490);
nand U221 (N_221,In_378,In_735);
or U222 (N_222,In_1027,In_151);
and U223 (N_223,In_315,In_1033);
or U224 (N_224,In_1542,In_1429);
nor U225 (N_225,In_1313,In_1703);
and U226 (N_226,In_1857,In_686);
nor U227 (N_227,In_1772,In_1054);
nand U228 (N_228,In_654,In_168);
or U229 (N_229,In_741,In_1895);
and U230 (N_230,In_1538,In_1609);
or U231 (N_231,In_1614,In_649);
nand U232 (N_232,In_440,In_1302);
and U233 (N_233,In_1518,In_1194);
and U234 (N_234,In_523,In_184);
nand U235 (N_235,In_1358,In_1603);
and U236 (N_236,In_697,In_1874);
nor U237 (N_237,In_1575,In_826);
nand U238 (N_238,In_448,In_1905);
nand U239 (N_239,In_1252,In_1776);
nand U240 (N_240,In_569,In_915);
and U241 (N_241,In_1572,In_169);
or U242 (N_242,In_115,In_438);
nor U243 (N_243,In_918,In_1474);
and U244 (N_244,In_607,In_819);
nand U245 (N_245,In_337,In_97);
and U246 (N_246,In_1125,In_104);
nor U247 (N_247,In_729,In_791);
nand U248 (N_248,In_288,In_1558);
xor U249 (N_249,In_1280,In_765);
and U250 (N_250,In_1426,In_468);
nand U251 (N_251,In_1548,In_1263);
nand U252 (N_252,In_1247,In_25);
nand U253 (N_253,In_1372,In_144);
and U254 (N_254,In_1201,In_1192);
nand U255 (N_255,In_433,In_745);
or U256 (N_256,In_1559,In_1418);
or U257 (N_257,In_96,In_1427);
nand U258 (N_258,In_947,In_1014);
nor U259 (N_259,In_1715,In_347);
nor U260 (N_260,In_1535,In_1393);
nand U261 (N_261,In_1847,In_1815);
nand U262 (N_262,In_611,In_653);
or U263 (N_263,In_1761,In_231);
nand U264 (N_264,In_1112,In_201);
or U265 (N_265,In_1514,In_1434);
nor U266 (N_266,In_978,In_1000);
and U267 (N_267,In_1896,In_1105);
nand U268 (N_268,In_1168,In_211);
nand U269 (N_269,In_1499,In_567);
and U270 (N_270,In_675,In_1193);
or U271 (N_271,In_1727,In_650);
and U272 (N_272,In_498,In_173);
nor U273 (N_273,In_950,In_1160);
and U274 (N_274,In_1348,In_1881);
nand U275 (N_275,In_137,In_1191);
or U276 (N_276,In_1562,In_1865);
nand U277 (N_277,In_332,In_810);
or U278 (N_278,In_1851,In_469);
or U279 (N_279,In_182,In_1786);
or U280 (N_280,In_1632,In_1659);
nor U281 (N_281,In_862,In_1750);
or U282 (N_282,In_684,In_679);
nor U283 (N_283,In_924,In_576);
nor U284 (N_284,In_126,In_548);
and U285 (N_285,In_743,In_1277);
or U286 (N_286,In_840,In_357);
and U287 (N_287,In_1141,In_111);
and U288 (N_288,In_1643,In_1974);
nand U289 (N_289,In_1079,In_1707);
nor U290 (N_290,In_1316,In_1417);
nand U291 (N_291,In_1352,In_267);
or U292 (N_292,In_1340,In_361);
or U293 (N_293,In_1732,In_1162);
or U294 (N_294,In_374,In_1940);
and U295 (N_295,In_843,In_1216);
nor U296 (N_296,In_617,In_683);
nor U297 (N_297,In_1777,In_1717);
nand U298 (N_298,In_1992,In_1177);
and U299 (N_299,In_88,In_1275);
or U300 (N_300,In_102,In_171);
and U301 (N_301,In_555,In_1869);
or U302 (N_302,In_1526,In_1481);
and U303 (N_303,In_196,In_1743);
nor U304 (N_304,In_798,In_139);
nand U305 (N_305,In_968,In_135);
nand U306 (N_306,In_1586,In_1297);
or U307 (N_307,In_1749,In_1966);
nor U308 (N_308,In_140,In_134);
or U309 (N_309,In_494,In_541);
nand U310 (N_310,In_1003,In_1121);
nor U311 (N_311,In_375,In_711);
and U312 (N_312,In_997,In_1272);
and U313 (N_313,In_983,In_1531);
nand U314 (N_314,In_583,In_853);
or U315 (N_315,In_1710,In_1910);
and U316 (N_316,In_676,In_106);
or U317 (N_317,In_1662,In_391);
or U318 (N_318,In_1164,In_294);
nor U319 (N_319,In_1924,In_1797);
or U320 (N_320,In_1600,In_935);
and U321 (N_321,In_1476,In_1638);
nand U322 (N_322,In_1330,In_1350);
and U323 (N_323,In_1695,In_1126);
or U324 (N_324,In_1008,In_91);
nand U325 (N_325,In_1241,In_333);
nand U326 (N_326,In_1253,In_794);
nand U327 (N_327,In_1889,In_596);
nand U328 (N_328,In_425,In_1202);
or U329 (N_329,In_586,In_1157);
and U330 (N_330,In_1987,In_865);
nor U331 (N_331,In_121,In_153);
and U332 (N_332,In_394,In_48);
and U333 (N_333,In_1299,In_352);
nand U334 (N_334,In_136,In_1206);
nand U335 (N_335,In_1229,In_483);
or U336 (N_336,In_277,In_71);
nand U337 (N_337,In_1294,In_1509);
nor U338 (N_338,In_786,In_1325);
and U339 (N_339,In_738,In_1366);
nand U340 (N_340,In_524,In_1913);
nor U341 (N_341,In_836,In_1689);
and U342 (N_342,In_354,In_750);
and U343 (N_343,In_299,In_1292);
nor U344 (N_344,In_412,In_801);
and U345 (N_345,In_176,In_472);
and U346 (N_346,In_610,In_365);
nor U347 (N_347,In_1696,In_1955);
nor U348 (N_348,In_23,In_1920);
or U349 (N_349,In_240,In_1856);
and U350 (N_350,In_317,In_1699);
and U351 (N_351,In_955,In_1849);
or U352 (N_352,In_291,In_1702);
and U353 (N_353,In_272,In_1485);
or U354 (N_354,In_871,In_1892);
nand U355 (N_355,In_626,In_1839);
nand U356 (N_356,In_1238,In_1595);
or U357 (N_357,In_1675,In_1718);
nand U358 (N_358,In_1219,In_1886);
xnor U359 (N_359,In_846,In_537);
nor U360 (N_360,In_521,In_1904);
nor U361 (N_361,In_1615,In_235);
nand U362 (N_362,In_1698,In_874);
nand U363 (N_363,In_1914,In_1315);
nand U364 (N_364,In_1467,In_129);
nand U365 (N_365,In_1812,In_485);
nand U366 (N_366,In_1731,In_251);
and U367 (N_367,In_35,In_951);
and U368 (N_368,In_1724,In_1273);
and U369 (N_369,In_1950,In_1947);
or U370 (N_370,In_673,In_1137);
nor U371 (N_371,In_700,In_258);
and U372 (N_372,In_1767,In_1285);
or U373 (N_373,In_712,In_212);
nor U374 (N_374,In_460,In_239);
and U375 (N_375,In_710,In_1502);
and U376 (N_376,In_1629,In_1818);
nand U377 (N_377,In_1553,In_228);
or U378 (N_378,In_1604,In_937);
and U379 (N_379,In_1808,In_1435);
nand U380 (N_380,In_268,In_1922);
nor U381 (N_381,In_195,In_706);
and U382 (N_382,In_1639,In_1667);
nor U383 (N_383,In_692,In_533);
nor U384 (N_384,In_330,In_1415);
nor U385 (N_385,In_1658,In_175);
nor U386 (N_386,In_1086,In_852);
or U387 (N_387,In_276,In_1071);
or U388 (N_388,In_519,In_306);
or U389 (N_389,In_1563,In_1375);
nand U390 (N_390,In_864,In_825);
and U391 (N_391,In_1399,In_680);
or U392 (N_392,In_1520,In_8);
nand U393 (N_393,In_248,In_298);
nor U394 (N_394,In_566,In_1006);
and U395 (N_395,In_1734,In_1532);
nor U396 (N_396,In_1544,In_1062);
and U397 (N_397,In_1622,In_270);
nand U398 (N_398,In_719,In_1533);
nand U399 (N_399,In_593,In_1317);
nor U400 (N_400,In_63,In_1420);
nand U401 (N_401,In_397,In_200);
nor U402 (N_402,In_1268,In_1962);
or U403 (N_403,In_1766,In_348);
nand U404 (N_404,In_477,In_1218);
xnor U405 (N_405,In_1721,In_1089);
nand U406 (N_406,In_1163,In_854);
nor U407 (N_407,In_418,In_1653);
nor U408 (N_408,In_619,In_1915);
nand U409 (N_409,In_1233,In_1577);
or U410 (N_410,In_934,In_486);
nand U411 (N_411,In_725,In_116);
and U412 (N_412,In_1369,In_94);
nand U413 (N_413,In_280,In_1276);
nor U414 (N_414,In_560,In_304);
and U415 (N_415,In_732,In_130);
nand U416 (N_416,In_1377,In_1396);
nand U417 (N_417,In_1154,In_1165);
nor U418 (N_418,In_1525,In_1780);
nand U419 (N_419,In_500,In_1303);
or U420 (N_420,In_977,In_1278);
or U421 (N_421,In_1136,In_1130);
or U422 (N_422,In_782,In_696);
and U423 (N_423,In_1344,In_1599);
nor U424 (N_424,In_1053,In_621);
or U425 (N_425,In_1444,In_1844);
nand U426 (N_426,In_648,In_1879);
nand U427 (N_427,In_154,In_1097);
nand U428 (N_428,In_841,In_582);
nor U429 (N_429,In_170,In_9);
nand U430 (N_430,In_589,In_811);
nor U431 (N_431,In_165,In_807);
nand U432 (N_432,In_1180,In_559);
and U433 (N_433,In_1537,In_770);
nand U434 (N_434,In_1934,In_1183);
or U435 (N_435,In_1064,In_1242);
or U436 (N_436,In_1389,In_892);
and U437 (N_437,In_1634,In_1414);
nor U438 (N_438,In_1708,In_1146);
nor U439 (N_439,In_38,In_192);
and U440 (N_440,In_764,In_746);
or U441 (N_441,In_1179,In_1416);
and U442 (N_442,In_704,In_538);
nand U443 (N_443,In_49,In_1981);
nand U444 (N_444,In_806,In_1582);
and U445 (N_445,In_1794,In_1020);
and U446 (N_446,In_731,In_671);
and U447 (N_447,In_831,In_1227);
and U448 (N_448,In_1331,In_1867);
nor U449 (N_449,In_1501,In_1998);
and U450 (N_450,In_1090,In_687);
nand U451 (N_451,In_1339,In_1909);
and U452 (N_452,In_241,In_1666);
or U453 (N_453,In_695,In_1770);
nor U454 (N_454,In_1436,In_578);
nor U455 (N_455,In_1468,In_969);
and U456 (N_456,In_736,In_190);
nor U457 (N_457,In_14,In_1825);
nand U458 (N_458,In_606,In_1588);
nand U459 (N_459,In_1309,In_131);
nor U460 (N_460,In_1866,In_1101);
and U461 (N_461,In_199,In_752);
nor U462 (N_462,In_166,In_1026);
nor U463 (N_463,In_534,In_149);
and U464 (N_464,In_156,In_322);
or U465 (N_465,In_1753,In_628);
and U466 (N_466,In_1805,In_338);
and U467 (N_467,In_656,In_1106);
or U468 (N_468,In_1212,In_1237);
and U469 (N_469,In_1013,In_1965);
nand U470 (N_470,In_113,In_145);
nor U471 (N_471,In_845,In_1832);
and U472 (N_472,In_442,In_247);
and U473 (N_473,In_1128,In_1084);
or U474 (N_474,In_1334,In_734);
nand U475 (N_475,In_393,In_645);
and U476 (N_476,In_1848,In_326);
nor U477 (N_477,In_1406,In_1534);
nand U478 (N_478,In_1230,In_1332);
nand U479 (N_479,In_237,In_1061);
nor U480 (N_480,In_1073,In_1295);
nor U481 (N_481,In_1561,In_1500);
or U482 (N_482,In_755,In_681);
nand U483 (N_483,In_1082,In_1868);
nor U484 (N_484,In_813,In_1826);
nand U485 (N_485,In_1058,In_1774);
nor U486 (N_486,In_1686,In_848);
and U487 (N_487,In_1283,In_161);
or U488 (N_488,In_920,In_463);
nor U489 (N_489,In_22,In_1755);
or U490 (N_490,In_1769,In_1536);
nor U491 (N_491,In_98,In_1827);
nand U492 (N_492,In_1453,In_60);
and U493 (N_493,In_209,In_405);
or U494 (N_494,In_1960,In_1075);
or U495 (N_495,In_1540,In_1077);
and U496 (N_496,In_401,In_763);
xor U497 (N_497,In_1254,In_835);
nor U498 (N_498,In_1005,In_219);
nand U499 (N_499,In_1232,In_866);
or U500 (N_500,In_1510,In_52);
or U501 (N_501,In_761,In_1597);
nor U502 (N_502,In_818,In_1859);
or U503 (N_503,In_363,In_327);
nand U504 (N_504,In_1447,In_1454);
nand U505 (N_505,In_1763,In_1907);
and U506 (N_506,In_1030,In_1438);
or U507 (N_507,In_309,In_1875);
nor U508 (N_508,In_620,In_451);
nor U509 (N_509,In_1871,In_1817);
nor U510 (N_510,In_1460,In_960);
and U511 (N_511,In_1694,In_1570);
nand U512 (N_512,In_1195,In_894);
or U513 (N_513,In_124,In_513);
nor U514 (N_514,In_571,In_629);
and U515 (N_515,In_1256,In_380);
or U516 (N_516,In_1988,In_625);
nand U517 (N_517,In_474,In_1382);
and U518 (N_518,In_870,In_1311);
nor U519 (N_519,In_85,In_1828);
nand U520 (N_520,In_562,In_1679);
or U521 (N_521,In_286,In_931);
or U522 (N_522,In_565,In_369);
or U523 (N_523,In_217,In_1007);
and U524 (N_524,In_1746,In_324);
and U525 (N_525,In_29,In_1419);
nand U526 (N_526,In_32,In_318);
nand U527 (N_527,In_503,In_1989);
and U528 (N_528,In_1182,In_1972);
and U529 (N_529,In_608,In_1939);
nor U530 (N_530,In_180,In_1517);
nor U531 (N_531,In_1961,In_584);
or U532 (N_532,In_499,In_344);
or U533 (N_533,In_827,In_1504);
and U534 (N_534,In_1487,In_428);
and U535 (N_535,In_21,In_1752);
or U536 (N_536,In_1764,In_563);
nor U537 (N_537,In_1370,In_1048);
nand U538 (N_538,In_1901,In_1221);
nand U539 (N_539,In_87,In_895);
nand U540 (N_540,In_1169,In_1361);
or U541 (N_541,In_1085,In_1713);
nor U542 (N_542,In_1759,In_863);
nand U543 (N_543,In_1994,In_1104);
nor U544 (N_544,In_998,In_123);
and U545 (N_545,In_416,In_1282);
and U546 (N_546,In_778,In_528);
nand U547 (N_547,In_441,In_313);
nor U548 (N_548,In_598,In_1873);
nor U549 (N_549,In_1087,In_342);
or U550 (N_550,In_899,In_221);
and U551 (N_551,In_945,In_108);
and U552 (N_552,In_1837,In_1050);
or U553 (N_553,In_1722,In_1834);
or U554 (N_554,In_1945,In_302);
and U555 (N_555,In_532,In_349);
or U556 (N_556,In_1804,In_1657);
nor U557 (N_557,In_747,In_62);
nand U558 (N_558,In_366,In_1069);
nor U559 (N_559,In_600,In_1425);
and U560 (N_560,In_1486,In_964);
or U561 (N_561,In_907,In_1646);
and U562 (N_562,In_1301,In_529);
nor U563 (N_563,In_672,In_114);
nand U564 (N_564,In_803,In_514);
nor U565 (N_565,In_1457,In_1475);
or U566 (N_566,In_1635,In_984);
and U567 (N_567,In_1654,In_698);
nor U568 (N_568,In_229,In_1305);
nor U569 (N_569,In_61,In_748);
nor U570 (N_570,In_1312,In_1991);
nand U571 (N_571,In_446,In_218);
xnor U572 (N_572,In_1779,In_101);
and U573 (N_573,In_1433,In_1637);
nor U574 (N_574,In_1935,In_857);
or U575 (N_575,In_967,In_1651);
nor U576 (N_576,In_585,In_1472);
and U577 (N_577,In_1190,In_975);
nor U578 (N_578,In_1959,In_254);
and U579 (N_579,In_1809,In_1685);
or U580 (N_580,In_1730,In_289);
nand U581 (N_581,In_249,In_622);
and U582 (N_582,In_92,In_449);
or U583 (N_583,In_1441,In_1709);
nand U584 (N_584,In_847,In_1001);
nand U585 (N_585,In_721,In_1140);
and U586 (N_586,In_404,In_1142);
and U587 (N_587,In_1880,In_64);
and U588 (N_588,In_186,In_44);
nor U589 (N_589,In_929,In_962);
or U590 (N_590,In_1576,In_1259);
or U591 (N_591,In_100,In_651);
nor U592 (N_592,In_1284,In_407);
and U593 (N_593,In_1336,In_545);
and U594 (N_594,In_284,In_490);
nand U595 (N_595,In_1421,In_1209);
nor U596 (N_596,In_552,In_1581);
nor U597 (N_597,In_1511,In_904);
nand U598 (N_598,In_885,In_595);
nor U599 (N_599,In_1785,In_1044);
nor U600 (N_600,In_829,In_643);
nor U601 (N_601,In_1365,In_897);
xnor U602 (N_602,In_1096,In_1757);
or U603 (N_603,In_949,In_282);
or U604 (N_604,In_805,In_1683);
nor U605 (N_605,In_718,In_808);
or U606 (N_606,In_1289,In_1933);
nor U607 (N_607,In_204,In_1956);
nand U608 (N_608,In_1899,In_1768);
and U609 (N_609,In_994,In_985);
and U610 (N_610,In_1158,In_1110);
nor U611 (N_611,In_1778,In_1024);
nor U612 (N_612,In_1705,In_635);
nand U613 (N_613,In_1953,In_995);
or U614 (N_614,In_216,In_1327);
nand U615 (N_615,In_632,In_336);
and U616 (N_616,In_678,In_75);
or U617 (N_617,In_1279,In_594);
nor U618 (N_618,In_867,In_403);
nor U619 (N_619,In_1872,In_467);
nand U620 (N_620,In_1067,In_1287);
or U621 (N_621,In_896,In_1621);
nand U622 (N_622,In_547,In_346);
and U623 (N_623,In_384,In_1204);
nand U624 (N_624,In_1028,In_1236);
nor U625 (N_625,In_259,In_93);
or U626 (N_626,In_1149,In_1134);
nand U627 (N_627,In_409,In_392);
nor U628 (N_628,In_222,In_990);
nor U629 (N_629,In_265,In_1918);
or U630 (N_630,In_1585,In_634);
and U631 (N_631,In_312,In_6);
and U632 (N_632,In_1144,In_1494);
nand U633 (N_633,In_283,In_162);
nand U634 (N_634,In_30,In_1373);
nor U635 (N_635,In_1300,In_1567);
or U636 (N_636,In_1555,In_501);
nand U637 (N_637,In_551,In_910);
and U638 (N_638,In_492,In_142);
nand U639 (N_639,In_1628,In_1841);
and U640 (N_640,In_717,In_1329);
and U641 (N_641,In_1298,In_41);
and U642 (N_642,In_1115,In_728);
or U643 (N_643,In_633,In_714);
nor U644 (N_644,In_1488,In_1409);
nor U645 (N_645,In_1095,In_1384);
and U646 (N_646,In_455,In_1004);
xnor U647 (N_647,In_148,In_1919);
or U648 (N_648,In_1528,In_1356);
nor U649 (N_649,In_1430,In_1245);
nand U650 (N_650,In_553,In_160);
nor U651 (N_651,In_759,In_1564);
nand U652 (N_652,In_1123,In_1941);
nor U653 (N_653,In_630,In_1250);
or U654 (N_654,In_1712,In_814);
and U655 (N_655,In_143,In_210);
and U656 (N_656,In_273,In_466);
and U657 (N_657,In_1573,In_689);
nor U658 (N_658,In_1251,In_480);
or U659 (N_659,In_766,In_1043);
and U660 (N_660,In_155,In_1930);
and U661 (N_661,In_128,In_615);
or U662 (N_662,In_1820,In_66);
and U663 (N_663,In_708,In_522);
or U664 (N_664,In_50,In_305);
nor U665 (N_665,In_912,In_58);
nor U666 (N_666,In_74,In_879);
nor U667 (N_667,In_1440,In_59);
nand U668 (N_668,In_1265,In_1065);
and U669 (N_669,In_1937,In_988);
and U670 (N_670,In_447,In_367);
xnor U671 (N_671,In_223,In_926);
or U672 (N_672,In_1072,In_971);
nor U673 (N_673,In_1213,In_1728);
and U674 (N_674,In_382,In_536);
and U675 (N_675,In_1748,In_1884);
or U676 (N_676,In_57,In_1723);
nand U677 (N_677,In_402,In_1187);
and U678 (N_678,In_214,In_1037);
or U679 (N_679,In_597,In_1156);
nor U680 (N_680,In_355,In_1648);
or U681 (N_681,In_1131,In_1337);
nor U682 (N_682,In_256,In_509);
or U683 (N_683,In_1210,In_657);
or U684 (N_684,In_1161,In_1976);
nand U685 (N_685,In_178,In_2);
and U686 (N_686,In_942,In_1607);
nand U687 (N_687,In_82,In_1644);
nor U688 (N_688,In_795,In_450);
and U689 (N_689,In_1482,In_1459);
and U690 (N_690,In_1368,In_1971);
nand U691 (N_691,In_1326,In_478);
nor U692 (N_692,In_1422,In_1954);
or U693 (N_693,In_187,In_1611);
or U694 (N_694,In_705,In_1047);
nor U695 (N_695,In_1449,In_3);
and U696 (N_696,In_1584,In_1690);
xnor U697 (N_697,In_373,In_1034);
and U698 (N_698,In_579,In_557);
and U699 (N_699,In_624,In_385);
or U700 (N_700,In_424,In_158);
nor U701 (N_701,In_172,In_793);
or U702 (N_702,In_1678,In_285);
nor U703 (N_703,In_1627,In_1590);
nand U704 (N_704,In_1470,In_1171);
nor U705 (N_705,In_1802,In_435);
nand U706 (N_706,In_1946,In_1813);
or U707 (N_707,In_771,In_257);
and U708 (N_708,In_850,In_444);
and U709 (N_709,In_1261,In_520);
nand U710 (N_710,In_506,In_1921);
and U711 (N_711,In_24,In_266);
nand U712 (N_712,In_262,In_1010);
xor U713 (N_713,In_922,In_1244);
and U714 (N_714,In_660,In_507);
nand U715 (N_715,In_1341,In_502);
nand U716 (N_716,In_1623,In_1152);
nand U717 (N_717,In_781,In_1568);
or U718 (N_718,In_1663,In_816);
nand U719 (N_719,In_1656,In_882);
or U720 (N_720,In_1290,In_1484);
and U721 (N_721,In_1853,In_1092);
or U722 (N_722,In_1345,In_1701);
or U723 (N_723,In_1636,In_627);
nor U724 (N_724,In_923,In_530);
and U725 (N_725,In_1258,In_609);
and U726 (N_726,In_674,In_1458);
and U727 (N_727,In_1973,In_1122);
and U728 (N_728,In_880,In_601);
nor U729 (N_729,In_452,In_1580);
nand U730 (N_730,In_544,In_163);
or U731 (N_731,In_1943,In_1758);
or U732 (N_732,In_132,In_542);
nor U733 (N_733,In_773,In_1512);
and U734 (N_734,In_255,In_351);
and U735 (N_735,In_1080,In_510);
nand U736 (N_736,In_1093,In_1545);
nor U737 (N_737,In_1451,In_1355);
nor U738 (N_738,In_42,In_278);
nand U739 (N_739,In_1594,In_602);
and U740 (N_740,In_944,In_1668);
or U741 (N_741,In_353,In_1111);
and U742 (N_742,In_512,In_389);
nand U743 (N_743,In_1068,In_1716);
nand U744 (N_744,In_1228,In_1932);
nand U745 (N_745,In_1226,In_465);
or U746 (N_746,In_1842,In_1819);
nand U747 (N_747,In_1351,In_390);
nand U748 (N_748,In_1016,In_105);
nand U749 (N_749,In_335,In_1359);
or U750 (N_750,In_1477,In_779);
and U751 (N_751,In_588,In_688);
or U752 (N_752,In_245,In_1736);
nor U753 (N_753,In_1997,In_395);
nor U754 (N_754,In_1811,In_462);
or U755 (N_755,In_445,In_638);
nand U756 (N_756,In_1114,In_376);
nor U757 (N_757,In_459,In_70);
nand U758 (N_758,In_1473,In_125);
and U759 (N_759,In_183,In_1017);
or U760 (N_760,In_1049,In_1843);
nor U761 (N_761,In_1605,In_1060);
nand U762 (N_762,In_1624,In_953);
nor U763 (N_763,In_1176,In_334);
nand U764 (N_764,In_1442,In_1032);
and U765 (N_765,In_1103,In_1952);
and U766 (N_766,In_1129,In_1035);
or U767 (N_767,In_1948,In_1625);
nand U768 (N_768,In_525,In_754);
nand U769 (N_769,In_1838,In_1830);
nand U770 (N_770,In_243,In_1401);
nand U771 (N_771,In_1944,In_1513);
nand U772 (N_772,In_573,In_271);
and U773 (N_773,In_1737,In_727);
or U774 (N_774,In_1633,In_84);
nor U775 (N_775,In_546,In_83);
and U776 (N_776,In_1342,In_1951);
and U777 (N_777,In_1491,In_613);
and U778 (N_778,In_1391,In_15);
nand U779 (N_779,In_417,In_691);
nand U780 (N_780,In_1610,In_799);
nand U781 (N_781,In_618,In_493);
and U782 (N_782,In_339,In_1719);
nor U783 (N_783,In_331,In_851);
or U784 (N_784,In_1493,In_796);
nor U785 (N_785,In_220,In_1480);
or U786 (N_786,In_1524,In_604);
or U787 (N_787,In_122,In_1380);
or U788 (N_788,In_481,In_138);
and U789 (N_789,In_133,In_1118);
nor U790 (N_790,In_1091,In_1109);
and U791 (N_791,In_1583,In_1552);
nor U792 (N_792,In_36,In_1387);
or U793 (N_793,In_1220,In_1682);
nand U794 (N_794,In_421,In_1108);
or U795 (N_795,In_1410,In_603);
nor U796 (N_796,In_709,In_45);
or U797 (N_797,In_193,In_1546);
nand U798 (N_798,In_1801,In_701);
and U799 (N_799,In_911,In_86);
nor U800 (N_800,In_946,In_1747);
and U801 (N_801,In_10,In_67);
and U802 (N_802,In_1357,In_1383);
nand U803 (N_803,In_43,In_1660);
nor U804 (N_804,In_1836,In_1446);
and U805 (N_805,In_1835,In_1367);
and U806 (N_806,In_320,In_1150);
or U807 (N_807,In_19,In_69);
and U808 (N_808,In_458,In_1455);
and U809 (N_809,In_1413,In_1056);
nor U810 (N_810,In_909,In_314);
nand U811 (N_811,In_1980,In_1439);
nand U812 (N_812,In_1408,In_823);
or U813 (N_813,In_1579,In_1985);
or U814 (N_814,In_1461,In_834);
and U815 (N_815,In_890,In_1412);
or U816 (N_816,In_1967,In_1281);
or U817 (N_817,In_1314,In_1432);
nor U818 (N_818,In_505,In_999);
xor U819 (N_819,In_762,In_1618);
and U820 (N_820,In_694,In_226);
or U821 (N_821,In_927,In_631);
nor U822 (N_822,In_1274,In_203);
nor U823 (N_823,In_1596,In_399);
nand U824 (N_824,In_1088,In_815);
nand U825 (N_825,In_1516,In_1845);
or U826 (N_826,In_1903,In_933);
and U827 (N_827,In_408,In_1234);
nor U828 (N_828,In_90,In_1405);
nand U829 (N_829,In_824,In_1557);
nor U830 (N_830,In_119,In_1688);
nand U831 (N_831,In_103,In_1178);
xor U832 (N_832,In_1665,In_749);
nor U833 (N_833,In_1074,In_868);
and U834 (N_834,In_1465,In_956);
and U835 (N_835,In_321,In_1173);
nand U836 (N_836,In_1902,In_1680);
nand U837 (N_837,In_191,In_888);
nor U838 (N_838,In_1464,In_1725);
or U839 (N_839,In_1246,In_238);
nor U840 (N_840,In_141,In_431);
nor U841 (N_841,In_1288,In_670);
and U842 (N_842,In_1645,In_215);
nand U843 (N_843,In_1335,In_981);
nand U844 (N_844,In_647,In_900);
nand U845 (N_845,In_1784,In_383);
nor U846 (N_846,In_1612,In_1549);
nand U847 (N_847,In_1620,In_1354);
nor U848 (N_848,In_539,In_1452);
or U849 (N_849,In_1673,In_1124);
xnor U850 (N_850,In_768,In_1207);
or U851 (N_851,In_561,In_362);
and U852 (N_852,In_740,In_1729);
and U853 (N_853,In_916,In_1565);
nor U854 (N_854,In_943,In_1787);
nor U855 (N_855,In_785,In_1174);
or U856 (N_856,In_1040,In_26);
and U857 (N_857,In_157,In_1205);
nor U858 (N_858,In_1821,In_1066);
nor U859 (N_859,In_1492,In_842);
and U860 (N_860,In_570,In_767);
or U861 (N_861,In_720,In_400);
or U862 (N_862,In_1015,In_37);
nor U863 (N_863,In_11,In_1269);
and U864 (N_864,In_110,In_112);
or U865 (N_865,In_1404,In_642);
nor U866 (N_866,In_556,In_18);
nand U867 (N_867,In_993,In_77);
or U868 (N_868,In_1248,In_360);
nor U869 (N_869,In_1507,In_461);
or U870 (N_870,In_1323,In_1906);
and U871 (N_871,In_1773,In_1496);
nor U872 (N_872,In_1019,In_1012);
or U873 (N_873,In_1649,In_487);
nand U874 (N_874,In_343,In_508);
nand U875 (N_875,In_1676,In_1890);
and U876 (N_876,In_358,In_1379);
nand U877 (N_877,In_760,In_51);
and U878 (N_878,In_1508,In_1497);
nand U879 (N_879,In_1984,In_484);
nor U880 (N_880,In_516,In_1554);
or U881 (N_881,In_861,In_1070);
and U882 (N_882,In_1116,In_1891);
and U883 (N_883,In_1293,In_1846);
nor U884 (N_884,In_1,In_1882);
or U885 (N_885,In_350,In_742);
nor U886 (N_886,In_511,In_1550);
nand U887 (N_887,In_1591,In_580);
or U888 (N_888,In_1022,In_568);
nand U889 (N_889,In_189,In_1928);
and U890 (N_890,In_1170,In_1495);
or U891 (N_891,In_550,In_274);
xnor U892 (N_892,In_68,In_1977);
nor U893 (N_893,In_1829,In_372);
nand U894 (N_894,In_777,In_1466);
or U895 (N_895,In_820,In_1215);
and U896 (N_896,In_667,In_388);
and U897 (N_897,In_47,In_652);
nand U898 (N_898,In_167,In_1893);
nor U899 (N_899,In_703,In_849);
and U900 (N_900,In_605,In_906);
nor U901 (N_901,In_1456,In_1539);
nand U902 (N_902,In_470,In_381);
and U903 (N_903,In_655,In_297);
or U904 (N_904,In_1424,In_12);
nand U905 (N_905,In_1002,In_1260);
and U906 (N_906,In_1400,In_1957);
and U907 (N_907,In_1917,In_797);
nand U908 (N_908,In_973,In_902);
nand U909 (N_909,In_328,In_1704);
and U910 (N_910,In_932,In_1411);
nor U911 (N_911,In_869,In_1592);
nand U912 (N_912,In_1885,In_89);
nand U913 (N_913,In_1908,In_1601);
or U914 (N_914,In_72,In_396);
nor U915 (N_915,In_860,In_31);
xor U916 (N_916,In_658,In_225);
or U917 (N_917,In_188,In_1319);
nand U918 (N_918,In_963,In_1135);
and U919 (N_919,In_1958,In_1741);
and U920 (N_920,In_877,In_475);
nand U921 (N_921,In_913,In_364);
xnor U922 (N_922,In_415,In_699);
nor U923 (N_923,In_930,In_1986);
nand U924 (N_924,In_325,In_1322);
and U925 (N_925,In_844,In_1257);
or U926 (N_926,In_1669,In_1691);
or U927 (N_927,In_1107,In_1318);
and U928 (N_928,In_1498,In_1664);
and U929 (N_929,In_822,In_1642);
nand U930 (N_930,In_1308,In_1083);
or U931 (N_931,In_833,In_1745);
or U932 (N_932,In_379,In_1598);
nor U933 (N_933,In_772,In_936);
nor U934 (N_934,In_702,In_1423);
and U935 (N_935,In_1291,In_1711);
xor U936 (N_936,In_1222,In_17);
nor U937 (N_937,In_479,In_1522);
or U938 (N_938,In_1796,In_341);
or U939 (N_939,In_1547,In_884);
or U940 (N_940,In_263,In_269);
and U941 (N_941,In_1018,In_1765);
and U942 (N_942,In_637,In_443);
and U943 (N_943,In_250,In_246);
nor U944 (N_944,In_1374,In_804);
nor U945 (N_945,In_437,In_1938);
and U946 (N_946,In_275,In_1324);
and U947 (N_947,In_1978,In_1990);
and U948 (N_948,In_1198,In_1840);
or U949 (N_949,In_1850,In_181);
and U950 (N_950,In_453,In_751);
nand U951 (N_951,In_1571,In_898);
nor U952 (N_952,In_1148,In_436);
nand U953 (N_953,In_1661,In_1613);
and U954 (N_954,In_1714,In_307);
and U955 (N_955,In_1782,In_1155);
and U956 (N_956,In_723,In_789);
and U957 (N_957,In_1671,In_1687);
nand U958 (N_958,In_1181,In_1863);
and U959 (N_959,In_1364,In_1057);
nor U960 (N_960,In_855,In_120);
and U961 (N_961,In_1530,In_1602);
and U962 (N_962,In_1999,In_290);
nand U963 (N_963,In_939,In_531);
or U964 (N_964,In_79,In_1995);
nand U965 (N_965,In_980,In_1754);
or U966 (N_966,In_724,In_208);
and U967 (N_967,In_891,In_1751);
nor U968 (N_968,In_1249,In_901);
nor U969 (N_969,In_599,In_370);
or U970 (N_970,In_821,In_1394);
nand U971 (N_971,In_1059,In_65);
or U972 (N_972,In_917,In_234);
nor U973 (N_973,In_310,In_558);
or U974 (N_974,In_572,In_1392);
and U975 (N_975,In_1036,In_1551);
and U976 (N_976,In_726,In_1793);
nand U977 (N_977,In_856,In_1078);
or U978 (N_978,In_1262,In_518);
or U979 (N_979,In_682,In_159);
and U980 (N_980,In_1927,In_1021);
nand U981 (N_981,In_1445,In_664);
nor U982 (N_982,In_661,In_1039);
and U983 (N_983,In_644,In_575);
nand U984 (N_984,In_413,In_1320);
xor U985 (N_985,In_780,In_1483);
nor U986 (N_986,In_1463,In_482);
nor U987 (N_987,In_1692,In_1102);
and U988 (N_988,In_1197,In_439);
or U989 (N_989,In_1431,In_316);
or U990 (N_990,In_991,In_1515);
or U991 (N_991,In_1009,In_1081);
or U992 (N_992,In_323,In_27);
nor U993 (N_993,In_1593,In_1652);
nand U994 (N_994,In_1479,In_13);
or U995 (N_995,In_1139,In_279);
and U996 (N_996,In_179,In_616);
nand U997 (N_997,In_757,In_287);
or U998 (N_998,In_883,In_1214);
nand U999 (N_999,In_473,In_227);
nor U1000 (N_1000,In_438,In_107);
nand U1001 (N_1001,In_948,In_1141);
and U1002 (N_1002,In_412,In_1161);
and U1003 (N_1003,In_879,In_1336);
or U1004 (N_1004,In_1378,In_494);
or U1005 (N_1005,In_1413,In_1903);
nor U1006 (N_1006,In_1014,In_1329);
nand U1007 (N_1007,In_1294,In_1821);
and U1008 (N_1008,In_580,In_225);
or U1009 (N_1009,In_1626,In_1600);
nand U1010 (N_1010,In_862,In_647);
nand U1011 (N_1011,In_139,In_1334);
and U1012 (N_1012,In_1720,In_987);
or U1013 (N_1013,In_505,In_211);
nand U1014 (N_1014,In_1133,In_1631);
nand U1015 (N_1015,In_1692,In_968);
or U1016 (N_1016,In_803,In_1930);
nor U1017 (N_1017,In_1040,In_1816);
nand U1018 (N_1018,In_383,In_418);
nor U1019 (N_1019,In_1805,In_1001);
nor U1020 (N_1020,In_1913,In_765);
or U1021 (N_1021,In_1870,In_425);
and U1022 (N_1022,In_695,In_552);
nand U1023 (N_1023,In_1277,In_423);
and U1024 (N_1024,In_1854,In_1728);
nand U1025 (N_1025,In_854,In_1701);
nand U1026 (N_1026,In_1594,In_642);
nor U1027 (N_1027,In_1541,In_579);
and U1028 (N_1028,In_1251,In_1218);
or U1029 (N_1029,In_1342,In_1860);
and U1030 (N_1030,In_299,In_1489);
nand U1031 (N_1031,In_1240,In_382);
and U1032 (N_1032,In_1005,In_633);
and U1033 (N_1033,In_819,In_862);
and U1034 (N_1034,In_10,In_1171);
nand U1035 (N_1035,In_492,In_1775);
and U1036 (N_1036,In_834,In_666);
nor U1037 (N_1037,In_1015,In_1064);
nor U1038 (N_1038,In_1920,In_1700);
and U1039 (N_1039,In_410,In_442);
and U1040 (N_1040,In_1821,In_79);
and U1041 (N_1041,In_114,In_835);
nor U1042 (N_1042,In_1406,In_811);
nor U1043 (N_1043,In_993,In_578);
nor U1044 (N_1044,In_570,In_124);
and U1045 (N_1045,In_1504,In_1350);
nor U1046 (N_1046,In_1198,In_331);
or U1047 (N_1047,In_893,In_1008);
nand U1048 (N_1048,In_1656,In_1179);
or U1049 (N_1049,In_1624,In_1465);
and U1050 (N_1050,In_140,In_760);
nand U1051 (N_1051,In_1568,In_231);
or U1052 (N_1052,In_1815,In_733);
or U1053 (N_1053,In_909,In_843);
or U1054 (N_1054,In_16,In_679);
or U1055 (N_1055,In_1798,In_103);
nand U1056 (N_1056,In_159,In_769);
or U1057 (N_1057,In_435,In_1709);
and U1058 (N_1058,In_1061,In_696);
and U1059 (N_1059,In_263,In_1495);
or U1060 (N_1060,In_1968,In_1510);
or U1061 (N_1061,In_1858,In_1442);
and U1062 (N_1062,In_1402,In_1926);
and U1063 (N_1063,In_1362,In_874);
and U1064 (N_1064,In_161,In_1379);
nand U1065 (N_1065,In_1356,In_1390);
or U1066 (N_1066,In_755,In_564);
nor U1067 (N_1067,In_1330,In_1742);
nand U1068 (N_1068,In_1862,In_1886);
or U1069 (N_1069,In_1307,In_1654);
nand U1070 (N_1070,In_625,In_751);
or U1071 (N_1071,In_667,In_1301);
nor U1072 (N_1072,In_817,In_1646);
nand U1073 (N_1073,In_70,In_373);
nand U1074 (N_1074,In_1131,In_776);
nand U1075 (N_1075,In_1963,In_1641);
and U1076 (N_1076,In_936,In_1846);
and U1077 (N_1077,In_678,In_1469);
and U1078 (N_1078,In_370,In_601);
or U1079 (N_1079,In_909,In_1087);
or U1080 (N_1080,In_1998,In_409);
nand U1081 (N_1081,In_1249,In_1160);
nor U1082 (N_1082,In_1050,In_1707);
or U1083 (N_1083,In_1356,In_1292);
nor U1084 (N_1084,In_460,In_1221);
nand U1085 (N_1085,In_652,In_1943);
nor U1086 (N_1086,In_222,In_817);
nand U1087 (N_1087,In_344,In_1236);
or U1088 (N_1088,In_1353,In_67);
nor U1089 (N_1089,In_905,In_310);
nor U1090 (N_1090,In_58,In_1222);
nand U1091 (N_1091,In_246,In_1246);
nor U1092 (N_1092,In_1689,In_726);
nor U1093 (N_1093,In_1942,In_1832);
nand U1094 (N_1094,In_700,In_975);
nor U1095 (N_1095,In_469,In_202);
and U1096 (N_1096,In_1223,In_801);
nor U1097 (N_1097,In_67,In_1968);
and U1098 (N_1098,In_729,In_1530);
nand U1099 (N_1099,In_857,In_442);
nor U1100 (N_1100,In_1007,In_164);
or U1101 (N_1101,In_1452,In_65);
nand U1102 (N_1102,In_7,In_11);
nor U1103 (N_1103,In_1234,In_97);
nor U1104 (N_1104,In_480,In_849);
nor U1105 (N_1105,In_46,In_1305);
and U1106 (N_1106,In_1900,In_1749);
nand U1107 (N_1107,In_1464,In_1610);
nor U1108 (N_1108,In_538,In_1811);
nor U1109 (N_1109,In_791,In_1887);
and U1110 (N_1110,In_1942,In_1687);
nand U1111 (N_1111,In_1839,In_414);
nor U1112 (N_1112,In_4,In_1534);
or U1113 (N_1113,In_1634,In_1674);
nand U1114 (N_1114,In_672,In_674);
nor U1115 (N_1115,In_391,In_200);
nor U1116 (N_1116,In_732,In_765);
nand U1117 (N_1117,In_937,In_1129);
or U1118 (N_1118,In_1956,In_193);
nand U1119 (N_1119,In_709,In_397);
nand U1120 (N_1120,In_376,In_513);
and U1121 (N_1121,In_26,In_454);
nand U1122 (N_1122,In_1336,In_1159);
and U1123 (N_1123,In_989,In_1476);
nor U1124 (N_1124,In_169,In_1355);
nor U1125 (N_1125,In_1348,In_1143);
nand U1126 (N_1126,In_1760,In_768);
and U1127 (N_1127,In_1656,In_391);
and U1128 (N_1128,In_1178,In_546);
and U1129 (N_1129,In_122,In_1479);
nand U1130 (N_1130,In_993,In_1147);
or U1131 (N_1131,In_723,In_685);
nand U1132 (N_1132,In_1536,In_1107);
nand U1133 (N_1133,In_756,In_1718);
and U1134 (N_1134,In_267,In_730);
nor U1135 (N_1135,In_729,In_193);
and U1136 (N_1136,In_697,In_871);
nand U1137 (N_1137,In_596,In_1603);
or U1138 (N_1138,In_1896,In_678);
nor U1139 (N_1139,In_854,In_242);
nor U1140 (N_1140,In_1592,In_503);
or U1141 (N_1141,In_1230,In_1456);
or U1142 (N_1142,In_1923,In_1261);
or U1143 (N_1143,In_542,In_730);
and U1144 (N_1144,In_821,In_1204);
nor U1145 (N_1145,In_956,In_1567);
or U1146 (N_1146,In_1749,In_1129);
and U1147 (N_1147,In_1349,In_1533);
and U1148 (N_1148,In_1968,In_1233);
or U1149 (N_1149,In_23,In_219);
nand U1150 (N_1150,In_1231,In_323);
and U1151 (N_1151,In_225,In_642);
nand U1152 (N_1152,In_1250,In_570);
nor U1153 (N_1153,In_1764,In_918);
nand U1154 (N_1154,In_351,In_911);
nand U1155 (N_1155,In_277,In_1423);
nand U1156 (N_1156,In_1279,In_1782);
or U1157 (N_1157,In_334,In_945);
or U1158 (N_1158,In_1999,In_1756);
nor U1159 (N_1159,In_1332,In_464);
and U1160 (N_1160,In_286,In_927);
or U1161 (N_1161,In_173,In_1315);
and U1162 (N_1162,In_1577,In_821);
and U1163 (N_1163,In_36,In_436);
or U1164 (N_1164,In_408,In_1462);
nor U1165 (N_1165,In_748,In_509);
nor U1166 (N_1166,In_110,In_35);
nand U1167 (N_1167,In_1063,In_1627);
or U1168 (N_1168,In_296,In_438);
or U1169 (N_1169,In_701,In_1762);
and U1170 (N_1170,In_1505,In_767);
nand U1171 (N_1171,In_371,In_1965);
nand U1172 (N_1172,In_1294,In_1566);
nand U1173 (N_1173,In_386,In_701);
and U1174 (N_1174,In_66,In_1291);
or U1175 (N_1175,In_1186,In_719);
and U1176 (N_1176,In_736,In_1074);
and U1177 (N_1177,In_1423,In_1863);
nor U1178 (N_1178,In_128,In_1190);
or U1179 (N_1179,In_1083,In_1284);
or U1180 (N_1180,In_1092,In_734);
nand U1181 (N_1181,In_1694,In_1268);
nor U1182 (N_1182,In_875,In_587);
xnor U1183 (N_1183,In_359,In_23);
or U1184 (N_1184,In_430,In_340);
and U1185 (N_1185,In_1877,In_1103);
or U1186 (N_1186,In_1202,In_15);
or U1187 (N_1187,In_447,In_1477);
or U1188 (N_1188,In_1769,In_620);
nand U1189 (N_1189,In_1739,In_1687);
nand U1190 (N_1190,In_1003,In_1497);
nand U1191 (N_1191,In_878,In_379);
nor U1192 (N_1192,In_518,In_988);
or U1193 (N_1193,In_416,In_644);
nor U1194 (N_1194,In_1439,In_1107);
nor U1195 (N_1195,In_571,In_948);
nand U1196 (N_1196,In_781,In_1289);
or U1197 (N_1197,In_1573,In_1458);
nand U1198 (N_1198,In_1254,In_700);
nand U1199 (N_1199,In_29,In_1799);
nor U1200 (N_1200,In_310,In_1628);
or U1201 (N_1201,In_652,In_343);
or U1202 (N_1202,In_1572,In_1839);
nor U1203 (N_1203,In_1185,In_220);
nor U1204 (N_1204,In_1513,In_1262);
nor U1205 (N_1205,In_30,In_1988);
nor U1206 (N_1206,In_1855,In_1947);
nand U1207 (N_1207,In_774,In_1775);
nand U1208 (N_1208,In_261,In_1523);
nand U1209 (N_1209,In_561,In_1650);
and U1210 (N_1210,In_1841,In_925);
or U1211 (N_1211,In_785,In_144);
or U1212 (N_1212,In_787,In_1780);
nor U1213 (N_1213,In_1790,In_618);
or U1214 (N_1214,In_1905,In_1962);
nor U1215 (N_1215,In_707,In_230);
nand U1216 (N_1216,In_1788,In_1871);
or U1217 (N_1217,In_472,In_286);
nand U1218 (N_1218,In_487,In_1272);
and U1219 (N_1219,In_836,In_1956);
nor U1220 (N_1220,In_325,In_794);
nor U1221 (N_1221,In_813,In_1348);
or U1222 (N_1222,In_988,In_248);
and U1223 (N_1223,In_1818,In_143);
or U1224 (N_1224,In_916,In_505);
or U1225 (N_1225,In_827,In_1429);
or U1226 (N_1226,In_107,In_1165);
nand U1227 (N_1227,In_1049,In_1348);
or U1228 (N_1228,In_1820,In_897);
nor U1229 (N_1229,In_760,In_1694);
nand U1230 (N_1230,In_1850,In_545);
or U1231 (N_1231,In_1042,In_1014);
or U1232 (N_1232,In_206,In_562);
nor U1233 (N_1233,In_735,In_1717);
or U1234 (N_1234,In_342,In_1058);
and U1235 (N_1235,In_1755,In_1794);
and U1236 (N_1236,In_222,In_1442);
or U1237 (N_1237,In_297,In_860);
nand U1238 (N_1238,In_1083,In_534);
nand U1239 (N_1239,In_1071,In_1452);
nand U1240 (N_1240,In_277,In_565);
nand U1241 (N_1241,In_1683,In_1524);
nand U1242 (N_1242,In_485,In_1819);
or U1243 (N_1243,In_469,In_42);
nand U1244 (N_1244,In_691,In_955);
or U1245 (N_1245,In_387,In_32);
nand U1246 (N_1246,In_1545,In_1513);
or U1247 (N_1247,In_946,In_830);
or U1248 (N_1248,In_204,In_646);
nand U1249 (N_1249,In_1528,In_3);
and U1250 (N_1250,In_958,In_1466);
and U1251 (N_1251,In_1918,In_468);
nand U1252 (N_1252,In_969,In_1418);
and U1253 (N_1253,In_61,In_47);
or U1254 (N_1254,In_172,In_1152);
nor U1255 (N_1255,In_1196,In_940);
nand U1256 (N_1256,In_718,In_194);
nand U1257 (N_1257,In_31,In_1763);
or U1258 (N_1258,In_452,In_1232);
nand U1259 (N_1259,In_906,In_873);
nor U1260 (N_1260,In_191,In_1822);
nand U1261 (N_1261,In_1580,In_263);
or U1262 (N_1262,In_461,In_1954);
and U1263 (N_1263,In_927,In_690);
and U1264 (N_1264,In_129,In_41);
or U1265 (N_1265,In_1274,In_1613);
nand U1266 (N_1266,In_278,In_1134);
or U1267 (N_1267,In_1360,In_1991);
nand U1268 (N_1268,In_687,In_59);
and U1269 (N_1269,In_1327,In_1901);
or U1270 (N_1270,In_1594,In_3);
nand U1271 (N_1271,In_502,In_568);
nand U1272 (N_1272,In_245,In_341);
nand U1273 (N_1273,In_928,In_54);
or U1274 (N_1274,In_565,In_1563);
or U1275 (N_1275,In_276,In_165);
nor U1276 (N_1276,In_1901,In_549);
nor U1277 (N_1277,In_1429,In_215);
or U1278 (N_1278,In_1583,In_1058);
and U1279 (N_1279,In_1646,In_794);
nand U1280 (N_1280,In_239,In_900);
nand U1281 (N_1281,In_1101,In_398);
and U1282 (N_1282,In_1073,In_400);
nand U1283 (N_1283,In_607,In_636);
and U1284 (N_1284,In_193,In_512);
or U1285 (N_1285,In_1607,In_1463);
or U1286 (N_1286,In_772,In_1077);
and U1287 (N_1287,In_1663,In_323);
and U1288 (N_1288,In_1943,In_531);
nor U1289 (N_1289,In_469,In_398);
nor U1290 (N_1290,In_1975,In_86);
nand U1291 (N_1291,In_1852,In_954);
or U1292 (N_1292,In_988,In_343);
nor U1293 (N_1293,In_1624,In_324);
or U1294 (N_1294,In_1357,In_1012);
nand U1295 (N_1295,In_453,In_1247);
nor U1296 (N_1296,In_1061,In_34);
nor U1297 (N_1297,In_942,In_711);
nand U1298 (N_1298,In_233,In_1271);
nand U1299 (N_1299,In_1335,In_253);
or U1300 (N_1300,In_1561,In_696);
or U1301 (N_1301,In_615,In_131);
xnor U1302 (N_1302,In_1955,In_1586);
and U1303 (N_1303,In_474,In_1244);
or U1304 (N_1304,In_1192,In_228);
nand U1305 (N_1305,In_1761,In_441);
and U1306 (N_1306,In_1029,In_357);
and U1307 (N_1307,In_133,In_1330);
or U1308 (N_1308,In_1914,In_493);
nand U1309 (N_1309,In_263,In_1793);
or U1310 (N_1310,In_166,In_1372);
or U1311 (N_1311,In_253,In_220);
nand U1312 (N_1312,In_219,In_186);
or U1313 (N_1313,In_681,In_781);
and U1314 (N_1314,In_983,In_978);
or U1315 (N_1315,In_538,In_1678);
nor U1316 (N_1316,In_1402,In_655);
and U1317 (N_1317,In_1188,In_290);
nand U1318 (N_1318,In_459,In_189);
nand U1319 (N_1319,In_1197,In_1554);
and U1320 (N_1320,In_1738,In_648);
and U1321 (N_1321,In_1433,In_1749);
nor U1322 (N_1322,In_1762,In_1604);
nor U1323 (N_1323,In_506,In_358);
nor U1324 (N_1324,In_109,In_1310);
nor U1325 (N_1325,In_1437,In_1624);
nand U1326 (N_1326,In_679,In_1278);
nor U1327 (N_1327,In_1608,In_166);
and U1328 (N_1328,In_1016,In_1292);
nor U1329 (N_1329,In_1345,In_1820);
and U1330 (N_1330,In_79,In_601);
or U1331 (N_1331,In_1141,In_566);
nor U1332 (N_1332,In_925,In_1914);
and U1333 (N_1333,In_1927,In_1245);
nand U1334 (N_1334,In_1151,In_599);
or U1335 (N_1335,In_1498,In_1367);
nand U1336 (N_1336,In_497,In_1588);
and U1337 (N_1337,In_1523,In_228);
nand U1338 (N_1338,In_1771,In_1331);
xor U1339 (N_1339,In_434,In_617);
nor U1340 (N_1340,In_885,In_1682);
nand U1341 (N_1341,In_511,In_715);
and U1342 (N_1342,In_1690,In_698);
nand U1343 (N_1343,In_1496,In_350);
nand U1344 (N_1344,In_1614,In_1684);
or U1345 (N_1345,In_164,In_1711);
and U1346 (N_1346,In_495,In_309);
nor U1347 (N_1347,In_940,In_1603);
and U1348 (N_1348,In_1675,In_1551);
nor U1349 (N_1349,In_166,In_1132);
nand U1350 (N_1350,In_226,In_1250);
nor U1351 (N_1351,In_34,In_1381);
and U1352 (N_1352,In_1767,In_56);
or U1353 (N_1353,In_1568,In_438);
nand U1354 (N_1354,In_517,In_1070);
and U1355 (N_1355,In_1802,In_393);
nor U1356 (N_1356,In_1194,In_1917);
nand U1357 (N_1357,In_1827,In_216);
and U1358 (N_1358,In_1291,In_1106);
nor U1359 (N_1359,In_164,In_448);
nor U1360 (N_1360,In_582,In_1401);
nand U1361 (N_1361,In_769,In_1191);
nand U1362 (N_1362,In_800,In_286);
nand U1363 (N_1363,In_442,In_1126);
nor U1364 (N_1364,In_969,In_1858);
or U1365 (N_1365,In_85,In_550);
and U1366 (N_1366,In_1368,In_1602);
and U1367 (N_1367,In_1427,In_166);
and U1368 (N_1368,In_1206,In_1707);
and U1369 (N_1369,In_140,In_111);
nor U1370 (N_1370,In_903,In_362);
and U1371 (N_1371,In_341,In_501);
and U1372 (N_1372,In_1634,In_777);
nor U1373 (N_1373,In_919,In_1194);
and U1374 (N_1374,In_290,In_1274);
nor U1375 (N_1375,In_826,In_517);
and U1376 (N_1376,In_42,In_1754);
nand U1377 (N_1377,In_722,In_190);
nand U1378 (N_1378,In_990,In_1867);
nor U1379 (N_1379,In_1584,In_1650);
nor U1380 (N_1380,In_1216,In_507);
or U1381 (N_1381,In_1757,In_1618);
nand U1382 (N_1382,In_768,In_762);
and U1383 (N_1383,In_45,In_275);
or U1384 (N_1384,In_532,In_1314);
nor U1385 (N_1385,In_820,In_1782);
nor U1386 (N_1386,In_579,In_29);
nand U1387 (N_1387,In_329,In_1992);
or U1388 (N_1388,In_918,In_1453);
nand U1389 (N_1389,In_1343,In_1509);
nand U1390 (N_1390,In_418,In_685);
nor U1391 (N_1391,In_1808,In_484);
or U1392 (N_1392,In_46,In_572);
nand U1393 (N_1393,In_771,In_1700);
nor U1394 (N_1394,In_1061,In_1377);
and U1395 (N_1395,In_253,In_1756);
or U1396 (N_1396,In_1698,In_1982);
nor U1397 (N_1397,In_603,In_354);
nor U1398 (N_1398,In_1751,In_462);
and U1399 (N_1399,In_1816,In_830);
and U1400 (N_1400,In_1704,In_1609);
nand U1401 (N_1401,In_1783,In_1118);
nand U1402 (N_1402,In_1524,In_1243);
nand U1403 (N_1403,In_705,In_16);
and U1404 (N_1404,In_659,In_327);
nor U1405 (N_1405,In_88,In_200);
nand U1406 (N_1406,In_640,In_477);
nand U1407 (N_1407,In_1792,In_1091);
or U1408 (N_1408,In_405,In_1437);
and U1409 (N_1409,In_376,In_1623);
nand U1410 (N_1410,In_1202,In_254);
and U1411 (N_1411,In_1844,In_1543);
nand U1412 (N_1412,In_1399,In_236);
and U1413 (N_1413,In_462,In_1285);
nor U1414 (N_1414,In_712,In_1737);
or U1415 (N_1415,In_1181,In_1807);
xor U1416 (N_1416,In_968,In_450);
nor U1417 (N_1417,In_799,In_798);
and U1418 (N_1418,In_1283,In_153);
or U1419 (N_1419,In_621,In_1409);
and U1420 (N_1420,In_1077,In_1502);
or U1421 (N_1421,In_78,In_612);
and U1422 (N_1422,In_1556,In_1950);
or U1423 (N_1423,In_1344,In_1203);
nor U1424 (N_1424,In_1123,In_1519);
or U1425 (N_1425,In_1719,In_1482);
or U1426 (N_1426,In_806,In_1146);
nor U1427 (N_1427,In_921,In_1031);
nor U1428 (N_1428,In_874,In_1916);
nand U1429 (N_1429,In_1430,In_698);
or U1430 (N_1430,In_920,In_1665);
or U1431 (N_1431,In_507,In_486);
and U1432 (N_1432,In_1742,In_182);
nor U1433 (N_1433,In_1527,In_820);
nor U1434 (N_1434,In_517,In_111);
nor U1435 (N_1435,In_712,In_536);
nand U1436 (N_1436,In_1251,In_1285);
and U1437 (N_1437,In_309,In_1684);
nor U1438 (N_1438,In_1715,In_1234);
nand U1439 (N_1439,In_952,In_740);
or U1440 (N_1440,In_511,In_810);
nor U1441 (N_1441,In_1765,In_874);
nor U1442 (N_1442,In_999,In_1963);
nand U1443 (N_1443,In_617,In_1938);
and U1444 (N_1444,In_1994,In_488);
or U1445 (N_1445,In_1783,In_329);
or U1446 (N_1446,In_1398,In_842);
and U1447 (N_1447,In_1626,In_1316);
or U1448 (N_1448,In_1461,In_734);
or U1449 (N_1449,In_923,In_266);
nand U1450 (N_1450,In_1568,In_715);
or U1451 (N_1451,In_1676,In_1496);
nand U1452 (N_1452,In_765,In_360);
and U1453 (N_1453,In_1069,In_1091);
nor U1454 (N_1454,In_1819,In_1082);
nand U1455 (N_1455,In_195,In_931);
nor U1456 (N_1456,In_1685,In_1344);
or U1457 (N_1457,In_1239,In_1279);
nand U1458 (N_1458,In_1057,In_424);
nand U1459 (N_1459,In_453,In_942);
nand U1460 (N_1460,In_727,In_1721);
nand U1461 (N_1461,In_413,In_1116);
and U1462 (N_1462,In_1033,In_387);
nor U1463 (N_1463,In_1315,In_1796);
or U1464 (N_1464,In_637,In_1506);
nor U1465 (N_1465,In_313,In_1360);
nand U1466 (N_1466,In_158,In_1993);
xnor U1467 (N_1467,In_1990,In_1437);
and U1468 (N_1468,In_675,In_912);
nand U1469 (N_1469,In_480,In_608);
or U1470 (N_1470,In_1067,In_96);
or U1471 (N_1471,In_879,In_705);
nor U1472 (N_1472,In_1492,In_1611);
nor U1473 (N_1473,In_826,In_1918);
nor U1474 (N_1474,In_1121,In_1957);
nand U1475 (N_1475,In_1941,In_409);
nand U1476 (N_1476,In_268,In_635);
and U1477 (N_1477,In_631,In_1046);
nor U1478 (N_1478,In_1700,In_1896);
and U1479 (N_1479,In_753,In_1914);
nand U1480 (N_1480,In_1517,In_1656);
nand U1481 (N_1481,In_62,In_1954);
or U1482 (N_1482,In_302,In_1080);
nand U1483 (N_1483,In_977,In_1226);
nand U1484 (N_1484,In_1442,In_1265);
or U1485 (N_1485,In_800,In_1586);
nor U1486 (N_1486,In_479,In_181);
xnor U1487 (N_1487,In_323,In_1545);
or U1488 (N_1488,In_790,In_1579);
nor U1489 (N_1489,In_1004,In_1503);
nand U1490 (N_1490,In_1231,In_403);
nand U1491 (N_1491,In_1576,In_1631);
nor U1492 (N_1492,In_692,In_1965);
nor U1493 (N_1493,In_469,In_319);
nand U1494 (N_1494,In_843,In_515);
nor U1495 (N_1495,In_1020,In_435);
nand U1496 (N_1496,In_123,In_1058);
or U1497 (N_1497,In_1006,In_712);
nand U1498 (N_1498,In_850,In_800);
nand U1499 (N_1499,In_841,In_1999);
nand U1500 (N_1500,In_1366,In_1337);
xor U1501 (N_1501,In_963,In_118);
nor U1502 (N_1502,In_1488,In_1200);
or U1503 (N_1503,In_1829,In_835);
nor U1504 (N_1504,In_1222,In_1051);
nand U1505 (N_1505,In_1406,In_1996);
or U1506 (N_1506,In_1312,In_160);
and U1507 (N_1507,In_720,In_1416);
nor U1508 (N_1508,In_1249,In_861);
nor U1509 (N_1509,In_1143,In_1798);
or U1510 (N_1510,In_1830,In_789);
or U1511 (N_1511,In_1105,In_44);
and U1512 (N_1512,In_75,In_937);
and U1513 (N_1513,In_924,In_699);
nor U1514 (N_1514,In_1885,In_985);
nor U1515 (N_1515,In_848,In_604);
or U1516 (N_1516,In_820,In_1211);
or U1517 (N_1517,In_1826,In_1550);
nand U1518 (N_1518,In_899,In_62);
nor U1519 (N_1519,In_1755,In_1778);
or U1520 (N_1520,In_1203,In_567);
and U1521 (N_1521,In_1062,In_956);
nor U1522 (N_1522,In_1834,In_1736);
and U1523 (N_1523,In_1617,In_1750);
or U1524 (N_1524,In_840,In_1737);
and U1525 (N_1525,In_1206,In_1309);
and U1526 (N_1526,In_497,In_174);
and U1527 (N_1527,In_1071,In_1001);
or U1528 (N_1528,In_138,In_273);
and U1529 (N_1529,In_1553,In_418);
nor U1530 (N_1530,In_398,In_486);
xnor U1531 (N_1531,In_1005,In_992);
nor U1532 (N_1532,In_539,In_81);
nand U1533 (N_1533,In_882,In_65);
or U1534 (N_1534,In_1022,In_1838);
or U1535 (N_1535,In_590,In_534);
nand U1536 (N_1536,In_1950,In_1513);
nand U1537 (N_1537,In_843,In_1584);
or U1538 (N_1538,In_930,In_309);
or U1539 (N_1539,In_277,In_825);
nor U1540 (N_1540,In_658,In_267);
nand U1541 (N_1541,In_1447,In_1152);
or U1542 (N_1542,In_1437,In_1486);
nor U1543 (N_1543,In_1469,In_1417);
nand U1544 (N_1544,In_906,In_519);
nand U1545 (N_1545,In_1885,In_1280);
nor U1546 (N_1546,In_1600,In_1614);
and U1547 (N_1547,In_565,In_544);
or U1548 (N_1548,In_854,In_58);
and U1549 (N_1549,In_590,In_41);
or U1550 (N_1550,In_944,In_838);
nor U1551 (N_1551,In_1734,In_455);
and U1552 (N_1552,In_438,In_1343);
nand U1553 (N_1553,In_1285,In_1700);
nand U1554 (N_1554,In_1217,In_1328);
nor U1555 (N_1555,In_54,In_721);
nor U1556 (N_1556,In_1621,In_905);
nand U1557 (N_1557,In_1149,In_1015);
nor U1558 (N_1558,In_789,In_1057);
or U1559 (N_1559,In_1352,In_1780);
and U1560 (N_1560,In_1247,In_1318);
or U1561 (N_1561,In_1271,In_1236);
nor U1562 (N_1562,In_1240,In_1705);
and U1563 (N_1563,In_464,In_366);
and U1564 (N_1564,In_1892,In_1510);
and U1565 (N_1565,In_1220,In_846);
nor U1566 (N_1566,In_199,In_1381);
or U1567 (N_1567,In_426,In_1370);
and U1568 (N_1568,In_99,In_144);
nor U1569 (N_1569,In_1984,In_1411);
or U1570 (N_1570,In_171,In_34);
or U1571 (N_1571,In_1507,In_941);
or U1572 (N_1572,In_769,In_1895);
nand U1573 (N_1573,In_652,In_1248);
nor U1574 (N_1574,In_252,In_944);
nor U1575 (N_1575,In_5,In_1259);
nor U1576 (N_1576,In_709,In_510);
or U1577 (N_1577,In_305,In_1290);
and U1578 (N_1578,In_1202,In_843);
and U1579 (N_1579,In_482,In_1474);
nand U1580 (N_1580,In_1021,In_1002);
nand U1581 (N_1581,In_1543,In_37);
nor U1582 (N_1582,In_181,In_539);
and U1583 (N_1583,In_265,In_1659);
and U1584 (N_1584,In_1426,In_284);
nand U1585 (N_1585,In_681,In_340);
or U1586 (N_1586,In_391,In_1901);
nand U1587 (N_1587,In_1333,In_341);
or U1588 (N_1588,In_1709,In_974);
and U1589 (N_1589,In_1626,In_1842);
nor U1590 (N_1590,In_1055,In_245);
or U1591 (N_1591,In_25,In_806);
nand U1592 (N_1592,In_21,In_1089);
nor U1593 (N_1593,In_607,In_1071);
or U1594 (N_1594,In_1507,In_125);
nand U1595 (N_1595,In_1383,In_707);
and U1596 (N_1596,In_1027,In_838);
nand U1597 (N_1597,In_113,In_344);
nand U1598 (N_1598,In_257,In_1648);
and U1599 (N_1599,In_1596,In_887);
nand U1600 (N_1600,In_958,In_142);
or U1601 (N_1601,In_1116,In_1334);
nand U1602 (N_1602,In_766,In_1788);
or U1603 (N_1603,In_396,In_1901);
and U1604 (N_1604,In_1640,In_1193);
nand U1605 (N_1605,In_131,In_1145);
nor U1606 (N_1606,In_789,In_1381);
nand U1607 (N_1607,In_546,In_599);
nand U1608 (N_1608,In_1461,In_904);
or U1609 (N_1609,In_459,In_1681);
and U1610 (N_1610,In_1966,In_743);
or U1611 (N_1611,In_1394,In_1006);
nand U1612 (N_1612,In_1690,In_1953);
nor U1613 (N_1613,In_528,In_1468);
and U1614 (N_1614,In_644,In_1221);
nand U1615 (N_1615,In_1090,In_809);
and U1616 (N_1616,In_173,In_352);
and U1617 (N_1617,In_475,In_927);
xnor U1618 (N_1618,In_598,In_852);
or U1619 (N_1619,In_148,In_1239);
nand U1620 (N_1620,In_178,In_1109);
nand U1621 (N_1621,In_1625,In_735);
nor U1622 (N_1622,In_935,In_1430);
nand U1623 (N_1623,In_1358,In_1250);
nand U1624 (N_1624,In_1415,In_380);
xnor U1625 (N_1625,In_967,In_1023);
or U1626 (N_1626,In_96,In_1086);
or U1627 (N_1627,In_1505,In_1577);
nor U1628 (N_1628,In_1303,In_1770);
or U1629 (N_1629,In_716,In_1252);
nand U1630 (N_1630,In_623,In_302);
nor U1631 (N_1631,In_492,In_906);
nor U1632 (N_1632,In_326,In_1332);
or U1633 (N_1633,In_822,In_669);
nor U1634 (N_1634,In_953,In_750);
nand U1635 (N_1635,In_656,In_916);
nand U1636 (N_1636,In_591,In_1567);
or U1637 (N_1637,In_1533,In_1311);
or U1638 (N_1638,In_1658,In_1146);
nand U1639 (N_1639,In_1293,In_1633);
nand U1640 (N_1640,In_1165,In_511);
and U1641 (N_1641,In_1514,In_1062);
nand U1642 (N_1642,In_1661,In_1596);
nor U1643 (N_1643,In_493,In_589);
or U1644 (N_1644,In_302,In_710);
nand U1645 (N_1645,In_1231,In_1148);
nand U1646 (N_1646,In_1586,In_1696);
and U1647 (N_1647,In_118,In_951);
or U1648 (N_1648,In_1430,In_1462);
and U1649 (N_1649,In_1106,In_591);
and U1650 (N_1650,In_1091,In_1898);
and U1651 (N_1651,In_1135,In_413);
nor U1652 (N_1652,In_802,In_396);
nand U1653 (N_1653,In_558,In_1416);
nand U1654 (N_1654,In_19,In_921);
nor U1655 (N_1655,In_815,In_1459);
nor U1656 (N_1656,In_1257,In_1613);
and U1657 (N_1657,In_1849,In_1457);
or U1658 (N_1658,In_629,In_1125);
or U1659 (N_1659,In_230,In_1622);
nand U1660 (N_1660,In_254,In_850);
nor U1661 (N_1661,In_299,In_1831);
xnor U1662 (N_1662,In_755,In_1832);
nor U1663 (N_1663,In_1439,In_2);
nand U1664 (N_1664,In_142,In_624);
and U1665 (N_1665,In_944,In_672);
nand U1666 (N_1666,In_841,In_1977);
or U1667 (N_1667,In_889,In_346);
or U1668 (N_1668,In_1818,In_571);
xnor U1669 (N_1669,In_468,In_782);
and U1670 (N_1670,In_396,In_1250);
and U1671 (N_1671,In_1778,In_1912);
nor U1672 (N_1672,In_1066,In_1664);
or U1673 (N_1673,In_966,In_1966);
or U1674 (N_1674,In_527,In_16);
nand U1675 (N_1675,In_1831,In_600);
or U1676 (N_1676,In_1569,In_1476);
nand U1677 (N_1677,In_304,In_1482);
nand U1678 (N_1678,In_538,In_596);
and U1679 (N_1679,In_797,In_321);
nor U1680 (N_1680,In_1645,In_413);
and U1681 (N_1681,In_1445,In_571);
or U1682 (N_1682,In_291,In_846);
nand U1683 (N_1683,In_1820,In_1754);
nor U1684 (N_1684,In_922,In_1238);
and U1685 (N_1685,In_1480,In_1386);
nand U1686 (N_1686,In_1456,In_1764);
nor U1687 (N_1687,In_1336,In_111);
nor U1688 (N_1688,In_1258,In_869);
or U1689 (N_1689,In_195,In_1174);
or U1690 (N_1690,In_149,In_1843);
nand U1691 (N_1691,In_1756,In_1981);
or U1692 (N_1692,In_573,In_521);
xor U1693 (N_1693,In_1950,In_1223);
and U1694 (N_1694,In_890,In_1881);
and U1695 (N_1695,In_172,In_1642);
nand U1696 (N_1696,In_947,In_1895);
or U1697 (N_1697,In_395,In_1244);
or U1698 (N_1698,In_398,In_1431);
or U1699 (N_1699,In_1920,In_1582);
and U1700 (N_1700,In_1260,In_572);
nor U1701 (N_1701,In_224,In_1440);
nand U1702 (N_1702,In_797,In_502);
nor U1703 (N_1703,In_961,In_1909);
nand U1704 (N_1704,In_772,In_604);
and U1705 (N_1705,In_59,In_1827);
nand U1706 (N_1706,In_1213,In_451);
or U1707 (N_1707,In_1799,In_426);
nand U1708 (N_1708,In_1499,In_265);
nand U1709 (N_1709,In_127,In_1327);
nor U1710 (N_1710,In_375,In_1825);
nand U1711 (N_1711,In_1893,In_865);
and U1712 (N_1712,In_1502,In_724);
nor U1713 (N_1713,In_1411,In_1661);
nand U1714 (N_1714,In_1279,In_1342);
nand U1715 (N_1715,In_441,In_1638);
and U1716 (N_1716,In_1229,In_53);
or U1717 (N_1717,In_950,In_1290);
or U1718 (N_1718,In_886,In_1443);
nor U1719 (N_1719,In_948,In_177);
nand U1720 (N_1720,In_326,In_1441);
or U1721 (N_1721,In_1383,In_1791);
and U1722 (N_1722,In_1220,In_1931);
nand U1723 (N_1723,In_1487,In_1205);
nand U1724 (N_1724,In_118,In_1708);
or U1725 (N_1725,In_257,In_98);
nand U1726 (N_1726,In_1806,In_1044);
nor U1727 (N_1727,In_1686,In_1851);
nand U1728 (N_1728,In_1595,In_440);
and U1729 (N_1729,In_1039,In_1308);
and U1730 (N_1730,In_172,In_132);
and U1731 (N_1731,In_962,In_516);
nor U1732 (N_1732,In_461,In_1244);
nand U1733 (N_1733,In_1841,In_529);
and U1734 (N_1734,In_740,In_149);
or U1735 (N_1735,In_149,In_123);
or U1736 (N_1736,In_743,In_1651);
and U1737 (N_1737,In_865,In_805);
xnor U1738 (N_1738,In_1851,In_142);
nor U1739 (N_1739,In_616,In_1902);
and U1740 (N_1740,In_264,In_893);
and U1741 (N_1741,In_547,In_1520);
or U1742 (N_1742,In_720,In_1840);
nand U1743 (N_1743,In_1733,In_912);
nor U1744 (N_1744,In_1626,In_111);
and U1745 (N_1745,In_917,In_597);
nor U1746 (N_1746,In_613,In_1459);
and U1747 (N_1747,In_1557,In_1860);
nand U1748 (N_1748,In_950,In_1544);
or U1749 (N_1749,In_1645,In_1683);
nor U1750 (N_1750,In_317,In_742);
nand U1751 (N_1751,In_705,In_144);
and U1752 (N_1752,In_1366,In_1681);
or U1753 (N_1753,In_1908,In_543);
nor U1754 (N_1754,In_774,In_1179);
nor U1755 (N_1755,In_875,In_414);
or U1756 (N_1756,In_1478,In_607);
nor U1757 (N_1757,In_1030,In_166);
and U1758 (N_1758,In_508,In_783);
and U1759 (N_1759,In_929,In_1826);
nor U1760 (N_1760,In_1030,In_1281);
nor U1761 (N_1761,In_1564,In_1521);
nor U1762 (N_1762,In_1800,In_1496);
xor U1763 (N_1763,In_1369,In_1567);
nor U1764 (N_1764,In_617,In_368);
xor U1765 (N_1765,In_1310,In_1120);
nand U1766 (N_1766,In_649,In_265);
and U1767 (N_1767,In_186,In_1053);
nand U1768 (N_1768,In_1877,In_191);
nand U1769 (N_1769,In_1542,In_1851);
and U1770 (N_1770,In_1443,In_93);
or U1771 (N_1771,In_605,In_466);
or U1772 (N_1772,In_1046,In_1496);
nor U1773 (N_1773,In_212,In_327);
or U1774 (N_1774,In_253,In_1484);
or U1775 (N_1775,In_1240,In_3);
and U1776 (N_1776,In_908,In_515);
nand U1777 (N_1777,In_1301,In_716);
nor U1778 (N_1778,In_771,In_1776);
nor U1779 (N_1779,In_1026,In_1824);
nor U1780 (N_1780,In_469,In_468);
or U1781 (N_1781,In_1014,In_837);
nor U1782 (N_1782,In_1011,In_1973);
nand U1783 (N_1783,In_1942,In_1871);
nor U1784 (N_1784,In_1120,In_926);
nor U1785 (N_1785,In_1033,In_872);
and U1786 (N_1786,In_893,In_1950);
or U1787 (N_1787,In_1761,In_237);
nor U1788 (N_1788,In_1838,In_7);
or U1789 (N_1789,In_1628,In_601);
or U1790 (N_1790,In_110,In_930);
or U1791 (N_1791,In_1537,In_634);
xnor U1792 (N_1792,In_848,In_375);
nand U1793 (N_1793,In_918,In_790);
xnor U1794 (N_1794,In_1079,In_1300);
nor U1795 (N_1795,In_817,In_1075);
nor U1796 (N_1796,In_235,In_424);
and U1797 (N_1797,In_1381,In_1330);
or U1798 (N_1798,In_1980,In_129);
nor U1799 (N_1799,In_1846,In_1159);
nor U1800 (N_1800,In_1490,In_1489);
nand U1801 (N_1801,In_1480,In_681);
and U1802 (N_1802,In_57,In_547);
nor U1803 (N_1803,In_862,In_1594);
and U1804 (N_1804,In_62,In_1683);
and U1805 (N_1805,In_1612,In_1017);
nor U1806 (N_1806,In_1332,In_99);
nor U1807 (N_1807,In_1404,In_441);
nor U1808 (N_1808,In_180,In_847);
and U1809 (N_1809,In_201,In_1761);
or U1810 (N_1810,In_1150,In_668);
nand U1811 (N_1811,In_259,In_1435);
and U1812 (N_1812,In_1358,In_1977);
nor U1813 (N_1813,In_1477,In_1871);
nor U1814 (N_1814,In_165,In_728);
nor U1815 (N_1815,In_444,In_321);
nand U1816 (N_1816,In_534,In_1502);
nand U1817 (N_1817,In_1949,In_878);
nand U1818 (N_1818,In_1921,In_812);
nor U1819 (N_1819,In_828,In_728);
nand U1820 (N_1820,In_1669,In_677);
or U1821 (N_1821,In_1189,In_1388);
nor U1822 (N_1822,In_667,In_427);
and U1823 (N_1823,In_112,In_1545);
and U1824 (N_1824,In_387,In_815);
and U1825 (N_1825,In_1477,In_1037);
and U1826 (N_1826,In_1097,In_281);
nor U1827 (N_1827,In_1820,In_1725);
nand U1828 (N_1828,In_1208,In_82);
and U1829 (N_1829,In_1252,In_745);
nor U1830 (N_1830,In_1898,In_859);
nand U1831 (N_1831,In_194,In_178);
or U1832 (N_1832,In_1943,In_1023);
nor U1833 (N_1833,In_1652,In_423);
nor U1834 (N_1834,In_515,In_64);
or U1835 (N_1835,In_337,In_281);
nand U1836 (N_1836,In_1627,In_1891);
nand U1837 (N_1837,In_1196,In_1646);
nand U1838 (N_1838,In_1590,In_1971);
or U1839 (N_1839,In_578,In_1873);
and U1840 (N_1840,In_351,In_1630);
and U1841 (N_1841,In_1789,In_614);
or U1842 (N_1842,In_385,In_1021);
and U1843 (N_1843,In_1976,In_1569);
nor U1844 (N_1844,In_721,In_120);
nand U1845 (N_1845,In_771,In_115);
nor U1846 (N_1846,In_1931,In_912);
nand U1847 (N_1847,In_705,In_484);
nand U1848 (N_1848,In_767,In_545);
or U1849 (N_1849,In_32,In_1386);
nor U1850 (N_1850,In_1246,In_75);
or U1851 (N_1851,In_566,In_1728);
or U1852 (N_1852,In_1156,In_865);
nand U1853 (N_1853,In_187,In_1543);
and U1854 (N_1854,In_1825,In_396);
and U1855 (N_1855,In_210,In_939);
nor U1856 (N_1856,In_635,In_1467);
or U1857 (N_1857,In_846,In_1708);
and U1858 (N_1858,In_1003,In_1053);
nor U1859 (N_1859,In_1190,In_251);
nor U1860 (N_1860,In_1896,In_402);
or U1861 (N_1861,In_1911,In_62);
or U1862 (N_1862,In_707,In_466);
or U1863 (N_1863,In_1648,In_186);
or U1864 (N_1864,In_471,In_1228);
and U1865 (N_1865,In_647,In_194);
or U1866 (N_1866,In_1546,In_1552);
or U1867 (N_1867,In_1012,In_360);
nand U1868 (N_1868,In_414,In_1119);
nand U1869 (N_1869,In_1522,In_1412);
nand U1870 (N_1870,In_1570,In_410);
nor U1871 (N_1871,In_643,In_783);
or U1872 (N_1872,In_846,In_46);
or U1873 (N_1873,In_924,In_310);
and U1874 (N_1874,In_1762,In_1519);
and U1875 (N_1875,In_826,In_1586);
and U1876 (N_1876,In_1825,In_1991);
and U1877 (N_1877,In_657,In_846);
or U1878 (N_1878,In_1837,In_828);
nor U1879 (N_1879,In_338,In_1701);
nor U1880 (N_1880,In_1560,In_1764);
nand U1881 (N_1881,In_1504,In_1276);
nand U1882 (N_1882,In_1484,In_587);
or U1883 (N_1883,In_1934,In_711);
nand U1884 (N_1884,In_1523,In_579);
nor U1885 (N_1885,In_192,In_221);
nand U1886 (N_1886,In_1731,In_1990);
nor U1887 (N_1887,In_1097,In_214);
or U1888 (N_1888,In_985,In_478);
or U1889 (N_1889,In_307,In_1169);
nand U1890 (N_1890,In_1436,In_440);
nand U1891 (N_1891,In_1052,In_120);
or U1892 (N_1892,In_850,In_550);
or U1893 (N_1893,In_709,In_1814);
and U1894 (N_1894,In_1713,In_356);
and U1895 (N_1895,In_412,In_139);
and U1896 (N_1896,In_584,In_609);
nor U1897 (N_1897,In_197,In_239);
nand U1898 (N_1898,In_372,In_773);
and U1899 (N_1899,In_1208,In_791);
and U1900 (N_1900,In_1832,In_1733);
and U1901 (N_1901,In_819,In_837);
and U1902 (N_1902,In_46,In_546);
nand U1903 (N_1903,In_1146,In_1528);
or U1904 (N_1904,In_409,In_1930);
or U1905 (N_1905,In_1840,In_906);
and U1906 (N_1906,In_1003,In_313);
nand U1907 (N_1907,In_1880,In_329);
and U1908 (N_1908,In_992,In_599);
and U1909 (N_1909,In_452,In_1718);
and U1910 (N_1910,In_1850,In_359);
and U1911 (N_1911,In_1987,In_421);
nand U1912 (N_1912,In_1021,In_467);
nand U1913 (N_1913,In_1526,In_1118);
nor U1914 (N_1914,In_473,In_1363);
nor U1915 (N_1915,In_496,In_22);
and U1916 (N_1916,In_1312,In_140);
nor U1917 (N_1917,In_1138,In_5);
or U1918 (N_1918,In_353,In_1305);
xnor U1919 (N_1919,In_16,In_754);
or U1920 (N_1920,In_1522,In_1318);
nand U1921 (N_1921,In_1906,In_1717);
and U1922 (N_1922,In_1515,In_97);
nor U1923 (N_1923,In_1144,In_363);
nor U1924 (N_1924,In_33,In_1881);
and U1925 (N_1925,In_18,In_357);
and U1926 (N_1926,In_333,In_1165);
or U1927 (N_1927,In_949,In_420);
or U1928 (N_1928,In_135,In_439);
nand U1929 (N_1929,In_1854,In_1216);
nand U1930 (N_1930,In_347,In_1607);
and U1931 (N_1931,In_434,In_981);
nor U1932 (N_1932,In_1611,In_1927);
nor U1933 (N_1933,In_480,In_753);
nand U1934 (N_1934,In_732,In_1957);
nand U1935 (N_1935,In_223,In_85);
nor U1936 (N_1936,In_1776,In_1971);
and U1937 (N_1937,In_1034,In_876);
nand U1938 (N_1938,In_685,In_553);
nand U1939 (N_1939,In_260,In_1331);
and U1940 (N_1940,In_1245,In_1233);
nand U1941 (N_1941,In_525,In_1321);
and U1942 (N_1942,In_576,In_876);
nor U1943 (N_1943,In_345,In_114);
nor U1944 (N_1944,In_1233,In_252);
nand U1945 (N_1945,In_442,In_1667);
nand U1946 (N_1946,In_444,In_1211);
nor U1947 (N_1947,In_1858,In_938);
and U1948 (N_1948,In_34,In_971);
or U1949 (N_1949,In_1120,In_658);
and U1950 (N_1950,In_187,In_850);
nand U1951 (N_1951,In_781,In_1525);
and U1952 (N_1952,In_529,In_399);
nor U1953 (N_1953,In_304,In_385);
or U1954 (N_1954,In_919,In_278);
nor U1955 (N_1955,In_1172,In_1683);
nor U1956 (N_1956,In_1181,In_1035);
and U1957 (N_1957,In_724,In_1090);
nor U1958 (N_1958,In_181,In_1251);
and U1959 (N_1959,In_1861,In_590);
or U1960 (N_1960,In_1507,In_272);
nor U1961 (N_1961,In_511,In_1135);
nand U1962 (N_1962,In_451,In_759);
or U1963 (N_1963,In_1345,In_1827);
nor U1964 (N_1964,In_1219,In_168);
and U1965 (N_1965,In_623,In_1620);
nor U1966 (N_1966,In_1311,In_1437);
nor U1967 (N_1967,In_1167,In_587);
nand U1968 (N_1968,In_1244,In_350);
nor U1969 (N_1969,In_388,In_325);
or U1970 (N_1970,In_842,In_674);
nor U1971 (N_1971,In_634,In_1402);
or U1972 (N_1972,In_607,In_1467);
nor U1973 (N_1973,In_1016,In_1384);
and U1974 (N_1974,In_749,In_961);
nand U1975 (N_1975,In_1616,In_1363);
or U1976 (N_1976,In_1765,In_1431);
nand U1977 (N_1977,In_376,In_1180);
nand U1978 (N_1978,In_1670,In_1930);
or U1979 (N_1979,In_1581,In_555);
nand U1980 (N_1980,In_1949,In_956);
or U1981 (N_1981,In_1711,In_165);
xor U1982 (N_1982,In_1561,In_396);
nor U1983 (N_1983,In_1298,In_904);
and U1984 (N_1984,In_630,In_303);
and U1985 (N_1985,In_731,In_831);
nand U1986 (N_1986,In_1897,In_1398);
and U1987 (N_1987,In_720,In_440);
or U1988 (N_1988,In_1047,In_362);
nand U1989 (N_1989,In_1198,In_996);
or U1990 (N_1990,In_58,In_495);
and U1991 (N_1991,In_1198,In_262);
and U1992 (N_1992,In_1895,In_1747);
nor U1993 (N_1993,In_1063,In_642);
and U1994 (N_1994,In_634,In_982);
nor U1995 (N_1995,In_847,In_760);
xor U1996 (N_1996,In_628,In_1632);
nor U1997 (N_1997,In_444,In_209);
and U1998 (N_1998,In_1965,In_1875);
nor U1999 (N_1999,In_972,In_1784);
nor U2000 (N_2000,In_1903,In_366);
and U2001 (N_2001,In_1733,In_575);
or U2002 (N_2002,In_1172,In_1701);
and U2003 (N_2003,In_1486,In_1462);
nor U2004 (N_2004,In_119,In_1503);
or U2005 (N_2005,In_1513,In_65);
and U2006 (N_2006,In_646,In_1712);
and U2007 (N_2007,In_658,In_646);
nand U2008 (N_2008,In_1001,In_1595);
nor U2009 (N_2009,In_842,In_1734);
nor U2010 (N_2010,In_1936,In_1141);
nand U2011 (N_2011,In_1296,In_1509);
nor U2012 (N_2012,In_1832,In_783);
nor U2013 (N_2013,In_1524,In_857);
nor U2014 (N_2014,In_1919,In_1179);
and U2015 (N_2015,In_1575,In_1524);
and U2016 (N_2016,In_544,In_672);
nand U2017 (N_2017,In_985,In_1647);
nor U2018 (N_2018,In_402,In_1582);
nand U2019 (N_2019,In_1590,In_95);
and U2020 (N_2020,In_1345,In_1783);
nand U2021 (N_2021,In_1477,In_1630);
or U2022 (N_2022,In_413,In_1646);
nand U2023 (N_2023,In_1326,In_284);
or U2024 (N_2024,In_157,In_705);
and U2025 (N_2025,In_1879,In_255);
or U2026 (N_2026,In_518,In_274);
or U2027 (N_2027,In_1095,In_295);
nor U2028 (N_2028,In_532,In_296);
or U2029 (N_2029,In_139,In_1531);
and U2030 (N_2030,In_758,In_897);
or U2031 (N_2031,In_13,In_297);
or U2032 (N_2032,In_601,In_465);
or U2033 (N_2033,In_291,In_1521);
nand U2034 (N_2034,In_1471,In_931);
or U2035 (N_2035,In_605,In_1516);
nand U2036 (N_2036,In_1408,In_1725);
nand U2037 (N_2037,In_736,In_285);
nand U2038 (N_2038,In_671,In_401);
and U2039 (N_2039,In_661,In_726);
and U2040 (N_2040,In_1534,In_503);
nand U2041 (N_2041,In_1145,In_98);
and U2042 (N_2042,In_1606,In_791);
nor U2043 (N_2043,In_1406,In_1664);
nand U2044 (N_2044,In_1839,In_1966);
and U2045 (N_2045,In_1441,In_700);
nand U2046 (N_2046,In_690,In_1044);
nand U2047 (N_2047,In_1930,In_1548);
nor U2048 (N_2048,In_66,In_146);
nor U2049 (N_2049,In_471,In_57);
and U2050 (N_2050,In_1502,In_311);
nor U2051 (N_2051,In_635,In_1742);
nand U2052 (N_2052,In_485,In_329);
and U2053 (N_2053,In_425,In_540);
and U2054 (N_2054,In_509,In_622);
nand U2055 (N_2055,In_179,In_794);
nand U2056 (N_2056,In_981,In_49);
or U2057 (N_2057,In_658,In_1595);
and U2058 (N_2058,In_461,In_134);
or U2059 (N_2059,In_1192,In_1474);
or U2060 (N_2060,In_38,In_1748);
and U2061 (N_2061,In_1382,In_49);
nor U2062 (N_2062,In_901,In_1626);
or U2063 (N_2063,In_399,In_1602);
and U2064 (N_2064,In_640,In_1424);
or U2065 (N_2065,In_1158,In_637);
nor U2066 (N_2066,In_1221,In_85);
nand U2067 (N_2067,In_1340,In_1942);
or U2068 (N_2068,In_454,In_897);
nor U2069 (N_2069,In_1493,In_978);
or U2070 (N_2070,In_337,In_1523);
nor U2071 (N_2071,In_1031,In_808);
nor U2072 (N_2072,In_795,In_1587);
or U2073 (N_2073,In_1705,In_915);
nand U2074 (N_2074,In_575,In_1015);
and U2075 (N_2075,In_1501,In_1853);
or U2076 (N_2076,In_123,In_1257);
nand U2077 (N_2077,In_1207,In_1901);
nand U2078 (N_2078,In_708,In_272);
nand U2079 (N_2079,In_63,In_55);
or U2080 (N_2080,In_1127,In_470);
nand U2081 (N_2081,In_711,In_1365);
nand U2082 (N_2082,In_1739,In_319);
and U2083 (N_2083,In_1184,In_830);
and U2084 (N_2084,In_487,In_1651);
or U2085 (N_2085,In_1410,In_556);
nand U2086 (N_2086,In_1712,In_730);
or U2087 (N_2087,In_1151,In_1109);
nor U2088 (N_2088,In_1892,In_1986);
or U2089 (N_2089,In_386,In_1506);
nand U2090 (N_2090,In_654,In_463);
and U2091 (N_2091,In_253,In_175);
nand U2092 (N_2092,In_1673,In_1434);
nand U2093 (N_2093,In_1785,In_633);
nand U2094 (N_2094,In_131,In_345);
nor U2095 (N_2095,In_153,In_115);
nand U2096 (N_2096,In_1992,In_1439);
and U2097 (N_2097,In_1195,In_36);
or U2098 (N_2098,In_784,In_1073);
nor U2099 (N_2099,In_288,In_218);
or U2100 (N_2100,In_1907,In_1096);
or U2101 (N_2101,In_739,In_121);
or U2102 (N_2102,In_145,In_756);
or U2103 (N_2103,In_1275,In_600);
nor U2104 (N_2104,In_1371,In_124);
nor U2105 (N_2105,In_809,In_995);
or U2106 (N_2106,In_1152,In_1220);
nor U2107 (N_2107,In_1385,In_1568);
nor U2108 (N_2108,In_475,In_1720);
or U2109 (N_2109,In_1785,In_8);
and U2110 (N_2110,In_1056,In_402);
nand U2111 (N_2111,In_964,In_317);
or U2112 (N_2112,In_731,In_1755);
and U2113 (N_2113,In_1796,In_1854);
nor U2114 (N_2114,In_1203,In_1151);
nand U2115 (N_2115,In_931,In_1213);
and U2116 (N_2116,In_1467,In_760);
and U2117 (N_2117,In_1193,In_1217);
nor U2118 (N_2118,In_1193,In_363);
nor U2119 (N_2119,In_763,In_991);
nor U2120 (N_2120,In_899,In_1350);
or U2121 (N_2121,In_1427,In_147);
nand U2122 (N_2122,In_1051,In_1043);
nand U2123 (N_2123,In_1010,In_1884);
nand U2124 (N_2124,In_494,In_1934);
or U2125 (N_2125,In_738,In_1974);
nor U2126 (N_2126,In_574,In_857);
or U2127 (N_2127,In_77,In_499);
nor U2128 (N_2128,In_1590,In_1778);
nand U2129 (N_2129,In_73,In_1378);
nand U2130 (N_2130,In_894,In_110);
nor U2131 (N_2131,In_1198,In_1066);
nand U2132 (N_2132,In_460,In_1727);
nand U2133 (N_2133,In_914,In_1243);
and U2134 (N_2134,In_162,In_548);
or U2135 (N_2135,In_628,In_1412);
or U2136 (N_2136,In_660,In_1672);
or U2137 (N_2137,In_1438,In_415);
or U2138 (N_2138,In_1845,In_1211);
or U2139 (N_2139,In_563,In_1529);
nand U2140 (N_2140,In_834,In_664);
or U2141 (N_2141,In_995,In_813);
nand U2142 (N_2142,In_1434,In_800);
nand U2143 (N_2143,In_411,In_1588);
or U2144 (N_2144,In_972,In_1844);
nand U2145 (N_2145,In_1524,In_1729);
nand U2146 (N_2146,In_1858,In_456);
or U2147 (N_2147,In_842,In_1708);
nand U2148 (N_2148,In_338,In_775);
and U2149 (N_2149,In_829,In_627);
or U2150 (N_2150,In_1267,In_1821);
or U2151 (N_2151,In_1465,In_699);
and U2152 (N_2152,In_69,In_1327);
or U2153 (N_2153,In_457,In_1016);
nor U2154 (N_2154,In_1555,In_1363);
or U2155 (N_2155,In_316,In_1749);
nand U2156 (N_2156,In_988,In_1811);
and U2157 (N_2157,In_1786,In_1341);
and U2158 (N_2158,In_1043,In_1937);
nand U2159 (N_2159,In_928,In_150);
or U2160 (N_2160,In_447,In_1188);
nor U2161 (N_2161,In_712,In_48);
nor U2162 (N_2162,In_135,In_1520);
nand U2163 (N_2163,In_1021,In_1483);
nor U2164 (N_2164,In_1835,In_1363);
nand U2165 (N_2165,In_871,In_1821);
or U2166 (N_2166,In_1394,In_1265);
and U2167 (N_2167,In_176,In_867);
nor U2168 (N_2168,In_1156,In_1811);
or U2169 (N_2169,In_1093,In_1736);
nor U2170 (N_2170,In_1964,In_1893);
or U2171 (N_2171,In_602,In_1745);
or U2172 (N_2172,In_631,In_1696);
nand U2173 (N_2173,In_266,In_166);
or U2174 (N_2174,In_120,In_737);
or U2175 (N_2175,In_1654,In_531);
nor U2176 (N_2176,In_1229,In_1665);
or U2177 (N_2177,In_1141,In_1);
or U2178 (N_2178,In_698,In_632);
and U2179 (N_2179,In_797,In_630);
and U2180 (N_2180,In_927,In_306);
and U2181 (N_2181,In_1846,In_710);
or U2182 (N_2182,In_1933,In_790);
or U2183 (N_2183,In_783,In_536);
nor U2184 (N_2184,In_554,In_607);
and U2185 (N_2185,In_137,In_1437);
or U2186 (N_2186,In_1756,In_742);
nor U2187 (N_2187,In_1530,In_30);
nand U2188 (N_2188,In_388,In_1023);
nand U2189 (N_2189,In_1892,In_792);
nand U2190 (N_2190,In_659,In_1218);
and U2191 (N_2191,In_38,In_1529);
and U2192 (N_2192,In_1478,In_151);
and U2193 (N_2193,In_1956,In_1451);
xnor U2194 (N_2194,In_735,In_943);
and U2195 (N_2195,In_462,In_652);
and U2196 (N_2196,In_367,In_538);
and U2197 (N_2197,In_59,In_516);
and U2198 (N_2198,In_1986,In_133);
nor U2199 (N_2199,In_989,In_1415);
and U2200 (N_2200,In_1694,In_731);
nor U2201 (N_2201,In_729,In_409);
nand U2202 (N_2202,In_1859,In_1816);
nor U2203 (N_2203,In_386,In_838);
or U2204 (N_2204,In_314,In_1063);
xnor U2205 (N_2205,In_834,In_1054);
nor U2206 (N_2206,In_1793,In_610);
or U2207 (N_2207,In_1411,In_369);
nand U2208 (N_2208,In_504,In_1508);
nor U2209 (N_2209,In_988,In_1883);
nand U2210 (N_2210,In_1759,In_1267);
nor U2211 (N_2211,In_1375,In_1191);
or U2212 (N_2212,In_1959,In_20);
xnor U2213 (N_2213,In_741,In_1576);
and U2214 (N_2214,In_701,In_431);
nand U2215 (N_2215,In_304,In_1891);
and U2216 (N_2216,In_114,In_557);
nor U2217 (N_2217,In_1497,In_1766);
nand U2218 (N_2218,In_358,In_1132);
nor U2219 (N_2219,In_1015,In_1713);
nand U2220 (N_2220,In_1458,In_731);
nor U2221 (N_2221,In_1788,In_1665);
or U2222 (N_2222,In_936,In_1099);
nand U2223 (N_2223,In_279,In_897);
nand U2224 (N_2224,In_1997,In_1167);
or U2225 (N_2225,In_922,In_928);
and U2226 (N_2226,In_234,In_1108);
or U2227 (N_2227,In_254,In_1532);
nor U2228 (N_2228,In_921,In_180);
nor U2229 (N_2229,In_1456,In_1345);
or U2230 (N_2230,In_1575,In_458);
nor U2231 (N_2231,In_1486,In_1807);
and U2232 (N_2232,In_114,In_1408);
nor U2233 (N_2233,In_1888,In_222);
nor U2234 (N_2234,In_1817,In_1593);
nand U2235 (N_2235,In_1960,In_247);
nor U2236 (N_2236,In_1669,In_689);
nand U2237 (N_2237,In_511,In_553);
or U2238 (N_2238,In_996,In_1134);
or U2239 (N_2239,In_1873,In_1798);
or U2240 (N_2240,In_497,In_510);
or U2241 (N_2241,In_1142,In_800);
and U2242 (N_2242,In_797,In_249);
or U2243 (N_2243,In_979,In_783);
and U2244 (N_2244,In_1950,In_1773);
or U2245 (N_2245,In_513,In_318);
nor U2246 (N_2246,In_1293,In_956);
nand U2247 (N_2247,In_1313,In_1901);
nor U2248 (N_2248,In_543,In_1375);
and U2249 (N_2249,In_1328,In_1993);
nand U2250 (N_2250,In_630,In_1083);
or U2251 (N_2251,In_1341,In_1950);
nand U2252 (N_2252,In_105,In_1045);
or U2253 (N_2253,In_1342,In_1776);
and U2254 (N_2254,In_1911,In_1627);
and U2255 (N_2255,In_1598,In_1367);
or U2256 (N_2256,In_1767,In_1696);
nand U2257 (N_2257,In_783,In_1449);
nor U2258 (N_2258,In_1536,In_398);
and U2259 (N_2259,In_1945,In_438);
nand U2260 (N_2260,In_982,In_1476);
nor U2261 (N_2261,In_718,In_1152);
nand U2262 (N_2262,In_1053,In_272);
and U2263 (N_2263,In_74,In_446);
nand U2264 (N_2264,In_1266,In_1471);
or U2265 (N_2265,In_1828,In_1265);
nand U2266 (N_2266,In_447,In_923);
nand U2267 (N_2267,In_1808,In_36);
or U2268 (N_2268,In_1909,In_652);
or U2269 (N_2269,In_1702,In_1351);
nand U2270 (N_2270,In_1087,In_1344);
nand U2271 (N_2271,In_305,In_754);
or U2272 (N_2272,In_387,In_46);
and U2273 (N_2273,In_685,In_388);
nor U2274 (N_2274,In_629,In_772);
and U2275 (N_2275,In_1347,In_1248);
or U2276 (N_2276,In_885,In_1056);
nand U2277 (N_2277,In_490,In_1278);
nor U2278 (N_2278,In_807,In_551);
or U2279 (N_2279,In_656,In_1099);
and U2280 (N_2280,In_1501,In_1874);
and U2281 (N_2281,In_535,In_1857);
or U2282 (N_2282,In_1555,In_1525);
and U2283 (N_2283,In_597,In_1718);
and U2284 (N_2284,In_1355,In_1936);
nor U2285 (N_2285,In_970,In_611);
nand U2286 (N_2286,In_888,In_1893);
or U2287 (N_2287,In_1371,In_110);
nand U2288 (N_2288,In_781,In_821);
or U2289 (N_2289,In_983,In_227);
and U2290 (N_2290,In_1935,In_560);
or U2291 (N_2291,In_560,In_1761);
or U2292 (N_2292,In_862,In_342);
or U2293 (N_2293,In_479,In_1312);
nand U2294 (N_2294,In_952,In_1744);
nor U2295 (N_2295,In_1275,In_468);
nor U2296 (N_2296,In_175,In_917);
nor U2297 (N_2297,In_752,In_1773);
and U2298 (N_2298,In_370,In_1709);
and U2299 (N_2299,In_1712,In_1876);
nand U2300 (N_2300,In_1657,In_124);
and U2301 (N_2301,In_36,In_1309);
nor U2302 (N_2302,In_885,In_1135);
and U2303 (N_2303,In_884,In_1898);
nand U2304 (N_2304,In_1128,In_1917);
and U2305 (N_2305,In_741,In_795);
nand U2306 (N_2306,In_1044,In_1135);
or U2307 (N_2307,In_491,In_41);
nand U2308 (N_2308,In_1367,In_1604);
nor U2309 (N_2309,In_186,In_311);
nor U2310 (N_2310,In_1633,In_423);
nor U2311 (N_2311,In_1812,In_1282);
and U2312 (N_2312,In_579,In_162);
and U2313 (N_2313,In_3,In_1364);
nor U2314 (N_2314,In_133,In_1145);
nor U2315 (N_2315,In_449,In_1174);
nand U2316 (N_2316,In_1511,In_1695);
nand U2317 (N_2317,In_690,In_1134);
nand U2318 (N_2318,In_1974,In_176);
nand U2319 (N_2319,In_1150,In_1295);
and U2320 (N_2320,In_1919,In_1639);
or U2321 (N_2321,In_1902,In_1107);
and U2322 (N_2322,In_838,In_424);
nand U2323 (N_2323,In_1295,In_1154);
or U2324 (N_2324,In_547,In_737);
nor U2325 (N_2325,In_938,In_1456);
xnor U2326 (N_2326,In_1131,In_1760);
and U2327 (N_2327,In_633,In_1943);
or U2328 (N_2328,In_285,In_232);
nor U2329 (N_2329,In_1865,In_1947);
nand U2330 (N_2330,In_433,In_1360);
nor U2331 (N_2331,In_1424,In_1167);
and U2332 (N_2332,In_354,In_1428);
nor U2333 (N_2333,In_1233,In_1897);
nand U2334 (N_2334,In_1046,In_1448);
nor U2335 (N_2335,In_964,In_1267);
or U2336 (N_2336,In_939,In_1536);
and U2337 (N_2337,In_1446,In_1431);
and U2338 (N_2338,In_269,In_948);
or U2339 (N_2339,In_649,In_433);
nand U2340 (N_2340,In_400,In_1939);
and U2341 (N_2341,In_1468,In_1559);
and U2342 (N_2342,In_1402,In_85);
nor U2343 (N_2343,In_1368,In_13);
nor U2344 (N_2344,In_1537,In_1692);
nand U2345 (N_2345,In_224,In_592);
and U2346 (N_2346,In_907,In_1239);
or U2347 (N_2347,In_975,In_875);
nor U2348 (N_2348,In_1935,In_46);
nor U2349 (N_2349,In_1056,In_220);
nor U2350 (N_2350,In_1984,In_924);
nand U2351 (N_2351,In_1148,In_740);
and U2352 (N_2352,In_1777,In_1727);
nor U2353 (N_2353,In_1586,In_372);
nand U2354 (N_2354,In_350,In_1850);
and U2355 (N_2355,In_50,In_426);
or U2356 (N_2356,In_1628,In_526);
or U2357 (N_2357,In_720,In_1499);
xor U2358 (N_2358,In_1269,In_134);
and U2359 (N_2359,In_1725,In_98);
or U2360 (N_2360,In_1940,In_1046);
nand U2361 (N_2361,In_917,In_1049);
nor U2362 (N_2362,In_809,In_740);
and U2363 (N_2363,In_1671,In_1870);
nor U2364 (N_2364,In_1371,In_1250);
nand U2365 (N_2365,In_188,In_482);
or U2366 (N_2366,In_1832,In_334);
and U2367 (N_2367,In_1549,In_1113);
nor U2368 (N_2368,In_49,In_498);
nand U2369 (N_2369,In_330,In_1404);
nor U2370 (N_2370,In_1408,In_1694);
or U2371 (N_2371,In_1769,In_1495);
and U2372 (N_2372,In_444,In_435);
nand U2373 (N_2373,In_101,In_371);
or U2374 (N_2374,In_811,In_1164);
nor U2375 (N_2375,In_678,In_1435);
nor U2376 (N_2376,In_439,In_566);
and U2377 (N_2377,In_391,In_1551);
nor U2378 (N_2378,In_1227,In_1317);
and U2379 (N_2379,In_1725,In_1898);
nand U2380 (N_2380,In_1289,In_1713);
or U2381 (N_2381,In_1600,In_1408);
or U2382 (N_2382,In_1920,In_289);
or U2383 (N_2383,In_212,In_1346);
or U2384 (N_2384,In_1832,In_957);
or U2385 (N_2385,In_279,In_223);
nor U2386 (N_2386,In_1660,In_1914);
nor U2387 (N_2387,In_1151,In_1);
or U2388 (N_2388,In_80,In_85);
nand U2389 (N_2389,In_650,In_863);
nand U2390 (N_2390,In_1202,In_1793);
or U2391 (N_2391,In_86,In_1229);
or U2392 (N_2392,In_1001,In_772);
and U2393 (N_2393,In_594,In_378);
or U2394 (N_2394,In_1435,In_1942);
nor U2395 (N_2395,In_756,In_1163);
and U2396 (N_2396,In_1387,In_1101);
nand U2397 (N_2397,In_141,In_1411);
and U2398 (N_2398,In_592,In_1999);
nor U2399 (N_2399,In_1633,In_506);
or U2400 (N_2400,In_679,In_1398);
or U2401 (N_2401,In_692,In_705);
nand U2402 (N_2402,In_1572,In_726);
or U2403 (N_2403,In_1409,In_1198);
or U2404 (N_2404,In_135,In_479);
nand U2405 (N_2405,In_215,In_809);
or U2406 (N_2406,In_1792,In_492);
nand U2407 (N_2407,In_769,In_794);
or U2408 (N_2408,In_1495,In_28);
nand U2409 (N_2409,In_1486,In_1635);
nor U2410 (N_2410,In_1140,In_1373);
nor U2411 (N_2411,In_1362,In_786);
nand U2412 (N_2412,In_1246,In_474);
nor U2413 (N_2413,In_125,In_240);
and U2414 (N_2414,In_315,In_363);
or U2415 (N_2415,In_1972,In_1593);
and U2416 (N_2416,In_1662,In_1088);
nand U2417 (N_2417,In_1407,In_2);
nor U2418 (N_2418,In_1617,In_603);
and U2419 (N_2419,In_243,In_652);
or U2420 (N_2420,In_537,In_1467);
nor U2421 (N_2421,In_1131,In_1441);
nor U2422 (N_2422,In_1590,In_632);
nor U2423 (N_2423,In_1914,In_129);
and U2424 (N_2424,In_160,In_1979);
nand U2425 (N_2425,In_99,In_1614);
and U2426 (N_2426,In_740,In_338);
nand U2427 (N_2427,In_370,In_910);
or U2428 (N_2428,In_95,In_626);
or U2429 (N_2429,In_1683,In_628);
and U2430 (N_2430,In_865,In_682);
or U2431 (N_2431,In_252,In_1899);
or U2432 (N_2432,In_674,In_669);
and U2433 (N_2433,In_493,In_836);
nor U2434 (N_2434,In_331,In_1734);
nand U2435 (N_2435,In_1960,In_115);
nand U2436 (N_2436,In_712,In_1280);
nor U2437 (N_2437,In_1250,In_1400);
or U2438 (N_2438,In_969,In_1347);
nor U2439 (N_2439,In_1171,In_316);
and U2440 (N_2440,In_1970,In_456);
nand U2441 (N_2441,In_369,In_1407);
nand U2442 (N_2442,In_471,In_220);
nand U2443 (N_2443,In_1312,In_790);
nand U2444 (N_2444,In_1997,In_1623);
nor U2445 (N_2445,In_1120,In_1982);
or U2446 (N_2446,In_211,In_1816);
xor U2447 (N_2447,In_801,In_1582);
or U2448 (N_2448,In_1922,In_390);
or U2449 (N_2449,In_512,In_353);
and U2450 (N_2450,In_1998,In_465);
and U2451 (N_2451,In_1853,In_636);
or U2452 (N_2452,In_494,In_322);
and U2453 (N_2453,In_412,In_686);
nor U2454 (N_2454,In_621,In_1736);
and U2455 (N_2455,In_1650,In_810);
and U2456 (N_2456,In_418,In_1625);
and U2457 (N_2457,In_1786,In_793);
or U2458 (N_2458,In_304,In_964);
and U2459 (N_2459,In_927,In_106);
nor U2460 (N_2460,In_1620,In_979);
and U2461 (N_2461,In_559,In_351);
nor U2462 (N_2462,In_1821,In_1651);
xnor U2463 (N_2463,In_896,In_250);
nand U2464 (N_2464,In_894,In_431);
nand U2465 (N_2465,In_36,In_664);
or U2466 (N_2466,In_241,In_16);
or U2467 (N_2467,In_1113,In_1347);
or U2468 (N_2468,In_1964,In_637);
or U2469 (N_2469,In_644,In_359);
xor U2470 (N_2470,In_1009,In_963);
nor U2471 (N_2471,In_558,In_1073);
or U2472 (N_2472,In_738,In_1084);
and U2473 (N_2473,In_667,In_1029);
and U2474 (N_2474,In_706,In_506);
nand U2475 (N_2475,In_760,In_280);
and U2476 (N_2476,In_1608,In_215);
nor U2477 (N_2477,In_1594,In_1803);
or U2478 (N_2478,In_1055,In_1797);
or U2479 (N_2479,In_1458,In_1412);
or U2480 (N_2480,In_538,In_192);
and U2481 (N_2481,In_629,In_1668);
nor U2482 (N_2482,In_1624,In_1087);
nor U2483 (N_2483,In_637,In_812);
and U2484 (N_2484,In_472,In_418);
nand U2485 (N_2485,In_691,In_1223);
or U2486 (N_2486,In_174,In_1472);
and U2487 (N_2487,In_1111,In_1672);
and U2488 (N_2488,In_211,In_0);
and U2489 (N_2489,In_918,In_1876);
or U2490 (N_2490,In_1542,In_1362);
nor U2491 (N_2491,In_783,In_796);
or U2492 (N_2492,In_1130,In_1009);
nor U2493 (N_2493,In_521,In_926);
or U2494 (N_2494,In_1635,In_727);
or U2495 (N_2495,In_1012,In_823);
nand U2496 (N_2496,In_262,In_1731);
nor U2497 (N_2497,In_231,In_927);
nor U2498 (N_2498,In_1038,In_1071);
nand U2499 (N_2499,In_234,In_933);
or U2500 (N_2500,In_386,In_1203);
and U2501 (N_2501,In_1351,In_298);
nand U2502 (N_2502,In_477,In_1687);
or U2503 (N_2503,In_179,In_859);
nor U2504 (N_2504,In_1427,In_1830);
or U2505 (N_2505,In_1502,In_1120);
nand U2506 (N_2506,In_1519,In_294);
and U2507 (N_2507,In_1871,In_1106);
and U2508 (N_2508,In_443,In_470);
and U2509 (N_2509,In_1352,In_1091);
or U2510 (N_2510,In_989,In_1963);
or U2511 (N_2511,In_1322,In_1071);
or U2512 (N_2512,In_386,In_83);
nor U2513 (N_2513,In_1475,In_1935);
nor U2514 (N_2514,In_589,In_1459);
or U2515 (N_2515,In_1685,In_64);
nand U2516 (N_2516,In_880,In_1956);
and U2517 (N_2517,In_492,In_1635);
nand U2518 (N_2518,In_1160,In_840);
nor U2519 (N_2519,In_521,In_1979);
and U2520 (N_2520,In_534,In_1397);
or U2521 (N_2521,In_1789,In_442);
nand U2522 (N_2522,In_515,In_1159);
or U2523 (N_2523,In_794,In_1580);
nand U2524 (N_2524,In_1156,In_1803);
and U2525 (N_2525,In_93,In_1962);
or U2526 (N_2526,In_789,In_1938);
nor U2527 (N_2527,In_836,In_715);
or U2528 (N_2528,In_1736,In_1733);
nor U2529 (N_2529,In_1724,In_420);
or U2530 (N_2530,In_1221,In_717);
nor U2531 (N_2531,In_381,In_97);
nor U2532 (N_2532,In_1562,In_1999);
and U2533 (N_2533,In_1045,In_199);
nor U2534 (N_2534,In_776,In_1081);
nor U2535 (N_2535,In_321,In_1397);
and U2536 (N_2536,In_1606,In_1109);
nor U2537 (N_2537,In_1716,In_1439);
nor U2538 (N_2538,In_778,In_667);
or U2539 (N_2539,In_1245,In_63);
and U2540 (N_2540,In_478,In_397);
nand U2541 (N_2541,In_1729,In_477);
and U2542 (N_2542,In_1760,In_529);
and U2543 (N_2543,In_779,In_1309);
and U2544 (N_2544,In_475,In_1079);
nand U2545 (N_2545,In_645,In_161);
and U2546 (N_2546,In_1503,In_1062);
and U2547 (N_2547,In_1389,In_639);
nand U2548 (N_2548,In_1374,In_1899);
and U2549 (N_2549,In_1986,In_1086);
or U2550 (N_2550,In_1988,In_660);
and U2551 (N_2551,In_814,In_428);
nand U2552 (N_2552,In_1088,In_1536);
nand U2553 (N_2553,In_491,In_413);
nand U2554 (N_2554,In_930,In_1888);
or U2555 (N_2555,In_839,In_323);
or U2556 (N_2556,In_322,In_458);
and U2557 (N_2557,In_1105,In_333);
or U2558 (N_2558,In_1359,In_81);
xnor U2559 (N_2559,In_448,In_666);
nand U2560 (N_2560,In_18,In_161);
nand U2561 (N_2561,In_359,In_806);
nand U2562 (N_2562,In_134,In_546);
and U2563 (N_2563,In_348,In_1768);
and U2564 (N_2564,In_364,In_1198);
and U2565 (N_2565,In_1872,In_259);
nor U2566 (N_2566,In_623,In_1052);
and U2567 (N_2567,In_135,In_7);
nor U2568 (N_2568,In_898,In_1383);
or U2569 (N_2569,In_887,In_1642);
nor U2570 (N_2570,In_1315,In_1540);
and U2571 (N_2571,In_1100,In_607);
nand U2572 (N_2572,In_384,In_1709);
nand U2573 (N_2573,In_383,In_983);
nand U2574 (N_2574,In_1382,In_354);
nor U2575 (N_2575,In_633,In_141);
nor U2576 (N_2576,In_334,In_1083);
nand U2577 (N_2577,In_1590,In_772);
nand U2578 (N_2578,In_432,In_1490);
nand U2579 (N_2579,In_357,In_1876);
nor U2580 (N_2580,In_14,In_644);
and U2581 (N_2581,In_1151,In_402);
nor U2582 (N_2582,In_588,In_320);
and U2583 (N_2583,In_867,In_1608);
or U2584 (N_2584,In_1223,In_158);
and U2585 (N_2585,In_306,In_1164);
nor U2586 (N_2586,In_937,In_1044);
nand U2587 (N_2587,In_711,In_338);
nor U2588 (N_2588,In_258,In_1485);
nor U2589 (N_2589,In_1196,In_1852);
nand U2590 (N_2590,In_1932,In_1258);
nor U2591 (N_2591,In_560,In_561);
nand U2592 (N_2592,In_1835,In_289);
nand U2593 (N_2593,In_765,In_187);
and U2594 (N_2594,In_593,In_123);
or U2595 (N_2595,In_1134,In_860);
nor U2596 (N_2596,In_1613,In_1089);
or U2597 (N_2597,In_63,In_603);
and U2598 (N_2598,In_1449,In_955);
nand U2599 (N_2599,In_1292,In_473);
or U2600 (N_2600,In_1226,In_1586);
xnor U2601 (N_2601,In_537,In_1468);
nand U2602 (N_2602,In_1137,In_1134);
nor U2603 (N_2603,In_527,In_1714);
nor U2604 (N_2604,In_979,In_1404);
nand U2605 (N_2605,In_1687,In_1361);
nor U2606 (N_2606,In_1982,In_592);
nand U2607 (N_2607,In_942,In_1296);
or U2608 (N_2608,In_345,In_1656);
nor U2609 (N_2609,In_373,In_709);
and U2610 (N_2610,In_914,In_1107);
nand U2611 (N_2611,In_647,In_649);
and U2612 (N_2612,In_472,In_615);
nand U2613 (N_2613,In_957,In_1414);
or U2614 (N_2614,In_534,In_787);
and U2615 (N_2615,In_1434,In_980);
and U2616 (N_2616,In_775,In_1683);
nand U2617 (N_2617,In_1959,In_1796);
and U2618 (N_2618,In_836,In_915);
nor U2619 (N_2619,In_397,In_665);
xor U2620 (N_2620,In_309,In_1159);
and U2621 (N_2621,In_1389,In_1994);
nand U2622 (N_2622,In_186,In_167);
nand U2623 (N_2623,In_1495,In_1585);
nand U2624 (N_2624,In_596,In_1498);
nor U2625 (N_2625,In_794,In_898);
or U2626 (N_2626,In_774,In_1766);
or U2627 (N_2627,In_1093,In_1698);
or U2628 (N_2628,In_1803,In_615);
nor U2629 (N_2629,In_1240,In_897);
nand U2630 (N_2630,In_1240,In_599);
or U2631 (N_2631,In_795,In_428);
or U2632 (N_2632,In_1375,In_1979);
or U2633 (N_2633,In_563,In_142);
and U2634 (N_2634,In_1336,In_1607);
and U2635 (N_2635,In_1316,In_1023);
and U2636 (N_2636,In_743,In_1507);
and U2637 (N_2637,In_1818,In_311);
nand U2638 (N_2638,In_123,In_1958);
and U2639 (N_2639,In_547,In_932);
nor U2640 (N_2640,In_1751,In_266);
nor U2641 (N_2641,In_1567,In_225);
and U2642 (N_2642,In_1842,In_244);
and U2643 (N_2643,In_1639,In_850);
and U2644 (N_2644,In_1726,In_753);
nand U2645 (N_2645,In_886,In_119);
nor U2646 (N_2646,In_637,In_1574);
or U2647 (N_2647,In_1185,In_80);
or U2648 (N_2648,In_1557,In_1748);
and U2649 (N_2649,In_964,In_1368);
nor U2650 (N_2650,In_805,In_1815);
or U2651 (N_2651,In_1259,In_1356);
nand U2652 (N_2652,In_87,In_1564);
and U2653 (N_2653,In_1588,In_576);
or U2654 (N_2654,In_985,In_1278);
nor U2655 (N_2655,In_947,In_1717);
nor U2656 (N_2656,In_481,In_546);
or U2657 (N_2657,In_278,In_1459);
nor U2658 (N_2658,In_1800,In_1434);
or U2659 (N_2659,In_157,In_229);
or U2660 (N_2660,In_448,In_1593);
or U2661 (N_2661,In_964,In_602);
or U2662 (N_2662,In_353,In_1682);
or U2663 (N_2663,In_663,In_1958);
or U2664 (N_2664,In_767,In_1842);
or U2665 (N_2665,In_540,In_1511);
nor U2666 (N_2666,In_964,In_496);
nand U2667 (N_2667,In_1024,In_900);
and U2668 (N_2668,In_1250,In_1533);
or U2669 (N_2669,In_1729,In_782);
or U2670 (N_2670,In_995,In_1940);
nand U2671 (N_2671,In_1130,In_173);
nor U2672 (N_2672,In_339,In_420);
or U2673 (N_2673,In_1753,In_1260);
or U2674 (N_2674,In_922,In_1750);
or U2675 (N_2675,In_1840,In_1658);
and U2676 (N_2676,In_34,In_1689);
or U2677 (N_2677,In_1536,In_1758);
and U2678 (N_2678,In_668,In_1761);
or U2679 (N_2679,In_400,In_1083);
nor U2680 (N_2680,In_652,In_1444);
nor U2681 (N_2681,In_354,In_1215);
nor U2682 (N_2682,In_482,In_1079);
and U2683 (N_2683,In_1876,In_447);
and U2684 (N_2684,In_829,In_1314);
nand U2685 (N_2685,In_1393,In_1885);
nor U2686 (N_2686,In_1895,In_1610);
nand U2687 (N_2687,In_475,In_1877);
nand U2688 (N_2688,In_1828,In_833);
nand U2689 (N_2689,In_456,In_663);
or U2690 (N_2690,In_895,In_1396);
nand U2691 (N_2691,In_271,In_579);
nor U2692 (N_2692,In_1616,In_1171);
or U2693 (N_2693,In_536,In_1897);
and U2694 (N_2694,In_1682,In_429);
and U2695 (N_2695,In_1309,In_671);
nor U2696 (N_2696,In_768,In_1539);
or U2697 (N_2697,In_314,In_437);
or U2698 (N_2698,In_614,In_341);
and U2699 (N_2699,In_44,In_1808);
nor U2700 (N_2700,In_1897,In_1654);
and U2701 (N_2701,In_769,In_416);
nand U2702 (N_2702,In_1199,In_1037);
or U2703 (N_2703,In_1845,In_1414);
and U2704 (N_2704,In_1216,In_1846);
or U2705 (N_2705,In_1410,In_170);
xor U2706 (N_2706,In_1212,In_1346);
and U2707 (N_2707,In_266,In_1470);
and U2708 (N_2708,In_319,In_1063);
and U2709 (N_2709,In_1180,In_1988);
or U2710 (N_2710,In_441,In_1416);
nor U2711 (N_2711,In_1559,In_1906);
nor U2712 (N_2712,In_521,In_1977);
or U2713 (N_2713,In_1466,In_1227);
and U2714 (N_2714,In_728,In_69);
and U2715 (N_2715,In_65,In_1293);
nor U2716 (N_2716,In_1640,In_1354);
nor U2717 (N_2717,In_91,In_216);
and U2718 (N_2718,In_698,In_1642);
nor U2719 (N_2719,In_33,In_48);
nand U2720 (N_2720,In_728,In_1699);
nand U2721 (N_2721,In_1808,In_29);
nor U2722 (N_2722,In_1248,In_988);
nand U2723 (N_2723,In_1265,In_1182);
nor U2724 (N_2724,In_1553,In_645);
nand U2725 (N_2725,In_729,In_1674);
nor U2726 (N_2726,In_1110,In_1906);
xor U2727 (N_2727,In_1351,In_1944);
nand U2728 (N_2728,In_1531,In_813);
and U2729 (N_2729,In_1917,In_621);
nand U2730 (N_2730,In_1216,In_597);
nor U2731 (N_2731,In_1090,In_1685);
and U2732 (N_2732,In_1431,In_1465);
nand U2733 (N_2733,In_423,In_559);
nor U2734 (N_2734,In_92,In_58);
xor U2735 (N_2735,In_1071,In_1102);
nor U2736 (N_2736,In_1573,In_907);
and U2737 (N_2737,In_291,In_1884);
and U2738 (N_2738,In_1550,In_808);
or U2739 (N_2739,In_1461,In_711);
or U2740 (N_2740,In_1017,In_25);
nand U2741 (N_2741,In_959,In_327);
nor U2742 (N_2742,In_1343,In_157);
and U2743 (N_2743,In_104,In_1227);
nor U2744 (N_2744,In_1688,In_957);
nand U2745 (N_2745,In_87,In_1625);
or U2746 (N_2746,In_759,In_104);
and U2747 (N_2747,In_1254,In_1688);
and U2748 (N_2748,In_571,In_1393);
nor U2749 (N_2749,In_819,In_1505);
and U2750 (N_2750,In_278,In_116);
or U2751 (N_2751,In_839,In_1898);
nand U2752 (N_2752,In_1601,In_1312);
nor U2753 (N_2753,In_440,In_629);
nor U2754 (N_2754,In_1192,In_909);
nand U2755 (N_2755,In_593,In_1960);
nand U2756 (N_2756,In_636,In_1959);
and U2757 (N_2757,In_502,In_1844);
or U2758 (N_2758,In_750,In_331);
or U2759 (N_2759,In_707,In_1476);
nor U2760 (N_2760,In_1065,In_495);
and U2761 (N_2761,In_604,In_1794);
and U2762 (N_2762,In_1722,In_1956);
nor U2763 (N_2763,In_1917,In_1446);
nor U2764 (N_2764,In_1488,In_77);
nand U2765 (N_2765,In_1969,In_140);
and U2766 (N_2766,In_1383,In_1040);
nand U2767 (N_2767,In_1998,In_954);
and U2768 (N_2768,In_1870,In_1961);
nand U2769 (N_2769,In_1690,In_1824);
and U2770 (N_2770,In_541,In_1598);
and U2771 (N_2771,In_1672,In_1480);
or U2772 (N_2772,In_651,In_1727);
nor U2773 (N_2773,In_994,In_1774);
and U2774 (N_2774,In_988,In_717);
or U2775 (N_2775,In_1569,In_1243);
nand U2776 (N_2776,In_1156,In_1605);
and U2777 (N_2777,In_1998,In_532);
nor U2778 (N_2778,In_249,In_305);
and U2779 (N_2779,In_288,In_1839);
nor U2780 (N_2780,In_1741,In_879);
and U2781 (N_2781,In_1406,In_184);
and U2782 (N_2782,In_1737,In_285);
or U2783 (N_2783,In_1056,In_1509);
nor U2784 (N_2784,In_1864,In_633);
nor U2785 (N_2785,In_809,In_430);
or U2786 (N_2786,In_805,In_1711);
nand U2787 (N_2787,In_784,In_1092);
nor U2788 (N_2788,In_918,In_987);
nand U2789 (N_2789,In_1061,In_1431);
and U2790 (N_2790,In_1276,In_1327);
and U2791 (N_2791,In_1294,In_714);
and U2792 (N_2792,In_1940,In_1639);
nand U2793 (N_2793,In_915,In_299);
or U2794 (N_2794,In_1,In_1921);
nand U2795 (N_2795,In_525,In_1347);
or U2796 (N_2796,In_1768,In_246);
nor U2797 (N_2797,In_1464,In_895);
or U2798 (N_2798,In_390,In_424);
nor U2799 (N_2799,In_1913,In_188);
or U2800 (N_2800,In_1935,In_1775);
or U2801 (N_2801,In_1386,In_510);
or U2802 (N_2802,In_1671,In_1237);
nand U2803 (N_2803,In_1602,In_1019);
nor U2804 (N_2804,In_211,In_1422);
or U2805 (N_2805,In_1129,In_664);
or U2806 (N_2806,In_44,In_1046);
and U2807 (N_2807,In_1505,In_941);
nor U2808 (N_2808,In_309,In_836);
nor U2809 (N_2809,In_1371,In_1477);
nor U2810 (N_2810,In_356,In_508);
or U2811 (N_2811,In_524,In_891);
or U2812 (N_2812,In_1142,In_1513);
or U2813 (N_2813,In_1100,In_1168);
and U2814 (N_2814,In_1381,In_229);
and U2815 (N_2815,In_137,In_1800);
and U2816 (N_2816,In_1611,In_1880);
and U2817 (N_2817,In_1700,In_94);
nor U2818 (N_2818,In_570,In_1220);
nand U2819 (N_2819,In_857,In_1693);
and U2820 (N_2820,In_1431,In_1280);
and U2821 (N_2821,In_1932,In_1624);
nor U2822 (N_2822,In_1005,In_1876);
nand U2823 (N_2823,In_67,In_38);
and U2824 (N_2824,In_1928,In_1779);
or U2825 (N_2825,In_1654,In_1754);
or U2826 (N_2826,In_1439,In_1750);
nor U2827 (N_2827,In_124,In_277);
nand U2828 (N_2828,In_319,In_809);
and U2829 (N_2829,In_1409,In_707);
or U2830 (N_2830,In_1645,In_569);
or U2831 (N_2831,In_1499,In_1958);
nor U2832 (N_2832,In_1050,In_1449);
nor U2833 (N_2833,In_817,In_1297);
or U2834 (N_2834,In_1172,In_1400);
nand U2835 (N_2835,In_1281,In_123);
or U2836 (N_2836,In_917,In_693);
or U2837 (N_2837,In_1905,In_1940);
or U2838 (N_2838,In_293,In_952);
and U2839 (N_2839,In_648,In_348);
and U2840 (N_2840,In_368,In_1163);
and U2841 (N_2841,In_272,In_24);
and U2842 (N_2842,In_1302,In_852);
nor U2843 (N_2843,In_1940,In_377);
nand U2844 (N_2844,In_467,In_416);
nor U2845 (N_2845,In_495,In_1911);
and U2846 (N_2846,In_1468,In_323);
nand U2847 (N_2847,In_1160,In_104);
nor U2848 (N_2848,In_1872,In_407);
or U2849 (N_2849,In_910,In_940);
xor U2850 (N_2850,In_813,In_1834);
or U2851 (N_2851,In_772,In_1492);
and U2852 (N_2852,In_644,In_1607);
nor U2853 (N_2853,In_1975,In_1806);
nand U2854 (N_2854,In_687,In_340);
nor U2855 (N_2855,In_977,In_1887);
or U2856 (N_2856,In_1055,In_488);
nor U2857 (N_2857,In_1373,In_1454);
nor U2858 (N_2858,In_396,In_1003);
nor U2859 (N_2859,In_1437,In_634);
or U2860 (N_2860,In_230,In_1316);
and U2861 (N_2861,In_46,In_1879);
nor U2862 (N_2862,In_1590,In_64);
nand U2863 (N_2863,In_388,In_1861);
nor U2864 (N_2864,In_370,In_527);
and U2865 (N_2865,In_1569,In_938);
nor U2866 (N_2866,In_1487,In_1165);
or U2867 (N_2867,In_1607,In_1195);
nor U2868 (N_2868,In_1333,In_330);
nor U2869 (N_2869,In_1306,In_93);
nand U2870 (N_2870,In_102,In_903);
nand U2871 (N_2871,In_163,In_1142);
or U2872 (N_2872,In_1891,In_1223);
or U2873 (N_2873,In_1402,In_1043);
or U2874 (N_2874,In_1226,In_897);
nor U2875 (N_2875,In_1754,In_496);
or U2876 (N_2876,In_133,In_882);
nand U2877 (N_2877,In_105,In_642);
and U2878 (N_2878,In_1741,In_656);
nand U2879 (N_2879,In_565,In_525);
or U2880 (N_2880,In_354,In_491);
or U2881 (N_2881,In_844,In_289);
nor U2882 (N_2882,In_1803,In_762);
nand U2883 (N_2883,In_1308,In_259);
nor U2884 (N_2884,In_810,In_1486);
nor U2885 (N_2885,In_176,In_387);
and U2886 (N_2886,In_172,In_523);
and U2887 (N_2887,In_1564,In_1085);
nor U2888 (N_2888,In_881,In_1852);
and U2889 (N_2889,In_1297,In_1566);
nand U2890 (N_2890,In_1635,In_902);
or U2891 (N_2891,In_1623,In_265);
nor U2892 (N_2892,In_1008,In_1006);
nand U2893 (N_2893,In_1656,In_1666);
and U2894 (N_2894,In_1740,In_36);
nor U2895 (N_2895,In_651,In_1753);
nor U2896 (N_2896,In_392,In_1857);
nor U2897 (N_2897,In_1566,In_270);
nand U2898 (N_2898,In_382,In_150);
nor U2899 (N_2899,In_19,In_1507);
nand U2900 (N_2900,In_943,In_1190);
or U2901 (N_2901,In_598,In_140);
nor U2902 (N_2902,In_633,In_1440);
nand U2903 (N_2903,In_1626,In_1821);
or U2904 (N_2904,In_1955,In_1513);
nor U2905 (N_2905,In_496,In_688);
and U2906 (N_2906,In_672,In_9);
or U2907 (N_2907,In_637,In_1052);
nor U2908 (N_2908,In_1465,In_94);
or U2909 (N_2909,In_1383,In_1393);
nor U2910 (N_2910,In_1089,In_424);
nand U2911 (N_2911,In_572,In_5);
and U2912 (N_2912,In_561,In_1866);
or U2913 (N_2913,In_1246,In_1856);
and U2914 (N_2914,In_1359,In_346);
and U2915 (N_2915,In_168,In_995);
and U2916 (N_2916,In_194,In_1255);
nand U2917 (N_2917,In_695,In_1402);
and U2918 (N_2918,In_1782,In_542);
or U2919 (N_2919,In_580,In_890);
nand U2920 (N_2920,In_1193,In_1268);
and U2921 (N_2921,In_737,In_1892);
and U2922 (N_2922,In_643,In_410);
or U2923 (N_2923,In_392,In_1343);
or U2924 (N_2924,In_1456,In_1873);
nand U2925 (N_2925,In_262,In_680);
and U2926 (N_2926,In_1890,In_1851);
and U2927 (N_2927,In_877,In_588);
nor U2928 (N_2928,In_1085,In_830);
and U2929 (N_2929,In_576,In_48);
or U2930 (N_2930,In_847,In_59);
nor U2931 (N_2931,In_1064,In_527);
nor U2932 (N_2932,In_1791,In_254);
and U2933 (N_2933,In_897,In_345);
and U2934 (N_2934,In_283,In_838);
nor U2935 (N_2935,In_696,In_1085);
or U2936 (N_2936,In_331,In_98);
nand U2937 (N_2937,In_915,In_1102);
or U2938 (N_2938,In_749,In_1449);
nor U2939 (N_2939,In_676,In_719);
xnor U2940 (N_2940,In_1965,In_1776);
nor U2941 (N_2941,In_1707,In_1778);
nand U2942 (N_2942,In_1783,In_613);
nand U2943 (N_2943,In_1839,In_27);
nor U2944 (N_2944,In_1967,In_398);
or U2945 (N_2945,In_240,In_356);
nor U2946 (N_2946,In_928,In_675);
and U2947 (N_2947,In_1312,In_336);
and U2948 (N_2948,In_180,In_878);
or U2949 (N_2949,In_1360,In_660);
and U2950 (N_2950,In_134,In_1595);
and U2951 (N_2951,In_856,In_1452);
nor U2952 (N_2952,In_1445,In_678);
and U2953 (N_2953,In_1977,In_994);
nand U2954 (N_2954,In_1617,In_1974);
or U2955 (N_2955,In_1340,In_1539);
and U2956 (N_2956,In_1176,In_769);
nand U2957 (N_2957,In_1129,In_1346);
nand U2958 (N_2958,In_326,In_902);
nand U2959 (N_2959,In_719,In_950);
or U2960 (N_2960,In_959,In_127);
and U2961 (N_2961,In_1030,In_395);
or U2962 (N_2962,In_291,In_1973);
nor U2963 (N_2963,In_1697,In_355);
or U2964 (N_2964,In_35,In_20);
nand U2965 (N_2965,In_1036,In_1266);
or U2966 (N_2966,In_394,In_1866);
nand U2967 (N_2967,In_1163,In_1410);
nand U2968 (N_2968,In_274,In_1859);
and U2969 (N_2969,In_1903,In_655);
nand U2970 (N_2970,In_1988,In_1478);
nor U2971 (N_2971,In_611,In_1493);
nand U2972 (N_2972,In_1069,In_934);
and U2973 (N_2973,In_1963,In_378);
nand U2974 (N_2974,In_1241,In_244);
nand U2975 (N_2975,In_699,In_293);
nor U2976 (N_2976,In_283,In_1407);
and U2977 (N_2977,In_979,In_777);
or U2978 (N_2978,In_941,In_799);
nor U2979 (N_2979,In_151,In_1733);
and U2980 (N_2980,In_683,In_800);
or U2981 (N_2981,In_1090,In_1226);
nor U2982 (N_2982,In_582,In_1482);
and U2983 (N_2983,In_1700,In_472);
and U2984 (N_2984,In_865,In_473);
nor U2985 (N_2985,In_1811,In_1450);
nor U2986 (N_2986,In_1278,In_472);
nand U2987 (N_2987,In_39,In_249);
or U2988 (N_2988,In_1610,In_230);
nor U2989 (N_2989,In_1449,In_1335);
nor U2990 (N_2990,In_938,In_1596);
and U2991 (N_2991,In_644,In_1957);
and U2992 (N_2992,In_1234,In_1436);
nor U2993 (N_2993,In_456,In_5);
or U2994 (N_2994,In_1291,In_605);
or U2995 (N_2995,In_1471,In_593);
nor U2996 (N_2996,In_1352,In_581);
nand U2997 (N_2997,In_729,In_1101);
or U2998 (N_2998,In_1618,In_1617);
nor U2999 (N_2999,In_1082,In_992);
nor U3000 (N_3000,In_1977,In_530);
nand U3001 (N_3001,In_1581,In_1511);
and U3002 (N_3002,In_856,In_1451);
nor U3003 (N_3003,In_1624,In_1900);
nor U3004 (N_3004,In_1042,In_939);
and U3005 (N_3005,In_310,In_650);
and U3006 (N_3006,In_402,In_1935);
or U3007 (N_3007,In_205,In_9);
nand U3008 (N_3008,In_105,In_208);
nand U3009 (N_3009,In_12,In_879);
or U3010 (N_3010,In_1838,In_1786);
nand U3011 (N_3011,In_1937,In_7);
or U3012 (N_3012,In_1448,In_970);
nand U3013 (N_3013,In_42,In_1163);
nand U3014 (N_3014,In_17,In_655);
nand U3015 (N_3015,In_176,In_651);
nor U3016 (N_3016,In_736,In_212);
nor U3017 (N_3017,In_1668,In_898);
and U3018 (N_3018,In_1130,In_403);
nand U3019 (N_3019,In_729,In_1780);
nand U3020 (N_3020,In_872,In_611);
and U3021 (N_3021,In_666,In_1065);
nand U3022 (N_3022,In_1337,In_931);
nor U3023 (N_3023,In_529,In_177);
nor U3024 (N_3024,In_791,In_784);
nor U3025 (N_3025,In_1427,In_885);
and U3026 (N_3026,In_136,In_466);
nand U3027 (N_3027,In_174,In_1996);
nand U3028 (N_3028,In_496,In_1563);
and U3029 (N_3029,In_201,In_27);
or U3030 (N_3030,In_1801,In_1237);
or U3031 (N_3031,In_1676,In_268);
nor U3032 (N_3032,In_1664,In_674);
nand U3033 (N_3033,In_251,In_440);
and U3034 (N_3034,In_47,In_440);
nor U3035 (N_3035,In_279,In_526);
or U3036 (N_3036,In_1354,In_929);
and U3037 (N_3037,In_4,In_593);
nand U3038 (N_3038,In_76,In_1506);
or U3039 (N_3039,In_160,In_1820);
and U3040 (N_3040,In_289,In_1663);
or U3041 (N_3041,In_671,In_468);
nor U3042 (N_3042,In_659,In_1092);
and U3043 (N_3043,In_959,In_20);
or U3044 (N_3044,In_1175,In_1211);
or U3045 (N_3045,In_976,In_1068);
or U3046 (N_3046,In_1216,In_619);
and U3047 (N_3047,In_1105,In_434);
and U3048 (N_3048,In_215,In_786);
nand U3049 (N_3049,In_1038,In_1785);
and U3050 (N_3050,In_1273,In_1605);
and U3051 (N_3051,In_69,In_26);
or U3052 (N_3052,In_883,In_1637);
or U3053 (N_3053,In_242,In_1393);
or U3054 (N_3054,In_943,In_861);
and U3055 (N_3055,In_1465,In_1487);
nor U3056 (N_3056,In_63,In_1822);
or U3057 (N_3057,In_1686,In_1241);
or U3058 (N_3058,In_1763,In_850);
or U3059 (N_3059,In_497,In_1240);
or U3060 (N_3060,In_1548,In_1462);
and U3061 (N_3061,In_1839,In_1730);
or U3062 (N_3062,In_1672,In_1839);
nor U3063 (N_3063,In_1929,In_1512);
or U3064 (N_3064,In_959,In_113);
nand U3065 (N_3065,In_1045,In_1333);
nor U3066 (N_3066,In_984,In_514);
nor U3067 (N_3067,In_623,In_457);
and U3068 (N_3068,In_1890,In_1886);
and U3069 (N_3069,In_592,In_83);
and U3070 (N_3070,In_621,In_1234);
nand U3071 (N_3071,In_1209,In_1629);
or U3072 (N_3072,In_1330,In_540);
nor U3073 (N_3073,In_952,In_1778);
nor U3074 (N_3074,In_84,In_1108);
and U3075 (N_3075,In_758,In_1537);
and U3076 (N_3076,In_1222,In_1719);
nor U3077 (N_3077,In_1624,In_1065);
or U3078 (N_3078,In_973,In_528);
nor U3079 (N_3079,In_405,In_1014);
nand U3080 (N_3080,In_1754,In_1566);
nand U3081 (N_3081,In_161,In_1258);
xor U3082 (N_3082,In_23,In_1841);
and U3083 (N_3083,In_202,In_1133);
xor U3084 (N_3084,In_426,In_540);
or U3085 (N_3085,In_1145,In_999);
or U3086 (N_3086,In_436,In_1484);
and U3087 (N_3087,In_1427,In_1080);
or U3088 (N_3088,In_793,In_527);
or U3089 (N_3089,In_1799,In_1168);
and U3090 (N_3090,In_136,In_1537);
or U3091 (N_3091,In_569,In_1334);
nor U3092 (N_3092,In_411,In_438);
nand U3093 (N_3093,In_565,In_1260);
nor U3094 (N_3094,In_672,In_712);
and U3095 (N_3095,In_1974,In_1123);
nor U3096 (N_3096,In_1878,In_1296);
or U3097 (N_3097,In_37,In_1398);
nor U3098 (N_3098,In_652,In_1933);
nand U3099 (N_3099,In_1115,In_218);
and U3100 (N_3100,In_1905,In_1130);
nand U3101 (N_3101,In_1708,In_87);
nand U3102 (N_3102,In_587,In_897);
nor U3103 (N_3103,In_626,In_279);
nand U3104 (N_3104,In_921,In_1794);
or U3105 (N_3105,In_1851,In_728);
nand U3106 (N_3106,In_31,In_1810);
nand U3107 (N_3107,In_961,In_1415);
nand U3108 (N_3108,In_914,In_403);
or U3109 (N_3109,In_890,In_619);
and U3110 (N_3110,In_1490,In_387);
or U3111 (N_3111,In_1591,In_540);
and U3112 (N_3112,In_24,In_889);
nand U3113 (N_3113,In_1664,In_1076);
nor U3114 (N_3114,In_370,In_1742);
or U3115 (N_3115,In_1886,In_1576);
nor U3116 (N_3116,In_1483,In_1199);
and U3117 (N_3117,In_32,In_394);
and U3118 (N_3118,In_1616,In_876);
nand U3119 (N_3119,In_962,In_55);
xor U3120 (N_3120,In_782,In_1614);
nor U3121 (N_3121,In_1232,In_197);
nor U3122 (N_3122,In_363,In_1380);
and U3123 (N_3123,In_1954,In_948);
nand U3124 (N_3124,In_546,In_1524);
nor U3125 (N_3125,In_1378,In_1940);
nand U3126 (N_3126,In_266,In_653);
or U3127 (N_3127,In_1028,In_1297);
and U3128 (N_3128,In_210,In_382);
and U3129 (N_3129,In_1724,In_1409);
and U3130 (N_3130,In_1741,In_1843);
and U3131 (N_3131,In_1823,In_543);
and U3132 (N_3132,In_107,In_768);
and U3133 (N_3133,In_1615,In_78);
and U3134 (N_3134,In_1120,In_1758);
and U3135 (N_3135,In_966,In_1711);
and U3136 (N_3136,In_1372,In_1669);
nor U3137 (N_3137,In_674,In_1743);
nor U3138 (N_3138,In_124,In_1002);
or U3139 (N_3139,In_1032,In_773);
nand U3140 (N_3140,In_1738,In_460);
nor U3141 (N_3141,In_164,In_431);
or U3142 (N_3142,In_814,In_518);
nor U3143 (N_3143,In_1585,In_1475);
or U3144 (N_3144,In_858,In_139);
xnor U3145 (N_3145,In_1663,In_1271);
nand U3146 (N_3146,In_784,In_507);
nand U3147 (N_3147,In_772,In_796);
nor U3148 (N_3148,In_441,In_295);
and U3149 (N_3149,In_1554,In_844);
and U3150 (N_3150,In_668,In_706);
and U3151 (N_3151,In_208,In_964);
nor U3152 (N_3152,In_735,In_1551);
and U3153 (N_3153,In_414,In_1506);
nand U3154 (N_3154,In_598,In_1524);
nor U3155 (N_3155,In_1354,In_0);
and U3156 (N_3156,In_238,In_1299);
nor U3157 (N_3157,In_1089,In_886);
nor U3158 (N_3158,In_291,In_729);
and U3159 (N_3159,In_1951,In_504);
and U3160 (N_3160,In_410,In_715);
or U3161 (N_3161,In_863,In_844);
and U3162 (N_3162,In_1796,In_142);
or U3163 (N_3163,In_1450,In_485);
nand U3164 (N_3164,In_1615,In_1456);
nor U3165 (N_3165,In_315,In_1453);
and U3166 (N_3166,In_331,In_1673);
or U3167 (N_3167,In_257,In_1329);
and U3168 (N_3168,In_1228,In_615);
nor U3169 (N_3169,In_1762,In_863);
nor U3170 (N_3170,In_1068,In_1495);
nor U3171 (N_3171,In_613,In_41);
or U3172 (N_3172,In_1951,In_1227);
nand U3173 (N_3173,In_1041,In_592);
or U3174 (N_3174,In_1353,In_983);
and U3175 (N_3175,In_1288,In_447);
nand U3176 (N_3176,In_1846,In_236);
nor U3177 (N_3177,In_948,In_1122);
and U3178 (N_3178,In_1498,In_1132);
and U3179 (N_3179,In_1488,In_635);
and U3180 (N_3180,In_102,In_540);
and U3181 (N_3181,In_681,In_1958);
nor U3182 (N_3182,In_704,In_1348);
or U3183 (N_3183,In_983,In_1266);
nand U3184 (N_3184,In_305,In_1226);
nor U3185 (N_3185,In_203,In_501);
and U3186 (N_3186,In_458,In_1192);
or U3187 (N_3187,In_1129,In_92);
or U3188 (N_3188,In_252,In_766);
or U3189 (N_3189,In_1104,In_303);
and U3190 (N_3190,In_873,In_1845);
nand U3191 (N_3191,In_984,In_1163);
and U3192 (N_3192,In_47,In_1141);
nor U3193 (N_3193,In_530,In_1790);
nor U3194 (N_3194,In_902,In_1801);
nand U3195 (N_3195,In_235,In_1719);
nor U3196 (N_3196,In_1425,In_1352);
xor U3197 (N_3197,In_1620,In_1652);
nand U3198 (N_3198,In_432,In_282);
nand U3199 (N_3199,In_1644,In_1909);
and U3200 (N_3200,In_1073,In_1908);
and U3201 (N_3201,In_376,In_1073);
nor U3202 (N_3202,In_1045,In_1461);
or U3203 (N_3203,In_1181,In_1997);
or U3204 (N_3204,In_870,In_1416);
nand U3205 (N_3205,In_1185,In_1105);
nor U3206 (N_3206,In_1101,In_141);
nand U3207 (N_3207,In_927,In_841);
and U3208 (N_3208,In_200,In_935);
xnor U3209 (N_3209,In_821,In_1021);
and U3210 (N_3210,In_712,In_308);
and U3211 (N_3211,In_1673,In_134);
nand U3212 (N_3212,In_1328,In_1451);
and U3213 (N_3213,In_1647,In_1535);
nand U3214 (N_3214,In_1721,In_557);
and U3215 (N_3215,In_473,In_1344);
or U3216 (N_3216,In_532,In_1667);
nor U3217 (N_3217,In_1733,In_872);
and U3218 (N_3218,In_27,In_726);
nor U3219 (N_3219,In_1590,In_1298);
or U3220 (N_3220,In_703,In_1873);
or U3221 (N_3221,In_932,In_802);
nand U3222 (N_3222,In_640,In_239);
or U3223 (N_3223,In_1358,In_1245);
or U3224 (N_3224,In_1568,In_1398);
nor U3225 (N_3225,In_558,In_1937);
nand U3226 (N_3226,In_1350,In_375);
and U3227 (N_3227,In_939,In_503);
or U3228 (N_3228,In_58,In_899);
or U3229 (N_3229,In_1144,In_1789);
nor U3230 (N_3230,In_1866,In_303);
or U3231 (N_3231,In_290,In_697);
or U3232 (N_3232,In_1780,In_1711);
or U3233 (N_3233,In_1243,In_1497);
and U3234 (N_3234,In_1417,In_817);
nand U3235 (N_3235,In_714,In_1257);
nor U3236 (N_3236,In_510,In_1881);
nor U3237 (N_3237,In_1985,In_1890);
and U3238 (N_3238,In_742,In_392);
nand U3239 (N_3239,In_1591,In_1589);
and U3240 (N_3240,In_187,In_1144);
or U3241 (N_3241,In_394,In_408);
and U3242 (N_3242,In_853,In_773);
xor U3243 (N_3243,In_530,In_987);
or U3244 (N_3244,In_1524,In_904);
nand U3245 (N_3245,In_50,In_198);
nor U3246 (N_3246,In_342,In_465);
nor U3247 (N_3247,In_388,In_504);
nand U3248 (N_3248,In_1873,In_1123);
nor U3249 (N_3249,In_461,In_1526);
nand U3250 (N_3250,In_413,In_539);
or U3251 (N_3251,In_1661,In_603);
nand U3252 (N_3252,In_996,In_586);
nand U3253 (N_3253,In_1252,In_384);
nand U3254 (N_3254,In_729,In_1222);
nand U3255 (N_3255,In_1938,In_107);
nor U3256 (N_3256,In_1192,In_989);
and U3257 (N_3257,In_1880,In_590);
or U3258 (N_3258,In_1495,In_645);
nor U3259 (N_3259,In_1955,In_136);
nand U3260 (N_3260,In_211,In_26);
and U3261 (N_3261,In_1788,In_647);
nor U3262 (N_3262,In_1331,In_1896);
and U3263 (N_3263,In_1011,In_342);
nand U3264 (N_3264,In_1233,In_662);
nand U3265 (N_3265,In_1077,In_212);
and U3266 (N_3266,In_1904,In_1951);
or U3267 (N_3267,In_165,In_948);
nand U3268 (N_3268,In_694,In_1846);
nand U3269 (N_3269,In_1120,In_974);
or U3270 (N_3270,In_322,In_520);
nor U3271 (N_3271,In_685,In_1846);
and U3272 (N_3272,In_700,In_1140);
or U3273 (N_3273,In_1118,In_1805);
or U3274 (N_3274,In_1269,In_1474);
nand U3275 (N_3275,In_251,In_616);
or U3276 (N_3276,In_282,In_644);
nor U3277 (N_3277,In_1284,In_135);
nand U3278 (N_3278,In_453,In_1022);
and U3279 (N_3279,In_1075,In_1116);
nand U3280 (N_3280,In_942,In_671);
and U3281 (N_3281,In_392,In_1324);
or U3282 (N_3282,In_723,In_1357);
or U3283 (N_3283,In_107,In_816);
or U3284 (N_3284,In_165,In_1276);
nand U3285 (N_3285,In_1231,In_1499);
and U3286 (N_3286,In_445,In_1602);
nor U3287 (N_3287,In_1070,In_1073);
or U3288 (N_3288,In_1675,In_585);
nand U3289 (N_3289,In_1223,In_383);
nor U3290 (N_3290,In_1569,In_159);
nor U3291 (N_3291,In_94,In_1375);
xnor U3292 (N_3292,In_167,In_679);
or U3293 (N_3293,In_1251,In_1086);
nand U3294 (N_3294,In_711,In_1410);
xor U3295 (N_3295,In_218,In_921);
or U3296 (N_3296,In_208,In_596);
or U3297 (N_3297,In_1248,In_1790);
nand U3298 (N_3298,In_489,In_1890);
and U3299 (N_3299,In_1592,In_379);
xor U3300 (N_3300,In_1323,In_576);
nor U3301 (N_3301,In_550,In_719);
nor U3302 (N_3302,In_1861,In_1246);
or U3303 (N_3303,In_1792,In_1162);
nor U3304 (N_3304,In_1790,In_484);
or U3305 (N_3305,In_1232,In_1683);
nand U3306 (N_3306,In_504,In_1578);
nor U3307 (N_3307,In_436,In_1552);
nand U3308 (N_3308,In_1710,In_1685);
nor U3309 (N_3309,In_760,In_1731);
nand U3310 (N_3310,In_1456,In_372);
nor U3311 (N_3311,In_683,In_977);
nand U3312 (N_3312,In_353,In_571);
or U3313 (N_3313,In_39,In_1255);
or U3314 (N_3314,In_1080,In_685);
nand U3315 (N_3315,In_1822,In_183);
or U3316 (N_3316,In_217,In_1059);
nand U3317 (N_3317,In_475,In_176);
and U3318 (N_3318,In_1640,In_117);
nor U3319 (N_3319,In_991,In_1495);
or U3320 (N_3320,In_42,In_1121);
nand U3321 (N_3321,In_63,In_1294);
or U3322 (N_3322,In_285,In_1897);
and U3323 (N_3323,In_1959,In_1299);
or U3324 (N_3324,In_783,In_850);
nand U3325 (N_3325,In_584,In_908);
and U3326 (N_3326,In_1816,In_999);
nor U3327 (N_3327,In_66,In_1610);
nor U3328 (N_3328,In_1998,In_1726);
nand U3329 (N_3329,In_952,In_861);
nor U3330 (N_3330,In_1204,In_596);
nand U3331 (N_3331,In_799,In_619);
nand U3332 (N_3332,In_1804,In_678);
or U3333 (N_3333,In_1563,In_1308);
nor U3334 (N_3334,In_1116,In_85);
nor U3335 (N_3335,In_1289,In_8);
nand U3336 (N_3336,In_1876,In_548);
and U3337 (N_3337,In_1982,In_1626);
and U3338 (N_3338,In_3,In_1380);
or U3339 (N_3339,In_203,In_1799);
nor U3340 (N_3340,In_1967,In_683);
or U3341 (N_3341,In_857,In_520);
and U3342 (N_3342,In_1420,In_736);
and U3343 (N_3343,In_1106,In_1905);
and U3344 (N_3344,In_380,In_593);
nor U3345 (N_3345,In_372,In_1138);
nand U3346 (N_3346,In_347,In_415);
or U3347 (N_3347,In_655,In_663);
and U3348 (N_3348,In_1196,In_1815);
nor U3349 (N_3349,In_418,In_1945);
nand U3350 (N_3350,In_834,In_1483);
nand U3351 (N_3351,In_1479,In_1297);
or U3352 (N_3352,In_1176,In_4);
and U3353 (N_3353,In_1256,In_862);
and U3354 (N_3354,In_660,In_748);
nor U3355 (N_3355,In_924,In_23);
nand U3356 (N_3356,In_699,In_1346);
nand U3357 (N_3357,In_1233,In_1223);
nand U3358 (N_3358,In_1673,In_78);
nand U3359 (N_3359,In_990,In_1577);
nor U3360 (N_3360,In_1511,In_1996);
and U3361 (N_3361,In_1927,In_1173);
or U3362 (N_3362,In_1318,In_260);
nand U3363 (N_3363,In_728,In_978);
nand U3364 (N_3364,In_1525,In_692);
or U3365 (N_3365,In_610,In_900);
or U3366 (N_3366,In_1724,In_543);
and U3367 (N_3367,In_1211,In_733);
or U3368 (N_3368,In_515,In_1692);
nor U3369 (N_3369,In_563,In_731);
nand U3370 (N_3370,In_1093,In_1843);
and U3371 (N_3371,In_667,In_941);
nor U3372 (N_3372,In_949,In_89);
nor U3373 (N_3373,In_1862,In_1725);
nor U3374 (N_3374,In_1139,In_1927);
and U3375 (N_3375,In_649,In_490);
or U3376 (N_3376,In_743,In_1234);
nor U3377 (N_3377,In_1994,In_1098);
or U3378 (N_3378,In_135,In_1161);
nand U3379 (N_3379,In_1322,In_1771);
nand U3380 (N_3380,In_776,In_1525);
or U3381 (N_3381,In_1531,In_1698);
nand U3382 (N_3382,In_159,In_787);
nand U3383 (N_3383,In_1428,In_81);
nand U3384 (N_3384,In_1357,In_1985);
nand U3385 (N_3385,In_1215,In_1700);
or U3386 (N_3386,In_448,In_1967);
or U3387 (N_3387,In_154,In_1313);
or U3388 (N_3388,In_1413,In_995);
nor U3389 (N_3389,In_1202,In_652);
nor U3390 (N_3390,In_1989,In_1847);
nand U3391 (N_3391,In_725,In_1929);
or U3392 (N_3392,In_479,In_409);
or U3393 (N_3393,In_1746,In_796);
and U3394 (N_3394,In_278,In_1144);
nand U3395 (N_3395,In_1930,In_1300);
or U3396 (N_3396,In_891,In_1211);
or U3397 (N_3397,In_936,In_1566);
nor U3398 (N_3398,In_1014,In_1533);
nand U3399 (N_3399,In_1484,In_16);
nor U3400 (N_3400,In_1104,In_1992);
and U3401 (N_3401,In_1215,In_1805);
nand U3402 (N_3402,In_956,In_1264);
or U3403 (N_3403,In_1095,In_1163);
and U3404 (N_3404,In_640,In_823);
xnor U3405 (N_3405,In_598,In_429);
xnor U3406 (N_3406,In_1339,In_293);
nand U3407 (N_3407,In_1573,In_1937);
or U3408 (N_3408,In_968,In_106);
or U3409 (N_3409,In_470,In_1717);
and U3410 (N_3410,In_1438,In_330);
or U3411 (N_3411,In_335,In_728);
and U3412 (N_3412,In_112,In_1356);
or U3413 (N_3413,In_935,In_604);
and U3414 (N_3414,In_1068,In_1607);
and U3415 (N_3415,In_1290,In_1565);
or U3416 (N_3416,In_1378,In_1077);
nor U3417 (N_3417,In_1178,In_1376);
or U3418 (N_3418,In_462,In_1076);
and U3419 (N_3419,In_1219,In_209);
nor U3420 (N_3420,In_1549,In_1862);
and U3421 (N_3421,In_852,In_1240);
nor U3422 (N_3422,In_122,In_356);
or U3423 (N_3423,In_1455,In_230);
or U3424 (N_3424,In_1772,In_1246);
nand U3425 (N_3425,In_1008,In_1943);
and U3426 (N_3426,In_154,In_812);
and U3427 (N_3427,In_1106,In_210);
nor U3428 (N_3428,In_1693,In_598);
nor U3429 (N_3429,In_227,In_150);
or U3430 (N_3430,In_1032,In_596);
nand U3431 (N_3431,In_818,In_596);
nand U3432 (N_3432,In_1910,In_1598);
or U3433 (N_3433,In_1520,In_1935);
nor U3434 (N_3434,In_189,In_1702);
and U3435 (N_3435,In_505,In_1985);
nor U3436 (N_3436,In_454,In_115);
or U3437 (N_3437,In_349,In_679);
nand U3438 (N_3438,In_1872,In_422);
nand U3439 (N_3439,In_1495,In_969);
nor U3440 (N_3440,In_207,In_1637);
or U3441 (N_3441,In_1018,In_1087);
and U3442 (N_3442,In_1544,In_1903);
nor U3443 (N_3443,In_1354,In_745);
or U3444 (N_3444,In_439,In_713);
nand U3445 (N_3445,In_639,In_169);
nand U3446 (N_3446,In_64,In_373);
nor U3447 (N_3447,In_1953,In_1862);
nor U3448 (N_3448,In_1554,In_909);
and U3449 (N_3449,In_185,In_847);
nor U3450 (N_3450,In_1785,In_141);
and U3451 (N_3451,In_31,In_434);
and U3452 (N_3452,In_374,In_979);
or U3453 (N_3453,In_896,In_212);
or U3454 (N_3454,In_898,In_514);
and U3455 (N_3455,In_1301,In_1246);
and U3456 (N_3456,In_1752,In_515);
nor U3457 (N_3457,In_575,In_56);
or U3458 (N_3458,In_1116,In_779);
and U3459 (N_3459,In_710,In_404);
nor U3460 (N_3460,In_1210,In_105);
and U3461 (N_3461,In_1474,In_1169);
nand U3462 (N_3462,In_1006,In_1799);
or U3463 (N_3463,In_1230,In_1502);
or U3464 (N_3464,In_1930,In_1475);
nor U3465 (N_3465,In_1232,In_599);
nor U3466 (N_3466,In_1071,In_371);
nand U3467 (N_3467,In_1917,In_1742);
nor U3468 (N_3468,In_296,In_644);
or U3469 (N_3469,In_1476,In_299);
and U3470 (N_3470,In_132,In_303);
or U3471 (N_3471,In_1412,In_1294);
nor U3472 (N_3472,In_1058,In_1542);
nor U3473 (N_3473,In_304,In_1710);
nor U3474 (N_3474,In_1085,In_4);
nand U3475 (N_3475,In_1227,In_1647);
nand U3476 (N_3476,In_971,In_1121);
nand U3477 (N_3477,In_697,In_491);
nand U3478 (N_3478,In_426,In_1933);
nor U3479 (N_3479,In_1554,In_1292);
and U3480 (N_3480,In_1326,In_1722);
and U3481 (N_3481,In_1040,In_609);
nor U3482 (N_3482,In_1490,In_7);
or U3483 (N_3483,In_1208,In_866);
or U3484 (N_3484,In_689,In_1214);
and U3485 (N_3485,In_589,In_267);
nand U3486 (N_3486,In_1650,In_1116);
and U3487 (N_3487,In_856,In_963);
nor U3488 (N_3488,In_1205,In_162);
or U3489 (N_3489,In_1416,In_328);
nor U3490 (N_3490,In_1482,In_903);
nor U3491 (N_3491,In_443,In_1157);
or U3492 (N_3492,In_1516,In_1006);
nor U3493 (N_3493,In_1785,In_1835);
or U3494 (N_3494,In_1685,In_1812);
nor U3495 (N_3495,In_379,In_134);
nor U3496 (N_3496,In_821,In_798);
or U3497 (N_3497,In_1284,In_1852);
nor U3498 (N_3498,In_1098,In_799);
nor U3499 (N_3499,In_387,In_1688);
nand U3500 (N_3500,In_677,In_591);
or U3501 (N_3501,In_182,In_1723);
or U3502 (N_3502,In_988,In_1665);
and U3503 (N_3503,In_473,In_919);
nand U3504 (N_3504,In_179,In_1126);
and U3505 (N_3505,In_648,In_904);
nor U3506 (N_3506,In_727,In_1194);
or U3507 (N_3507,In_1017,In_1437);
and U3508 (N_3508,In_1563,In_1739);
or U3509 (N_3509,In_923,In_1283);
nor U3510 (N_3510,In_1128,In_1912);
nor U3511 (N_3511,In_1569,In_1322);
nand U3512 (N_3512,In_336,In_1992);
and U3513 (N_3513,In_1401,In_1321);
nand U3514 (N_3514,In_1377,In_924);
nand U3515 (N_3515,In_1512,In_1565);
or U3516 (N_3516,In_1849,In_88);
and U3517 (N_3517,In_870,In_118);
and U3518 (N_3518,In_598,In_1694);
or U3519 (N_3519,In_1419,In_1598);
nor U3520 (N_3520,In_1899,In_170);
nand U3521 (N_3521,In_1129,In_205);
or U3522 (N_3522,In_1402,In_1027);
or U3523 (N_3523,In_914,In_306);
nor U3524 (N_3524,In_1317,In_94);
and U3525 (N_3525,In_729,In_1614);
nand U3526 (N_3526,In_1181,In_1058);
nor U3527 (N_3527,In_78,In_417);
and U3528 (N_3528,In_685,In_642);
nor U3529 (N_3529,In_596,In_173);
nor U3530 (N_3530,In_1786,In_509);
and U3531 (N_3531,In_1006,In_784);
and U3532 (N_3532,In_1583,In_598);
and U3533 (N_3533,In_847,In_270);
nor U3534 (N_3534,In_1731,In_246);
nand U3535 (N_3535,In_452,In_112);
nor U3536 (N_3536,In_1563,In_310);
and U3537 (N_3537,In_1036,In_658);
nand U3538 (N_3538,In_1317,In_387);
or U3539 (N_3539,In_1333,In_1796);
nor U3540 (N_3540,In_1268,In_1297);
or U3541 (N_3541,In_1402,In_1549);
and U3542 (N_3542,In_108,In_1030);
or U3543 (N_3543,In_837,In_1447);
nand U3544 (N_3544,In_1103,In_1095);
and U3545 (N_3545,In_1622,In_1403);
nor U3546 (N_3546,In_1743,In_444);
or U3547 (N_3547,In_138,In_272);
nand U3548 (N_3548,In_780,In_750);
nor U3549 (N_3549,In_1682,In_463);
and U3550 (N_3550,In_1589,In_1502);
nand U3551 (N_3551,In_1920,In_1847);
nand U3552 (N_3552,In_1271,In_98);
and U3553 (N_3553,In_323,In_75);
or U3554 (N_3554,In_63,In_307);
and U3555 (N_3555,In_1174,In_63);
or U3556 (N_3556,In_1048,In_1293);
nand U3557 (N_3557,In_637,In_673);
or U3558 (N_3558,In_184,In_40);
xnor U3559 (N_3559,In_1199,In_10);
nor U3560 (N_3560,In_214,In_1234);
and U3561 (N_3561,In_1860,In_1588);
xnor U3562 (N_3562,In_1338,In_209);
and U3563 (N_3563,In_1074,In_153);
or U3564 (N_3564,In_443,In_902);
nand U3565 (N_3565,In_953,In_1890);
nor U3566 (N_3566,In_666,In_1727);
nand U3567 (N_3567,In_1721,In_1943);
and U3568 (N_3568,In_1064,In_909);
or U3569 (N_3569,In_652,In_1317);
nor U3570 (N_3570,In_1728,In_300);
nand U3571 (N_3571,In_1250,In_1276);
nand U3572 (N_3572,In_1583,In_636);
nor U3573 (N_3573,In_709,In_446);
nor U3574 (N_3574,In_380,In_441);
and U3575 (N_3575,In_958,In_436);
nor U3576 (N_3576,In_849,In_263);
and U3577 (N_3577,In_1291,In_121);
and U3578 (N_3578,In_949,In_1279);
or U3579 (N_3579,In_342,In_380);
and U3580 (N_3580,In_435,In_359);
nand U3581 (N_3581,In_1173,In_1289);
nand U3582 (N_3582,In_1792,In_928);
or U3583 (N_3583,In_1407,In_1329);
nor U3584 (N_3584,In_665,In_77);
and U3585 (N_3585,In_665,In_934);
nor U3586 (N_3586,In_1837,In_1949);
nand U3587 (N_3587,In_1969,In_1308);
or U3588 (N_3588,In_1696,In_1282);
nor U3589 (N_3589,In_1092,In_1397);
or U3590 (N_3590,In_446,In_678);
nand U3591 (N_3591,In_219,In_1102);
nand U3592 (N_3592,In_715,In_182);
and U3593 (N_3593,In_1039,In_301);
or U3594 (N_3594,In_720,In_1015);
or U3595 (N_3595,In_1089,In_97);
or U3596 (N_3596,In_1425,In_1062);
or U3597 (N_3597,In_655,In_1404);
and U3598 (N_3598,In_1139,In_1001);
nand U3599 (N_3599,In_1579,In_1620);
nand U3600 (N_3600,In_1223,In_1515);
or U3601 (N_3601,In_479,In_112);
or U3602 (N_3602,In_1440,In_1287);
nand U3603 (N_3603,In_70,In_1746);
and U3604 (N_3604,In_1272,In_1539);
nor U3605 (N_3605,In_871,In_1575);
or U3606 (N_3606,In_1684,In_973);
nand U3607 (N_3607,In_1286,In_729);
nand U3608 (N_3608,In_1978,In_18);
nor U3609 (N_3609,In_778,In_831);
nand U3610 (N_3610,In_1505,In_530);
or U3611 (N_3611,In_558,In_1953);
nand U3612 (N_3612,In_500,In_1017);
or U3613 (N_3613,In_1722,In_1500);
or U3614 (N_3614,In_1092,In_126);
nor U3615 (N_3615,In_913,In_1342);
nand U3616 (N_3616,In_881,In_1290);
nand U3617 (N_3617,In_897,In_415);
and U3618 (N_3618,In_748,In_105);
or U3619 (N_3619,In_790,In_223);
nand U3620 (N_3620,In_574,In_1624);
xnor U3621 (N_3621,In_290,In_212);
nor U3622 (N_3622,In_260,In_601);
nand U3623 (N_3623,In_1701,In_1486);
nand U3624 (N_3624,In_549,In_1547);
or U3625 (N_3625,In_1908,In_1328);
and U3626 (N_3626,In_728,In_1162);
nor U3627 (N_3627,In_1421,In_1533);
or U3628 (N_3628,In_506,In_1640);
or U3629 (N_3629,In_1552,In_913);
or U3630 (N_3630,In_833,In_1422);
and U3631 (N_3631,In_376,In_481);
and U3632 (N_3632,In_447,In_510);
or U3633 (N_3633,In_1493,In_1080);
nand U3634 (N_3634,In_1868,In_606);
nand U3635 (N_3635,In_886,In_1469);
nand U3636 (N_3636,In_1351,In_431);
nand U3637 (N_3637,In_21,In_685);
and U3638 (N_3638,In_928,In_1154);
nand U3639 (N_3639,In_319,In_1398);
and U3640 (N_3640,In_491,In_1912);
and U3641 (N_3641,In_930,In_1792);
and U3642 (N_3642,In_680,In_1171);
xor U3643 (N_3643,In_1736,In_1610);
and U3644 (N_3644,In_213,In_807);
or U3645 (N_3645,In_1163,In_1409);
nand U3646 (N_3646,In_499,In_1780);
nor U3647 (N_3647,In_1965,In_1716);
nand U3648 (N_3648,In_1872,In_1286);
nand U3649 (N_3649,In_1662,In_839);
or U3650 (N_3650,In_1646,In_1776);
and U3651 (N_3651,In_1119,In_231);
and U3652 (N_3652,In_161,In_1482);
or U3653 (N_3653,In_394,In_1900);
and U3654 (N_3654,In_1278,In_1442);
xnor U3655 (N_3655,In_968,In_153);
nand U3656 (N_3656,In_1296,In_1969);
and U3657 (N_3657,In_114,In_1913);
nor U3658 (N_3658,In_379,In_1789);
xnor U3659 (N_3659,In_1947,In_278);
nand U3660 (N_3660,In_1189,In_1174);
nor U3661 (N_3661,In_995,In_1377);
and U3662 (N_3662,In_1364,In_285);
nand U3663 (N_3663,In_64,In_1592);
or U3664 (N_3664,In_252,In_1916);
nor U3665 (N_3665,In_872,In_1325);
nand U3666 (N_3666,In_1512,In_1940);
and U3667 (N_3667,In_845,In_958);
and U3668 (N_3668,In_1358,In_1027);
xnor U3669 (N_3669,In_1221,In_1714);
nor U3670 (N_3670,In_1753,In_1100);
nand U3671 (N_3671,In_1377,In_1112);
nor U3672 (N_3672,In_729,In_115);
or U3673 (N_3673,In_1547,In_1738);
nor U3674 (N_3674,In_301,In_163);
nor U3675 (N_3675,In_527,In_328);
or U3676 (N_3676,In_1014,In_482);
and U3677 (N_3677,In_41,In_1357);
or U3678 (N_3678,In_1880,In_705);
and U3679 (N_3679,In_1478,In_448);
nand U3680 (N_3680,In_616,In_958);
or U3681 (N_3681,In_1101,In_1355);
nand U3682 (N_3682,In_1367,In_98);
or U3683 (N_3683,In_1912,In_395);
nand U3684 (N_3684,In_187,In_746);
and U3685 (N_3685,In_289,In_263);
and U3686 (N_3686,In_1307,In_532);
nand U3687 (N_3687,In_717,In_1670);
nand U3688 (N_3688,In_1621,In_595);
nand U3689 (N_3689,In_1798,In_122);
nand U3690 (N_3690,In_937,In_77);
nand U3691 (N_3691,In_742,In_668);
or U3692 (N_3692,In_1176,In_1288);
and U3693 (N_3693,In_1839,In_1036);
nor U3694 (N_3694,In_1663,In_1471);
and U3695 (N_3695,In_745,In_1513);
nor U3696 (N_3696,In_1585,In_1971);
nor U3697 (N_3697,In_1116,In_1958);
and U3698 (N_3698,In_728,In_1686);
nor U3699 (N_3699,In_659,In_1168);
or U3700 (N_3700,In_824,In_1596);
and U3701 (N_3701,In_614,In_1475);
and U3702 (N_3702,In_473,In_142);
nor U3703 (N_3703,In_179,In_876);
nor U3704 (N_3704,In_1812,In_1988);
or U3705 (N_3705,In_826,In_1845);
nand U3706 (N_3706,In_1643,In_654);
and U3707 (N_3707,In_205,In_995);
nand U3708 (N_3708,In_462,In_1391);
nor U3709 (N_3709,In_429,In_1233);
nand U3710 (N_3710,In_1734,In_876);
nor U3711 (N_3711,In_1094,In_328);
nor U3712 (N_3712,In_575,In_59);
nor U3713 (N_3713,In_326,In_1049);
nor U3714 (N_3714,In_1600,In_1628);
and U3715 (N_3715,In_926,In_1370);
and U3716 (N_3716,In_307,In_679);
nand U3717 (N_3717,In_347,In_444);
nor U3718 (N_3718,In_586,In_101);
nor U3719 (N_3719,In_376,In_818);
and U3720 (N_3720,In_856,In_445);
or U3721 (N_3721,In_924,In_920);
xor U3722 (N_3722,In_1493,In_1397);
and U3723 (N_3723,In_427,In_572);
or U3724 (N_3724,In_874,In_781);
nand U3725 (N_3725,In_429,In_1979);
nor U3726 (N_3726,In_642,In_1278);
and U3727 (N_3727,In_265,In_109);
or U3728 (N_3728,In_1148,In_1976);
and U3729 (N_3729,In_315,In_691);
nand U3730 (N_3730,In_616,In_408);
nor U3731 (N_3731,In_1244,In_29);
and U3732 (N_3732,In_1900,In_383);
and U3733 (N_3733,In_1985,In_156);
nor U3734 (N_3734,In_1345,In_1193);
and U3735 (N_3735,In_826,In_477);
or U3736 (N_3736,In_1869,In_1455);
and U3737 (N_3737,In_1792,In_1557);
nand U3738 (N_3738,In_161,In_1187);
and U3739 (N_3739,In_1495,In_648);
or U3740 (N_3740,In_1773,In_25);
nor U3741 (N_3741,In_779,In_1044);
or U3742 (N_3742,In_791,In_1922);
and U3743 (N_3743,In_168,In_906);
nor U3744 (N_3744,In_1734,In_1434);
or U3745 (N_3745,In_735,In_1152);
or U3746 (N_3746,In_81,In_1286);
or U3747 (N_3747,In_1298,In_1565);
nand U3748 (N_3748,In_494,In_1518);
nor U3749 (N_3749,In_1407,In_1693);
nand U3750 (N_3750,In_90,In_849);
nor U3751 (N_3751,In_1206,In_1373);
nor U3752 (N_3752,In_141,In_1389);
or U3753 (N_3753,In_1634,In_752);
nand U3754 (N_3754,In_174,In_64);
nor U3755 (N_3755,In_1335,In_267);
and U3756 (N_3756,In_1213,In_1926);
and U3757 (N_3757,In_1081,In_712);
nand U3758 (N_3758,In_936,In_1988);
nand U3759 (N_3759,In_654,In_1609);
or U3760 (N_3760,In_1697,In_980);
nor U3761 (N_3761,In_966,In_1815);
nand U3762 (N_3762,In_1563,In_833);
and U3763 (N_3763,In_1380,In_1195);
or U3764 (N_3764,In_1493,In_391);
or U3765 (N_3765,In_1260,In_935);
or U3766 (N_3766,In_1323,In_327);
and U3767 (N_3767,In_1344,In_1901);
nand U3768 (N_3768,In_735,In_1585);
nor U3769 (N_3769,In_1250,In_875);
or U3770 (N_3770,In_1257,In_1300);
or U3771 (N_3771,In_731,In_284);
nand U3772 (N_3772,In_1300,In_1023);
and U3773 (N_3773,In_711,In_1385);
xor U3774 (N_3774,In_1158,In_65);
or U3775 (N_3775,In_472,In_1070);
or U3776 (N_3776,In_1159,In_611);
nor U3777 (N_3777,In_1220,In_281);
and U3778 (N_3778,In_1748,In_280);
nor U3779 (N_3779,In_1027,In_645);
or U3780 (N_3780,In_1494,In_933);
or U3781 (N_3781,In_1074,In_1979);
nor U3782 (N_3782,In_1428,In_266);
nor U3783 (N_3783,In_1717,In_1910);
nand U3784 (N_3784,In_625,In_324);
nor U3785 (N_3785,In_1595,In_976);
nor U3786 (N_3786,In_1541,In_1680);
nand U3787 (N_3787,In_889,In_1546);
or U3788 (N_3788,In_1431,In_422);
and U3789 (N_3789,In_710,In_1541);
or U3790 (N_3790,In_582,In_29);
nor U3791 (N_3791,In_1623,In_576);
nand U3792 (N_3792,In_291,In_85);
nor U3793 (N_3793,In_1271,In_983);
nor U3794 (N_3794,In_1272,In_831);
or U3795 (N_3795,In_1111,In_611);
nand U3796 (N_3796,In_32,In_1845);
or U3797 (N_3797,In_1162,In_5);
nor U3798 (N_3798,In_1182,In_162);
nand U3799 (N_3799,In_1870,In_1952);
nand U3800 (N_3800,In_635,In_202);
nand U3801 (N_3801,In_718,In_1836);
nand U3802 (N_3802,In_693,In_463);
or U3803 (N_3803,In_1467,In_369);
and U3804 (N_3804,In_1694,In_1014);
and U3805 (N_3805,In_1131,In_508);
nand U3806 (N_3806,In_805,In_1766);
or U3807 (N_3807,In_572,In_1082);
and U3808 (N_3808,In_1919,In_1665);
or U3809 (N_3809,In_525,In_1718);
and U3810 (N_3810,In_267,In_1515);
nor U3811 (N_3811,In_682,In_1485);
and U3812 (N_3812,In_1494,In_1747);
xnor U3813 (N_3813,In_810,In_647);
xor U3814 (N_3814,In_1416,In_566);
nand U3815 (N_3815,In_1598,In_1593);
and U3816 (N_3816,In_1823,In_1019);
nand U3817 (N_3817,In_543,In_1340);
nor U3818 (N_3818,In_286,In_1123);
nand U3819 (N_3819,In_1300,In_1836);
nor U3820 (N_3820,In_1227,In_717);
nand U3821 (N_3821,In_229,In_958);
or U3822 (N_3822,In_1652,In_1017);
and U3823 (N_3823,In_787,In_1898);
nand U3824 (N_3824,In_508,In_265);
nand U3825 (N_3825,In_227,In_1462);
or U3826 (N_3826,In_1004,In_1631);
and U3827 (N_3827,In_395,In_1949);
and U3828 (N_3828,In_1977,In_239);
and U3829 (N_3829,In_664,In_583);
or U3830 (N_3830,In_1266,In_604);
nand U3831 (N_3831,In_1416,In_1033);
and U3832 (N_3832,In_1328,In_564);
nor U3833 (N_3833,In_1608,In_884);
nor U3834 (N_3834,In_1543,In_377);
nor U3835 (N_3835,In_359,In_1566);
or U3836 (N_3836,In_1137,In_1176);
and U3837 (N_3837,In_981,In_410);
and U3838 (N_3838,In_1165,In_1782);
nor U3839 (N_3839,In_144,In_1490);
and U3840 (N_3840,In_813,In_1183);
or U3841 (N_3841,In_714,In_1890);
nor U3842 (N_3842,In_95,In_705);
or U3843 (N_3843,In_1945,In_1853);
nand U3844 (N_3844,In_930,In_1425);
nor U3845 (N_3845,In_1958,In_1746);
nand U3846 (N_3846,In_1146,In_965);
nand U3847 (N_3847,In_91,In_399);
nand U3848 (N_3848,In_761,In_639);
and U3849 (N_3849,In_1656,In_1263);
and U3850 (N_3850,In_394,In_571);
and U3851 (N_3851,In_1473,In_818);
nor U3852 (N_3852,In_679,In_327);
and U3853 (N_3853,In_459,In_1750);
and U3854 (N_3854,In_1272,In_9);
and U3855 (N_3855,In_862,In_1150);
nand U3856 (N_3856,In_1506,In_691);
and U3857 (N_3857,In_742,In_801);
nor U3858 (N_3858,In_485,In_573);
nand U3859 (N_3859,In_767,In_1241);
nand U3860 (N_3860,In_1407,In_1274);
nor U3861 (N_3861,In_628,In_1956);
nor U3862 (N_3862,In_1290,In_1017);
nand U3863 (N_3863,In_1259,In_1729);
nand U3864 (N_3864,In_762,In_1989);
and U3865 (N_3865,In_1997,In_1244);
or U3866 (N_3866,In_1763,In_1581);
and U3867 (N_3867,In_991,In_1578);
nor U3868 (N_3868,In_978,In_1007);
nor U3869 (N_3869,In_170,In_1949);
or U3870 (N_3870,In_1346,In_56);
and U3871 (N_3871,In_1269,In_899);
nor U3872 (N_3872,In_664,In_1682);
nand U3873 (N_3873,In_874,In_1047);
nor U3874 (N_3874,In_336,In_1786);
nand U3875 (N_3875,In_469,In_803);
nand U3876 (N_3876,In_296,In_1768);
or U3877 (N_3877,In_268,In_653);
nor U3878 (N_3878,In_984,In_705);
nor U3879 (N_3879,In_1125,In_689);
nand U3880 (N_3880,In_469,In_1391);
nand U3881 (N_3881,In_139,In_1638);
xor U3882 (N_3882,In_414,In_1140);
nand U3883 (N_3883,In_1552,In_1523);
nor U3884 (N_3884,In_1869,In_1983);
and U3885 (N_3885,In_697,In_76);
or U3886 (N_3886,In_1039,In_26);
nand U3887 (N_3887,In_681,In_1853);
and U3888 (N_3888,In_1265,In_1477);
and U3889 (N_3889,In_468,In_173);
nand U3890 (N_3890,In_94,In_643);
nand U3891 (N_3891,In_570,In_1680);
and U3892 (N_3892,In_664,In_712);
nor U3893 (N_3893,In_177,In_1712);
and U3894 (N_3894,In_1326,In_1287);
or U3895 (N_3895,In_1896,In_983);
nand U3896 (N_3896,In_395,In_907);
nand U3897 (N_3897,In_1912,In_1380);
nor U3898 (N_3898,In_1195,In_575);
nand U3899 (N_3899,In_1372,In_1308);
nor U3900 (N_3900,In_520,In_1144);
nor U3901 (N_3901,In_251,In_1471);
or U3902 (N_3902,In_969,In_817);
nor U3903 (N_3903,In_303,In_1628);
nand U3904 (N_3904,In_877,In_1613);
or U3905 (N_3905,In_449,In_523);
nor U3906 (N_3906,In_1163,In_348);
or U3907 (N_3907,In_1658,In_527);
nor U3908 (N_3908,In_367,In_534);
nor U3909 (N_3909,In_1677,In_537);
and U3910 (N_3910,In_984,In_1385);
nand U3911 (N_3911,In_447,In_243);
and U3912 (N_3912,In_235,In_845);
nand U3913 (N_3913,In_825,In_1746);
nand U3914 (N_3914,In_383,In_679);
nand U3915 (N_3915,In_1650,In_28);
or U3916 (N_3916,In_381,In_1639);
or U3917 (N_3917,In_1432,In_1923);
or U3918 (N_3918,In_1292,In_862);
and U3919 (N_3919,In_263,In_1568);
or U3920 (N_3920,In_857,In_918);
or U3921 (N_3921,In_1411,In_1752);
or U3922 (N_3922,In_186,In_1639);
or U3923 (N_3923,In_1636,In_1962);
and U3924 (N_3924,In_1838,In_1123);
nand U3925 (N_3925,In_319,In_67);
and U3926 (N_3926,In_1677,In_507);
xor U3927 (N_3927,In_400,In_33);
or U3928 (N_3928,In_864,In_1066);
nand U3929 (N_3929,In_1048,In_557);
and U3930 (N_3930,In_494,In_1068);
and U3931 (N_3931,In_583,In_1);
or U3932 (N_3932,In_603,In_1449);
and U3933 (N_3933,In_882,In_994);
and U3934 (N_3934,In_1720,In_1656);
or U3935 (N_3935,In_1347,In_1886);
and U3936 (N_3936,In_239,In_1310);
nor U3937 (N_3937,In_355,In_615);
nor U3938 (N_3938,In_1033,In_74);
nor U3939 (N_3939,In_518,In_388);
nand U3940 (N_3940,In_1406,In_964);
nor U3941 (N_3941,In_12,In_1031);
and U3942 (N_3942,In_863,In_1417);
and U3943 (N_3943,In_1414,In_578);
nor U3944 (N_3944,In_1326,In_1710);
nand U3945 (N_3945,In_1451,In_566);
and U3946 (N_3946,In_1589,In_1322);
nand U3947 (N_3947,In_690,In_1719);
or U3948 (N_3948,In_1561,In_924);
and U3949 (N_3949,In_6,In_1652);
nand U3950 (N_3950,In_1483,In_124);
and U3951 (N_3951,In_593,In_780);
nand U3952 (N_3952,In_420,In_938);
nand U3953 (N_3953,In_599,In_45);
and U3954 (N_3954,In_700,In_1667);
nor U3955 (N_3955,In_996,In_1982);
or U3956 (N_3956,In_673,In_1620);
nor U3957 (N_3957,In_1233,In_198);
nor U3958 (N_3958,In_1328,In_949);
nand U3959 (N_3959,In_600,In_974);
or U3960 (N_3960,In_1068,In_1290);
and U3961 (N_3961,In_1999,In_1633);
nor U3962 (N_3962,In_1523,In_416);
and U3963 (N_3963,In_1697,In_1692);
or U3964 (N_3964,In_134,In_1555);
nand U3965 (N_3965,In_115,In_1274);
and U3966 (N_3966,In_1235,In_1166);
or U3967 (N_3967,In_817,In_360);
nand U3968 (N_3968,In_177,In_1732);
nand U3969 (N_3969,In_754,In_582);
nor U3970 (N_3970,In_842,In_1137);
nand U3971 (N_3971,In_143,In_213);
nor U3972 (N_3972,In_759,In_588);
nor U3973 (N_3973,In_1432,In_48);
and U3974 (N_3974,In_834,In_1720);
nand U3975 (N_3975,In_1672,In_615);
or U3976 (N_3976,In_1481,In_279);
or U3977 (N_3977,In_115,In_1127);
and U3978 (N_3978,In_509,In_1804);
and U3979 (N_3979,In_1758,In_1612);
and U3980 (N_3980,In_249,In_1869);
nor U3981 (N_3981,In_1912,In_366);
and U3982 (N_3982,In_792,In_160);
nand U3983 (N_3983,In_1685,In_1226);
nand U3984 (N_3984,In_514,In_1895);
nor U3985 (N_3985,In_1324,In_798);
nand U3986 (N_3986,In_229,In_574);
or U3987 (N_3987,In_783,In_114);
and U3988 (N_3988,In_103,In_1960);
and U3989 (N_3989,In_912,In_1196);
nand U3990 (N_3990,In_1406,In_774);
nand U3991 (N_3991,In_757,In_369);
and U3992 (N_3992,In_1577,In_1275);
and U3993 (N_3993,In_1487,In_897);
and U3994 (N_3994,In_1892,In_1118);
or U3995 (N_3995,In_1586,In_1269);
nand U3996 (N_3996,In_1426,In_1360);
nor U3997 (N_3997,In_855,In_754);
or U3998 (N_3998,In_249,In_1359);
nand U3999 (N_3999,In_196,In_1974);
nand U4000 (N_4000,N_2161,N_1800);
and U4001 (N_4001,N_2823,N_1738);
nor U4002 (N_4002,N_3850,N_3876);
nor U4003 (N_4003,N_3866,N_2553);
and U4004 (N_4004,N_370,N_35);
nand U4005 (N_4005,N_2583,N_3751);
and U4006 (N_4006,N_3321,N_1246);
nor U4007 (N_4007,N_3326,N_3402);
or U4008 (N_4008,N_2192,N_956);
nor U4009 (N_4009,N_3291,N_1520);
nor U4010 (N_4010,N_110,N_2969);
or U4011 (N_4011,N_1216,N_768);
and U4012 (N_4012,N_856,N_954);
or U4013 (N_4013,N_3968,N_375);
or U4014 (N_4014,N_3969,N_1480);
and U4015 (N_4015,N_2370,N_484);
nand U4016 (N_4016,N_2475,N_3363);
or U4017 (N_4017,N_355,N_1045);
nor U4018 (N_4018,N_3693,N_3043);
and U4019 (N_4019,N_2171,N_1046);
nand U4020 (N_4020,N_70,N_518);
or U4021 (N_4021,N_2247,N_1065);
and U4022 (N_4022,N_3952,N_1871);
nor U4023 (N_4023,N_3209,N_2907);
and U4024 (N_4024,N_2094,N_1845);
nand U4025 (N_4025,N_174,N_3373);
nand U4026 (N_4026,N_2374,N_3914);
or U4027 (N_4027,N_1115,N_1126);
nor U4028 (N_4028,N_3390,N_3022);
or U4029 (N_4029,N_1359,N_3051);
nor U4030 (N_4030,N_2088,N_1863);
and U4031 (N_4031,N_1828,N_11);
xor U4032 (N_4032,N_2024,N_2238);
nor U4033 (N_4033,N_1457,N_3251);
nor U4034 (N_4034,N_1164,N_520);
nor U4035 (N_4035,N_3995,N_1456);
nor U4036 (N_4036,N_1025,N_794);
and U4037 (N_4037,N_604,N_148);
and U4038 (N_4038,N_2599,N_2114);
nor U4039 (N_4039,N_1669,N_2209);
nor U4040 (N_4040,N_1004,N_17);
or U4041 (N_4041,N_8,N_3989);
or U4042 (N_4042,N_2998,N_2637);
and U4043 (N_4043,N_1764,N_1125);
nand U4044 (N_4044,N_1847,N_1124);
or U4045 (N_4045,N_1439,N_466);
nand U4046 (N_4046,N_987,N_3240);
nand U4047 (N_4047,N_2430,N_1498);
or U4048 (N_4048,N_2232,N_932);
or U4049 (N_4049,N_599,N_2841);
and U4050 (N_4050,N_3613,N_2139);
and U4051 (N_4051,N_2741,N_879);
nor U4052 (N_4052,N_2473,N_742);
nand U4053 (N_4053,N_2158,N_246);
nand U4054 (N_4054,N_480,N_2331);
and U4055 (N_4055,N_3197,N_711);
nor U4056 (N_4056,N_57,N_44);
or U4057 (N_4057,N_1763,N_2235);
or U4058 (N_4058,N_2421,N_3011);
or U4059 (N_4059,N_313,N_493);
or U4060 (N_4060,N_30,N_1588);
nor U4061 (N_4061,N_426,N_1695);
nor U4062 (N_4062,N_1191,N_1467);
or U4063 (N_4063,N_3708,N_2979);
xor U4064 (N_4064,N_2973,N_94);
nor U4065 (N_4065,N_3211,N_1628);
xnor U4066 (N_4066,N_1374,N_1469);
or U4067 (N_4067,N_1364,N_3726);
nand U4068 (N_4068,N_1114,N_3109);
nand U4069 (N_4069,N_3714,N_1265);
nand U4070 (N_4070,N_736,N_1597);
or U4071 (N_4071,N_412,N_42);
and U4072 (N_4072,N_430,N_1454);
nor U4073 (N_4073,N_1809,N_1227);
nand U4074 (N_4074,N_2575,N_1591);
or U4075 (N_4075,N_1721,N_3340);
nand U4076 (N_4076,N_2497,N_2211);
and U4077 (N_4077,N_3210,N_238);
nor U4078 (N_4078,N_239,N_1388);
or U4079 (N_4079,N_380,N_114);
and U4080 (N_4080,N_559,N_3981);
and U4081 (N_4081,N_1733,N_1404);
or U4082 (N_4082,N_2526,N_2483);
nor U4083 (N_4083,N_2154,N_3806);
nor U4084 (N_4084,N_1602,N_3165);
nor U4085 (N_4085,N_1250,N_15);
nor U4086 (N_4086,N_801,N_131);
nor U4087 (N_4087,N_2103,N_1200);
and U4088 (N_4088,N_1236,N_1130);
xor U4089 (N_4089,N_2491,N_339);
nand U4090 (N_4090,N_846,N_1482);
and U4091 (N_4091,N_3136,N_1245);
or U4092 (N_4092,N_968,N_2166);
nor U4093 (N_4093,N_1251,N_660);
nor U4094 (N_4094,N_3830,N_2809);
nor U4095 (N_4095,N_2332,N_969);
nor U4096 (N_4096,N_2182,N_1709);
nand U4097 (N_4097,N_2616,N_3488);
or U4098 (N_4098,N_2866,N_3563);
nor U4099 (N_4099,N_3848,N_2359);
and U4100 (N_4100,N_860,N_404);
and U4101 (N_4101,N_2535,N_2002);
nand U4102 (N_4102,N_2673,N_3031);
xor U4103 (N_4103,N_3319,N_2034);
nor U4104 (N_4104,N_1116,N_3976);
and U4105 (N_4105,N_3464,N_1710);
and U4106 (N_4106,N_3865,N_2576);
nor U4107 (N_4107,N_1321,N_1765);
and U4108 (N_4108,N_3010,N_2444);
nand U4109 (N_4109,N_912,N_658);
or U4110 (N_4110,N_1197,N_3840);
nor U4111 (N_4111,N_3451,N_2302);
nor U4112 (N_4112,N_1948,N_1749);
or U4113 (N_4113,N_903,N_3349);
and U4114 (N_4114,N_2684,N_3843);
and U4115 (N_4115,N_2419,N_3379);
nand U4116 (N_4116,N_1564,N_2469);
nor U4117 (N_4117,N_391,N_2360);
or U4118 (N_4118,N_1899,N_3455);
nand U4119 (N_4119,N_883,N_245);
nor U4120 (N_4120,N_728,N_2791);
and U4121 (N_4121,N_612,N_1018);
nand U4122 (N_4122,N_920,N_3772);
nand U4123 (N_4123,N_3869,N_31);
or U4124 (N_4124,N_3584,N_820);
nor U4125 (N_4125,N_1458,N_3334);
nor U4126 (N_4126,N_3965,N_970);
nor U4127 (N_4127,N_309,N_3044);
nand U4128 (N_4128,N_368,N_1965);
or U4129 (N_4129,N_457,N_3424);
and U4130 (N_4130,N_1335,N_2005);
nand U4131 (N_4131,N_137,N_3318);
or U4132 (N_4132,N_282,N_2521);
nor U4133 (N_4133,N_2168,N_2717);
nor U4134 (N_4134,N_3774,N_3337);
nor U4135 (N_4135,N_1147,N_1796);
nand U4136 (N_4136,N_390,N_881);
nand U4137 (N_4137,N_2722,N_402);
nor U4138 (N_4138,N_3588,N_1425);
and U4139 (N_4139,N_2536,N_964);
nor U4140 (N_4140,N_3870,N_2325);
nand U4141 (N_4141,N_2733,N_598);
nand U4142 (N_4142,N_3554,N_3753);
and U4143 (N_4143,N_1369,N_3308);
nor U4144 (N_4144,N_3875,N_2932);
nand U4145 (N_4145,N_1553,N_3208);
nand U4146 (N_4146,N_2726,N_3019);
nand U4147 (N_4147,N_387,N_2015);
xnor U4148 (N_4148,N_3648,N_3028);
and U4149 (N_4149,N_2495,N_2128);
nand U4150 (N_4150,N_696,N_1746);
nor U4151 (N_4151,N_1193,N_2357);
nor U4152 (N_4152,N_2311,N_3509);
or U4153 (N_4153,N_385,N_1032);
nand U4154 (N_4154,N_2762,N_1473);
nor U4155 (N_4155,N_2819,N_806);
and U4156 (N_4156,N_3395,N_1795);
or U4157 (N_4157,N_2222,N_1515);
or U4158 (N_4158,N_3645,N_1692);
nand U4159 (N_4159,N_3361,N_588);
nand U4160 (N_4160,N_1451,N_3632);
nor U4161 (N_4161,N_3024,N_1519);
nor U4162 (N_4162,N_3570,N_2178);
nand U4163 (N_4163,N_720,N_2920);
nor U4164 (N_4164,N_1638,N_1403);
nor U4165 (N_4165,N_3264,N_914);
or U4166 (N_4166,N_3184,N_470);
or U4167 (N_4167,N_3078,N_2763);
nor U4168 (N_4168,N_3892,N_3545);
nor U4169 (N_4169,N_611,N_310);
nor U4170 (N_4170,N_1743,N_1975);
nand U4171 (N_4171,N_2615,N_1180);
and U4172 (N_4172,N_170,N_3769);
xnor U4173 (N_4173,N_2348,N_3482);
and U4174 (N_4174,N_804,N_2265);
nor U4175 (N_4175,N_469,N_550);
and U4176 (N_4176,N_3335,N_789);
or U4177 (N_4177,N_1323,N_1850);
or U4178 (N_4178,N_1900,N_1254);
nand U4179 (N_4179,N_3489,N_1481);
or U4180 (N_4180,N_3516,N_1605);
or U4181 (N_4181,N_3532,N_3849);
nand U4182 (N_4182,N_3822,N_3872);
nor U4183 (N_4183,N_281,N_1230);
nand U4184 (N_4184,N_2793,N_224);
nand U4185 (N_4185,N_1044,N_250);
or U4186 (N_4186,N_756,N_837);
and U4187 (N_4187,N_1675,N_3261);
or U4188 (N_4188,N_369,N_993);
nand U4189 (N_4189,N_304,N_88);
nor U4190 (N_4190,N_2596,N_894);
nor U4191 (N_4191,N_2938,N_3137);
nor U4192 (N_4192,N_3069,N_3504);
and U4193 (N_4193,N_3433,N_3606);
nor U4194 (N_4194,N_2046,N_1437);
nand U4195 (N_4195,N_3441,N_2428);
nand U4196 (N_4196,N_2507,N_2636);
or U4197 (N_4197,N_2287,N_3320);
nand U4198 (N_4198,N_775,N_121);
nor U4199 (N_4199,N_1702,N_2062);
nor U4200 (N_4200,N_1433,N_3375);
or U4201 (N_4201,N_3317,N_3686);
and U4202 (N_4202,N_691,N_2860);
nand U4203 (N_4203,N_529,N_1257);
or U4204 (N_4204,N_2908,N_2591);
and U4205 (N_4205,N_1214,N_396);
or U4206 (N_4206,N_188,N_2987);
nor U4207 (N_4207,N_3752,N_2692);
and U4208 (N_4208,N_2167,N_3634);
nor U4209 (N_4209,N_3707,N_1258);
nand U4210 (N_4210,N_3717,N_346);
and U4211 (N_4211,N_2269,N_2709);
nor U4212 (N_4212,N_1993,N_584);
or U4213 (N_4213,N_1831,N_3877);
or U4214 (N_4214,N_1249,N_2785);
or U4215 (N_4215,N_2886,N_1056);
and U4216 (N_4216,N_189,N_1677);
or U4217 (N_4217,N_3053,N_917);
nand U4218 (N_4218,N_3583,N_3585);
and U4219 (N_4219,N_3470,N_1579);
and U4220 (N_4220,N_365,N_592);
nor U4221 (N_4221,N_2163,N_1483);
nor U4222 (N_4222,N_3980,N_2669);
nor U4223 (N_4223,N_144,N_2858);
nor U4224 (N_4224,N_2116,N_3163);
and U4225 (N_4225,N_1646,N_2060);
nor U4226 (N_4226,N_2997,N_3512);
nand U4227 (N_4227,N_2658,N_1842);
and U4228 (N_4228,N_1362,N_1219);
nor U4229 (N_4229,N_3644,N_3819);
nor U4230 (N_4230,N_164,N_1274);
nor U4231 (N_4231,N_3929,N_2652);
or U4232 (N_4232,N_3192,N_74);
nor U4233 (N_4233,N_938,N_274);
or U4234 (N_4234,N_1931,N_3797);
nor U4235 (N_4235,N_2778,N_3421);
nor U4236 (N_4236,N_1512,N_2079);
or U4237 (N_4237,N_3151,N_1912);
and U4238 (N_4238,N_1231,N_3382);
or U4239 (N_4239,N_1853,N_3500);
nand U4240 (N_4240,N_474,N_1587);
or U4241 (N_4241,N_659,N_7);
nor U4242 (N_4242,N_1953,N_2445);
nand U4243 (N_4243,N_428,N_3802);
or U4244 (N_4244,N_3546,N_3612);
nand U4245 (N_4245,N_2234,N_294);
or U4246 (N_4246,N_3073,N_1021);
nor U4247 (N_4247,N_2050,N_1228);
nor U4248 (N_4248,N_3637,N_1547);
nor U4249 (N_4249,N_3032,N_3659);
or U4250 (N_4250,N_982,N_26);
or U4251 (N_4251,N_438,N_578);
nor U4252 (N_4252,N_1781,N_2217);
nor U4253 (N_4253,N_2693,N_679);
nor U4254 (N_4254,N_1140,N_3205);
or U4255 (N_4255,N_2057,N_1063);
and U4256 (N_4256,N_3267,N_3993);
and U4257 (N_4257,N_939,N_1492);
nand U4258 (N_4258,N_2423,N_2565);
and U4259 (N_4259,N_3037,N_1070);
or U4260 (N_4260,N_2221,N_1291);
nor U4261 (N_4261,N_3782,N_3131);
and U4262 (N_4262,N_3089,N_2623);
nand U4263 (N_4263,N_730,N_2665);
or U4264 (N_4264,N_3913,N_2329);
or U4265 (N_4265,N_82,N_3219);
nand U4266 (N_4266,N_3780,N_1616);
and U4267 (N_4267,N_1752,N_3573);
nor U4268 (N_4268,N_1969,N_1067);
nor U4269 (N_4269,N_947,N_877);
or U4270 (N_4270,N_2533,N_1460);
nand U4271 (N_4271,N_3496,N_1058);
nor U4272 (N_4272,N_1143,N_2455);
nor U4273 (N_4273,N_143,N_1664);
nand U4274 (N_4274,N_1570,N_741);
nand U4275 (N_4275,N_1431,N_2670);
or U4276 (N_4276,N_3933,N_2552);
and U4277 (N_4277,N_3878,N_1536);
nor U4278 (N_4278,N_2147,N_3419);
nor U4279 (N_4279,N_3936,N_467);
or U4280 (N_4280,N_2208,N_3156);
nor U4281 (N_4281,N_504,N_115);
or U4282 (N_4282,N_3259,N_924);
or U4283 (N_4283,N_2694,N_2939);
or U4284 (N_4284,N_576,N_3403);
nand U4285 (N_4285,N_360,N_1598);
nor U4286 (N_4286,N_999,N_3890);
and U4287 (N_4287,N_3578,N_107);
nand U4288 (N_4288,N_3345,N_1356);
nor U4289 (N_4289,N_1865,N_420);
and U4290 (N_4290,N_2316,N_2082);
nor U4291 (N_4291,N_1872,N_1332);
and U4292 (N_4292,N_3786,N_1340);
and U4293 (N_4293,N_198,N_1509);
or U4294 (N_4294,N_891,N_3443);
or U4295 (N_4295,N_2914,N_2405);
or U4296 (N_4296,N_297,N_3930);
nand U4297 (N_4297,N_1019,N_6);
nor U4298 (N_4298,N_1484,N_2951);
or U4299 (N_4299,N_171,N_3873);
nor U4300 (N_4300,N_1844,N_2981);
and U4301 (N_4301,N_610,N_434);
nor U4302 (N_4302,N_1833,N_2980);
or U4303 (N_4303,N_2011,N_2032);
nor U4304 (N_4304,N_2634,N_1317);
and U4305 (N_4305,N_1131,N_686);
nor U4306 (N_4306,N_3541,N_3339);
nor U4307 (N_4307,N_3127,N_2874);
nand U4308 (N_4308,N_76,N_1855);
nor U4309 (N_4309,N_3795,N_2344);
or U4310 (N_4310,N_2889,N_1626);
nand U4311 (N_4311,N_413,N_307);
nor U4312 (N_4312,N_1017,N_3682);
nor U4313 (N_4313,N_1946,N_3939);
nand U4314 (N_4314,N_2558,N_2897);
nor U4315 (N_4315,N_2365,N_1665);
or U4316 (N_4316,N_1778,N_431);
nor U4317 (N_4317,N_3486,N_3364);
or U4318 (N_4318,N_1555,N_178);
or U4319 (N_4319,N_1790,N_613);
or U4320 (N_4320,N_996,N_2283);
nand U4321 (N_4321,N_3766,N_3549);
nor U4322 (N_4322,N_3166,N_1703);
nor U4323 (N_4323,N_1732,N_2108);
and U4324 (N_4324,N_1985,N_2417);
nor U4325 (N_4325,N_2878,N_2856);
nand U4326 (N_4326,N_1128,N_1939);
nor U4327 (N_4327,N_1071,N_564);
nand U4328 (N_4328,N_895,N_96);
nand U4329 (N_4329,N_3323,N_1687);
and U4330 (N_4330,N_2508,N_1905);
nand U4331 (N_4331,N_3255,N_2572);
nor U4332 (N_4332,N_1206,N_1590);
nor U4333 (N_4333,N_2194,N_3428);
or U4334 (N_4334,N_3738,N_3749);
nor U4335 (N_4335,N_1455,N_196);
nor U4336 (N_4336,N_2440,N_347);
nor U4337 (N_4337,N_487,N_3005);
nor U4338 (N_4338,N_3773,N_3760);
and U4339 (N_4339,N_3330,N_3108);
nor U4340 (N_4340,N_482,N_2790);
nand U4341 (N_4341,N_2853,N_1613);
nand U4342 (N_4342,N_2100,N_2227);
nand U4343 (N_4343,N_754,N_244);
nand U4344 (N_4344,N_1154,N_3423);
nand U4345 (N_4345,N_650,N_2281);
nand U4346 (N_4346,N_1755,N_1312);
and U4347 (N_4347,N_3017,N_3880);
or U4348 (N_4348,N_1366,N_2934);
nand U4349 (N_4349,N_3799,N_2952);
xor U4350 (N_4350,N_2319,N_2277);
or U4351 (N_4351,N_2588,N_2604);
or U4352 (N_4352,N_928,N_1138);
nand U4353 (N_4353,N_71,N_3139);
and U4354 (N_4354,N_959,N_326);
nor U4355 (N_4355,N_4,N_2102);
or U4356 (N_4356,N_111,N_2321);
and U4357 (N_4357,N_834,N_436);
nor U4358 (N_4358,N_528,N_1995);
nor U4359 (N_4359,N_1997,N_859);
or U4360 (N_4360,N_1575,N_135);
nor U4361 (N_4361,N_3539,N_3172);
nor U4362 (N_4362,N_3391,N_701);
xnor U4363 (N_4363,N_2600,N_1052);
and U4364 (N_4364,N_2725,N_278);
or U4365 (N_4365,N_880,N_3857);
nand U4366 (N_4366,N_3133,N_2447);
and U4367 (N_4367,N_1854,N_3737);
nor U4368 (N_4368,N_3485,N_2869);
or U4369 (N_4369,N_853,N_2891);
nand U4370 (N_4370,N_3919,N_2944);
nand U4371 (N_4371,N_3860,N_39);
nand U4372 (N_4372,N_721,N_3847);
and U4373 (N_4373,N_875,N_887);
or U4374 (N_4374,N_454,N_1714);
or U4375 (N_4375,N_2774,N_1040);
and U4376 (N_4376,N_3275,N_481);
and U4377 (N_4377,N_2931,N_957);
nor U4378 (N_4378,N_3220,N_2561);
or U4379 (N_4379,N_1479,N_955);
nor U4380 (N_4380,N_544,N_2230);
xnor U4381 (N_4381,N_2191,N_718);
and U4382 (N_4382,N_2342,N_2481);
nand U4383 (N_4383,N_1622,N_2160);
or U4384 (N_4384,N_3503,N_2551);
and U4385 (N_4385,N_502,N_483);
nand U4386 (N_4386,N_3007,N_1525);
nor U4387 (N_4387,N_3371,N_2775);
nor U4388 (N_4388,N_722,N_1859);
nand U4389 (N_4389,N_2894,N_3125);
and U4390 (N_4390,N_2426,N_288);
nand U4391 (N_4391,N_3740,N_795);
nand U4392 (N_4392,N_3378,N_3915);
and U4393 (N_4393,N_2272,N_3864);
nand U4394 (N_4394,N_3805,N_3761);
nand U4395 (N_4395,N_3091,N_1630);
nand U4396 (N_4396,N_2511,N_1252);
nor U4397 (N_4397,N_3954,N_733);
and U4398 (N_4398,N_509,N_2040);
nor U4399 (N_4399,N_60,N_348);
or U4400 (N_4400,N_3609,N_2493);
nor U4401 (N_4401,N_336,N_2383);
nor U4402 (N_4402,N_3181,N_2314);
nor U4403 (N_4403,N_1401,N_745);
or U4404 (N_4404,N_3577,N_1267);
nor U4405 (N_4405,N_3683,N_2564);
or U4406 (N_4406,N_739,N_2095);
nand U4407 (N_4407,N_2346,N_324);
and U4408 (N_4408,N_2366,N_1350);
nand U4409 (N_4409,N_399,N_1843);
or U4410 (N_4410,N_442,N_3757);
nand U4411 (N_4411,N_2458,N_3076);
or U4412 (N_4412,N_2186,N_958);
and U4413 (N_4413,N_1827,N_1349);
nor U4414 (N_4414,N_1820,N_748);
or U4415 (N_4415,N_2259,N_2524);
nor U4416 (N_4416,N_565,N_2412);
and U4417 (N_4417,N_3800,N_2459);
nor U4418 (N_4418,N_1314,N_854);
nand U4419 (N_4419,N_3863,N_2584);
nand U4420 (N_4420,N_2685,N_285);
and U4421 (N_4421,N_862,N_1560);
and U4422 (N_4422,N_991,N_3359);
nand U4423 (N_4423,N_1650,N_3654);
nor U4424 (N_4424,N_3353,N_343);
nor U4425 (N_4425,N_3083,N_1717);
nor U4426 (N_4426,N_3506,N_2590);
and U4427 (N_4427,N_2449,N_203);
nor U4428 (N_4428,N_3288,N_3346);
nand U4429 (N_4429,N_3140,N_3234);
nand U4430 (N_4430,N_1806,N_2753);
nand U4431 (N_4431,N_3107,N_3587);
or U4432 (N_4432,N_1099,N_1508);
and U4433 (N_4433,N_2305,N_2832);
or U4434 (N_4434,N_433,N_1829);
nor U4435 (N_4435,N_2432,N_663);
or U4436 (N_4436,N_2683,N_1857);
and U4437 (N_4437,N_3104,N_3979);
nand U4438 (N_4438,N_3175,N_2334);
or U4439 (N_4439,N_717,N_253);
and U4440 (N_4440,N_1725,N_2004);
and U4441 (N_4441,N_1719,N_800);
or U4442 (N_4442,N_1470,N_423);
or U4443 (N_4443,N_3605,N_1033);
or U4444 (N_4444,N_1619,N_2164);
nand U4445 (N_4445,N_777,N_587);
nor U4446 (N_4446,N_3653,N_3960);
nand U4447 (N_4447,N_1452,N_3871);
and U4448 (N_4448,N_1450,N_1610);
and U4449 (N_4449,N_429,N_1060);
and U4450 (N_4450,N_3988,N_583);
nor U4451 (N_4451,N_1448,N_2156);
and U4452 (N_4452,N_2420,N_2863);
and U4453 (N_4453,N_1976,N_2345);
or U4454 (N_4454,N_1756,N_2755);
nand U4455 (N_4455,N_2077,N_1649);
nand U4456 (N_4456,N_1101,N_1290);
nand U4457 (N_4457,N_1566,N_1625);
and U4458 (N_4458,N_427,N_2971);
and U4459 (N_4459,N_1916,N_3491);
and U4460 (N_4460,N_3299,N_3484);
nand U4461 (N_4461,N_1208,N_1438);
nor U4462 (N_4462,N_1270,N_3307);
nor U4463 (N_4463,N_2900,N_1313);
or U4464 (N_4464,N_1989,N_3001);
nor U4465 (N_4465,N_1540,N_3972);
and U4466 (N_4466,N_1218,N_2946);
and U4467 (N_4467,N_3056,N_1851);
and U4468 (N_4468,N_2566,N_3305);
or U4469 (N_4469,N_2547,N_829);
and U4470 (N_4470,N_965,N_1959);
nand U4471 (N_4471,N_3216,N_2075);
nor U4472 (N_4472,N_361,N_1468);
nand U4473 (N_4473,N_275,N_931);
or U4474 (N_4474,N_3789,N_1426);
nand U4475 (N_4475,N_2361,N_2326);
and U4476 (N_4476,N_217,N_2000);
or U4477 (N_4477,N_2715,N_119);
or U4478 (N_4478,N_3457,N_2834);
and U4479 (N_4479,N_523,N_835);
and U4480 (N_4480,N_2245,N_828);
or U4481 (N_4481,N_120,N_3967);
and U4482 (N_4482,N_2390,N_1495);
or U4483 (N_4483,N_1656,N_619);
nand U4484 (N_4484,N_2389,N_439);
or U4485 (N_4485,N_3592,N_2610);
nor U4486 (N_4486,N_2527,N_3668);
and U4487 (N_4487,N_2068,N_3884);
and U4488 (N_4488,N_3164,N_1574);
nand U4489 (N_4489,N_3560,N_3018);
nand U4490 (N_4490,N_1557,N_2628);
nor U4491 (N_4491,N_2422,N_651);
nand U4492 (N_4492,N_3096,N_734);
and U4493 (N_4493,N_1594,N_2396);
and U4494 (N_4494,N_1760,N_1518);
and U4495 (N_4495,N_802,N_1963);
and U4496 (N_4496,N_2810,N_642);
nor U4497 (N_4497,N_1647,N_3452);
or U4498 (N_4498,N_2700,N_750);
nor U4499 (N_4499,N_3436,N_1996);
nand U4500 (N_4500,N_625,N_2736);
and U4501 (N_4501,N_3315,N_329);
nor U4502 (N_4502,N_3077,N_3372);
nor U4503 (N_4503,N_2789,N_3568);
or U4504 (N_4504,N_791,N_3710);
or U4505 (N_4505,N_3669,N_1632);
nand U4506 (N_4506,N_940,N_3505);
or U4507 (N_4507,N_476,N_1176);
nor U4508 (N_4508,N_126,N_3700);
or U4509 (N_4509,N_3312,N_3727);
nand U4510 (N_4510,N_2587,N_3273);
nand U4511 (N_4511,N_3343,N_2732);
nand U4512 (N_4512,N_868,N_3879);
nand U4513 (N_4513,N_644,N_590);
or U4514 (N_4514,N_2391,N_3134);
and U4515 (N_4515,N_3111,N_1260);
and U4516 (N_4516,N_1223,N_661);
or U4517 (N_4517,N_3442,N_142);
and U4518 (N_4518,N_2697,N_1173);
nand U4519 (N_4519,N_1648,N_3515);
nor U4520 (N_4520,N_3129,N_1165);
xor U4521 (N_4521,N_3818,N_549);
or U4522 (N_4522,N_2003,N_532);
and U4523 (N_4523,N_1973,N_944);
and U4524 (N_4524,N_827,N_3049);
nor U4525 (N_4525,N_2418,N_1885);
nor U4526 (N_4526,N_715,N_1586);
or U4527 (N_4527,N_3257,N_1023);
nand U4528 (N_4528,N_3713,N_494);
nor U4529 (N_4529,N_377,N_374);
nand U4530 (N_4530,N_1264,N_2795);
nand U4531 (N_4531,N_3511,N_3651);
nand U4532 (N_4532,N_735,N_2734);
nand U4533 (N_4533,N_3286,N_444);
and U4534 (N_4534,N_1041,N_1753);
nand U4535 (N_4535,N_2532,N_208);
nand U4536 (N_4536,N_595,N_1888);
nand U4537 (N_4537,N_3928,N_2993);
nand U4538 (N_4538,N_1798,N_1097);
nand U4539 (N_4539,N_2905,N_89);
nor U4540 (N_4540,N_1676,N_3271);
nand U4541 (N_4541,N_1053,N_2876);
nor U4542 (N_4542,N_2070,N_3697);
or U4543 (N_4543,N_3694,N_786);
and U4544 (N_4544,N_1834,N_2594);
or U4545 (N_4545,N_3723,N_3425);
nor U4546 (N_4546,N_749,N_2974);
or U4547 (N_4547,N_140,N_3638);
and U4548 (N_4548,N_2090,N_2065);
or U4549 (N_4549,N_2701,N_3762);
or U4550 (N_4550,N_2398,N_1668);
nand U4551 (N_4551,N_2620,N_1416);
nand U4552 (N_4552,N_2892,N_1920);
nor U4553 (N_4553,N_1705,N_477);
or U4554 (N_4554,N_3206,N_1195);
nand U4555 (N_4555,N_3739,N_1330);
and U4556 (N_4556,N_418,N_1292);
nand U4557 (N_4557,N_1672,N_552);
nand U4558 (N_4558,N_3828,N_3063);
and U4559 (N_4559,N_1381,N_50);
or U4560 (N_4560,N_1375,N_3026);
and U4561 (N_4561,N_3896,N_3962);
nand U4562 (N_4562,N_1029,N_3183);
or U4563 (N_4563,N_1242,N_2196);
or U4564 (N_4564,N_1568,N_1861);
nand U4565 (N_4565,N_1783,N_3189);
and U4566 (N_4566,N_2923,N_3118);
or U4567 (N_4567,N_1136,N_724);
or U4568 (N_4568,N_2279,N_1110);
nand U4569 (N_4569,N_3394,N_490);
and U4570 (N_4570,N_3322,N_2667);
and U4571 (N_4571,N_3122,N_3987);
nor U4572 (N_4572,N_545,N_819);
nand U4573 (N_4573,N_3327,N_1137);
nand U4574 (N_4574,N_75,N_3473);
nand U4575 (N_4575,N_112,N_150);
and U4576 (N_4576,N_1471,N_2586);
nor U4577 (N_4577,N_1127,N_283);
nor U4578 (N_4578,N_3961,N_2007);
and U4579 (N_4579,N_3833,N_972);
or U4580 (N_4580,N_3852,N_2833);
nand U4581 (N_4581,N_496,N_1205);
or U4582 (N_4582,N_2746,N_3179);
nand U4583 (N_4583,N_3071,N_1226);
or U4584 (N_4584,N_2339,N_1550);
nor U4585 (N_4585,N_247,N_3925);
and U4586 (N_4586,N_2071,N_1036);
and U4587 (N_4587,N_521,N_1713);
nor U4588 (N_4588,N_2001,N_124);
and U4589 (N_4589,N_3177,N_479);
nor U4590 (N_4590,N_2333,N_3365);
nand U4591 (N_4591,N_1624,N_1529);
and U4592 (N_4592,N_173,N_1870);
or U4593 (N_4593,N_1322,N_3298);
and U4594 (N_4594,N_976,N_3100);
nand U4595 (N_4595,N_2513,N_1024);
nand U4596 (N_4596,N_3661,N_424);
and U4597 (N_4597,N_1802,N_77);
and U4598 (N_4598,N_617,N_746);
and U4599 (N_4599,N_1734,N_2848);
nand U4600 (N_4600,N_416,N_3949);
nand U4601 (N_4601,N_1561,N_2078);
and U4602 (N_4602,N_3050,N_2373);
xnor U4603 (N_4603,N_472,N_252);
and U4604 (N_4604,N_2101,N_488);
or U4605 (N_4605,N_367,N_1892);
nand U4606 (N_4606,N_2385,N_3589);
and U4607 (N_4607,N_2274,N_3012);
and U4608 (N_4608,N_386,N_1813);
nand U4609 (N_4609,N_784,N_184);
nand U4610 (N_4610,N_3158,N_2772);
and U4611 (N_4611,N_2503,N_692);
nor U4612 (N_4612,N_3985,N_3947);
and U4613 (N_4613,N_3266,N_2461);
and U4614 (N_4614,N_3374,N_3622);
or U4615 (N_4615,N_2155,N_1031);
or U4616 (N_4616,N_857,N_738);
or U4617 (N_4617,N_1447,N_378);
or U4618 (N_4618,N_3520,N_2084);
nor U4619 (N_4619,N_3688,N_2237);
nor U4620 (N_4620,N_3767,N_1373);
or U4621 (N_4621,N_762,N_656);
and U4622 (N_4622,N_2133,N_1463);
or U4623 (N_4623,N_1810,N_1237);
nor U4624 (N_4624,N_3923,N_162);
nand U4625 (N_4625,N_2462,N_3845);
xor U4626 (N_4626,N_3788,N_539);
and U4627 (N_4627,N_3282,N_2335);
nand U4628 (N_4628,N_1100,N_1192);
nor U4629 (N_4629,N_1659,N_1316);
and U4630 (N_4630,N_3831,N_1670);
and U4631 (N_4631,N_1609,N_1567);
nand U4632 (N_4632,N_3709,N_1990);
or U4633 (N_4633,N_966,N_838);
nor U4634 (N_4634,N_3296,N_3676);
and U4635 (N_4635,N_1503,N_1690);
or U4636 (N_4636,N_906,N_2786);
and U4637 (N_4637,N_2153,N_2782);
nor U4638 (N_4638,N_3973,N_3008);
nand U4639 (N_4639,N_602,N_3047);
and U4640 (N_4640,N_2750,N_2355);
nor U4641 (N_4641,N_2215,N_2253);
and U4642 (N_4642,N_2119,N_269);
and U4643 (N_4643,N_1992,N_3030);
and U4644 (N_4644,N_1917,N_2142);
or U4645 (N_4645,N_1122,N_3499);
or U4646 (N_4646,N_3775,N_1222);
nand U4647 (N_4647,N_1506,N_3029);
or U4648 (N_4648,N_2143,N_3200);
nand U4649 (N_4649,N_2567,N_2047);
and U4650 (N_4650,N_175,N_2067);
nor U4651 (N_4651,N_2268,N_3674);
and U4652 (N_4652,N_177,N_3121);
nand U4653 (N_4653,N_3405,N_2251);
nor U4654 (N_4654,N_3883,N_2206);
and U4655 (N_4655,N_3791,N_2045);
nand U4656 (N_4656,N_554,N_2985);
nor U4657 (N_4657,N_344,N_2557);
and U4658 (N_4658,N_312,N_2443);
or U4659 (N_4659,N_3715,N_3841);
xor U4660 (N_4660,N_93,N_2482);
nor U4661 (N_4661,N_3430,N_1149);
nand U4662 (N_4662,N_681,N_3983);
or U4663 (N_4663,N_1633,N_852);
or U4664 (N_4664,N_2541,N_130);
and U4665 (N_4665,N_2677,N_1098);
nand U4666 (N_4666,N_195,N_1740);
xor U4667 (N_4667,N_1421,N_1611);
and U4668 (N_4668,N_92,N_971);
or U4669 (N_4669,N_716,N_2804);
nor U4670 (N_4670,N_287,N_757);
nand U4671 (N_4671,N_3075,N_2127);
and U4672 (N_4672,N_2500,N_759);
nand U4673 (N_4673,N_1277,N_3438);
nor U4674 (N_4674,N_52,N_1837);
nor U4675 (N_4675,N_1129,N_787);
or U4676 (N_4676,N_2766,N_2059);
or U4677 (N_4677,N_1824,N_645);
xor U4678 (N_4678,N_305,N_1879);
and U4679 (N_4679,N_2574,N_2330);
or U4680 (N_4680,N_364,N_2777);
nand U4681 (N_4681,N_2427,N_2976);
nand U4682 (N_4682,N_21,N_3734);
nand U4683 (N_4683,N_3639,N_761);
and U4684 (N_4684,N_1631,N_1935);
nor U4685 (N_4685,N_2120,N_1583);
nand U4686 (N_4686,N_394,N_3905);
nand U4687 (N_4687,N_505,N_2801);
or U4688 (N_4688,N_3141,N_446);
nor U4689 (N_4689,N_3497,N_1394);
and U4690 (N_4690,N_3437,N_1510);
and U4691 (N_4691,N_3755,N_901);
and U4692 (N_4692,N_1343,N_2528);
and U4693 (N_4693,N_2960,N_2903);
nor U4694 (N_4694,N_593,N_2170);
nand U4695 (N_4695,N_1476,N_3630);
nor U4696 (N_4696,N_3039,N_580);
nor U4697 (N_4697,N_3268,N_1535);
nor U4698 (N_4698,N_3994,N_3193);
nor U4699 (N_4699,N_1042,N_1177);
or U4700 (N_4700,N_376,N_2220);
nand U4701 (N_4701,N_2214,N_1822);
and U4702 (N_4702,N_2861,N_513);
or U4703 (N_4703,N_2195,N_2608);
and U4704 (N_4704,N_2376,N_2606);
nor U4705 (N_4705,N_3931,N_1107);
and U4706 (N_4706,N_3202,N_54);
or U4707 (N_4707,N_3918,N_1396);
nor U4708 (N_4708,N_1663,N_1516);
nor U4709 (N_4709,N_1901,N_3675);
nand U4710 (N_4710,N_641,N_330);
nand U4711 (N_4711,N_2674,N_2118);
nand U4712 (N_4712,N_3553,N_2712);
nor U4713 (N_4713,N_3218,N_1720);
and U4714 (N_4714,N_2761,N_1729);
nor U4715 (N_4715,N_236,N_271);
nand U4716 (N_4716,N_1701,N_3445);
nand U4717 (N_4717,N_3508,N_1696);
or U4718 (N_4718,N_2307,N_2436);
nor U4719 (N_4719,N_2501,N_2463);
nand U4720 (N_4720,N_2924,N_2883);
nand U4721 (N_4721,N_2957,N_713);
or U4722 (N_4722,N_1545,N_3106);
nand U4723 (N_4723,N_945,N_3025);
and U4724 (N_4724,N_2852,N_2431);
nand U4725 (N_4725,N_2505,N_1889);
and U4726 (N_4726,N_3997,N_1694);
nand U4727 (N_4727,N_2288,N_1166);
or U4728 (N_4728,N_3957,N_3538);
or U4729 (N_4729,N_2991,N_1262);
and U4730 (N_4730,N_3416,N_1980);
or U4731 (N_4731,N_3518,N_83);
or U4732 (N_4732,N_694,N_202);
nand U4733 (N_4733,N_2241,N_3564);
nand U4734 (N_4734,N_3617,N_905);
nand U4735 (N_4735,N_1298,N_2913);
or U4736 (N_4736,N_1420,N_2687);
or U4737 (N_4737,N_1679,N_3274);
nand U4738 (N_4738,N_2956,N_676);
or U4739 (N_4739,N_1918,N_1397);
nor U4740 (N_4740,N_1848,N_664);
nor U4741 (N_4741,N_3784,N_1096);
or U4742 (N_4742,N_3474,N_501);
nor U4743 (N_4743,N_2893,N_1247);
and U4744 (N_4744,N_3458,N_3493);
nand U4745 (N_4745,N_1315,N_435);
nand U4746 (N_4746,N_1662,N_1442);
nand U4747 (N_4747,N_3746,N_2486);
nor U4748 (N_4748,N_5,N_463);
and U4749 (N_4749,N_2271,N_2631);
nor U4750 (N_4750,N_280,N_3842);
and U4751 (N_4751,N_631,N_3471);
or U4752 (N_4752,N_395,N_2571);
or U4753 (N_4753,N_3519,N_1748);
and U4754 (N_4754,N_2854,N_2613);
nand U4755 (N_4755,N_2593,N_1534);
nand U4756 (N_4756,N_1414,N_2977);
or U4757 (N_4757,N_1273,N_2758);
nor U4758 (N_4758,N_3524,N_2515);
nor U4759 (N_4759,N_3839,N_2134);
and U4760 (N_4760,N_2747,N_2918);
and U4761 (N_4761,N_3358,N_2087);
nor U4762 (N_4762,N_1325,N_1085);
nor U4763 (N_4763,N_3556,N_946);
and U4764 (N_4764,N_13,N_1329);
or U4765 (N_4765,N_522,N_2506);
and U4766 (N_4766,N_485,N_465);
and U4767 (N_4767,N_1599,N_3874);
nor U4768 (N_4768,N_3376,N_1064);
nand U4769 (N_4769,N_432,N_2783);
or U4770 (N_4770,N_1794,N_3277);
nor U4771 (N_4771,N_3745,N_586);
nand U4772 (N_4772,N_3702,N_3594);
and U4773 (N_4773,N_1121,N_3858);
or U4774 (N_4774,N_1938,N_186);
and U4775 (N_4775,N_653,N_2017);
nor U4776 (N_4776,N_1440,N_2621);
nor U4777 (N_4777,N_3641,N_1123);
and U4778 (N_4778,N_3623,N_1982);
and U4779 (N_4779,N_279,N_3704);
nand U4780 (N_4780,N_108,N_1741);
or U4781 (N_4781,N_296,N_258);
nor U4782 (N_4782,N_2708,N_1275);
or U4783 (N_4783,N_3383,N_2009);
nor U4784 (N_4784,N_2409,N_3649);
nand U4785 (N_4785,N_191,N_194);
nand U4786 (N_4786,N_3064,N_3329);
and U4787 (N_4787,N_3671,N_425);
nand U4788 (N_4788,N_2146,N_833);
or U4789 (N_4789,N_1849,N_86);
or U4790 (N_4790,N_1637,N_902);
or U4791 (N_4791,N_3033,N_1187);
xnor U4792 (N_4792,N_1788,N_421);
nand U4793 (N_4793,N_0,N_366);
or U4794 (N_4794,N_1776,N_678);
and U4795 (N_4795,N_1148,N_3174);
or U4796 (N_4796,N_3730,N_2570);
nand U4797 (N_4797,N_899,N_363);
and U4798 (N_4798,N_2180,N_2464);
nor U4799 (N_4799,N_1907,N_3851);
and U4800 (N_4800,N_2585,N_3432);
or U4801 (N_4801,N_2203,N_1139);
and U4802 (N_4802,N_3945,N_1947);
and U4803 (N_4803,N_2996,N_1814);
and U4804 (N_4804,N_2554,N_1202);
nor U4805 (N_4805,N_2499,N_1062);
nor U4806 (N_4806,N_890,N_3814);
nand U4807 (N_4807,N_2239,N_3357);
nand U4808 (N_4808,N_1288,N_3581);
nand U4809 (N_4809,N_411,N_2661);
xnor U4810 (N_4810,N_2959,N_2818);
and U4811 (N_4811,N_2984,N_113);
and U4812 (N_4812,N_1168,N_2165);
nand U4813 (N_4813,N_2560,N_2144);
nor U4814 (N_4814,N_1429,N_608);
nand U4815 (N_4815,N_2131,N_1673);
or U4816 (N_4816,N_2053,N_2954);
nor U4817 (N_4817,N_1157,N_1392);
nor U4818 (N_4818,N_1612,N_2796);
or U4819 (N_4819,N_2243,N_889);
nor U4820 (N_4820,N_3909,N_3054);
nand U4821 (N_4821,N_2290,N_1759);
and U4822 (N_4822,N_1897,N_2051);
or U4823 (N_4823,N_3820,N_102);
or U4824 (N_4824,N_2740,N_2113);
nor U4825 (N_4825,N_1235,N_1689);
nor U4826 (N_4826,N_1576,N_536);
nor U4827 (N_4827,N_3227,N_2104);
and U4828 (N_4828,N_916,N_58);
and U4829 (N_4829,N_2825,N_2990);
nand U4830 (N_4830,N_3105,N_3042);
and U4831 (N_4831,N_1183,N_3698);
nand U4832 (N_4832,N_1327,N_49);
and U4833 (N_4833,N_712,N_3514);
or U4834 (N_4834,N_2964,N_3048);
nand U4835 (N_4835,N_556,N_1867);
nand U4836 (N_4836,N_1181,N_963);
and U4837 (N_4837,N_630,N_2025);
and U4838 (N_4838,N_125,N_320);
or U4839 (N_4839,N_3195,N_3341);
nand U4840 (N_4840,N_155,N_621);
or U4841 (N_4841,N_2441,N_867);
or U4842 (N_4842,N_2713,N_337);
nor U4843 (N_4843,N_1234,N_3369);
nor U4844 (N_4844,N_2019,N_910);
nor U4845 (N_4845,N_1651,N_241);
nor U4846 (N_4846,N_2364,N_1944);
nand U4847 (N_4847,N_2072,N_3236);
or U4848 (N_4848,N_193,N_1078);
and U4849 (N_4849,N_3162,N_2926);
and U4850 (N_4850,N_2308,N_3510);
or U4851 (N_4851,N_508,N_109);
nand U4852 (N_4852,N_1823,N_3920);
or U4853 (N_4853,N_2320,N_2555);
and U4854 (N_4854,N_1039,N_1000);
nand U4855 (N_4855,N_1028,N_1384);
nor U4856 (N_4856,N_805,N_2757);
or U4857 (N_4857,N_1528,N_3169);
and U4858 (N_4858,N_1009,N_567);
or U4859 (N_4859,N_1977,N_409);
nand U4860 (N_4860,N_1511,N_2136);
nor U4861 (N_4861,N_1789,N_1715);
nor U4862 (N_4862,N_3922,N_2812);
or U4863 (N_4863,N_3336,N_3072);
and U4864 (N_4864,N_1300,N_2703);
and U4865 (N_4865,N_2061,N_2837);
or U4866 (N_4866,N_1419,N_915);
and U4867 (N_4867,N_1391,N_1502);
and U4868 (N_4868,N_3492,N_2830);
or U4869 (N_4869,N_277,N_3910);
or U4870 (N_4870,N_2680,N_2972);
and U4871 (N_4871,N_2556,N_3978);
and U4872 (N_4872,N_3558,N_1770);
nor U4873 (N_4873,N_1109,N_2888);
or U4874 (N_4874,N_1441,N_3304);
nor U4875 (N_4875,N_3422,N_3355);
nor U4876 (N_4876,N_2205,N_551);
or U4877 (N_4877,N_3098,N_468);
nor U4878 (N_4878,N_1209,N_1059);
nand U4879 (N_4879,N_1395,N_221);
and U4880 (N_4880,N_2476,N_1604);
or U4881 (N_4881,N_1546,N_157);
nand U4882 (N_4882,N_3817,N_3706);
nand U4883 (N_4883,N_2442,N_3916);
nor U4884 (N_4884,N_316,N_1285);
nor U4885 (N_4885,N_3477,N_3387);
nand U4886 (N_4886,N_2967,N_1606);
and U4887 (N_4887,N_3625,N_677);
nand U4888 (N_4888,N_1531,N_1652);
and U4889 (N_4889,N_2484,N_1805);
or U4890 (N_4890,N_3908,N_1999);
nand U4891 (N_4891,N_790,N_3897);
xor U4892 (N_4892,N_2159,N_3113);
nand U4893 (N_4893,N_1818,N_807);
or U4894 (N_4894,N_2640,N_1517);
and U4895 (N_4895,N_232,N_2306);
nand U4896 (N_4896,N_1514,N_704);
or U4897 (N_4897,N_497,N_3170);
nand U4898 (N_4898,N_3217,N_3821);
nor U4899 (N_4899,N_937,N_654);
or U4900 (N_4900,N_1875,N_3690);
nor U4901 (N_4901,N_1681,N_220);
or U4902 (N_4902,N_2173,N_2614);
nand U4903 (N_4903,N_1960,N_3176);
or U4904 (N_4904,N_689,N_3417);
nand U4905 (N_4905,N_3178,N_1986);
xor U4906 (N_4906,N_1500,N_2759);
nand U4907 (N_4907,N_1758,N_3971);
nor U4908 (N_4908,N_3130,N_66);
nand U4909 (N_4909,N_810,N_574);
or U4910 (N_4910,N_2368,N_2262);
nand U4911 (N_4911,N_3191,N_2919);
nor U4912 (N_4912,N_359,N_872);
and U4913 (N_4913,N_3647,N_858);
nor U4914 (N_4914,N_3450,N_674);
nor U4915 (N_4915,N_1621,N_1532);
and U4916 (N_4916,N_925,N_95);
nor U4917 (N_4917,N_3935,N_3314);
nand U4918 (N_4918,N_2207,N_2219);
and U4919 (N_4919,N_3475,N_298);
or U4920 (N_4920,N_3629,N_471);
nand U4921 (N_4921,N_1043,N_871);
nor U4922 (N_4922,N_2965,N_3633);
or U4923 (N_4923,N_535,N_3526);
or U4924 (N_4924,N_695,N_1987);
or U4925 (N_4925,N_743,N_1432);
or U4926 (N_4926,N_2577,N_3941);
and U4927 (N_4927,N_1910,N_2132);
or U4928 (N_4928,N_2707,N_2729);
nand U4929 (N_4929,N_2935,N_2915);
or U4930 (N_4930,N_2612,N_2641);
nand U4931 (N_4931,N_63,N_254);
nand U4932 (N_4932,N_1486,N_1302);
nand U4933 (N_4933,N_579,N_1768);
or U4934 (N_4934,N_1083,N_655);
nor U4935 (N_4935,N_2927,N_3348);
nor U4936 (N_4936,N_1803,N_400);
and U4937 (N_4937,N_785,N_2664);
nand U4938 (N_4938,N_2814,N_1667);
and U4939 (N_4939,N_2768,N_1608);
and U4940 (N_4940,N_2936,N_3720);
nor U4941 (N_4941,N_1263,N_1241);
or U4942 (N_4942,N_2433,N_1580);
nand U4943 (N_4943,N_2369,N_128);
and U4944 (N_4944,N_2027,N_3014);
or U4945 (N_4945,N_2656,N_2912);
and U4946 (N_4946,N_2358,N_1887);
and U4947 (N_4947,N_1422,N_3190);
nor U4948 (N_4948,N_995,N_2714);
nand U4949 (N_4949,N_373,N_2792);
or U4950 (N_4950,N_99,N_813);
or U4951 (N_4951,N_327,N_101);
nand U4952 (N_4952,N_441,N_1466);
nand U4953 (N_4953,N_1011,N_1991);
and U4954 (N_4954,N_3600,N_3393);
or U4955 (N_4955,N_832,N_1658);
or U4956 (N_4956,N_1449,N_3311);
and U4957 (N_4957,N_2474,N_2172);
nand U4958 (N_4958,N_3885,N_2679);
or U4959 (N_4959,N_3370,N_2438);
nand U4960 (N_4960,N_2603,N_34);
nand U4961 (N_4961,N_2666,N_2520);
nor U4962 (N_4962,N_516,N_372);
nand U4963 (N_4963,N_3783,N_1864);
nand U4964 (N_4964,N_2994,N_2968);
nand U4965 (N_4965,N_2468,N_2543);
or U4966 (N_4966,N_3119,N_1413);
or U4967 (N_4967,N_290,N_1217);
nor U4968 (N_4968,N_922,N_3367);
and U4969 (N_4969,N_2504,N_199);
nor U4970 (N_4970,N_2091,N_1475);
and U4971 (N_4971,N_1411,N_149);
and U4972 (N_4972,N_473,N_1666);
and U4973 (N_4973,N_3061,N_1337);
nand U4974 (N_4974,N_2231,N_3853);
or U4975 (N_4975,N_3620,N_3447);
nand U4976 (N_4976,N_2244,N_2945);
and U4977 (N_4977,N_685,N_893);
nand U4978 (N_4978,N_1906,N_2393);
nand U4979 (N_4979,N_2408,N_1835);
or U4980 (N_4980,N_512,N_2270);
nor U4981 (N_4981,N_1784,N_3354);
nor U4982 (N_4982,N_3110,N_2816);
and U4983 (N_4983,N_2313,N_1142);
nand U4984 (N_4984,N_3085,N_3284);
nor U4985 (N_4985,N_1001,N_2902);
nand U4986 (N_4986,N_3938,N_2026);
nand U4987 (N_4987,N_3917,N_3565);
nor U4988 (N_4988,N_1541,N_1572);
or U4989 (N_4989,N_1026,N_3812);
or U4990 (N_4990,N_242,N_2568);
and U4991 (N_4991,N_3934,N_158);
and U4992 (N_4992,N_2843,N_3895);
or U4993 (N_4993,N_1928,N_1324);
or U4994 (N_4994,N_798,N_874);
nor U4995 (N_4995,N_869,N_2257);
nand U4996 (N_4996,N_1210,N_3530);
or U4997 (N_4997,N_3002,N_1582);
nand U4998 (N_4998,N_2049,N_849);
and U4999 (N_4999,N_2151,N_2479);
nor U5000 (N_5000,N_687,N_2776);
or U5001 (N_5001,N_601,N_3868);
and U5002 (N_5002,N_3759,N_3404);
or U5003 (N_5003,N_2054,N_3270);
nor U5004 (N_5004,N_753,N_2517);
or U5005 (N_5005,N_2873,N_1757);
and U5006 (N_5006,N_1051,N_2605);
nor U5007 (N_5007,N_2911,N_3461);
nand U5008 (N_5008,N_732,N_3124);
nand U5009 (N_5009,N_3289,N_219);
and U5010 (N_5010,N_1908,N_2092);
and U5011 (N_5011,N_541,N_3185);
and U5012 (N_5012,N_3628,N_2030);
nand U5013 (N_5013,N_3813,N_2872);
nand U5014 (N_5014,N_980,N_2898);
nor U5015 (N_5015,N_2828,N_990);
xnor U5016 (N_5016,N_1342,N_1955);
nor U5017 (N_5017,N_816,N_1896);
nand U5018 (N_5018,N_3087,N_1494);
nor U5019 (N_5019,N_265,N_2716);
nor U5020 (N_5020,N_1400,N_1636);
nand U5021 (N_5021,N_3758,N_3481);
or U5022 (N_5022,N_582,N_234);
nand U5023 (N_5023,N_499,N_2016);
or U5024 (N_5024,N_2573,N_3894);
nand U5025 (N_5025,N_1921,N_152);
or U5026 (N_5026,N_769,N_172);
nor U5027 (N_5027,N_3295,N_2839);
nor U5028 (N_5028,N_3034,N_2105);
and U5029 (N_5029,N_2371,N_864);
and U5030 (N_5030,N_2705,N_1762);
or U5031 (N_5031,N_2377,N_1978);
or U5032 (N_5032,N_2644,N_2548);
nor U5033 (N_5033,N_3229,N_1119);
and U5034 (N_5034,N_3590,N_176);
and U5035 (N_5035,N_2322,N_1090);
or U5036 (N_5036,N_2719,N_256);
and U5037 (N_5037,N_1198,N_3602);
nor U5038 (N_5038,N_1683,N_897);
or U5039 (N_5039,N_2111,N_3953);
nor U5040 (N_5040,N_3533,N_185);
or U5041 (N_5041,N_2749,N_3642);
and U5042 (N_5042,N_1932,N_2958);
xor U5043 (N_5043,N_397,N_921);
nand U5044 (N_5044,N_475,N_1376);
nor U5045 (N_5045,N_1868,N_1159);
nor U5046 (N_5046,N_331,N_1962);
nor U5047 (N_5047,N_1711,N_627);
nor U5048 (N_5048,N_3380,N_1461);
nand U5049 (N_5049,N_646,N_3547);
or U5050 (N_5050,N_1601,N_577);
nand U5051 (N_5051,N_763,N_2831);
or U5052 (N_5052,N_45,N_216);
nand U5053 (N_5053,N_2838,N_2356);
nor U5054 (N_5054,N_1779,N_2662);
and U5055 (N_5055,N_2249,N_2706);
or U5056 (N_5056,N_3670,N_14);
and U5057 (N_5057,N_138,N_1286);
nor U5058 (N_5058,N_3787,N_2174);
xor U5059 (N_5059,N_2323,N_3431);
nand U5060 (N_5060,N_2298,N_2882);
and U5061 (N_5061,N_2185,N_1348);
or U5062 (N_5062,N_2530,N_626);
nor U5063 (N_5063,N_1745,N_2602);
nand U5064 (N_5064,N_3984,N_3964);
nor U5065 (N_5065,N_2672,N_342);
nor U5066 (N_5066,N_1489,N_638);
or U5067 (N_5067,N_3912,N_2188);
and U5068 (N_5068,N_2328,N_1444);
and U5069 (N_5069,N_3368,N_388);
or U5070 (N_5070,N_3186,N_1390);
or U5071 (N_5071,N_451,N_1417);
and U5072 (N_5072,N_2502,N_896);
nor U5073 (N_5073,N_2415,N_3435);
nand U5074 (N_5074,N_3381,N_1792);
nand U5075 (N_5075,N_1927,N_100);
nand U5076 (N_5076,N_3215,N_3586);
and U5077 (N_5077,N_3467,N_985);
and U5078 (N_5078,N_614,N_1878);
or U5079 (N_5079,N_1894,N_1728);
nand U5080 (N_5080,N_2906,N_2042);
nor U5081 (N_5081,N_1581,N_2589);
nand U5082 (N_5082,N_2917,N_2388);
and U5083 (N_5083,N_752,N_2986);
nor U5084 (N_5084,N_3253,N_1537);
nor U5085 (N_5085,N_3744,N_2970);
nand U5086 (N_5086,N_3180,N_2689);
and U5087 (N_5087,N_2121,N_3837);
nand U5088 (N_5088,N_3529,N_1722);
nand U5089 (N_5089,N_2315,N_1956);
or U5090 (N_5090,N_850,N_1739);
and U5091 (N_5091,N_3582,N_262);
nor U5092 (N_5092,N_46,N_1015);
nor U5093 (N_5093,N_2404,N_973);
and U5094 (N_5094,N_51,N_2267);
nand U5095 (N_5095,N_2414,N_3279);
nand U5096 (N_5096,N_1408,N_3456);
and U5097 (N_5097,N_3212,N_79);
and U5098 (N_5098,N_2450,N_2940);
or U5099 (N_5099,N_511,N_1377);
or U5100 (N_5100,N_2829,N_815);
or U5101 (N_5101,N_3242,N_1856);
and U5102 (N_5102,N_2836,N_2864);
and U5103 (N_5103,N_2299,N_353);
and U5104 (N_5104,N_898,N_3689);
and U5105 (N_5105,N_3576,N_3555);
nor U5106 (N_5106,N_3408,N_2738);
or U5107 (N_5107,N_212,N_2250);
nand U5108 (N_5108,N_2048,N_3898);
and U5109 (N_5109,N_1357,N_2542);
nor U5110 (N_5110,N_1595,N_918);
nor U5111 (N_5111,N_2699,N_2340);
or U5112 (N_5112,N_719,N_1255);
xor U5113 (N_5113,N_2800,N_248);
or U5114 (N_5114,N_2779,N_1490);
nor U5115 (N_5115,N_38,N_3265);
nand U5116 (N_5116,N_1428,N_3115);
nor U5117 (N_5117,N_2611,N_1521);
nand U5118 (N_5118,N_3148,N_1108);
nor U5119 (N_5119,N_506,N_1685);
and U5120 (N_5120,N_141,N_190);
nand U5121 (N_5121,N_2149,N_2805);
or U5122 (N_5122,N_3942,N_2538);
nand U5123 (N_5123,N_1141,N_585);
and U5124 (N_5124,N_117,N_2663);
or U5125 (N_5125,N_3235,N_863);
or U5126 (N_5126,N_2437,N_1306);
or U5127 (N_5127,N_652,N_1079);
nor U5128 (N_5128,N_165,N_3414);
and U5129 (N_5129,N_276,N_2629);
nor U5130 (N_5130,N_2721,N_1016);
and U5131 (N_5131,N_3867,N_2115);
and U5132 (N_5132,N_2654,N_3834);
or U5133 (N_5133,N_1775,N_2252);
nor U5134 (N_5134,N_2681,N_3472);
and U5135 (N_5135,N_1761,N_136);
and U5136 (N_5136,N_1554,N_2941);
nor U5137 (N_5137,N_3460,N_3347);
nor U5138 (N_5138,N_3794,N_3650);
nand U5139 (N_5139,N_1640,N_2140);
and U5140 (N_5140,N_3815,N_2386);
and U5141 (N_5141,N_3278,N_3237);
or U5142 (N_5142,N_1346,N_2434);
nor U5143 (N_5143,N_3951,N_3655);
and U5144 (N_5144,N_2767,N_2248);
or U5145 (N_5145,N_2582,N_1551);
or U5146 (N_5146,N_3611,N_1387);
nand U5147 (N_5147,N_2199,N_909);
and U5148 (N_5148,N_3469,N_2452);
and U5149 (N_5149,N_3711,N_1207);
nor U5150 (N_5150,N_1190,N_2480);
and U5151 (N_5151,N_2337,N_2815);
nor U5152 (N_5152,N_2563,N_2006);
and U5153 (N_5153,N_1472,N_1840);
nor U5154 (N_5154,N_384,N_2218);
nand U5155 (N_5155,N_1248,N_3453);
nand U5156 (N_5156,N_3055,N_1189);
and U5157 (N_5157,N_2787,N_1945);
or U5158 (N_5158,N_332,N_2887);
or U5159 (N_5159,N_793,N_1913);
and U5160 (N_5160,N_1133,N_2300);
and U5161 (N_5161,N_3059,N_2794);
nor U5162 (N_5162,N_3309,N_1003);
nor U5163 (N_5163,N_118,N_1704);
nand U5164 (N_5164,N_3899,N_2855);
or U5165 (N_5165,N_808,N_2201);
nand U5166 (N_5166,N_2294,N_3695);
and U5167 (N_5167,N_1094,N_2630);
or U5168 (N_5168,N_2350,N_1295);
nand U5169 (N_5169,N_773,N_437);
and U5170 (N_5170,N_447,N_1354);
nor U5171 (N_5171,N_930,N_1355);
and U5172 (N_5172,N_2451,N_1968);
nand U5173 (N_5173,N_448,N_3132);
and U5174 (N_5174,N_3400,N_2537);
nor U5175 (N_5175,N_765,N_1446);
nor U5176 (N_5176,N_1797,N_1172);
nand U5177 (N_5177,N_3067,N_2933);
and U5178 (N_5178,N_3226,N_1984);
nand U5179 (N_5179,N_553,N_3771);
and U5180 (N_5180,N_3982,N_2803);
nand U5181 (N_5181,N_725,N_3777);
and U5182 (N_5182,N_2138,N_1882);
or U5183 (N_5183,N_1435,N_2953);
nand U5184 (N_5184,N_3692,N_2516);
nor U5185 (N_5185,N_3593,N_462);
and U5186 (N_5186,N_3827,N_1727);
or U5187 (N_5187,N_41,N_1895);
or U5188 (N_5188,N_2546,N_2731);
nand U5189 (N_5189,N_2073,N_3377);
nand U5190 (N_5190,N_3463,N_240);
and U5191 (N_5191,N_338,N_3816);
or U5192 (N_5192,N_1886,N_1700);
nor U5193 (N_5193,N_766,N_1807);
nor U5194 (N_5194,N_3747,N_284);
nand U5195 (N_5195,N_3901,N_2813);
or U5196 (N_5196,N_1318,N_2756);
nand U5197 (N_5197,N_3803,N_414);
nand U5198 (N_5198,N_2525,N_670);
nor U5199 (N_5199,N_2727,N_1607);
nand U5200 (N_5200,N_2539,N_2216);
and U5201 (N_5201,N_1418,N_2058);
or U5202 (N_5202,N_1478,N_29);
and U5203 (N_5203,N_3006,N_1186);
nand U5204 (N_5204,N_1069,N_1578);
and U5205 (N_5205,N_1,N_3232);
nand U5206 (N_5206,N_3718,N_2961);
nand U5207 (N_5207,N_3665,N_3287);
nand U5208 (N_5208,N_24,N_2695);
nor U5209 (N_5209,N_2407,N_321);
or U5210 (N_5210,N_2943,N_187);
and U5211 (N_5211,N_3911,N_1937);
and U5212 (N_5212,N_491,N_2292);
and U5213 (N_5213,N_1293,N_2471);
or U5214 (N_5214,N_3306,N_2126);
nand U5215 (N_5215,N_206,N_2177);
and U5216 (N_5216,N_2372,N_1360);
or U5217 (N_5217,N_371,N_2871);
and U5218 (N_5218,N_3281,N_607);
or U5219 (N_5219,N_560,N_266);
nor U5220 (N_5220,N_2397,N_2978);
nand U5221 (N_5221,N_98,N_3490);
nand U5222 (N_5222,N_201,N_2282);
nor U5223 (N_5223,N_2764,N_3926);
or U5224 (N_5224,N_1530,N_1880);
nor U5225 (N_5225,N_2744,N_1006);
nand U5226 (N_5226,N_1858,N_3862);
or U5227 (N_5227,N_3207,N_345);
nor U5228 (N_5228,N_3103,N_3350);
nand U5229 (N_5229,N_10,N_2928);
nor U5230 (N_5230,N_1372,N_975);
and U5231 (N_5231,N_405,N_2760);
and U5232 (N_5232,N_1409,N_2702);
nand U5233 (N_5233,N_48,N_3685);
or U5234 (N_5234,N_3523,N_1577);
nor U5235 (N_5235,N_226,N_988);
or U5236 (N_5236,N_1459,N_2098);
and U5237 (N_5237,N_1559,N_1152);
and U5238 (N_5238,N_3150,N_3328);
and U5239 (N_5239,N_967,N_3244);
or U5240 (N_5240,N_2318,N_2737);
or U5241 (N_5241,N_2487,N_1949);
or U5242 (N_5242,N_3750,N_1105);
nor U5243 (N_5243,N_2148,N_69);
or U5244 (N_5244,N_886,N_213);
or U5245 (N_5245,N_1817,N_146);
or U5246 (N_5246,N_1940,N_1661);
nand U5247 (N_5247,N_3292,N_147);
nor U5248 (N_5248,N_2179,N_3114);
nor U5249 (N_5249,N_3084,N_1135);
or U5250 (N_5250,N_3561,N_997);
or U5251 (N_5251,N_1603,N_3389);
or U5252 (N_5252,N_1884,N_3384);
nand U5253 (N_5253,N_1936,N_1744);
nor U5254 (N_5254,N_2044,N_570);
nor U5255 (N_5255,N_1923,N_153);
nand U5256 (N_5256,N_1787,N_778);
or U5257 (N_5257,N_672,N_2921);
and U5258 (N_5258,N_639,N_3677);
or U5259 (N_5259,N_450,N_2896);
or U5260 (N_5260,N_1035,N_1751);
or U5261 (N_5261,N_291,N_1179);
nand U5262 (N_5262,N_458,N_888);
nand U5263 (N_5263,N_1077,N_293);
nand U5264 (N_5264,N_151,N_3093);
or U5265 (N_5265,N_1294,N_1642);
and U5266 (N_5266,N_1780,N_3102);
nand U5267 (N_5267,N_2728,N_2089);
nand U5268 (N_5268,N_594,N_986);
or U5269 (N_5269,N_1027,N_2363);
or U5270 (N_5270,N_2200,N_3932);
nor U5271 (N_5271,N_776,N_1596);
or U5272 (N_5272,N_3060,N_1902);
and U5273 (N_5273,N_3635,N_1076);
nand U5274 (N_5274,N_90,N_314);
nand U5275 (N_5275,N_211,N_2688);
or U5276 (N_5276,N_1382,N_933);
and U5277 (N_5277,N_2798,N_1393);
nand U5278 (N_5278,N_3741,N_515);
or U5279 (N_5279,N_3534,N_3479);
nor U5280 (N_5280,N_2788,N_249);
and U5281 (N_5281,N_2754,N_260);
xnor U5282 (N_5282,N_2338,N_495);
or U5283 (N_5283,N_538,N_2189);
or U5284 (N_5284,N_2124,N_3621);
and U5285 (N_5285,N_977,N_72);
or U5286 (N_5286,N_2353,N_2099);
nor U5287 (N_5287,N_2922,N_566);
nor U5288 (N_5288,N_3608,N_628);
and U5289 (N_5289,N_1766,N_2901);
or U5290 (N_5290,N_1614,N_2293);
and U5291 (N_5291,N_222,N_3537);
nor U5292 (N_5292,N_1682,N_1972);
or U5293 (N_5293,N_1057,N_1163);
and U5294 (N_5294,N_3691,N_1983);
and U5295 (N_5295,N_855,N_1548);
and U5296 (N_5296,N_563,N_747);
and U5297 (N_5297,N_3846,N_2276);
or U5298 (N_5298,N_351,N_700);
nand U5299 (N_5299,N_740,N_3092);
or U5300 (N_5300,N_2982,N_3020);
nand U5301 (N_5301,N_1268,N_3480);
nand U5302 (N_5302,N_3603,N_3664);
nand U5303 (N_5303,N_243,N_1522);
and U5304 (N_5304,N_831,N_3301);
and U5305 (N_5305,N_843,N_1203);
nand U5306 (N_5306,N_2229,N_1465);
or U5307 (N_5307,N_3778,N_3793);
and U5308 (N_5308,N_3615,N_261);
nor U5309 (N_5309,N_233,N_319);
and U5310 (N_5310,N_1132,N_2523);
nand U5311 (N_5311,N_3411,N_214);
and U5312 (N_5312,N_3239,N_3667);
and U5313 (N_5313,N_3966,N_455);
nand U5314 (N_5314,N_2352,N_1615);
and U5315 (N_5315,N_64,N_2107);
nor U5316 (N_5316,N_3882,N_379);
or U5317 (N_5317,N_3599,N_273);
or U5318 (N_5318,N_981,N_3597);
and U5319 (N_5319,N_333,N_2106);
and U5320 (N_5320,N_3646,N_2097);
nor U5321 (N_5321,N_1086,N_1150);
and U5322 (N_5322,N_1073,N_2975);
or U5323 (N_5323,N_2012,N_3058);
nor U5324 (N_5324,N_809,N_1038);
and U5325 (N_5325,N_2963,N_3959);
or U5326 (N_5326,N_3859,N_941);
and U5327 (N_5327,N_3944,N_684);
and U5328 (N_5328,N_3052,N_1926);
or U5329 (N_5329,N_2223,N_2635);
or U5330 (N_5330,N_2597,N_3352);
nor U5331 (N_5331,N_486,N_19);
nor U5332 (N_5332,N_1924,N_1891);
nor U5333 (N_5333,N_3907,N_3728);
or U5334 (N_5334,N_3955,N_3388);
or U5335 (N_5335,N_540,N_3399);
nand U5336 (N_5336,N_3095,N_97);
and U5337 (N_5337,N_572,N_2454);
nand U5338 (N_5338,N_2846,N_78);
or U5339 (N_5339,N_1922,N_3601);
and U5340 (N_5340,N_2802,N_3153);
or U5341 (N_5341,N_1368,N_1684);
nor U5342 (N_5342,N_2765,N_1430);
and U5343 (N_5343,N_2351,N_575);
or U5344 (N_5344,N_779,N_3699);
and U5345 (N_5345,N_3036,N_3658);
or U5346 (N_5346,N_962,N_1487);
nand U5347 (N_5347,N_3631,N_3426);
nand U5348 (N_5348,N_527,N_3887);
nand U5349 (N_5349,N_2890,N_2512);
and U5350 (N_5350,N_3903,N_861);
nand U5351 (N_5351,N_2296,N_3465);
nand U5352 (N_5352,N_389,N_299);
or U5353 (N_5353,N_842,N_1398);
and U5354 (N_5354,N_1385,N_1240);
or U5355 (N_5355,N_3294,N_1423);
nor U5356 (N_5356,N_772,N_680);
nand U5357 (N_5357,N_2509,N_1215);
or U5358 (N_5358,N_3086,N_3616);
nor U5359 (N_5359,N_3763,N_354);
nand U5360 (N_5360,N_1623,N_2123);
and U5361 (N_5361,N_3886,N_3807);
and U5362 (N_5362,N_2569,N_3854);
nand U5363 (N_5363,N_492,N_2880);
or U5364 (N_5364,N_318,N_2842);
or U5365 (N_5365,N_2752,N_2645);
nor U5366 (N_5366,N_2799,N_1134);
nand U5367 (N_5367,N_824,N_237);
and U5368 (N_5368,N_3768,N_1497);
xor U5369 (N_5369,N_949,N_876);
or U5370 (N_5370,N_180,N_1092);
or U5371 (N_5371,N_3495,N_1386);
or U5372 (N_5372,N_1378,N_3525);
nor U5373 (N_5373,N_2291,N_797);
nand U5374 (N_5374,N_2425,N_2157);
or U5375 (N_5375,N_3660,N_2137);
and U5376 (N_5376,N_3198,N_1365);
or U5377 (N_5377,N_1196,N_817);
nand U5378 (N_5378,N_23,N_3254);
or U5379 (N_5379,N_2028,N_1427);
nand U5380 (N_5380,N_1220,N_1405);
nand U5381 (N_5381,N_3798,N_2074);
nor U5382 (N_5382,N_2827,N_200);
nand U5383 (N_5383,N_3776,N_1272);
nor U5384 (N_5384,N_3410,N_705);
or U5385 (N_5385,N_1904,N_3250);
nand U5386 (N_5386,N_3351,N_3362);
nor U5387 (N_5387,N_3407,N_340);
and U5388 (N_5388,N_900,N_1261);
nor U5389 (N_5389,N_1627,N_1367);
and U5390 (N_5390,N_3160,N_1988);
and U5391 (N_5391,N_688,N_3861);
or U5392 (N_5392,N_3147,N_961);
nor U5393 (N_5393,N_2336,N_3356);
nor U5394 (N_5394,N_1653,N_2210);
and U5395 (N_5395,N_1336,N_1238);
nor U5396 (N_5396,N_818,N_3856);
nand U5397 (N_5397,N_537,N_145);
and U5398 (N_5398,N_1767,N_3015);
nand U5399 (N_5399,N_315,N_1309);
nand U5400 (N_5400,N_603,N_662);
xor U5401 (N_5401,N_2349,N_760);
nand U5402 (N_5402,N_2742,N_3213);
and U5403 (N_5403,N_878,N_2110);
nor U5404 (N_5404,N_885,N_3906);
and U5405 (N_5405,N_62,N_3146);
nand U5406 (N_5406,N_1304,N_1688);
nand U5407 (N_5407,N_984,N_3144);
and U5408 (N_5408,N_3300,N_406);
nor U5409 (N_5409,N_2014,N_3562);
or U5410 (N_5410,N_456,N_1543);
and U5411 (N_5411,N_3194,N_1269);
and U5412 (N_5412,N_3157,N_1331);
or U5413 (N_5413,N_3575,N_12);
xnor U5414 (N_5414,N_669,N_3487);
or U5415 (N_5415,N_306,N_2650);
or U5416 (N_5416,N_3468,N_2008);
and U5417 (N_5417,N_2424,N_671);
nor U5418 (N_5418,N_1194,N_1464);
and U5419 (N_5419,N_935,N_1010);
nand U5420 (N_5420,N_1054,N_65);
nand U5421 (N_5421,N_2743,N_3684);
and U5422 (N_5422,N_3090,N_3168);
nor U5423 (N_5423,N_104,N_2198);
nand U5424 (N_5424,N_2492,N_36);
nor U5425 (N_5425,N_1311,N_2379);
nor U5426 (N_5426,N_758,N_623);
and U5427 (N_5427,N_156,N_3551);
or U5428 (N_5428,N_445,N_1730);
nand U5429 (N_5429,N_510,N_3439);
or U5430 (N_5430,N_1145,N_3990);
or U5431 (N_5431,N_1524,N_3188);
or U5432 (N_5432,N_974,N_771);
nand U5433 (N_5433,N_3829,N_3155);
nand U5434 (N_5434,N_3543,N_3081);
nand U5435 (N_5435,N_3574,N_3027);
nor U5436 (N_5436,N_3297,N_1002);
nand U5437 (N_5437,N_43,N_3881);
nor U5438 (N_5438,N_1020,N_3998);
or U5439 (N_5439,N_690,N_2929);
nand U5440 (N_5440,N_417,N_3810);
or U5441 (N_5441,N_2518,N_2735);
or U5442 (N_5442,N_1925,N_1320);
and U5443 (N_5443,N_3360,N_3542);
or U5444 (N_5444,N_2122,N_600);
nor U5445 (N_5445,N_3950,N_3618);
nand U5446 (N_5446,N_2022,N_3214);
and U5447 (N_5447,N_2152,N_1866);
nand U5448 (N_5448,N_782,N_657);
and U5449 (N_5449,N_2076,N_1301);
or U5450 (N_5450,N_2465,N_1641);
and U5451 (N_5451,N_3992,N_3904);
and U5452 (N_5452,N_3513,N_3449);
nor U5453 (N_5453,N_1178,N_3228);
nand U5454 (N_5454,N_2242,N_2877);
or U5455 (N_5455,N_792,N_334);
and U5456 (N_5456,N_2909,N_3201);
or U5457 (N_5457,N_605,N_1552);
and U5458 (N_5458,N_3080,N_615);
nor U5459 (N_5459,N_3567,N_1777);
and U5460 (N_5460,N_1724,N_1162);
and U5461 (N_5461,N_209,N_1563);
or U5462 (N_5462,N_322,N_2857);
nor U5463 (N_5463,N_2285,N_3657);
and U5464 (N_5464,N_2682,N_3187);
nor U5465 (N_5465,N_1934,N_534);
and U5466 (N_5466,N_3610,N_3057);
and U5467 (N_5467,N_1699,N_3070);
nor U5468 (N_5468,N_1389,N_2999);
nand U5469 (N_5469,N_2845,N_1812);
xnor U5470 (N_5470,N_268,N_723);
and U5471 (N_5471,N_3943,N_3066);
nor U5472 (N_5472,N_1022,N_1326);
nor U5473 (N_5473,N_3790,N_2490);
nor U5474 (N_5474,N_1158,N_2317);
or U5475 (N_5475,N_822,N_2041);
and U5476 (N_5476,N_3434,N_1281);
nand U5477 (N_5477,N_865,N_163);
nand U5478 (N_5478,N_2439,N_1095);
nand U5479 (N_5479,N_40,N_3580);
and U5480 (N_5480,N_2236,N_3280);
and U5481 (N_5481,N_3152,N_1873);
nand U5482 (N_5482,N_3579,N_3182);
and U5483 (N_5483,N_767,N_948);
and U5484 (N_5484,N_1296,N_1253);
or U5485 (N_5485,N_3681,N_2730);
or U5486 (N_5486,N_3596,N_2510);
nand U5487 (N_5487,N_1723,N_1462);
and U5488 (N_5488,N_978,N_3527);
and U5489 (N_5489,N_2212,N_1341);
and U5490 (N_5490,N_3316,N_2748);
nand U5491 (N_5491,N_2711,N_2607);
and U5492 (N_5492,N_3332,N_317);
nand U5493 (N_5493,N_811,N_1799);
nand U5494 (N_5494,N_3900,N_2225);
and U5495 (N_5495,N_1282,N_382);
nor U5496 (N_5496,N_1731,N_823);
or U5497 (N_5497,N_517,N_989);
nor U5498 (N_5498,N_3501,N_3835);
and U5499 (N_5499,N_2826,N_2822);
nor U5500 (N_5500,N_2948,N_1287);
or U5501 (N_5501,N_1008,N_803);
nor U5502 (N_5502,N_3116,N_459);
nor U5503 (N_5503,N_2559,N_1617);
or U5504 (N_5504,N_667,N_2275);
nor U5505 (N_5505,N_489,N_1860);
nor U5506 (N_5506,N_1013,N_1144);
or U5507 (N_5507,N_2489,N_3948);
or U5508 (N_5508,N_3041,N_2676);
or U5509 (N_5509,N_3062,N_620);
or U5510 (N_5510,N_2021,N_3126);
nand U5511 (N_5511,N_911,N_1120);
or U5512 (N_5512,N_2303,N_2406);
and U5513 (N_5513,N_1584,N_1081);
or U5514 (N_5514,N_1911,N_2083);
nand U5515 (N_5515,N_3855,N_3498);
or U5516 (N_5516,N_1954,N_204);
nor U5517 (N_5517,N_3705,N_1089);
nand U5518 (N_5518,N_37,N_22);
and U5519 (N_5519,N_3342,N_192);
and U5520 (N_5520,N_2429,N_1087);
and U5521 (N_5521,N_710,N_825);
nor U5522 (N_5522,N_358,N_1527);
and U5523 (N_5523,N_3446,N_123);
nor U5524 (N_5524,N_2686,N_1406);
or U5525 (N_5525,N_1966,N_2130);
or U5526 (N_5526,N_2494,N_3808);
and U5527 (N_5527,N_1244,N_1161);
nor U5528 (N_5528,N_530,N_2966);
xnor U5529 (N_5529,N_1846,N_1155);
nor U5530 (N_5530,N_1333,N_675);
nor U5531 (N_5531,N_3135,N_3991);
nand U5532 (N_5532,N_323,N_629);
nand U5533 (N_5533,N_2327,N_2175);
nand U5534 (N_5534,N_2183,N_1898);
and U5535 (N_5535,N_1841,N_3544);
and U5536 (N_5536,N_228,N_3409);
nor U5537 (N_5537,N_1493,N_3940);
nand U5538 (N_5538,N_2,N_2184);
or U5539 (N_5539,N_2678,N_2204);
and U5540 (N_5540,N_2169,N_1998);
and U5541 (N_5541,N_1061,N_2817);
or U5542 (N_5542,N_1111,N_1305);
or U5543 (N_5543,N_3566,N_1825);
or U5544 (N_5544,N_1957,N_2657);
nor U5545 (N_5545,N_1971,N_3262);
nor U5546 (N_5546,N_215,N_731);
or U5547 (N_5547,N_2925,N_2875);
and U5548 (N_5548,N_1542,N_2691);
and U5549 (N_5549,N_543,N_2619);
or U5550 (N_5550,N_2895,N_449);
nor U5551 (N_5551,N_9,N_979);
nand U5552 (N_5552,N_2035,N_1585);
or U5553 (N_5553,N_2400,N_2129);
and U5554 (N_5554,N_2544,N_561);
nand U5555 (N_5555,N_3735,N_3824);
nand U5556 (N_5556,N_3719,N_2578);
or U5557 (N_5557,N_697,N_3809);
nor U5558 (N_5558,N_2519,N_3572);
nor U5559 (N_5559,N_1229,N_453);
nand U5560 (N_5560,N_1890,N_992);
and U5561 (N_5561,N_2381,N_1074);
nor U5562 (N_5562,N_3893,N_264);
xnor U5563 (N_5563,N_302,N_478);
or U5564 (N_5564,N_568,N_1289);
or U5565 (N_5565,N_3143,N_1151);
or U5566 (N_5566,N_3765,N_3785);
or U5567 (N_5567,N_1942,N_2806);
or U5568 (N_5568,N_461,N_3598);
and U5569 (N_5569,N_3742,N_2531);
nand U5570 (N_5570,N_1600,N_1499);
or U5571 (N_5571,N_665,N_618);
nand U5572 (N_5572,N_1146,N_2534);
nor U5573 (N_5573,N_2096,N_3958);
nand U5574 (N_5574,N_1118,N_183);
and U5575 (N_5575,N_73,N_1278);
and U5576 (N_5576,N_272,N_3401);
or U5577 (N_5577,N_160,N_2301);
nand U5578 (N_5578,N_1066,N_1204);
or U5579 (N_5579,N_1279,N_1629);
and U5580 (N_5580,N_709,N_2562);
nor U5581 (N_5581,N_2983,N_2807);
nand U5582 (N_5582,N_2739,N_2745);
nand U5583 (N_5583,N_2496,N_1224);
or U5584 (N_5584,N_1708,N_2950);
nor U5585 (N_5585,N_1526,N_1686);
nor U5586 (N_5586,N_1852,N_683);
nand U5587 (N_5587,N_3283,N_845);
and U5588 (N_5588,N_3673,N_589);
nor U5589 (N_5589,N_503,N_3247);
or U5590 (N_5590,N_2595,N_507);
or U5591 (N_5591,N_3231,N_2642);
nor U5592 (N_5592,N_2549,N_1211);
nor U5593 (N_5593,N_668,N_3724);
nor U5594 (N_5594,N_2367,N_3977);
nand U5595 (N_5595,N_3021,N_3406);
or U5596 (N_5596,N_2865,N_525);
nand U5597 (N_5597,N_547,N_3836);
nor U5598 (N_5598,N_923,N_1338);
or U5599 (N_5599,N_2648,N_2392);
or U5600 (N_5600,N_1979,N_1838);
nand U5601 (N_5601,N_2653,N_415);
nor U5602 (N_5602,N_546,N_352);
or U5603 (N_5603,N_103,N_632);
nand U5604 (N_5604,N_33,N_292);
nor U5605 (N_5605,N_3068,N_1399);
or U5606 (N_5606,N_1958,N_2470);
nand U5607 (N_5607,N_1380,N_2655);
nor U5608 (N_5608,N_951,N_2904);
or U5609 (N_5609,N_3550,N_2466);
nor U5610 (N_5610,N_3591,N_116);
or U5611 (N_5611,N_1075,N_3832);
nand U5612 (N_5612,N_2617,N_2310);
and U5613 (N_5613,N_3094,N_2284);
nand U5614 (N_5614,N_2341,N_2069);
and U5615 (N_5615,N_2273,N_2529);
nand U5616 (N_5616,N_2266,N_2514);
nand U5617 (N_5617,N_3999,N_1351);
and U5618 (N_5618,N_1943,N_2675);
nand U5619 (N_5619,N_1153,N_1562);
and U5620 (N_5620,N_707,N_2080);
nor U5621 (N_5621,N_812,N_3531);
nor U5622 (N_5622,N_422,N_1950);
nand U5623 (N_5623,N_557,N_1014);
and U5624 (N_5624,N_3412,N_3770);
nand U5625 (N_5625,N_3440,N_1276);
or U5626 (N_5626,N_2309,N_3825);
nor U5627 (N_5627,N_1674,N_2176);
nand U5628 (N_5628,N_3729,N_3224);
or U5629 (N_5629,N_1769,N_2646);
or U5630 (N_5630,N_32,N_666);
or U5631 (N_5631,N_3796,N_2835);
or U5632 (N_5632,N_2660,N_2580);
nand U5633 (N_5633,N_392,N_934);
or U5634 (N_5634,N_635,N_498);
nor U5635 (N_5635,N_2820,N_3569);
nand U5636 (N_5636,N_643,N_2633);
nor U5637 (N_5637,N_1544,N_3652);
and U5638 (N_5638,N_356,N_3732);
nor U5639 (N_5639,N_3494,N_726);
and U5640 (N_5640,N_3703,N_2135);
or U5641 (N_5641,N_3117,N_134);
or U5642 (N_5642,N_1877,N_3619);
nand U5643 (N_5643,N_1952,N_1961);
nand U5644 (N_5644,N_1909,N_3722);
nor U5645 (N_5645,N_1697,N_960);
nor U5646 (N_5646,N_3678,N_1112);
nor U5647 (N_5647,N_55,N_2258);
nor U5648 (N_5648,N_2162,N_2618);
nand U5649 (N_5649,N_381,N_2598);
nand U5650 (N_5650,N_2649,N_3392);
nor U5651 (N_5651,N_2647,N_2867);
nand U5652 (N_5652,N_2781,N_3792);
and U5653 (N_5653,N_362,N_3256);
nor U5654 (N_5654,N_3396,N_2478);
or U5655 (N_5655,N_637,N_2375);
nand U5656 (N_5656,N_311,N_1571);
nand U5657 (N_5657,N_2401,N_1082);
nor U5658 (N_5658,N_1453,N_3663);
or U5659 (N_5659,N_1303,N_1774);
nand U5660 (N_5660,N_3303,N_1232);
nand U5661 (N_5661,N_1410,N_81);
nand U5662 (N_5662,N_403,N_1201);
nor U5663 (N_5663,N_913,N_737);
and U5664 (N_5664,N_1271,N_2226);
nor U5665 (N_5665,N_3046,N_1772);
or U5666 (N_5666,N_1088,N_2399);
nand U5667 (N_5667,N_1050,N_1436);
and U5668 (N_5668,N_1068,N_1742);
or U5669 (N_5669,N_3324,N_3427);
nand U5670 (N_5670,N_1660,N_2840);
or U5671 (N_5671,N_1007,N_3230);
or U5672 (N_5672,N_2718,N_2622);
or U5673 (N_5673,N_3065,N_1919);
nor U5674 (N_5674,N_2910,N_1407);
nor U5675 (N_5675,N_2193,N_393);
and U5676 (N_5676,N_2190,N_3413);
and U5677 (N_5677,N_2304,N_1639);
nor U5678 (N_5678,N_3528,N_693);
or U5679 (N_5679,N_2467,N_2202);
or U5680 (N_5680,N_3571,N_1160);
or U5681 (N_5681,N_127,N_1169);
nand U5682 (N_5682,N_2031,N_440);
nor U5683 (N_5683,N_2246,N_1569);
nand U5684 (N_5684,N_2181,N_3975);
or U5685 (N_5685,N_866,N_2472);
nor U5686 (N_5686,N_3483,N_1712);
nor U5687 (N_5687,N_3397,N_2639);
nand U5688 (N_5688,N_1726,N_3656);
nand U5689 (N_5689,N_1785,N_1654);
nor U5690 (N_5690,N_179,N_1345);
and U5691 (N_5691,N_182,N_3996);
nand U5692 (N_5692,N_1307,N_3756);
and U5693 (N_5693,N_3263,N_851);
or U5694 (N_5694,N_3902,N_3238);
nor U5695 (N_5695,N_3721,N_698);
and U5696 (N_5696,N_1634,N_1037);
nand U5697 (N_5697,N_2029,N_3418);
nand U5698 (N_5698,N_2579,N_936);
nor U5699 (N_5699,N_25,N_3);
nor U5700 (N_5700,N_1754,N_706);
nand U5701 (N_5701,N_3459,N_56);
nand U5702 (N_5702,N_3252,N_2811);
nor U5703 (N_5703,N_2942,N_2930);
nand U5704 (N_5704,N_2394,N_3013);
and U5705 (N_5705,N_3420,N_3045);
nand U5706 (N_5706,N_2770,N_1474);
and U5707 (N_5707,N_169,N_18);
nand U5708 (N_5708,N_1371,N_443);
nor U5709 (N_5709,N_2632,N_2347);
and U5710 (N_5710,N_3640,N_573);
nand U5711 (N_5711,N_1951,N_907);
nand U5712 (N_5712,N_1914,N_1443);
nor U5713 (N_5713,N_3344,N_1175);
or U5714 (N_5714,N_3285,N_1718);
nor U5715 (N_5715,N_218,N_591);
nor U5716 (N_5716,N_3173,N_1735);
nor U5717 (N_5717,N_882,N_3145);
nor U5718 (N_5718,N_1819,N_53);
and U5719 (N_5719,N_870,N_3986);
and U5720 (N_5720,N_1259,N_783);
or U5721 (N_5721,N_1412,N_1113);
nor U5722 (N_5722,N_1212,N_519);
and U5723 (N_5723,N_407,N_1816);
or U5724 (N_5724,N_2995,N_383);
and U5725 (N_5725,N_1698,N_1941);
nor U5726 (N_5726,N_84,N_2378);
and U5727 (N_5727,N_1221,N_1930);
nand U5728 (N_5728,N_770,N_3624);
nor U5729 (N_5729,N_3112,N_1876);
nand U5730 (N_5730,N_2213,N_2773);
nand U5731 (N_5731,N_1334,N_3838);
nor U5732 (N_5732,N_2638,N_1030);
nand U5733 (N_5733,N_2624,N_1496);
or U5734 (N_5734,N_1513,N_3921);
or U5735 (N_5735,N_1488,N_634);
or U5736 (N_5736,N_1821,N_1370);
and U5737 (N_5737,N_3293,N_500);
and U5738 (N_5738,N_1970,N_640);
or U5739 (N_5739,N_2881,N_251);
or U5740 (N_5740,N_3366,N_1383);
and U5741 (N_5741,N_609,N_1485);
and U5742 (N_5742,N_1635,N_2899);
nand U5743 (N_5743,N_2036,N_2085);
nand U5744 (N_5744,N_2228,N_3385);
nand U5745 (N_5745,N_2821,N_27);
or U5746 (N_5746,N_3607,N_727);
nor U5747 (N_5747,N_3079,N_3074);
and U5748 (N_5748,N_3559,N_3325);
and U5749 (N_5749,N_349,N_20);
nand U5750 (N_5750,N_2851,N_1424);
and U5751 (N_5751,N_235,N_61);
or U5752 (N_5752,N_2720,N_780);
and U5753 (N_5753,N_2380,N_1167);
nor U5754 (N_5754,N_2224,N_2413);
nor U5755 (N_5755,N_2297,N_3733);
and U5756 (N_5756,N_1280,N_1328);
and U5757 (N_5757,N_1102,N_3891);
and U5758 (N_5758,N_3743,N_1266);
and U5759 (N_5759,N_3004,N_1786);
nand U5760 (N_5760,N_3517,N_3243);
nand U5761 (N_5761,N_2064,N_3023);
nand U5762 (N_5762,N_1549,N_3823);
and U5763 (N_5763,N_1538,N_47);
and U5764 (N_5764,N_3333,N_1239);
and U5765 (N_5765,N_2485,N_2625);
nand U5766 (N_5766,N_2289,N_3246);
nor U5767 (N_5767,N_633,N_1589);
nor U5768 (N_5768,N_826,N_1225);
nand U5769 (N_5769,N_1655,N_2150);
nor U5770 (N_5770,N_1593,N_2255);
nand U5771 (N_5771,N_2550,N_2522);
nand U5772 (N_5772,N_1750,N_1504);
or U5773 (N_5773,N_255,N_2384);
nand U5774 (N_5774,N_983,N_1862);
and U5775 (N_5775,N_223,N_3040);
nor U5776 (N_5776,N_1434,N_569);
nand U5777 (N_5777,N_230,N_1188);
and U5778 (N_5778,N_2751,N_873);
and U5779 (N_5779,N_3154,N_1903);
nor U5780 (N_5780,N_328,N_3731);
nand U5781 (N_5781,N_2312,N_649);
nor U5782 (N_5782,N_729,N_2043);
or U5783 (N_5783,N_2962,N_1707);
and U5784 (N_5784,N_205,N_2055);
nor U5785 (N_5785,N_3204,N_2592);
nor U5786 (N_5786,N_1310,N_159);
nor U5787 (N_5787,N_231,N_2039);
nand U5788 (N_5788,N_952,N_3779);
or U5789 (N_5789,N_2112,N_3502);
or U5790 (N_5790,N_2690,N_1184);
nand U5791 (N_5791,N_1174,N_132);
or U5792 (N_5792,N_3016,N_3142);
nor U5793 (N_5793,N_788,N_1893);
or U5794 (N_5794,N_129,N_2847);
nand U5795 (N_5795,N_2668,N_452);
nand U5796 (N_5796,N_596,N_3222);
or U5797 (N_5797,N_919,N_3454);
or U5798 (N_5798,N_308,N_3223);
and U5799 (N_5799,N_1691,N_229);
nor U5800 (N_5800,N_3696,N_950);
and U5801 (N_5801,N_3038,N_548);
nor U5802 (N_5802,N_2278,N_526);
and U5803 (N_5803,N_3970,N_3444);
nand U5804 (N_5804,N_2696,N_1618);
and U5805 (N_5805,N_2033,N_2324);
or U5806 (N_5806,N_2671,N_1106);
nand U5807 (N_5807,N_1592,N_714);
nor U5808 (N_5808,N_408,N_3088);
or U5809 (N_5809,N_2264,N_3302);
or U5810 (N_5810,N_2992,N_3120);
nor U5811 (N_5811,N_1881,N_3003);
nand U5812 (N_5812,N_1933,N_1156);
or U5813 (N_5813,N_764,N_270);
or U5814 (N_5814,N_1915,N_210);
nand U5815 (N_5815,N_844,N_998);
or U5816 (N_5816,N_2498,N_3429);
nand U5817 (N_5817,N_1299,N_994);
and U5818 (N_5818,N_3035,N_796);
or U5819 (N_5819,N_1213,N_139);
nand U5820 (N_5820,N_1243,N_2916);
or U5821 (N_5821,N_1644,N_1671);
nor U5822 (N_5822,N_3000,N_884);
nand U5823 (N_5823,N_350,N_3386);
and U5824 (N_5824,N_1256,N_1558);
or U5825 (N_5825,N_2862,N_839);
or U5826 (N_5826,N_2263,N_3099);
nand U5827 (N_5827,N_2197,N_703);
or U5828 (N_5828,N_2233,N_1773);
or U5829 (N_5829,N_571,N_2018);
nor U5830 (N_5830,N_1836,N_814);
or U5831 (N_5831,N_3687,N_1363);
nor U5832 (N_5832,N_1319,N_2260);
nand U5833 (N_5833,N_1055,N_3249);
nand U5834 (N_5834,N_106,N_2020);
and U5835 (N_5835,N_3974,N_3101);
and U5836 (N_5836,N_2280,N_3754);
nand U5837 (N_5837,N_3889,N_3826);
and U5838 (N_5838,N_1170,N_2949);
nor U5839 (N_5839,N_3701,N_1964);
nor U5840 (N_5840,N_181,N_1693);
nand U5841 (N_5841,N_1308,N_531);
or U5842 (N_5842,N_335,N_1353);
and U5843 (N_5843,N_682,N_3536);
or U5844 (N_5844,N_2448,N_2240);
or U5845 (N_5845,N_1379,N_1034);
nor U5846 (N_5846,N_1736,N_2037);
and U5847 (N_5847,N_1012,N_410);
nor U5848 (N_5848,N_122,N_154);
or U5849 (N_5849,N_533,N_3937);
nand U5850 (N_5850,N_3557,N_1103);
nor U5851 (N_5851,N_3248,N_3415);
or U5852 (N_5852,N_1782,N_821);
nand U5853 (N_5853,N_1839,N_289);
nand U5854 (N_5854,N_1361,N_2797);
nand U5855 (N_5855,N_1505,N_2354);
nand U5856 (N_5856,N_1539,N_295);
or U5857 (N_5857,N_1477,N_781);
nor U5858 (N_5858,N_1801,N_2456);
nor U5859 (N_5859,N_2117,N_3522);
and U5860 (N_5860,N_3233,N_836);
and U5861 (N_5861,N_1104,N_2187);
and U5862 (N_5862,N_3725,N_558);
or U5863 (N_5863,N_357,N_3679);
nand U5864 (N_5864,N_1678,N_3128);
and U5865 (N_5865,N_1974,N_636);
and U5866 (N_5866,N_1533,N_2477);
nor U5867 (N_5867,N_1091,N_755);
and U5868 (N_5868,N_300,N_1680);
or U5869 (N_5869,N_1832,N_1657);
nand U5870 (N_5870,N_3398,N_3614);
nor U5871 (N_5871,N_2704,N_616);
nor U5872 (N_5872,N_2723,N_1874);
or U5873 (N_5873,N_3764,N_59);
or U5874 (N_5874,N_2261,N_1491);
or U5875 (N_5875,N_3123,N_1339);
nor U5876 (N_5876,N_166,N_892);
and U5877 (N_5877,N_2013,N_702);
nand U5878 (N_5878,N_1445,N_1352);
or U5879 (N_5879,N_2435,N_2540);
or U5880 (N_5880,N_942,N_2879);
nand U5881 (N_5881,N_3196,N_1048);
nor U5882 (N_5882,N_744,N_3888);
or U5883 (N_5883,N_2446,N_3462);
or U5884 (N_5884,N_1981,N_3507);
nand U5885 (N_5885,N_647,N_2601);
and U5886 (N_5886,N_2609,N_648);
or U5887 (N_5887,N_2086,N_1182);
or U5888 (N_5888,N_3245,N_167);
or U5889 (N_5889,N_2410,N_1811);
nor U5890 (N_5890,N_87,N_67);
or U5891 (N_5891,N_1344,N_2141);
nand U5892 (N_5892,N_1706,N_2824);
and U5893 (N_5893,N_91,N_3338);
or U5894 (N_5894,N_751,N_1716);
or U5895 (N_5895,N_3009,N_3290);
and U5896 (N_5896,N_2859,N_581);
or U5897 (N_5897,N_3272,N_943);
and U5898 (N_5898,N_1072,N_3736);
nor U5899 (N_5899,N_2947,N_80);
and U5900 (N_5900,N_1771,N_2626);
nand U5901 (N_5901,N_1507,N_708);
and U5902 (N_5902,N_16,N_2453);
or U5903 (N_5903,N_848,N_908);
nand U5904 (N_5904,N_673,N_133);
nand U5905 (N_5905,N_2724,N_257);
nand U5906 (N_5906,N_3167,N_2063);
and U5907 (N_5907,N_1791,N_2460);
nand U5908 (N_5908,N_1804,N_325);
nand U5909 (N_5909,N_2784,N_267);
nor U5910 (N_5910,N_799,N_847);
nand U5911 (N_5911,N_3680,N_3662);
nor U5912 (N_5912,N_2295,N_2343);
or U5913 (N_5913,N_3225,N_3203);
or U5914 (N_5914,N_460,N_2710);
nand U5915 (N_5915,N_3221,N_840);
or U5916 (N_5916,N_2093,N_2254);
nand U5917 (N_5917,N_2109,N_1402);
nand U5918 (N_5918,N_2387,N_2651);
and U5919 (N_5919,N_3331,N_2808);
nand U5920 (N_5920,N_3844,N_2844);
and U5921 (N_5921,N_3666,N_904);
nand U5922 (N_5922,N_105,N_419);
nand U5923 (N_5923,N_3927,N_3626);
and U5924 (N_5924,N_3924,N_2850);
and U5925 (N_5925,N_3595,N_263);
nand U5926 (N_5926,N_68,N_259);
and U5927 (N_5927,N_3269,N_161);
nor U5928 (N_5928,N_3310,N_3548);
or U5929 (N_5929,N_1620,N_2698);
nor U5930 (N_5930,N_953,N_2769);
or U5931 (N_5931,N_774,N_3082);
or U5932 (N_5932,N_830,N_1994);
nor U5933 (N_5933,N_3963,N_3171);
nor U5934 (N_5934,N_3478,N_464);
nand U5935 (N_5935,N_2488,N_3636);
nand U5936 (N_5936,N_1523,N_3672);
and U5937 (N_5937,N_3258,N_2145);
nor U5938 (N_5938,N_1358,N_2457);
nor U5939 (N_5939,N_1005,N_3804);
nor U5940 (N_5940,N_514,N_1080);
nor U5941 (N_5941,N_1929,N_398);
or U5942 (N_5942,N_225,N_1093);
nand U5943 (N_5943,N_3097,N_3643);
or U5944 (N_5944,N_3149,N_2659);
xnor U5945 (N_5945,N_2023,N_1284);
nand U5946 (N_5946,N_1233,N_1556);
nand U5947 (N_5947,N_85,N_197);
nand U5948 (N_5948,N_207,N_2038);
and U5949 (N_5949,N_1171,N_3161);
or U5950 (N_5950,N_1793,N_1883);
nand U5951 (N_5951,N_926,N_3260);
or U5952 (N_5952,N_2056,N_301);
and U5953 (N_5953,N_3276,N_1117);
or U5954 (N_5954,N_2066,N_2403);
or U5955 (N_5955,N_562,N_2382);
and U5956 (N_5956,N_555,N_286);
and U5957 (N_5957,N_3801,N_3521);
nand U5958 (N_5958,N_542,N_1826);
or U5959 (N_5959,N_1501,N_624);
and U5960 (N_5960,N_1645,N_2411);
or U5961 (N_5961,N_2955,N_2870);
or U5962 (N_5962,N_168,N_2052);
nand U5963 (N_5963,N_1049,N_3627);
nor U5964 (N_5964,N_2849,N_927);
nand U5965 (N_5965,N_1297,N_3748);
or U5966 (N_5966,N_841,N_1643);
and U5967 (N_5967,N_3712,N_2771);
nand U5968 (N_5968,N_2780,N_28);
nor U5969 (N_5969,N_1047,N_2937);
or U5970 (N_5970,N_1347,N_606);
nand U5971 (N_5971,N_2868,N_2395);
or U5972 (N_5972,N_2125,N_2643);
or U5973 (N_5973,N_929,N_2256);
or U5974 (N_5974,N_3604,N_3811);
nand U5975 (N_5975,N_1573,N_303);
nand U5976 (N_5976,N_401,N_1084);
xnor U5977 (N_5977,N_1185,N_1747);
nand U5978 (N_5978,N_1737,N_3476);
nand U5979 (N_5979,N_524,N_1283);
or U5980 (N_5980,N_3540,N_3313);
nor U5981 (N_5981,N_2286,N_3448);
nand U5982 (N_5982,N_227,N_622);
nor U5983 (N_5983,N_1199,N_1869);
and U5984 (N_5984,N_3716,N_3466);
or U5985 (N_5985,N_2081,N_3781);
or U5986 (N_5986,N_699,N_1815);
nand U5987 (N_5987,N_2402,N_1808);
nand U5988 (N_5988,N_1967,N_3159);
nor U5989 (N_5989,N_3956,N_2416);
and U5990 (N_5990,N_3138,N_1830);
nand U5991 (N_5991,N_341,N_1565);
or U5992 (N_5992,N_1415,N_3552);
nand U5993 (N_5993,N_2627,N_2884);
nand U5994 (N_5994,N_2010,N_3535);
and U5995 (N_5995,N_2989,N_2885);
nand U5996 (N_5996,N_2362,N_2581);
nand U5997 (N_5997,N_3241,N_3199);
nor U5998 (N_5998,N_3946,N_597);
or U5999 (N_5999,N_2988,N_2545);
or U6000 (N_6000,N_2730,N_2746);
and U6001 (N_6001,N_1914,N_267);
and U6002 (N_6002,N_297,N_41);
nor U6003 (N_6003,N_279,N_3600);
and U6004 (N_6004,N_3696,N_3740);
nand U6005 (N_6005,N_3047,N_1015);
or U6006 (N_6006,N_3621,N_451);
and U6007 (N_6007,N_3190,N_1863);
nor U6008 (N_6008,N_1817,N_1027);
nand U6009 (N_6009,N_93,N_60);
and U6010 (N_6010,N_1605,N_1661);
or U6011 (N_6011,N_3423,N_3690);
nand U6012 (N_6012,N_2925,N_569);
and U6013 (N_6013,N_1060,N_3240);
xnor U6014 (N_6014,N_737,N_2877);
nand U6015 (N_6015,N_3427,N_2192);
nor U6016 (N_6016,N_3447,N_1331);
and U6017 (N_6017,N_3188,N_3568);
or U6018 (N_6018,N_2628,N_1610);
or U6019 (N_6019,N_1057,N_2514);
and U6020 (N_6020,N_1588,N_1390);
nor U6021 (N_6021,N_257,N_2166);
nand U6022 (N_6022,N_738,N_3247);
or U6023 (N_6023,N_588,N_428);
nand U6024 (N_6024,N_3908,N_2793);
nor U6025 (N_6025,N_2300,N_2728);
and U6026 (N_6026,N_3064,N_298);
nor U6027 (N_6027,N_846,N_1460);
nand U6028 (N_6028,N_1811,N_2733);
nand U6029 (N_6029,N_2344,N_3504);
and U6030 (N_6030,N_482,N_270);
nand U6031 (N_6031,N_846,N_810);
nor U6032 (N_6032,N_3233,N_2504);
nor U6033 (N_6033,N_1294,N_945);
nor U6034 (N_6034,N_2871,N_2908);
nor U6035 (N_6035,N_429,N_1199);
and U6036 (N_6036,N_3339,N_3070);
and U6037 (N_6037,N_2120,N_3117);
nor U6038 (N_6038,N_1044,N_238);
nor U6039 (N_6039,N_3088,N_2468);
nor U6040 (N_6040,N_2554,N_674);
and U6041 (N_6041,N_1613,N_2136);
nand U6042 (N_6042,N_3029,N_424);
and U6043 (N_6043,N_1474,N_1322);
or U6044 (N_6044,N_3399,N_2161);
nand U6045 (N_6045,N_3972,N_2123);
nand U6046 (N_6046,N_1143,N_2508);
nor U6047 (N_6047,N_686,N_2389);
or U6048 (N_6048,N_2455,N_2556);
nor U6049 (N_6049,N_718,N_220);
nor U6050 (N_6050,N_1536,N_1656);
or U6051 (N_6051,N_1094,N_3226);
and U6052 (N_6052,N_2921,N_3970);
nand U6053 (N_6053,N_593,N_588);
nand U6054 (N_6054,N_3506,N_3744);
nand U6055 (N_6055,N_102,N_3855);
xnor U6056 (N_6056,N_2383,N_1957);
nor U6057 (N_6057,N_3891,N_659);
or U6058 (N_6058,N_3494,N_1744);
nor U6059 (N_6059,N_3885,N_1610);
and U6060 (N_6060,N_2968,N_877);
nand U6061 (N_6061,N_1143,N_1614);
or U6062 (N_6062,N_1953,N_3387);
nand U6063 (N_6063,N_565,N_1919);
nor U6064 (N_6064,N_2543,N_2134);
nor U6065 (N_6065,N_1699,N_3654);
nand U6066 (N_6066,N_296,N_3551);
or U6067 (N_6067,N_2034,N_2506);
or U6068 (N_6068,N_3075,N_1287);
or U6069 (N_6069,N_869,N_617);
nor U6070 (N_6070,N_2178,N_2039);
nand U6071 (N_6071,N_3604,N_1873);
nor U6072 (N_6072,N_1123,N_2178);
and U6073 (N_6073,N_2034,N_2085);
or U6074 (N_6074,N_1792,N_2458);
nor U6075 (N_6075,N_2026,N_1334);
or U6076 (N_6076,N_3456,N_927);
and U6077 (N_6077,N_3503,N_3328);
nand U6078 (N_6078,N_351,N_1399);
nor U6079 (N_6079,N_728,N_744);
or U6080 (N_6080,N_2520,N_1076);
nor U6081 (N_6081,N_635,N_2980);
or U6082 (N_6082,N_3684,N_2821);
nor U6083 (N_6083,N_3664,N_2992);
and U6084 (N_6084,N_1622,N_341);
or U6085 (N_6085,N_401,N_1842);
and U6086 (N_6086,N_3354,N_1812);
and U6087 (N_6087,N_846,N_2045);
or U6088 (N_6088,N_2506,N_2060);
nor U6089 (N_6089,N_2176,N_1246);
nand U6090 (N_6090,N_2572,N_1968);
nor U6091 (N_6091,N_449,N_2179);
and U6092 (N_6092,N_387,N_1850);
and U6093 (N_6093,N_489,N_3886);
or U6094 (N_6094,N_1432,N_2221);
nand U6095 (N_6095,N_1479,N_3403);
nor U6096 (N_6096,N_3040,N_39);
and U6097 (N_6097,N_784,N_686);
nand U6098 (N_6098,N_3054,N_1764);
or U6099 (N_6099,N_3587,N_3322);
and U6100 (N_6100,N_2141,N_3865);
nand U6101 (N_6101,N_2857,N_1967);
nor U6102 (N_6102,N_1360,N_3309);
and U6103 (N_6103,N_3759,N_2206);
and U6104 (N_6104,N_3036,N_129);
nand U6105 (N_6105,N_1670,N_948);
nand U6106 (N_6106,N_567,N_3451);
nor U6107 (N_6107,N_1652,N_227);
nand U6108 (N_6108,N_1635,N_1411);
and U6109 (N_6109,N_878,N_3542);
and U6110 (N_6110,N_1113,N_329);
or U6111 (N_6111,N_110,N_3814);
and U6112 (N_6112,N_1878,N_2231);
nand U6113 (N_6113,N_3070,N_3294);
nand U6114 (N_6114,N_3115,N_2864);
and U6115 (N_6115,N_1401,N_583);
nor U6116 (N_6116,N_3477,N_1533);
or U6117 (N_6117,N_3084,N_11);
or U6118 (N_6118,N_1191,N_3549);
and U6119 (N_6119,N_2560,N_2423);
or U6120 (N_6120,N_2468,N_2028);
nor U6121 (N_6121,N_2024,N_670);
nor U6122 (N_6122,N_1701,N_2768);
nor U6123 (N_6123,N_979,N_2087);
nor U6124 (N_6124,N_2589,N_2593);
or U6125 (N_6125,N_804,N_2190);
or U6126 (N_6126,N_697,N_2990);
nand U6127 (N_6127,N_3708,N_2427);
nand U6128 (N_6128,N_3449,N_2995);
nand U6129 (N_6129,N_820,N_1968);
and U6130 (N_6130,N_3507,N_3942);
or U6131 (N_6131,N_987,N_2741);
nor U6132 (N_6132,N_997,N_1178);
or U6133 (N_6133,N_642,N_1138);
nand U6134 (N_6134,N_3331,N_2898);
and U6135 (N_6135,N_37,N_389);
and U6136 (N_6136,N_3450,N_3079);
or U6137 (N_6137,N_258,N_1024);
nand U6138 (N_6138,N_516,N_3371);
xor U6139 (N_6139,N_973,N_731);
nand U6140 (N_6140,N_2028,N_2841);
and U6141 (N_6141,N_3966,N_2866);
and U6142 (N_6142,N_907,N_2617);
nand U6143 (N_6143,N_50,N_1838);
or U6144 (N_6144,N_1742,N_3662);
and U6145 (N_6145,N_1195,N_2455);
or U6146 (N_6146,N_3899,N_311);
nand U6147 (N_6147,N_3768,N_2429);
and U6148 (N_6148,N_559,N_889);
nor U6149 (N_6149,N_687,N_3067);
or U6150 (N_6150,N_168,N_874);
nand U6151 (N_6151,N_1049,N_2825);
and U6152 (N_6152,N_3797,N_3506);
and U6153 (N_6153,N_332,N_3134);
and U6154 (N_6154,N_3915,N_3504);
and U6155 (N_6155,N_2269,N_25);
nor U6156 (N_6156,N_1642,N_3616);
nand U6157 (N_6157,N_1813,N_3083);
or U6158 (N_6158,N_3141,N_1039);
or U6159 (N_6159,N_761,N_1090);
nor U6160 (N_6160,N_1765,N_2369);
nor U6161 (N_6161,N_537,N_1903);
nor U6162 (N_6162,N_2719,N_1269);
nand U6163 (N_6163,N_3570,N_784);
xor U6164 (N_6164,N_616,N_1358);
or U6165 (N_6165,N_2799,N_3610);
and U6166 (N_6166,N_3812,N_3106);
nand U6167 (N_6167,N_3821,N_2383);
nor U6168 (N_6168,N_1631,N_1410);
nor U6169 (N_6169,N_644,N_3314);
or U6170 (N_6170,N_3868,N_78);
or U6171 (N_6171,N_2158,N_898);
nor U6172 (N_6172,N_3818,N_1368);
or U6173 (N_6173,N_2668,N_3889);
or U6174 (N_6174,N_2927,N_939);
nor U6175 (N_6175,N_1873,N_2640);
nand U6176 (N_6176,N_3222,N_3190);
nand U6177 (N_6177,N_800,N_1468);
or U6178 (N_6178,N_3537,N_961);
nor U6179 (N_6179,N_273,N_2095);
nand U6180 (N_6180,N_1638,N_2680);
or U6181 (N_6181,N_1082,N_3037);
nor U6182 (N_6182,N_1221,N_3959);
nand U6183 (N_6183,N_857,N_2566);
or U6184 (N_6184,N_3809,N_341);
nor U6185 (N_6185,N_3561,N_2726);
nor U6186 (N_6186,N_145,N_2688);
nor U6187 (N_6187,N_1505,N_1303);
nor U6188 (N_6188,N_395,N_2677);
nor U6189 (N_6189,N_1521,N_2312);
nand U6190 (N_6190,N_1072,N_858);
or U6191 (N_6191,N_1373,N_3032);
nor U6192 (N_6192,N_251,N_2633);
nor U6193 (N_6193,N_1187,N_509);
and U6194 (N_6194,N_163,N_1963);
nor U6195 (N_6195,N_867,N_809);
xnor U6196 (N_6196,N_17,N_620);
or U6197 (N_6197,N_1464,N_1415);
nor U6198 (N_6198,N_156,N_3389);
nand U6199 (N_6199,N_3914,N_3540);
and U6200 (N_6200,N_3787,N_3706);
nand U6201 (N_6201,N_1003,N_3086);
nor U6202 (N_6202,N_90,N_3911);
nand U6203 (N_6203,N_1381,N_369);
or U6204 (N_6204,N_2346,N_3183);
nor U6205 (N_6205,N_191,N_1346);
and U6206 (N_6206,N_720,N_2806);
and U6207 (N_6207,N_2825,N_3002);
nor U6208 (N_6208,N_1935,N_1849);
and U6209 (N_6209,N_2076,N_7);
or U6210 (N_6210,N_2806,N_3245);
and U6211 (N_6211,N_3291,N_2294);
nand U6212 (N_6212,N_3849,N_1842);
nor U6213 (N_6213,N_379,N_2387);
or U6214 (N_6214,N_2939,N_1654);
and U6215 (N_6215,N_3694,N_2646);
or U6216 (N_6216,N_228,N_3548);
or U6217 (N_6217,N_2024,N_2411);
nand U6218 (N_6218,N_3417,N_1329);
nor U6219 (N_6219,N_2534,N_1);
or U6220 (N_6220,N_3568,N_3166);
or U6221 (N_6221,N_1610,N_2624);
or U6222 (N_6222,N_2609,N_3162);
nand U6223 (N_6223,N_2903,N_1302);
or U6224 (N_6224,N_534,N_2870);
or U6225 (N_6225,N_2551,N_3824);
or U6226 (N_6226,N_2653,N_3789);
nor U6227 (N_6227,N_1205,N_3111);
nand U6228 (N_6228,N_1311,N_1901);
and U6229 (N_6229,N_1208,N_3520);
and U6230 (N_6230,N_2047,N_2570);
nand U6231 (N_6231,N_3570,N_589);
or U6232 (N_6232,N_574,N_1252);
and U6233 (N_6233,N_25,N_861);
and U6234 (N_6234,N_2581,N_131);
nor U6235 (N_6235,N_1195,N_3909);
nand U6236 (N_6236,N_1597,N_352);
nor U6237 (N_6237,N_2602,N_2280);
nand U6238 (N_6238,N_1706,N_955);
and U6239 (N_6239,N_1026,N_86);
or U6240 (N_6240,N_1002,N_2172);
and U6241 (N_6241,N_1982,N_1043);
or U6242 (N_6242,N_3379,N_73);
nor U6243 (N_6243,N_2709,N_3131);
nor U6244 (N_6244,N_2243,N_3580);
nor U6245 (N_6245,N_1645,N_2513);
or U6246 (N_6246,N_2503,N_3990);
and U6247 (N_6247,N_3495,N_1409);
nor U6248 (N_6248,N_1617,N_3550);
and U6249 (N_6249,N_1960,N_2309);
nand U6250 (N_6250,N_2310,N_2576);
and U6251 (N_6251,N_1439,N_1364);
nand U6252 (N_6252,N_840,N_2141);
and U6253 (N_6253,N_967,N_1608);
nand U6254 (N_6254,N_1587,N_934);
or U6255 (N_6255,N_3239,N_2345);
and U6256 (N_6256,N_2613,N_389);
and U6257 (N_6257,N_672,N_1746);
nand U6258 (N_6258,N_2816,N_2597);
nor U6259 (N_6259,N_3931,N_1265);
and U6260 (N_6260,N_2379,N_424);
nor U6261 (N_6261,N_3612,N_985);
and U6262 (N_6262,N_676,N_101);
nand U6263 (N_6263,N_441,N_1252);
and U6264 (N_6264,N_3368,N_2197);
or U6265 (N_6265,N_962,N_1113);
nand U6266 (N_6266,N_1646,N_997);
and U6267 (N_6267,N_2921,N_845);
xnor U6268 (N_6268,N_3748,N_2805);
and U6269 (N_6269,N_1018,N_1028);
and U6270 (N_6270,N_349,N_3104);
and U6271 (N_6271,N_1114,N_3544);
nor U6272 (N_6272,N_1407,N_3634);
nor U6273 (N_6273,N_2209,N_1495);
or U6274 (N_6274,N_1791,N_2386);
and U6275 (N_6275,N_1007,N_2880);
and U6276 (N_6276,N_1166,N_3446);
nor U6277 (N_6277,N_1765,N_1069);
and U6278 (N_6278,N_2231,N_3315);
or U6279 (N_6279,N_2687,N_2972);
and U6280 (N_6280,N_653,N_476);
nand U6281 (N_6281,N_74,N_1590);
nand U6282 (N_6282,N_3284,N_3252);
and U6283 (N_6283,N_309,N_1031);
nor U6284 (N_6284,N_693,N_3966);
and U6285 (N_6285,N_2369,N_2990);
or U6286 (N_6286,N_450,N_877);
nor U6287 (N_6287,N_2498,N_1709);
or U6288 (N_6288,N_3955,N_2136);
nand U6289 (N_6289,N_1647,N_3786);
or U6290 (N_6290,N_2838,N_2259);
and U6291 (N_6291,N_1566,N_2822);
xor U6292 (N_6292,N_3808,N_2961);
nand U6293 (N_6293,N_2685,N_2953);
and U6294 (N_6294,N_3813,N_1265);
nand U6295 (N_6295,N_2580,N_219);
nand U6296 (N_6296,N_1332,N_3916);
nor U6297 (N_6297,N_2818,N_1293);
and U6298 (N_6298,N_2371,N_278);
or U6299 (N_6299,N_2244,N_2093);
nor U6300 (N_6300,N_784,N_1707);
nor U6301 (N_6301,N_1209,N_1370);
nand U6302 (N_6302,N_2306,N_332);
nor U6303 (N_6303,N_2828,N_3397);
or U6304 (N_6304,N_2452,N_2358);
or U6305 (N_6305,N_673,N_1638);
nand U6306 (N_6306,N_93,N_1206);
nand U6307 (N_6307,N_937,N_3759);
or U6308 (N_6308,N_3388,N_3866);
and U6309 (N_6309,N_1237,N_1028);
nand U6310 (N_6310,N_828,N_3389);
nand U6311 (N_6311,N_435,N_799);
nor U6312 (N_6312,N_1779,N_138);
nor U6313 (N_6313,N_1154,N_787);
nor U6314 (N_6314,N_3823,N_3250);
and U6315 (N_6315,N_755,N_757);
and U6316 (N_6316,N_734,N_412);
or U6317 (N_6317,N_3497,N_3129);
nor U6318 (N_6318,N_1991,N_21);
or U6319 (N_6319,N_165,N_3327);
or U6320 (N_6320,N_1124,N_2965);
or U6321 (N_6321,N_3024,N_2642);
nor U6322 (N_6322,N_1822,N_3487);
or U6323 (N_6323,N_3856,N_1250);
nand U6324 (N_6324,N_3211,N_3993);
nor U6325 (N_6325,N_2459,N_1037);
nand U6326 (N_6326,N_3540,N_1874);
or U6327 (N_6327,N_941,N_3254);
nand U6328 (N_6328,N_2933,N_3143);
nor U6329 (N_6329,N_796,N_505);
or U6330 (N_6330,N_3508,N_3424);
nand U6331 (N_6331,N_370,N_176);
nand U6332 (N_6332,N_2028,N_1003);
nand U6333 (N_6333,N_3581,N_2633);
and U6334 (N_6334,N_3870,N_908);
or U6335 (N_6335,N_1075,N_2212);
or U6336 (N_6336,N_3907,N_2612);
nand U6337 (N_6337,N_2567,N_2598);
nand U6338 (N_6338,N_1737,N_426);
and U6339 (N_6339,N_1096,N_1753);
nor U6340 (N_6340,N_3209,N_1528);
and U6341 (N_6341,N_3650,N_1105);
nand U6342 (N_6342,N_2229,N_2108);
nor U6343 (N_6343,N_41,N_3153);
or U6344 (N_6344,N_1922,N_2722);
nand U6345 (N_6345,N_1445,N_3085);
or U6346 (N_6346,N_1083,N_943);
nand U6347 (N_6347,N_3842,N_3244);
and U6348 (N_6348,N_1801,N_240);
or U6349 (N_6349,N_104,N_713);
and U6350 (N_6350,N_3948,N_3868);
and U6351 (N_6351,N_686,N_2030);
nand U6352 (N_6352,N_164,N_2411);
nor U6353 (N_6353,N_907,N_2086);
or U6354 (N_6354,N_3325,N_512);
nor U6355 (N_6355,N_663,N_922);
nor U6356 (N_6356,N_3995,N_933);
nand U6357 (N_6357,N_2030,N_3080);
nor U6358 (N_6358,N_680,N_1899);
nand U6359 (N_6359,N_266,N_3091);
and U6360 (N_6360,N_238,N_1561);
nand U6361 (N_6361,N_767,N_1085);
and U6362 (N_6362,N_1757,N_326);
or U6363 (N_6363,N_1088,N_3593);
and U6364 (N_6364,N_3756,N_3918);
nor U6365 (N_6365,N_1586,N_2502);
nor U6366 (N_6366,N_3656,N_3702);
nor U6367 (N_6367,N_529,N_1988);
xor U6368 (N_6368,N_3545,N_2446);
nor U6369 (N_6369,N_1105,N_245);
and U6370 (N_6370,N_516,N_3275);
nor U6371 (N_6371,N_3712,N_2438);
nand U6372 (N_6372,N_1184,N_1975);
or U6373 (N_6373,N_3243,N_2301);
and U6374 (N_6374,N_122,N_3564);
nand U6375 (N_6375,N_892,N_303);
or U6376 (N_6376,N_621,N_1408);
and U6377 (N_6377,N_1021,N_1912);
and U6378 (N_6378,N_3367,N_2738);
nand U6379 (N_6379,N_2098,N_2329);
nor U6380 (N_6380,N_3113,N_3162);
nor U6381 (N_6381,N_1840,N_381);
nand U6382 (N_6382,N_2271,N_3605);
nand U6383 (N_6383,N_367,N_562);
and U6384 (N_6384,N_3969,N_1366);
and U6385 (N_6385,N_792,N_3190);
nand U6386 (N_6386,N_2360,N_2385);
nor U6387 (N_6387,N_905,N_3132);
nand U6388 (N_6388,N_3264,N_3291);
or U6389 (N_6389,N_1239,N_1465);
or U6390 (N_6390,N_373,N_2098);
and U6391 (N_6391,N_1586,N_3386);
or U6392 (N_6392,N_1963,N_3320);
and U6393 (N_6393,N_361,N_1862);
xnor U6394 (N_6394,N_2830,N_2034);
and U6395 (N_6395,N_1507,N_3716);
or U6396 (N_6396,N_2485,N_3010);
or U6397 (N_6397,N_380,N_747);
or U6398 (N_6398,N_2767,N_2610);
nor U6399 (N_6399,N_2109,N_698);
nor U6400 (N_6400,N_1672,N_3634);
and U6401 (N_6401,N_2835,N_2105);
nand U6402 (N_6402,N_2233,N_1670);
nor U6403 (N_6403,N_3527,N_1584);
and U6404 (N_6404,N_1684,N_672);
or U6405 (N_6405,N_3100,N_622);
nand U6406 (N_6406,N_1162,N_2475);
and U6407 (N_6407,N_2131,N_1964);
xnor U6408 (N_6408,N_1442,N_1580);
or U6409 (N_6409,N_2407,N_3793);
or U6410 (N_6410,N_3373,N_2398);
or U6411 (N_6411,N_3854,N_1768);
nand U6412 (N_6412,N_1820,N_10);
nor U6413 (N_6413,N_2021,N_1786);
nor U6414 (N_6414,N_1904,N_2628);
nand U6415 (N_6415,N_1813,N_3318);
nand U6416 (N_6416,N_1541,N_2443);
or U6417 (N_6417,N_47,N_1536);
nor U6418 (N_6418,N_568,N_1381);
or U6419 (N_6419,N_1596,N_68);
or U6420 (N_6420,N_3171,N_162);
xnor U6421 (N_6421,N_3562,N_2398);
nand U6422 (N_6422,N_2542,N_2103);
or U6423 (N_6423,N_1590,N_1846);
and U6424 (N_6424,N_340,N_793);
and U6425 (N_6425,N_3535,N_2651);
nor U6426 (N_6426,N_3571,N_1143);
nand U6427 (N_6427,N_2023,N_909);
nor U6428 (N_6428,N_3558,N_1821);
nand U6429 (N_6429,N_3742,N_2239);
xor U6430 (N_6430,N_2938,N_3727);
and U6431 (N_6431,N_3292,N_2989);
or U6432 (N_6432,N_1569,N_2549);
nor U6433 (N_6433,N_2815,N_2177);
nand U6434 (N_6434,N_3250,N_1370);
nand U6435 (N_6435,N_217,N_1343);
nand U6436 (N_6436,N_674,N_2404);
nand U6437 (N_6437,N_2250,N_3035);
and U6438 (N_6438,N_120,N_2291);
nor U6439 (N_6439,N_3104,N_3527);
nor U6440 (N_6440,N_2834,N_3297);
nand U6441 (N_6441,N_3833,N_721);
and U6442 (N_6442,N_62,N_1428);
and U6443 (N_6443,N_3037,N_3455);
and U6444 (N_6444,N_1524,N_1348);
and U6445 (N_6445,N_3810,N_1971);
nor U6446 (N_6446,N_1250,N_2598);
nor U6447 (N_6447,N_2707,N_3998);
or U6448 (N_6448,N_2327,N_837);
nand U6449 (N_6449,N_2929,N_3890);
nor U6450 (N_6450,N_3058,N_3737);
nand U6451 (N_6451,N_2783,N_665);
nand U6452 (N_6452,N_2339,N_3189);
and U6453 (N_6453,N_3606,N_3468);
nor U6454 (N_6454,N_3882,N_3778);
and U6455 (N_6455,N_527,N_115);
nand U6456 (N_6456,N_3682,N_905);
or U6457 (N_6457,N_718,N_466);
nand U6458 (N_6458,N_1525,N_2184);
and U6459 (N_6459,N_1046,N_1183);
nor U6460 (N_6460,N_277,N_3109);
and U6461 (N_6461,N_1093,N_2055);
and U6462 (N_6462,N_3663,N_390);
nor U6463 (N_6463,N_3654,N_2742);
nor U6464 (N_6464,N_2925,N_3360);
nand U6465 (N_6465,N_957,N_2351);
and U6466 (N_6466,N_2469,N_997);
xnor U6467 (N_6467,N_1428,N_2224);
and U6468 (N_6468,N_2613,N_786);
nand U6469 (N_6469,N_1711,N_3962);
xor U6470 (N_6470,N_1006,N_2632);
and U6471 (N_6471,N_2767,N_890);
or U6472 (N_6472,N_125,N_1744);
nor U6473 (N_6473,N_1464,N_1260);
and U6474 (N_6474,N_1835,N_629);
nand U6475 (N_6475,N_2096,N_2482);
nand U6476 (N_6476,N_1844,N_2691);
nand U6477 (N_6477,N_3158,N_2112);
and U6478 (N_6478,N_2846,N_1602);
or U6479 (N_6479,N_1654,N_2168);
nand U6480 (N_6480,N_3426,N_651);
and U6481 (N_6481,N_3255,N_2007);
and U6482 (N_6482,N_2831,N_1097);
and U6483 (N_6483,N_1813,N_105);
nor U6484 (N_6484,N_3611,N_3419);
nor U6485 (N_6485,N_3224,N_1223);
nor U6486 (N_6486,N_3821,N_1998);
or U6487 (N_6487,N_3741,N_1276);
nor U6488 (N_6488,N_1616,N_1796);
nand U6489 (N_6489,N_1025,N_379);
nand U6490 (N_6490,N_2090,N_6);
and U6491 (N_6491,N_1405,N_1358);
or U6492 (N_6492,N_2902,N_1076);
or U6493 (N_6493,N_3370,N_1217);
or U6494 (N_6494,N_3682,N_44);
nor U6495 (N_6495,N_2669,N_2213);
nor U6496 (N_6496,N_2996,N_3442);
nand U6497 (N_6497,N_1591,N_369);
and U6498 (N_6498,N_2303,N_1969);
and U6499 (N_6499,N_2952,N_1895);
nor U6500 (N_6500,N_531,N_542);
or U6501 (N_6501,N_164,N_531);
or U6502 (N_6502,N_444,N_2115);
nand U6503 (N_6503,N_3173,N_911);
nand U6504 (N_6504,N_137,N_456);
nand U6505 (N_6505,N_2626,N_2672);
and U6506 (N_6506,N_3605,N_3845);
or U6507 (N_6507,N_1913,N_1865);
or U6508 (N_6508,N_3502,N_1103);
or U6509 (N_6509,N_940,N_2760);
or U6510 (N_6510,N_3590,N_2353);
or U6511 (N_6511,N_776,N_2338);
nor U6512 (N_6512,N_3278,N_897);
or U6513 (N_6513,N_3643,N_72);
or U6514 (N_6514,N_2529,N_201);
or U6515 (N_6515,N_502,N_1050);
or U6516 (N_6516,N_2153,N_2360);
nor U6517 (N_6517,N_3999,N_2253);
and U6518 (N_6518,N_2067,N_92);
or U6519 (N_6519,N_2637,N_3648);
nor U6520 (N_6520,N_67,N_1519);
or U6521 (N_6521,N_1908,N_1404);
nand U6522 (N_6522,N_2175,N_179);
or U6523 (N_6523,N_570,N_659);
and U6524 (N_6524,N_3625,N_599);
nor U6525 (N_6525,N_2738,N_3559);
or U6526 (N_6526,N_3116,N_2895);
nand U6527 (N_6527,N_2243,N_1312);
nor U6528 (N_6528,N_2102,N_2096);
and U6529 (N_6529,N_2626,N_3871);
or U6530 (N_6530,N_1548,N_245);
nand U6531 (N_6531,N_2637,N_3953);
or U6532 (N_6532,N_1679,N_2313);
or U6533 (N_6533,N_2655,N_3436);
or U6534 (N_6534,N_3481,N_1158);
or U6535 (N_6535,N_3789,N_2376);
xnor U6536 (N_6536,N_1013,N_1481);
xnor U6537 (N_6537,N_325,N_3232);
nand U6538 (N_6538,N_1956,N_999);
nand U6539 (N_6539,N_2857,N_1803);
or U6540 (N_6540,N_245,N_3447);
or U6541 (N_6541,N_610,N_3176);
or U6542 (N_6542,N_962,N_2725);
or U6543 (N_6543,N_2408,N_3066);
nor U6544 (N_6544,N_1589,N_3573);
nand U6545 (N_6545,N_1776,N_3966);
nor U6546 (N_6546,N_2008,N_2212);
or U6547 (N_6547,N_3391,N_330);
nand U6548 (N_6548,N_948,N_2147);
nand U6549 (N_6549,N_3530,N_3811);
nand U6550 (N_6550,N_1917,N_1890);
and U6551 (N_6551,N_1645,N_982);
nand U6552 (N_6552,N_134,N_3828);
or U6553 (N_6553,N_977,N_113);
nand U6554 (N_6554,N_1438,N_3769);
nand U6555 (N_6555,N_372,N_2633);
or U6556 (N_6556,N_3183,N_1112);
nor U6557 (N_6557,N_3000,N_1913);
nor U6558 (N_6558,N_845,N_1347);
nor U6559 (N_6559,N_1837,N_1571);
nor U6560 (N_6560,N_2783,N_3271);
and U6561 (N_6561,N_162,N_3849);
or U6562 (N_6562,N_2210,N_1433);
and U6563 (N_6563,N_1091,N_3400);
nand U6564 (N_6564,N_3210,N_1941);
nor U6565 (N_6565,N_1170,N_69);
or U6566 (N_6566,N_2989,N_1070);
or U6567 (N_6567,N_1121,N_3602);
or U6568 (N_6568,N_2051,N_2707);
and U6569 (N_6569,N_3047,N_1124);
or U6570 (N_6570,N_1598,N_3175);
or U6571 (N_6571,N_1929,N_1642);
and U6572 (N_6572,N_3829,N_2043);
or U6573 (N_6573,N_1392,N_3631);
or U6574 (N_6574,N_2452,N_727);
or U6575 (N_6575,N_3263,N_1355);
and U6576 (N_6576,N_3924,N_304);
or U6577 (N_6577,N_164,N_796);
or U6578 (N_6578,N_2252,N_53);
or U6579 (N_6579,N_1889,N_2749);
and U6580 (N_6580,N_1664,N_2710);
xnor U6581 (N_6581,N_2708,N_2130);
nor U6582 (N_6582,N_741,N_1654);
or U6583 (N_6583,N_2187,N_2249);
and U6584 (N_6584,N_3046,N_2340);
nor U6585 (N_6585,N_3842,N_1832);
xnor U6586 (N_6586,N_1103,N_3045);
and U6587 (N_6587,N_1100,N_1530);
or U6588 (N_6588,N_3003,N_3331);
nor U6589 (N_6589,N_2671,N_1002);
nand U6590 (N_6590,N_3640,N_2327);
nor U6591 (N_6591,N_800,N_3746);
nand U6592 (N_6592,N_151,N_476);
nand U6593 (N_6593,N_1575,N_3713);
and U6594 (N_6594,N_1776,N_3303);
nor U6595 (N_6595,N_3983,N_694);
nand U6596 (N_6596,N_2672,N_2440);
and U6597 (N_6597,N_3224,N_2361);
and U6598 (N_6598,N_415,N_2320);
nor U6599 (N_6599,N_763,N_730);
or U6600 (N_6600,N_3379,N_1262);
nand U6601 (N_6601,N_394,N_1617);
and U6602 (N_6602,N_2397,N_3234);
nor U6603 (N_6603,N_1558,N_3320);
and U6604 (N_6604,N_3308,N_3413);
nor U6605 (N_6605,N_1179,N_2293);
nor U6606 (N_6606,N_593,N_2568);
nor U6607 (N_6607,N_2850,N_1419);
nand U6608 (N_6608,N_2900,N_1083);
nand U6609 (N_6609,N_3755,N_1546);
and U6610 (N_6610,N_2074,N_199);
nor U6611 (N_6611,N_3397,N_2970);
or U6612 (N_6612,N_224,N_3375);
and U6613 (N_6613,N_3371,N_1128);
or U6614 (N_6614,N_2414,N_2773);
nor U6615 (N_6615,N_3283,N_906);
nor U6616 (N_6616,N_2071,N_2519);
nand U6617 (N_6617,N_1242,N_3713);
nand U6618 (N_6618,N_3604,N_1150);
or U6619 (N_6619,N_3853,N_1738);
and U6620 (N_6620,N_2167,N_774);
and U6621 (N_6621,N_659,N_62);
or U6622 (N_6622,N_2771,N_495);
or U6623 (N_6623,N_1443,N_3353);
nand U6624 (N_6624,N_3017,N_606);
or U6625 (N_6625,N_819,N_3511);
or U6626 (N_6626,N_1978,N_373);
nand U6627 (N_6627,N_3643,N_3424);
nand U6628 (N_6628,N_1593,N_266);
or U6629 (N_6629,N_3068,N_3543);
and U6630 (N_6630,N_1398,N_3249);
nand U6631 (N_6631,N_2991,N_3538);
nor U6632 (N_6632,N_3617,N_1926);
or U6633 (N_6633,N_2168,N_225);
nand U6634 (N_6634,N_2980,N_1953);
nand U6635 (N_6635,N_1275,N_2579);
or U6636 (N_6636,N_2329,N_2350);
or U6637 (N_6637,N_1707,N_1365);
and U6638 (N_6638,N_3299,N_65);
nand U6639 (N_6639,N_215,N_3267);
and U6640 (N_6640,N_1393,N_3656);
nand U6641 (N_6641,N_3592,N_1515);
nand U6642 (N_6642,N_3744,N_1607);
nand U6643 (N_6643,N_749,N_3016);
nor U6644 (N_6644,N_2056,N_3752);
nand U6645 (N_6645,N_799,N_378);
nand U6646 (N_6646,N_1838,N_3990);
nor U6647 (N_6647,N_1140,N_643);
or U6648 (N_6648,N_1576,N_2926);
or U6649 (N_6649,N_2536,N_2277);
or U6650 (N_6650,N_583,N_2457);
or U6651 (N_6651,N_1425,N_2220);
or U6652 (N_6652,N_2727,N_842);
or U6653 (N_6653,N_3,N_395);
or U6654 (N_6654,N_2044,N_3491);
nand U6655 (N_6655,N_3558,N_1918);
nand U6656 (N_6656,N_1959,N_1699);
or U6657 (N_6657,N_2351,N_3416);
nand U6658 (N_6658,N_2181,N_1337);
nor U6659 (N_6659,N_1273,N_3970);
nor U6660 (N_6660,N_2442,N_859);
and U6661 (N_6661,N_3758,N_3628);
and U6662 (N_6662,N_2504,N_1675);
nand U6663 (N_6663,N_589,N_1169);
and U6664 (N_6664,N_3033,N_3994);
nor U6665 (N_6665,N_2149,N_3927);
nor U6666 (N_6666,N_3468,N_2816);
or U6667 (N_6667,N_2513,N_3520);
and U6668 (N_6668,N_2044,N_1802);
nor U6669 (N_6669,N_1975,N_2157);
or U6670 (N_6670,N_3080,N_891);
nand U6671 (N_6671,N_2954,N_3354);
nand U6672 (N_6672,N_3634,N_3250);
and U6673 (N_6673,N_1428,N_1579);
nand U6674 (N_6674,N_3171,N_3517);
nor U6675 (N_6675,N_309,N_2618);
or U6676 (N_6676,N_3271,N_873);
and U6677 (N_6677,N_2209,N_2556);
and U6678 (N_6678,N_1646,N_2509);
nand U6679 (N_6679,N_1475,N_2598);
and U6680 (N_6680,N_3952,N_472);
nor U6681 (N_6681,N_32,N_2560);
nand U6682 (N_6682,N_1682,N_276);
or U6683 (N_6683,N_554,N_3680);
and U6684 (N_6684,N_141,N_3642);
nor U6685 (N_6685,N_3138,N_2224);
nand U6686 (N_6686,N_3982,N_2656);
or U6687 (N_6687,N_2188,N_1936);
and U6688 (N_6688,N_2410,N_1469);
or U6689 (N_6689,N_2891,N_2724);
and U6690 (N_6690,N_421,N_27);
nor U6691 (N_6691,N_3274,N_2946);
nand U6692 (N_6692,N_2049,N_3979);
nand U6693 (N_6693,N_3744,N_1827);
and U6694 (N_6694,N_825,N_1745);
nor U6695 (N_6695,N_226,N_3975);
nand U6696 (N_6696,N_13,N_3046);
nor U6697 (N_6697,N_1172,N_398);
nand U6698 (N_6698,N_876,N_1501);
and U6699 (N_6699,N_245,N_931);
nor U6700 (N_6700,N_541,N_2724);
nand U6701 (N_6701,N_348,N_3333);
nand U6702 (N_6702,N_768,N_2565);
and U6703 (N_6703,N_1283,N_2558);
nor U6704 (N_6704,N_1994,N_871);
or U6705 (N_6705,N_3283,N_1483);
nor U6706 (N_6706,N_2191,N_3809);
and U6707 (N_6707,N_3473,N_2463);
or U6708 (N_6708,N_3845,N_1625);
nor U6709 (N_6709,N_2534,N_2716);
or U6710 (N_6710,N_98,N_1281);
and U6711 (N_6711,N_2465,N_2004);
nor U6712 (N_6712,N_3666,N_3712);
nand U6713 (N_6713,N_2507,N_1813);
and U6714 (N_6714,N_2464,N_520);
nor U6715 (N_6715,N_2881,N_1673);
or U6716 (N_6716,N_2694,N_1865);
nor U6717 (N_6717,N_487,N_856);
nor U6718 (N_6718,N_3867,N_8);
and U6719 (N_6719,N_2347,N_3916);
nor U6720 (N_6720,N_993,N_1342);
or U6721 (N_6721,N_1759,N_514);
nand U6722 (N_6722,N_2634,N_2502);
or U6723 (N_6723,N_1604,N_3414);
and U6724 (N_6724,N_3259,N_1411);
and U6725 (N_6725,N_3574,N_0);
and U6726 (N_6726,N_156,N_73);
or U6727 (N_6727,N_3077,N_3907);
nand U6728 (N_6728,N_1607,N_3411);
and U6729 (N_6729,N_653,N_298);
and U6730 (N_6730,N_214,N_313);
nor U6731 (N_6731,N_788,N_3690);
nor U6732 (N_6732,N_1215,N_1530);
nand U6733 (N_6733,N_2040,N_424);
and U6734 (N_6734,N_3476,N_609);
nand U6735 (N_6735,N_3917,N_2637);
nand U6736 (N_6736,N_1546,N_2585);
nor U6737 (N_6737,N_652,N_2359);
nand U6738 (N_6738,N_3552,N_1794);
or U6739 (N_6739,N_2628,N_2490);
xnor U6740 (N_6740,N_2418,N_3177);
nand U6741 (N_6741,N_1821,N_3060);
and U6742 (N_6742,N_488,N_60);
and U6743 (N_6743,N_738,N_2803);
and U6744 (N_6744,N_3637,N_1465);
nand U6745 (N_6745,N_3709,N_3358);
and U6746 (N_6746,N_2609,N_3879);
and U6747 (N_6747,N_444,N_818);
nor U6748 (N_6748,N_118,N_3138);
and U6749 (N_6749,N_3363,N_2404);
or U6750 (N_6750,N_1266,N_1849);
and U6751 (N_6751,N_3233,N_3209);
and U6752 (N_6752,N_838,N_3913);
or U6753 (N_6753,N_1331,N_418);
nor U6754 (N_6754,N_276,N_1675);
and U6755 (N_6755,N_2555,N_3232);
and U6756 (N_6756,N_2779,N_2302);
nand U6757 (N_6757,N_2188,N_1164);
and U6758 (N_6758,N_3302,N_3304);
nand U6759 (N_6759,N_3978,N_1182);
nor U6760 (N_6760,N_1480,N_1794);
nand U6761 (N_6761,N_2003,N_2);
or U6762 (N_6762,N_940,N_3838);
nand U6763 (N_6763,N_2127,N_1914);
nand U6764 (N_6764,N_2170,N_1486);
and U6765 (N_6765,N_2857,N_3060);
and U6766 (N_6766,N_123,N_476);
and U6767 (N_6767,N_2563,N_481);
nor U6768 (N_6768,N_3565,N_2590);
nor U6769 (N_6769,N_1866,N_2345);
or U6770 (N_6770,N_73,N_3321);
and U6771 (N_6771,N_2087,N_287);
or U6772 (N_6772,N_3050,N_1560);
nand U6773 (N_6773,N_170,N_998);
or U6774 (N_6774,N_3404,N_406);
or U6775 (N_6775,N_1842,N_3941);
or U6776 (N_6776,N_1728,N_3676);
nand U6777 (N_6777,N_1931,N_185);
nand U6778 (N_6778,N_1034,N_3230);
nor U6779 (N_6779,N_470,N_3124);
or U6780 (N_6780,N_2855,N_1117);
nand U6781 (N_6781,N_1475,N_2244);
and U6782 (N_6782,N_2983,N_2340);
nor U6783 (N_6783,N_1517,N_2392);
or U6784 (N_6784,N_2715,N_1380);
or U6785 (N_6785,N_1546,N_2399);
and U6786 (N_6786,N_2723,N_646);
or U6787 (N_6787,N_144,N_596);
or U6788 (N_6788,N_2801,N_2584);
nor U6789 (N_6789,N_1844,N_1824);
or U6790 (N_6790,N_3211,N_1271);
nand U6791 (N_6791,N_3237,N_3481);
or U6792 (N_6792,N_3335,N_334);
nor U6793 (N_6793,N_3547,N_3240);
or U6794 (N_6794,N_3213,N_956);
nand U6795 (N_6795,N_2831,N_1706);
nand U6796 (N_6796,N_1396,N_2333);
or U6797 (N_6797,N_829,N_2203);
nand U6798 (N_6798,N_589,N_100);
and U6799 (N_6799,N_3597,N_3219);
nand U6800 (N_6800,N_1465,N_3507);
or U6801 (N_6801,N_1074,N_2455);
or U6802 (N_6802,N_824,N_786);
or U6803 (N_6803,N_64,N_2248);
nor U6804 (N_6804,N_2939,N_354);
or U6805 (N_6805,N_602,N_1640);
and U6806 (N_6806,N_1418,N_1042);
or U6807 (N_6807,N_738,N_2348);
nand U6808 (N_6808,N_92,N_3638);
nor U6809 (N_6809,N_214,N_2772);
nor U6810 (N_6810,N_3727,N_2024);
nor U6811 (N_6811,N_2485,N_2804);
and U6812 (N_6812,N_3745,N_324);
nor U6813 (N_6813,N_3279,N_3842);
or U6814 (N_6814,N_2988,N_1761);
nor U6815 (N_6815,N_1103,N_1794);
nor U6816 (N_6816,N_2414,N_1928);
nand U6817 (N_6817,N_3739,N_1897);
or U6818 (N_6818,N_1729,N_1273);
or U6819 (N_6819,N_306,N_2821);
and U6820 (N_6820,N_309,N_2486);
and U6821 (N_6821,N_1138,N_2645);
and U6822 (N_6822,N_261,N_1161);
nor U6823 (N_6823,N_361,N_849);
nand U6824 (N_6824,N_3804,N_109);
or U6825 (N_6825,N_3658,N_2706);
and U6826 (N_6826,N_1888,N_2367);
and U6827 (N_6827,N_1260,N_365);
or U6828 (N_6828,N_1026,N_3800);
or U6829 (N_6829,N_376,N_516);
nor U6830 (N_6830,N_1072,N_2276);
nand U6831 (N_6831,N_3037,N_2904);
or U6832 (N_6832,N_2826,N_155);
and U6833 (N_6833,N_3521,N_3190);
and U6834 (N_6834,N_3706,N_1698);
nand U6835 (N_6835,N_251,N_3765);
nor U6836 (N_6836,N_1114,N_143);
xor U6837 (N_6837,N_633,N_3720);
nand U6838 (N_6838,N_143,N_220);
nand U6839 (N_6839,N_3263,N_3883);
nor U6840 (N_6840,N_3383,N_3106);
or U6841 (N_6841,N_1745,N_3906);
or U6842 (N_6842,N_3283,N_641);
and U6843 (N_6843,N_1076,N_1291);
nand U6844 (N_6844,N_2578,N_3246);
or U6845 (N_6845,N_366,N_3824);
nor U6846 (N_6846,N_3236,N_2892);
and U6847 (N_6847,N_2127,N_2803);
nor U6848 (N_6848,N_1875,N_2915);
or U6849 (N_6849,N_3821,N_2804);
and U6850 (N_6850,N_759,N_469);
nand U6851 (N_6851,N_2540,N_1798);
nand U6852 (N_6852,N_3593,N_3605);
nor U6853 (N_6853,N_3153,N_176);
and U6854 (N_6854,N_3456,N_1478);
or U6855 (N_6855,N_887,N_391);
nor U6856 (N_6856,N_2949,N_542);
nand U6857 (N_6857,N_405,N_2862);
nor U6858 (N_6858,N_61,N_873);
and U6859 (N_6859,N_3773,N_2061);
xor U6860 (N_6860,N_963,N_3452);
nand U6861 (N_6861,N_147,N_416);
nand U6862 (N_6862,N_301,N_618);
and U6863 (N_6863,N_3858,N_1367);
nor U6864 (N_6864,N_3408,N_2098);
nand U6865 (N_6865,N_108,N_3251);
and U6866 (N_6866,N_737,N_2753);
or U6867 (N_6867,N_3156,N_2846);
nand U6868 (N_6868,N_3377,N_3367);
or U6869 (N_6869,N_3655,N_1091);
and U6870 (N_6870,N_3532,N_639);
and U6871 (N_6871,N_2461,N_1857);
nor U6872 (N_6872,N_1945,N_353);
and U6873 (N_6873,N_3752,N_3321);
and U6874 (N_6874,N_2819,N_1078);
nand U6875 (N_6875,N_3034,N_1763);
nand U6876 (N_6876,N_94,N_3448);
nor U6877 (N_6877,N_1187,N_2599);
and U6878 (N_6878,N_2360,N_1489);
and U6879 (N_6879,N_2492,N_173);
and U6880 (N_6880,N_320,N_3697);
nor U6881 (N_6881,N_1822,N_2519);
nand U6882 (N_6882,N_988,N_3804);
nor U6883 (N_6883,N_3461,N_922);
or U6884 (N_6884,N_2776,N_1442);
nor U6885 (N_6885,N_2273,N_1284);
and U6886 (N_6886,N_154,N_3958);
and U6887 (N_6887,N_755,N_1914);
nand U6888 (N_6888,N_2963,N_1100);
nand U6889 (N_6889,N_3374,N_3815);
nor U6890 (N_6890,N_695,N_1992);
and U6891 (N_6891,N_3373,N_1932);
and U6892 (N_6892,N_1215,N_1454);
and U6893 (N_6893,N_2744,N_3268);
and U6894 (N_6894,N_2448,N_49);
and U6895 (N_6895,N_3854,N_3952);
and U6896 (N_6896,N_606,N_3365);
or U6897 (N_6897,N_1462,N_3467);
and U6898 (N_6898,N_1876,N_3339);
nor U6899 (N_6899,N_1696,N_146);
nand U6900 (N_6900,N_755,N_3788);
nand U6901 (N_6901,N_2111,N_3745);
and U6902 (N_6902,N_2498,N_2288);
nor U6903 (N_6903,N_1384,N_2332);
nor U6904 (N_6904,N_2335,N_3458);
nand U6905 (N_6905,N_3273,N_3214);
and U6906 (N_6906,N_873,N_3219);
nand U6907 (N_6907,N_3346,N_2650);
nand U6908 (N_6908,N_1030,N_2889);
and U6909 (N_6909,N_1914,N_2295);
nand U6910 (N_6910,N_2067,N_2770);
nor U6911 (N_6911,N_3713,N_473);
nor U6912 (N_6912,N_1825,N_73);
nor U6913 (N_6913,N_3735,N_2963);
or U6914 (N_6914,N_2473,N_2014);
nor U6915 (N_6915,N_1329,N_2192);
and U6916 (N_6916,N_2498,N_930);
nand U6917 (N_6917,N_1315,N_1097);
and U6918 (N_6918,N_1906,N_2576);
nand U6919 (N_6919,N_441,N_132);
nand U6920 (N_6920,N_2624,N_1697);
and U6921 (N_6921,N_2928,N_974);
nand U6922 (N_6922,N_1805,N_7);
and U6923 (N_6923,N_2602,N_3718);
nor U6924 (N_6924,N_3845,N_1380);
nor U6925 (N_6925,N_1342,N_2635);
or U6926 (N_6926,N_1675,N_2473);
and U6927 (N_6927,N_140,N_3163);
nand U6928 (N_6928,N_161,N_2731);
nand U6929 (N_6929,N_1954,N_118);
and U6930 (N_6930,N_492,N_2436);
and U6931 (N_6931,N_3623,N_964);
nand U6932 (N_6932,N_2731,N_3258);
or U6933 (N_6933,N_2180,N_2342);
nor U6934 (N_6934,N_3405,N_2046);
nor U6935 (N_6935,N_3453,N_5);
nor U6936 (N_6936,N_2283,N_515);
nor U6937 (N_6937,N_804,N_282);
nor U6938 (N_6938,N_2893,N_2768);
and U6939 (N_6939,N_3307,N_3736);
and U6940 (N_6940,N_2430,N_1194);
nand U6941 (N_6941,N_1173,N_2180);
nor U6942 (N_6942,N_1422,N_3742);
or U6943 (N_6943,N_891,N_117);
nand U6944 (N_6944,N_2136,N_1025);
and U6945 (N_6945,N_191,N_612);
nand U6946 (N_6946,N_2932,N_848);
and U6947 (N_6947,N_1851,N_1810);
or U6948 (N_6948,N_609,N_1627);
or U6949 (N_6949,N_841,N_2438);
and U6950 (N_6950,N_2023,N_1398);
or U6951 (N_6951,N_773,N_1739);
nand U6952 (N_6952,N_620,N_2106);
or U6953 (N_6953,N_1262,N_1371);
nor U6954 (N_6954,N_1301,N_671);
nor U6955 (N_6955,N_128,N_3375);
and U6956 (N_6956,N_432,N_3168);
nand U6957 (N_6957,N_843,N_3739);
or U6958 (N_6958,N_3917,N_309);
nand U6959 (N_6959,N_3932,N_1435);
nor U6960 (N_6960,N_3801,N_3206);
and U6961 (N_6961,N_1876,N_3350);
or U6962 (N_6962,N_3586,N_2239);
nand U6963 (N_6963,N_3320,N_1928);
or U6964 (N_6964,N_1524,N_2624);
nor U6965 (N_6965,N_2969,N_1764);
and U6966 (N_6966,N_3449,N_2226);
and U6967 (N_6967,N_2421,N_3964);
or U6968 (N_6968,N_1750,N_1417);
or U6969 (N_6969,N_3247,N_2443);
nor U6970 (N_6970,N_1669,N_2068);
and U6971 (N_6971,N_2286,N_3224);
nand U6972 (N_6972,N_2176,N_424);
or U6973 (N_6973,N_2751,N_1192);
or U6974 (N_6974,N_954,N_3317);
and U6975 (N_6975,N_2752,N_2687);
and U6976 (N_6976,N_2081,N_871);
nor U6977 (N_6977,N_143,N_1966);
and U6978 (N_6978,N_1162,N_1631);
or U6979 (N_6979,N_3958,N_515);
or U6980 (N_6980,N_1780,N_2469);
or U6981 (N_6981,N_1513,N_814);
nor U6982 (N_6982,N_392,N_2630);
nor U6983 (N_6983,N_2696,N_3647);
nand U6984 (N_6984,N_3306,N_680);
and U6985 (N_6985,N_512,N_1615);
and U6986 (N_6986,N_32,N_3262);
and U6987 (N_6987,N_3247,N_907);
or U6988 (N_6988,N_2453,N_218);
and U6989 (N_6989,N_2580,N_3168);
nor U6990 (N_6990,N_3231,N_338);
and U6991 (N_6991,N_3034,N_627);
or U6992 (N_6992,N_3798,N_3200);
nand U6993 (N_6993,N_3722,N_1683);
nand U6994 (N_6994,N_1373,N_706);
nor U6995 (N_6995,N_170,N_2782);
nor U6996 (N_6996,N_3152,N_1285);
nor U6997 (N_6997,N_3966,N_2244);
nand U6998 (N_6998,N_2241,N_1963);
or U6999 (N_6999,N_2162,N_1056);
or U7000 (N_7000,N_1270,N_1660);
or U7001 (N_7001,N_3284,N_3816);
nor U7002 (N_7002,N_3774,N_644);
and U7003 (N_7003,N_2127,N_1586);
and U7004 (N_7004,N_807,N_2122);
nor U7005 (N_7005,N_822,N_1158);
nand U7006 (N_7006,N_1951,N_2820);
and U7007 (N_7007,N_1661,N_2479);
and U7008 (N_7008,N_3369,N_1567);
or U7009 (N_7009,N_173,N_1170);
and U7010 (N_7010,N_2927,N_2759);
nand U7011 (N_7011,N_149,N_2258);
nor U7012 (N_7012,N_1148,N_3121);
and U7013 (N_7013,N_2033,N_3229);
nand U7014 (N_7014,N_3159,N_2370);
or U7015 (N_7015,N_1064,N_3347);
nand U7016 (N_7016,N_3255,N_1422);
and U7017 (N_7017,N_1323,N_1152);
or U7018 (N_7018,N_519,N_1643);
nand U7019 (N_7019,N_1304,N_3965);
or U7020 (N_7020,N_1824,N_1308);
nor U7021 (N_7021,N_565,N_1807);
nand U7022 (N_7022,N_736,N_2554);
nor U7023 (N_7023,N_3721,N_1926);
nand U7024 (N_7024,N_1816,N_1351);
nor U7025 (N_7025,N_421,N_905);
nand U7026 (N_7026,N_2820,N_86);
or U7027 (N_7027,N_3968,N_69);
or U7028 (N_7028,N_3058,N_756);
nor U7029 (N_7029,N_106,N_3399);
or U7030 (N_7030,N_1736,N_1001);
nand U7031 (N_7031,N_896,N_1944);
and U7032 (N_7032,N_2112,N_1547);
nor U7033 (N_7033,N_3743,N_2250);
nor U7034 (N_7034,N_3344,N_2197);
or U7035 (N_7035,N_2206,N_2933);
or U7036 (N_7036,N_1064,N_421);
or U7037 (N_7037,N_2773,N_1904);
or U7038 (N_7038,N_3349,N_218);
nand U7039 (N_7039,N_2605,N_291);
nand U7040 (N_7040,N_3926,N_1977);
nand U7041 (N_7041,N_3467,N_3989);
or U7042 (N_7042,N_2734,N_2215);
nand U7043 (N_7043,N_1682,N_606);
nand U7044 (N_7044,N_354,N_200);
nor U7045 (N_7045,N_2156,N_1856);
xor U7046 (N_7046,N_1953,N_911);
nand U7047 (N_7047,N_2030,N_745);
nor U7048 (N_7048,N_2424,N_3708);
and U7049 (N_7049,N_1404,N_3520);
or U7050 (N_7050,N_775,N_1758);
and U7051 (N_7051,N_3948,N_1350);
or U7052 (N_7052,N_1998,N_1270);
nor U7053 (N_7053,N_980,N_912);
or U7054 (N_7054,N_3797,N_2953);
nand U7055 (N_7055,N_216,N_3674);
or U7056 (N_7056,N_3618,N_548);
xnor U7057 (N_7057,N_2067,N_3582);
and U7058 (N_7058,N_3607,N_3525);
and U7059 (N_7059,N_1779,N_1446);
nor U7060 (N_7060,N_789,N_3328);
nand U7061 (N_7061,N_3223,N_326);
nand U7062 (N_7062,N_3257,N_764);
xor U7063 (N_7063,N_2391,N_1515);
and U7064 (N_7064,N_1360,N_209);
or U7065 (N_7065,N_3413,N_3216);
nor U7066 (N_7066,N_2815,N_3812);
and U7067 (N_7067,N_640,N_2405);
and U7068 (N_7068,N_3188,N_2623);
nor U7069 (N_7069,N_520,N_3822);
or U7070 (N_7070,N_2276,N_1603);
or U7071 (N_7071,N_321,N_1764);
nor U7072 (N_7072,N_1187,N_854);
and U7073 (N_7073,N_3310,N_3283);
and U7074 (N_7074,N_1668,N_1132);
nand U7075 (N_7075,N_687,N_2983);
or U7076 (N_7076,N_1175,N_3042);
and U7077 (N_7077,N_2860,N_1317);
nor U7078 (N_7078,N_475,N_3163);
and U7079 (N_7079,N_1717,N_1706);
nand U7080 (N_7080,N_1377,N_1683);
and U7081 (N_7081,N_2693,N_1663);
and U7082 (N_7082,N_609,N_192);
nand U7083 (N_7083,N_2510,N_299);
and U7084 (N_7084,N_1207,N_615);
or U7085 (N_7085,N_2167,N_1228);
or U7086 (N_7086,N_1668,N_342);
and U7087 (N_7087,N_864,N_1631);
or U7088 (N_7088,N_2683,N_3171);
nor U7089 (N_7089,N_2578,N_3336);
nor U7090 (N_7090,N_1082,N_1615);
nand U7091 (N_7091,N_3035,N_3881);
and U7092 (N_7092,N_3418,N_819);
nor U7093 (N_7093,N_1331,N_3893);
or U7094 (N_7094,N_741,N_241);
nor U7095 (N_7095,N_3787,N_2458);
and U7096 (N_7096,N_3863,N_2128);
and U7097 (N_7097,N_3125,N_1648);
and U7098 (N_7098,N_3179,N_968);
and U7099 (N_7099,N_2541,N_3202);
and U7100 (N_7100,N_3184,N_3750);
nor U7101 (N_7101,N_1562,N_1959);
and U7102 (N_7102,N_311,N_3671);
nor U7103 (N_7103,N_2554,N_1187);
or U7104 (N_7104,N_1797,N_1448);
nor U7105 (N_7105,N_2516,N_1150);
nor U7106 (N_7106,N_3469,N_1758);
nor U7107 (N_7107,N_2284,N_3053);
and U7108 (N_7108,N_2787,N_2401);
and U7109 (N_7109,N_1339,N_2315);
or U7110 (N_7110,N_1632,N_2549);
and U7111 (N_7111,N_882,N_2469);
or U7112 (N_7112,N_1680,N_1964);
nor U7113 (N_7113,N_3784,N_2728);
nor U7114 (N_7114,N_1394,N_2025);
or U7115 (N_7115,N_1336,N_2867);
nand U7116 (N_7116,N_3665,N_448);
nor U7117 (N_7117,N_2657,N_2827);
and U7118 (N_7118,N_3746,N_2958);
nor U7119 (N_7119,N_1861,N_3717);
and U7120 (N_7120,N_1986,N_445);
and U7121 (N_7121,N_2203,N_547);
and U7122 (N_7122,N_1858,N_171);
or U7123 (N_7123,N_2774,N_3362);
nand U7124 (N_7124,N_2405,N_2520);
nor U7125 (N_7125,N_54,N_800);
nor U7126 (N_7126,N_2821,N_2496);
and U7127 (N_7127,N_1495,N_2217);
and U7128 (N_7128,N_159,N_2844);
or U7129 (N_7129,N_1168,N_1713);
or U7130 (N_7130,N_3618,N_2368);
or U7131 (N_7131,N_2713,N_2006);
nand U7132 (N_7132,N_2493,N_3629);
nand U7133 (N_7133,N_939,N_1795);
or U7134 (N_7134,N_3686,N_2033);
and U7135 (N_7135,N_1915,N_1557);
nor U7136 (N_7136,N_3542,N_2506);
or U7137 (N_7137,N_2374,N_3647);
nand U7138 (N_7138,N_3544,N_3006);
and U7139 (N_7139,N_2323,N_2584);
and U7140 (N_7140,N_362,N_2077);
nand U7141 (N_7141,N_631,N_3408);
and U7142 (N_7142,N_2660,N_2625);
or U7143 (N_7143,N_103,N_2397);
and U7144 (N_7144,N_1994,N_2196);
or U7145 (N_7145,N_721,N_3882);
and U7146 (N_7146,N_2834,N_1429);
nor U7147 (N_7147,N_625,N_3547);
nor U7148 (N_7148,N_2291,N_17);
or U7149 (N_7149,N_1263,N_1973);
nand U7150 (N_7150,N_3127,N_3196);
or U7151 (N_7151,N_1039,N_1302);
nand U7152 (N_7152,N_2949,N_908);
or U7153 (N_7153,N_2154,N_2422);
nand U7154 (N_7154,N_2487,N_2326);
or U7155 (N_7155,N_3321,N_869);
nor U7156 (N_7156,N_315,N_3789);
or U7157 (N_7157,N_1671,N_1209);
nor U7158 (N_7158,N_3589,N_2713);
and U7159 (N_7159,N_95,N_426);
nor U7160 (N_7160,N_2773,N_1365);
and U7161 (N_7161,N_3218,N_1378);
and U7162 (N_7162,N_635,N_1761);
nor U7163 (N_7163,N_3145,N_2792);
and U7164 (N_7164,N_2209,N_2015);
or U7165 (N_7165,N_627,N_3478);
or U7166 (N_7166,N_3151,N_438);
nor U7167 (N_7167,N_568,N_3005);
nand U7168 (N_7168,N_1336,N_3058);
nor U7169 (N_7169,N_408,N_129);
nand U7170 (N_7170,N_2743,N_3320);
xnor U7171 (N_7171,N_2828,N_3000);
nand U7172 (N_7172,N_3732,N_2703);
or U7173 (N_7173,N_3464,N_1128);
or U7174 (N_7174,N_2021,N_2671);
or U7175 (N_7175,N_1644,N_797);
nand U7176 (N_7176,N_3594,N_839);
nand U7177 (N_7177,N_1220,N_2006);
and U7178 (N_7178,N_1332,N_1224);
nand U7179 (N_7179,N_1310,N_386);
nor U7180 (N_7180,N_3568,N_1885);
nor U7181 (N_7181,N_2256,N_2463);
and U7182 (N_7182,N_3771,N_1061);
or U7183 (N_7183,N_1296,N_541);
nor U7184 (N_7184,N_2050,N_2679);
nand U7185 (N_7185,N_1373,N_2507);
nor U7186 (N_7186,N_31,N_1036);
or U7187 (N_7187,N_3097,N_1548);
nor U7188 (N_7188,N_1378,N_575);
nor U7189 (N_7189,N_2958,N_902);
nand U7190 (N_7190,N_2344,N_2446);
nor U7191 (N_7191,N_1291,N_1737);
and U7192 (N_7192,N_764,N_106);
and U7193 (N_7193,N_740,N_2020);
nor U7194 (N_7194,N_3475,N_2989);
and U7195 (N_7195,N_176,N_3468);
nor U7196 (N_7196,N_2053,N_1803);
and U7197 (N_7197,N_2685,N_1168);
nand U7198 (N_7198,N_1219,N_3854);
nand U7199 (N_7199,N_1158,N_1958);
or U7200 (N_7200,N_1479,N_1447);
nor U7201 (N_7201,N_2132,N_136);
nand U7202 (N_7202,N_3270,N_2751);
nand U7203 (N_7203,N_3063,N_3344);
or U7204 (N_7204,N_750,N_1188);
or U7205 (N_7205,N_3435,N_1778);
nor U7206 (N_7206,N_2142,N_1144);
nor U7207 (N_7207,N_3849,N_3751);
nand U7208 (N_7208,N_465,N_777);
nor U7209 (N_7209,N_3811,N_451);
nand U7210 (N_7210,N_2334,N_107);
and U7211 (N_7211,N_3910,N_1548);
nor U7212 (N_7212,N_1758,N_3002);
or U7213 (N_7213,N_3579,N_3172);
nand U7214 (N_7214,N_2506,N_1033);
nor U7215 (N_7215,N_2505,N_2250);
nor U7216 (N_7216,N_104,N_188);
or U7217 (N_7217,N_1082,N_1837);
nor U7218 (N_7218,N_2347,N_190);
and U7219 (N_7219,N_2612,N_666);
nor U7220 (N_7220,N_2325,N_822);
or U7221 (N_7221,N_3066,N_2373);
and U7222 (N_7222,N_1229,N_1993);
or U7223 (N_7223,N_3748,N_2407);
or U7224 (N_7224,N_2791,N_2019);
and U7225 (N_7225,N_1376,N_2643);
and U7226 (N_7226,N_563,N_3645);
or U7227 (N_7227,N_1637,N_3248);
and U7228 (N_7228,N_3079,N_2206);
or U7229 (N_7229,N_1036,N_73);
nand U7230 (N_7230,N_1941,N_671);
nand U7231 (N_7231,N_660,N_407);
nand U7232 (N_7232,N_1377,N_480);
nand U7233 (N_7233,N_3454,N_2655);
or U7234 (N_7234,N_634,N_3452);
nor U7235 (N_7235,N_991,N_3815);
xor U7236 (N_7236,N_2076,N_1480);
and U7237 (N_7237,N_3573,N_58);
or U7238 (N_7238,N_2370,N_3337);
nor U7239 (N_7239,N_2488,N_3707);
or U7240 (N_7240,N_696,N_3101);
nand U7241 (N_7241,N_3506,N_1113);
nor U7242 (N_7242,N_1410,N_2470);
and U7243 (N_7243,N_1950,N_2745);
and U7244 (N_7244,N_267,N_672);
and U7245 (N_7245,N_946,N_1097);
nand U7246 (N_7246,N_2213,N_1089);
nor U7247 (N_7247,N_3393,N_3736);
and U7248 (N_7248,N_3351,N_2581);
and U7249 (N_7249,N_2993,N_2726);
and U7250 (N_7250,N_2180,N_2677);
or U7251 (N_7251,N_3008,N_3172);
nor U7252 (N_7252,N_3316,N_137);
or U7253 (N_7253,N_2880,N_2686);
nand U7254 (N_7254,N_598,N_277);
nor U7255 (N_7255,N_1748,N_3707);
and U7256 (N_7256,N_93,N_2497);
nor U7257 (N_7257,N_3910,N_3269);
nor U7258 (N_7258,N_1279,N_72);
nand U7259 (N_7259,N_2728,N_3375);
nand U7260 (N_7260,N_2714,N_2822);
nor U7261 (N_7261,N_1687,N_3667);
or U7262 (N_7262,N_2717,N_1003);
nand U7263 (N_7263,N_279,N_2551);
nand U7264 (N_7264,N_704,N_592);
or U7265 (N_7265,N_3736,N_1084);
nor U7266 (N_7266,N_3217,N_2197);
or U7267 (N_7267,N_3525,N_2201);
nor U7268 (N_7268,N_1708,N_1149);
nand U7269 (N_7269,N_965,N_3247);
nand U7270 (N_7270,N_525,N_1674);
or U7271 (N_7271,N_3703,N_1849);
or U7272 (N_7272,N_2348,N_1903);
nand U7273 (N_7273,N_3297,N_2048);
or U7274 (N_7274,N_390,N_175);
nor U7275 (N_7275,N_1585,N_3117);
xor U7276 (N_7276,N_3894,N_2239);
and U7277 (N_7277,N_1694,N_2470);
nand U7278 (N_7278,N_128,N_3777);
and U7279 (N_7279,N_1313,N_460);
nor U7280 (N_7280,N_3113,N_246);
nand U7281 (N_7281,N_3294,N_3257);
or U7282 (N_7282,N_2258,N_3273);
nand U7283 (N_7283,N_3579,N_9);
nand U7284 (N_7284,N_886,N_3137);
nor U7285 (N_7285,N_3517,N_1013);
nand U7286 (N_7286,N_3306,N_3858);
or U7287 (N_7287,N_178,N_2705);
nand U7288 (N_7288,N_222,N_367);
nand U7289 (N_7289,N_1010,N_2911);
nand U7290 (N_7290,N_3425,N_3460);
and U7291 (N_7291,N_3602,N_3141);
nor U7292 (N_7292,N_2611,N_101);
and U7293 (N_7293,N_93,N_1901);
or U7294 (N_7294,N_2917,N_1248);
nand U7295 (N_7295,N_309,N_3038);
nor U7296 (N_7296,N_2266,N_1539);
and U7297 (N_7297,N_2199,N_1375);
nand U7298 (N_7298,N_2513,N_3394);
nand U7299 (N_7299,N_1704,N_3161);
or U7300 (N_7300,N_1262,N_3765);
nor U7301 (N_7301,N_3366,N_3403);
nand U7302 (N_7302,N_1686,N_1060);
or U7303 (N_7303,N_1874,N_1488);
nor U7304 (N_7304,N_199,N_1856);
nor U7305 (N_7305,N_1260,N_3251);
or U7306 (N_7306,N_1276,N_2849);
and U7307 (N_7307,N_2370,N_3218);
nor U7308 (N_7308,N_671,N_1659);
and U7309 (N_7309,N_1536,N_981);
and U7310 (N_7310,N_478,N_2555);
or U7311 (N_7311,N_1534,N_1465);
or U7312 (N_7312,N_1347,N_2895);
or U7313 (N_7313,N_3473,N_1601);
or U7314 (N_7314,N_163,N_2639);
or U7315 (N_7315,N_1337,N_2428);
nor U7316 (N_7316,N_133,N_89);
or U7317 (N_7317,N_2334,N_2786);
nand U7318 (N_7318,N_3113,N_1907);
nand U7319 (N_7319,N_2922,N_587);
nor U7320 (N_7320,N_3492,N_2261);
nor U7321 (N_7321,N_3695,N_3648);
and U7322 (N_7322,N_1374,N_3671);
and U7323 (N_7323,N_1492,N_1028);
nand U7324 (N_7324,N_1466,N_635);
nand U7325 (N_7325,N_1274,N_3074);
nand U7326 (N_7326,N_1167,N_1174);
nand U7327 (N_7327,N_306,N_1698);
or U7328 (N_7328,N_1995,N_3016);
and U7329 (N_7329,N_1153,N_1912);
and U7330 (N_7330,N_3889,N_2381);
and U7331 (N_7331,N_2991,N_945);
nand U7332 (N_7332,N_3871,N_1458);
or U7333 (N_7333,N_2021,N_2659);
and U7334 (N_7334,N_251,N_250);
nor U7335 (N_7335,N_2298,N_65);
nor U7336 (N_7336,N_2258,N_3908);
nor U7337 (N_7337,N_1249,N_3790);
nand U7338 (N_7338,N_2085,N_2755);
nor U7339 (N_7339,N_3949,N_626);
nand U7340 (N_7340,N_660,N_1396);
and U7341 (N_7341,N_3329,N_549);
and U7342 (N_7342,N_1271,N_1430);
nand U7343 (N_7343,N_1805,N_2891);
or U7344 (N_7344,N_1904,N_756);
and U7345 (N_7345,N_3913,N_2983);
nand U7346 (N_7346,N_2276,N_2252);
nand U7347 (N_7347,N_2865,N_3967);
nand U7348 (N_7348,N_3693,N_1917);
and U7349 (N_7349,N_1776,N_3491);
and U7350 (N_7350,N_3892,N_1332);
nor U7351 (N_7351,N_2955,N_562);
or U7352 (N_7352,N_1339,N_2959);
or U7353 (N_7353,N_2350,N_891);
nor U7354 (N_7354,N_1713,N_3384);
and U7355 (N_7355,N_3955,N_2760);
or U7356 (N_7356,N_3018,N_1033);
or U7357 (N_7357,N_3585,N_2799);
nand U7358 (N_7358,N_318,N_2993);
or U7359 (N_7359,N_2744,N_624);
or U7360 (N_7360,N_1825,N_2285);
nand U7361 (N_7361,N_2126,N_2308);
nor U7362 (N_7362,N_3578,N_1129);
and U7363 (N_7363,N_2439,N_1373);
or U7364 (N_7364,N_2534,N_840);
or U7365 (N_7365,N_2152,N_3112);
nand U7366 (N_7366,N_1067,N_846);
xnor U7367 (N_7367,N_1541,N_3155);
nand U7368 (N_7368,N_1432,N_3784);
nor U7369 (N_7369,N_2529,N_1987);
or U7370 (N_7370,N_3675,N_882);
and U7371 (N_7371,N_347,N_3549);
and U7372 (N_7372,N_3136,N_982);
or U7373 (N_7373,N_2922,N_1378);
and U7374 (N_7374,N_101,N_429);
nor U7375 (N_7375,N_1977,N_831);
or U7376 (N_7376,N_1201,N_3653);
or U7377 (N_7377,N_1130,N_1255);
nor U7378 (N_7378,N_687,N_2797);
and U7379 (N_7379,N_2754,N_1957);
nor U7380 (N_7380,N_2198,N_3586);
or U7381 (N_7381,N_2708,N_3736);
and U7382 (N_7382,N_1131,N_3998);
nor U7383 (N_7383,N_1678,N_832);
nand U7384 (N_7384,N_2016,N_1366);
nand U7385 (N_7385,N_3152,N_41);
nand U7386 (N_7386,N_3743,N_1657);
nor U7387 (N_7387,N_1620,N_3045);
nor U7388 (N_7388,N_3042,N_2476);
nor U7389 (N_7389,N_3141,N_3956);
and U7390 (N_7390,N_3342,N_1294);
or U7391 (N_7391,N_3140,N_3491);
nor U7392 (N_7392,N_411,N_3618);
or U7393 (N_7393,N_1379,N_568);
nor U7394 (N_7394,N_3757,N_2324);
nand U7395 (N_7395,N_530,N_660);
nor U7396 (N_7396,N_1283,N_1646);
nor U7397 (N_7397,N_989,N_476);
nand U7398 (N_7398,N_3457,N_981);
nor U7399 (N_7399,N_1349,N_1596);
nand U7400 (N_7400,N_3150,N_2010);
nor U7401 (N_7401,N_3801,N_1804);
nand U7402 (N_7402,N_625,N_733);
or U7403 (N_7403,N_2447,N_332);
or U7404 (N_7404,N_2810,N_2908);
nand U7405 (N_7405,N_2832,N_786);
and U7406 (N_7406,N_3688,N_3799);
or U7407 (N_7407,N_889,N_244);
nand U7408 (N_7408,N_189,N_1194);
and U7409 (N_7409,N_3617,N_3442);
nand U7410 (N_7410,N_839,N_2739);
or U7411 (N_7411,N_2843,N_2395);
and U7412 (N_7412,N_2933,N_1034);
nor U7413 (N_7413,N_227,N_2426);
nor U7414 (N_7414,N_2768,N_2336);
nand U7415 (N_7415,N_3925,N_2871);
and U7416 (N_7416,N_613,N_3098);
nor U7417 (N_7417,N_1089,N_689);
or U7418 (N_7418,N_1223,N_944);
and U7419 (N_7419,N_3168,N_2928);
or U7420 (N_7420,N_2573,N_1288);
nor U7421 (N_7421,N_2694,N_1486);
nor U7422 (N_7422,N_2751,N_2517);
or U7423 (N_7423,N_1489,N_315);
nand U7424 (N_7424,N_1961,N_2740);
nand U7425 (N_7425,N_2974,N_2886);
and U7426 (N_7426,N_1601,N_2713);
nand U7427 (N_7427,N_2663,N_2968);
and U7428 (N_7428,N_3045,N_2411);
or U7429 (N_7429,N_1225,N_1158);
nand U7430 (N_7430,N_2472,N_2679);
or U7431 (N_7431,N_364,N_87);
and U7432 (N_7432,N_2909,N_885);
nor U7433 (N_7433,N_1068,N_3150);
or U7434 (N_7434,N_1643,N_3599);
or U7435 (N_7435,N_3124,N_2304);
and U7436 (N_7436,N_1463,N_3367);
or U7437 (N_7437,N_532,N_996);
and U7438 (N_7438,N_3447,N_983);
nor U7439 (N_7439,N_1706,N_452);
and U7440 (N_7440,N_3948,N_3883);
nand U7441 (N_7441,N_1992,N_2427);
nor U7442 (N_7442,N_877,N_1335);
nor U7443 (N_7443,N_1469,N_793);
nor U7444 (N_7444,N_3220,N_1924);
and U7445 (N_7445,N_1627,N_183);
nor U7446 (N_7446,N_3578,N_961);
nand U7447 (N_7447,N_1683,N_460);
nand U7448 (N_7448,N_38,N_1957);
and U7449 (N_7449,N_2114,N_3764);
or U7450 (N_7450,N_52,N_3806);
nor U7451 (N_7451,N_2484,N_2651);
and U7452 (N_7452,N_774,N_617);
or U7453 (N_7453,N_2380,N_1625);
or U7454 (N_7454,N_3313,N_1859);
or U7455 (N_7455,N_545,N_2398);
or U7456 (N_7456,N_2166,N_3439);
nor U7457 (N_7457,N_3117,N_2745);
nor U7458 (N_7458,N_1023,N_2916);
nand U7459 (N_7459,N_1274,N_886);
and U7460 (N_7460,N_2604,N_495);
or U7461 (N_7461,N_2810,N_89);
nand U7462 (N_7462,N_2598,N_2105);
nand U7463 (N_7463,N_1159,N_1402);
nor U7464 (N_7464,N_2188,N_1001);
nand U7465 (N_7465,N_3813,N_2622);
nor U7466 (N_7466,N_977,N_3262);
and U7467 (N_7467,N_1299,N_2016);
or U7468 (N_7468,N_3914,N_3768);
nand U7469 (N_7469,N_2140,N_2734);
nand U7470 (N_7470,N_1721,N_957);
nand U7471 (N_7471,N_3905,N_2480);
or U7472 (N_7472,N_3117,N_16);
or U7473 (N_7473,N_1319,N_3822);
nand U7474 (N_7474,N_3364,N_3407);
nand U7475 (N_7475,N_183,N_539);
nor U7476 (N_7476,N_3833,N_2939);
nand U7477 (N_7477,N_3119,N_438);
nand U7478 (N_7478,N_3490,N_1835);
nor U7479 (N_7479,N_3042,N_443);
and U7480 (N_7480,N_3334,N_2907);
nand U7481 (N_7481,N_1541,N_3758);
nand U7482 (N_7482,N_1519,N_246);
nor U7483 (N_7483,N_2685,N_1721);
or U7484 (N_7484,N_3131,N_582);
or U7485 (N_7485,N_2778,N_999);
and U7486 (N_7486,N_3852,N_2315);
nand U7487 (N_7487,N_2058,N_53);
nor U7488 (N_7488,N_1410,N_1221);
and U7489 (N_7489,N_1633,N_32);
nor U7490 (N_7490,N_455,N_836);
or U7491 (N_7491,N_149,N_3716);
nand U7492 (N_7492,N_2889,N_3695);
xnor U7493 (N_7493,N_2735,N_1636);
nand U7494 (N_7494,N_3413,N_3132);
nand U7495 (N_7495,N_412,N_3614);
and U7496 (N_7496,N_2971,N_2395);
xor U7497 (N_7497,N_1181,N_3808);
or U7498 (N_7498,N_2364,N_3905);
nand U7499 (N_7499,N_2341,N_3869);
nor U7500 (N_7500,N_736,N_3628);
or U7501 (N_7501,N_2486,N_878);
nand U7502 (N_7502,N_2516,N_90);
or U7503 (N_7503,N_2599,N_1095);
or U7504 (N_7504,N_1141,N_3498);
and U7505 (N_7505,N_2549,N_2212);
and U7506 (N_7506,N_1686,N_2674);
nor U7507 (N_7507,N_1422,N_3219);
nand U7508 (N_7508,N_3769,N_3258);
nand U7509 (N_7509,N_228,N_1925);
nor U7510 (N_7510,N_2055,N_1710);
and U7511 (N_7511,N_2698,N_2152);
nand U7512 (N_7512,N_2365,N_1577);
and U7513 (N_7513,N_2693,N_3203);
nor U7514 (N_7514,N_2226,N_1697);
nand U7515 (N_7515,N_2602,N_1200);
or U7516 (N_7516,N_1643,N_992);
xor U7517 (N_7517,N_3862,N_2323);
nor U7518 (N_7518,N_265,N_2574);
and U7519 (N_7519,N_2266,N_1687);
or U7520 (N_7520,N_59,N_1641);
and U7521 (N_7521,N_1591,N_76);
or U7522 (N_7522,N_1659,N_1664);
and U7523 (N_7523,N_492,N_1683);
nor U7524 (N_7524,N_3756,N_354);
nand U7525 (N_7525,N_1619,N_2547);
and U7526 (N_7526,N_248,N_1260);
and U7527 (N_7527,N_3410,N_166);
and U7528 (N_7528,N_1087,N_3989);
nor U7529 (N_7529,N_3278,N_3882);
nand U7530 (N_7530,N_3656,N_1031);
and U7531 (N_7531,N_3129,N_2825);
and U7532 (N_7532,N_1776,N_2926);
nor U7533 (N_7533,N_917,N_2513);
nor U7534 (N_7534,N_3733,N_2101);
or U7535 (N_7535,N_3404,N_804);
and U7536 (N_7536,N_1712,N_1337);
or U7537 (N_7537,N_3718,N_2903);
nand U7538 (N_7538,N_3457,N_203);
and U7539 (N_7539,N_3763,N_2874);
nor U7540 (N_7540,N_1353,N_2076);
nor U7541 (N_7541,N_2284,N_1099);
nand U7542 (N_7542,N_2391,N_1236);
nand U7543 (N_7543,N_2114,N_610);
nand U7544 (N_7544,N_1231,N_352);
or U7545 (N_7545,N_1799,N_3186);
nor U7546 (N_7546,N_635,N_2571);
nor U7547 (N_7547,N_3294,N_723);
or U7548 (N_7548,N_3215,N_421);
and U7549 (N_7549,N_1753,N_3398);
nor U7550 (N_7550,N_3072,N_1844);
nor U7551 (N_7551,N_1832,N_3797);
or U7552 (N_7552,N_1881,N_1498);
or U7553 (N_7553,N_2687,N_2285);
nand U7554 (N_7554,N_1211,N_1529);
nand U7555 (N_7555,N_1082,N_2254);
and U7556 (N_7556,N_3578,N_1685);
nand U7557 (N_7557,N_1535,N_719);
nand U7558 (N_7558,N_2455,N_2291);
and U7559 (N_7559,N_2444,N_3894);
or U7560 (N_7560,N_2273,N_0);
nor U7561 (N_7561,N_774,N_3490);
and U7562 (N_7562,N_3771,N_608);
and U7563 (N_7563,N_3932,N_893);
or U7564 (N_7564,N_2016,N_664);
nand U7565 (N_7565,N_765,N_2688);
nand U7566 (N_7566,N_2265,N_3910);
nand U7567 (N_7567,N_2346,N_3626);
nand U7568 (N_7568,N_3118,N_191);
or U7569 (N_7569,N_455,N_2256);
or U7570 (N_7570,N_1644,N_3540);
nor U7571 (N_7571,N_3060,N_1168);
nor U7572 (N_7572,N_1558,N_1302);
and U7573 (N_7573,N_3490,N_2321);
and U7574 (N_7574,N_227,N_1018);
or U7575 (N_7575,N_2232,N_1246);
nor U7576 (N_7576,N_2697,N_404);
nor U7577 (N_7577,N_3355,N_441);
nand U7578 (N_7578,N_55,N_2447);
nor U7579 (N_7579,N_2206,N_3196);
nor U7580 (N_7580,N_151,N_469);
nand U7581 (N_7581,N_587,N_210);
nor U7582 (N_7582,N_538,N_424);
nor U7583 (N_7583,N_720,N_1748);
or U7584 (N_7584,N_1834,N_3824);
nor U7585 (N_7585,N_2737,N_2185);
or U7586 (N_7586,N_3339,N_3679);
nand U7587 (N_7587,N_3608,N_2496);
nor U7588 (N_7588,N_2971,N_1799);
nor U7589 (N_7589,N_1665,N_1817);
or U7590 (N_7590,N_1227,N_2553);
or U7591 (N_7591,N_1281,N_2637);
and U7592 (N_7592,N_420,N_641);
nor U7593 (N_7593,N_1950,N_1865);
or U7594 (N_7594,N_888,N_1306);
and U7595 (N_7595,N_3196,N_2082);
nor U7596 (N_7596,N_1211,N_3605);
and U7597 (N_7597,N_361,N_1709);
nand U7598 (N_7598,N_1115,N_2452);
nor U7599 (N_7599,N_2096,N_2991);
or U7600 (N_7600,N_2000,N_2751);
or U7601 (N_7601,N_3654,N_1253);
nand U7602 (N_7602,N_2225,N_809);
nand U7603 (N_7603,N_3509,N_3932);
or U7604 (N_7604,N_2474,N_3186);
and U7605 (N_7605,N_1398,N_824);
nor U7606 (N_7606,N_1840,N_280);
or U7607 (N_7607,N_3856,N_1582);
nand U7608 (N_7608,N_1507,N_1376);
or U7609 (N_7609,N_1217,N_2657);
and U7610 (N_7610,N_2622,N_330);
or U7611 (N_7611,N_373,N_1864);
nand U7612 (N_7612,N_1311,N_669);
or U7613 (N_7613,N_1149,N_1195);
nand U7614 (N_7614,N_3602,N_2328);
or U7615 (N_7615,N_2063,N_1268);
nand U7616 (N_7616,N_3111,N_1040);
nor U7617 (N_7617,N_1596,N_2151);
or U7618 (N_7618,N_3171,N_679);
nand U7619 (N_7619,N_659,N_79);
nand U7620 (N_7620,N_3432,N_2440);
nor U7621 (N_7621,N_86,N_1036);
nor U7622 (N_7622,N_148,N_2187);
and U7623 (N_7623,N_704,N_1293);
and U7624 (N_7624,N_620,N_3256);
nand U7625 (N_7625,N_2258,N_3996);
or U7626 (N_7626,N_2630,N_470);
nand U7627 (N_7627,N_3865,N_3737);
and U7628 (N_7628,N_2496,N_3414);
or U7629 (N_7629,N_2420,N_489);
or U7630 (N_7630,N_3419,N_1338);
or U7631 (N_7631,N_1708,N_2668);
and U7632 (N_7632,N_408,N_1345);
and U7633 (N_7633,N_2930,N_1850);
nand U7634 (N_7634,N_2463,N_2596);
nor U7635 (N_7635,N_934,N_754);
and U7636 (N_7636,N_2911,N_904);
nand U7637 (N_7637,N_2552,N_3454);
or U7638 (N_7638,N_2065,N_1014);
and U7639 (N_7639,N_725,N_3012);
and U7640 (N_7640,N_3388,N_3804);
xor U7641 (N_7641,N_2482,N_3275);
nor U7642 (N_7642,N_1105,N_409);
and U7643 (N_7643,N_3148,N_2826);
or U7644 (N_7644,N_1149,N_3033);
and U7645 (N_7645,N_3113,N_3702);
or U7646 (N_7646,N_1886,N_773);
or U7647 (N_7647,N_402,N_3533);
and U7648 (N_7648,N_2528,N_3817);
nor U7649 (N_7649,N_2335,N_2488);
and U7650 (N_7650,N_3259,N_734);
or U7651 (N_7651,N_2040,N_1781);
nand U7652 (N_7652,N_860,N_3147);
nand U7653 (N_7653,N_3652,N_2083);
nor U7654 (N_7654,N_593,N_861);
xnor U7655 (N_7655,N_727,N_741);
nand U7656 (N_7656,N_3796,N_3724);
or U7657 (N_7657,N_1492,N_3618);
and U7658 (N_7658,N_734,N_3638);
and U7659 (N_7659,N_3673,N_3119);
nor U7660 (N_7660,N_687,N_2223);
and U7661 (N_7661,N_1255,N_2831);
nor U7662 (N_7662,N_2476,N_559);
or U7663 (N_7663,N_1654,N_3132);
nor U7664 (N_7664,N_2389,N_2243);
nand U7665 (N_7665,N_1937,N_2027);
or U7666 (N_7666,N_592,N_3411);
and U7667 (N_7667,N_1248,N_772);
nand U7668 (N_7668,N_754,N_1015);
and U7669 (N_7669,N_645,N_2053);
and U7670 (N_7670,N_410,N_229);
or U7671 (N_7671,N_1508,N_3055);
and U7672 (N_7672,N_2553,N_2527);
and U7673 (N_7673,N_358,N_3771);
or U7674 (N_7674,N_1630,N_1129);
or U7675 (N_7675,N_1820,N_410);
and U7676 (N_7676,N_937,N_3964);
and U7677 (N_7677,N_2730,N_2101);
nor U7678 (N_7678,N_3435,N_193);
and U7679 (N_7679,N_2417,N_3428);
nand U7680 (N_7680,N_2652,N_3069);
nor U7681 (N_7681,N_1375,N_3066);
and U7682 (N_7682,N_3535,N_133);
nor U7683 (N_7683,N_892,N_514);
nand U7684 (N_7684,N_2782,N_3737);
nor U7685 (N_7685,N_2258,N_1817);
nand U7686 (N_7686,N_2284,N_3589);
nand U7687 (N_7687,N_3907,N_941);
and U7688 (N_7688,N_3147,N_959);
nand U7689 (N_7689,N_38,N_3897);
nor U7690 (N_7690,N_66,N_1370);
nand U7691 (N_7691,N_1367,N_2977);
nor U7692 (N_7692,N_1171,N_3641);
xor U7693 (N_7693,N_150,N_580);
and U7694 (N_7694,N_1845,N_2773);
and U7695 (N_7695,N_412,N_979);
nand U7696 (N_7696,N_2131,N_2530);
or U7697 (N_7697,N_1897,N_2520);
nor U7698 (N_7698,N_3941,N_3679);
xor U7699 (N_7699,N_2250,N_1327);
nor U7700 (N_7700,N_1161,N_2819);
nor U7701 (N_7701,N_2132,N_1096);
or U7702 (N_7702,N_3609,N_3497);
xnor U7703 (N_7703,N_3566,N_3232);
nand U7704 (N_7704,N_851,N_2889);
nand U7705 (N_7705,N_1349,N_2656);
nor U7706 (N_7706,N_2746,N_970);
nor U7707 (N_7707,N_3902,N_3964);
nand U7708 (N_7708,N_440,N_375);
nor U7709 (N_7709,N_3322,N_1947);
and U7710 (N_7710,N_2671,N_971);
nor U7711 (N_7711,N_1250,N_2575);
xnor U7712 (N_7712,N_3399,N_345);
or U7713 (N_7713,N_1488,N_3240);
or U7714 (N_7714,N_1873,N_244);
or U7715 (N_7715,N_3981,N_3934);
nor U7716 (N_7716,N_1544,N_671);
or U7717 (N_7717,N_1039,N_1801);
nor U7718 (N_7718,N_3958,N_2976);
nand U7719 (N_7719,N_250,N_2728);
nor U7720 (N_7720,N_3146,N_3050);
or U7721 (N_7721,N_360,N_1014);
nand U7722 (N_7722,N_3031,N_2445);
nand U7723 (N_7723,N_1795,N_2882);
and U7724 (N_7724,N_2332,N_1747);
nor U7725 (N_7725,N_1570,N_528);
nor U7726 (N_7726,N_1400,N_2716);
and U7727 (N_7727,N_1856,N_459);
nor U7728 (N_7728,N_1326,N_541);
and U7729 (N_7729,N_755,N_448);
nand U7730 (N_7730,N_2599,N_292);
and U7731 (N_7731,N_3317,N_2040);
and U7732 (N_7732,N_194,N_1031);
nor U7733 (N_7733,N_827,N_852);
xnor U7734 (N_7734,N_313,N_3450);
or U7735 (N_7735,N_1166,N_2434);
nor U7736 (N_7736,N_3299,N_2482);
or U7737 (N_7737,N_1760,N_2376);
nor U7738 (N_7738,N_631,N_3918);
nor U7739 (N_7739,N_2271,N_3020);
nand U7740 (N_7740,N_1995,N_248);
or U7741 (N_7741,N_2393,N_1540);
nor U7742 (N_7742,N_1300,N_3639);
nor U7743 (N_7743,N_1504,N_1118);
and U7744 (N_7744,N_34,N_3781);
nand U7745 (N_7745,N_667,N_2696);
or U7746 (N_7746,N_3078,N_1831);
and U7747 (N_7747,N_3693,N_959);
nand U7748 (N_7748,N_1627,N_1758);
nand U7749 (N_7749,N_1837,N_1469);
or U7750 (N_7750,N_3621,N_3762);
nand U7751 (N_7751,N_3938,N_1211);
nand U7752 (N_7752,N_3688,N_557);
nor U7753 (N_7753,N_3035,N_2307);
or U7754 (N_7754,N_2685,N_2148);
nand U7755 (N_7755,N_1371,N_3504);
and U7756 (N_7756,N_3817,N_826);
and U7757 (N_7757,N_3688,N_3449);
nand U7758 (N_7758,N_1929,N_3310);
or U7759 (N_7759,N_2601,N_3393);
nor U7760 (N_7760,N_1356,N_3641);
or U7761 (N_7761,N_2410,N_438);
nor U7762 (N_7762,N_2193,N_448);
xnor U7763 (N_7763,N_3158,N_2890);
and U7764 (N_7764,N_2581,N_2542);
or U7765 (N_7765,N_1692,N_2799);
and U7766 (N_7766,N_2158,N_2296);
nand U7767 (N_7767,N_2524,N_992);
or U7768 (N_7768,N_787,N_470);
nand U7769 (N_7769,N_2364,N_1818);
nor U7770 (N_7770,N_1692,N_1021);
nor U7771 (N_7771,N_1196,N_3538);
and U7772 (N_7772,N_3471,N_156);
nor U7773 (N_7773,N_2287,N_2784);
nand U7774 (N_7774,N_1157,N_116);
nand U7775 (N_7775,N_2296,N_1366);
nor U7776 (N_7776,N_1909,N_394);
or U7777 (N_7777,N_1598,N_2008);
and U7778 (N_7778,N_2400,N_2372);
or U7779 (N_7779,N_3902,N_9);
and U7780 (N_7780,N_1446,N_1931);
and U7781 (N_7781,N_1058,N_753);
nor U7782 (N_7782,N_2132,N_1768);
or U7783 (N_7783,N_3592,N_345);
or U7784 (N_7784,N_3193,N_23);
nand U7785 (N_7785,N_2440,N_1403);
nand U7786 (N_7786,N_510,N_3478);
nor U7787 (N_7787,N_185,N_3290);
nand U7788 (N_7788,N_785,N_1558);
and U7789 (N_7789,N_1391,N_2028);
and U7790 (N_7790,N_1347,N_928);
nand U7791 (N_7791,N_665,N_299);
nand U7792 (N_7792,N_692,N_1230);
and U7793 (N_7793,N_3276,N_3688);
and U7794 (N_7794,N_984,N_739);
or U7795 (N_7795,N_1360,N_2309);
and U7796 (N_7796,N_3216,N_1519);
or U7797 (N_7797,N_653,N_2819);
and U7798 (N_7798,N_455,N_2457);
nor U7799 (N_7799,N_2828,N_1337);
nand U7800 (N_7800,N_1848,N_2439);
or U7801 (N_7801,N_1093,N_2219);
and U7802 (N_7802,N_516,N_1819);
and U7803 (N_7803,N_3720,N_2675);
nand U7804 (N_7804,N_889,N_2379);
nand U7805 (N_7805,N_1931,N_1905);
nor U7806 (N_7806,N_2476,N_1166);
nand U7807 (N_7807,N_2229,N_2324);
and U7808 (N_7808,N_3109,N_3125);
nand U7809 (N_7809,N_3675,N_483);
and U7810 (N_7810,N_3284,N_1487);
and U7811 (N_7811,N_3975,N_19);
and U7812 (N_7812,N_771,N_3789);
nand U7813 (N_7813,N_1023,N_730);
and U7814 (N_7814,N_3887,N_3917);
and U7815 (N_7815,N_1958,N_1696);
nand U7816 (N_7816,N_3479,N_3977);
nand U7817 (N_7817,N_2971,N_318);
nor U7818 (N_7818,N_580,N_2575);
or U7819 (N_7819,N_2647,N_3132);
or U7820 (N_7820,N_3185,N_246);
nor U7821 (N_7821,N_928,N_3188);
xor U7822 (N_7822,N_3982,N_2709);
nand U7823 (N_7823,N_1850,N_2435);
or U7824 (N_7824,N_3468,N_612);
nor U7825 (N_7825,N_199,N_3096);
or U7826 (N_7826,N_3841,N_653);
nor U7827 (N_7827,N_2262,N_2568);
nand U7828 (N_7828,N_2464,N_3543);
or U7829 (N_7829,N_579,N_719);
or U7830 (N_7830,N_1107,N_3489);
or U7831 (N_7831,N_787,N_2228);
or U7832 (N_7832,N_238,N_3637);
nand U7833 (N_7833,N_139,N_3863);
or U7834 (N_7834,N_1528,N_3921);
nand U7835 (N_7835,N_644,N_1595);
nand U7836 (N_7836,N_3801,N_815);
nand U7837 (N_7837,N_1001,N_140);
or U7838 (N_7838,N_1415,N_2467);
nor U7839 (N_7839,N_3356,N_3719);
or U7840 (N_7840,N_706,N_120);
or U7841 (N_7841,N_3843,N_3992);
or U7842 (N_7842,N_1256,N_387);
nor U7843 (N_7843,N_1465,N_2034);
nand U7844 (N_7844,N_3981,N_331);
nand U7845 (N_7845,N_927,N_2567);
nand U7846 (N_7846,N_3689,N_3146);
or U7847 (N_7847,N_1378,N_3334);
and U7848 (N_7848,N_925,N_387);
or U7849 (N_7849,N_64,N_2281);
or U7850 (N_7850,N_1399,N_92);
nor U7851 (N_7851,N_3164,N_3629);
or U7852 (N_7852,N_3699,N_147);
nor U7853 (N_7853,N_3694,N_2882);
and U7854 (N_7854,N_1759,N_3240);
or U7855 (N_7855,N_3421,N_460);
nor U7856 (N_7856,N_1180,N_3115);
nand U7857 (N_7857,N_1402,N_1921);
nor U7858 (N_7858,N_3453,N_3056);
nor U7859 (N_7859,N_679,N_2190);
and U7860 (N_7860,N_3530,N_1664);
and U7861 (N_7861,N_3526,N_2388);
or U7862 (N_7862,N_1443,N_3200);
nand U7863 (N_7863,N_3329,N_1201);
and U7864 (N_7864,N_3053,N_3918);
nand U7865 (N_7865,N_1854,N_1893);
nor U7866 (N_7866,N_2463,N_1477);
or U7867 (N_7867,N_1221,N_1163);
or U7868 (N_7868,N_654,N_3377);
or U7869 (N_7869,N_2561,N_1748);
nor U7870 (N_7870,N_2489,N_1768);
nand U7871 (N_7871,N_3776,N_1148);
nand U7872 (N_7872,N_930,N_3598);
nor U7873 (N_7873,N_1010,N_1424);
nor U7874 (N_7874,N_923,N_1815);
or U7875 (N_7875,N_988,N_1953);
or U7876 (N_7876,N_1754,N_2445);
nor U7877 (N_7877,N_2524,N_704);
or U7878 (N_7878,N_1256,N_3899);
and U7879 (N_7879,N_291,N_2879);
nand U7880 (N_7880,N_3154,N_3872);
nor U7881 (N_7881,N_1819,N_1536);
nor U7882 (N_7882,N_2069,N_1851);
nor U7883 (N_7883,N_1711,N_121);
nand U7884 (N_7884,N_2538,N_570);
and U7885 (N_7885,N_575,N_215);
nor U7886 (N_7886,N_2520,N_1499);
and U7887 (N_7887,N_3063,N_73);
nand U7888 (N_7888,N_1105,N_526);
or U7889 (N_7889,N_2737,N_2771);
nor U7890 (N_7890,N_2131,N_2921);
nor U7891 (N_7891,N_2930,N_2566);
or U7892 (N_7892,N_2007,N_1676);
nand U7893 (N_7893,N_301,N_2333);
or U7894 (N_7894,N_1685,N_1922);
or U7895 (N_7895,N_1590,N_3890);
or U7896 (N_7896,N_2834,N_2052);
nor U7897 (N_7897,N_1950,N_2902);
nor U7898 (N_7898,N_3511,N_886);
nor U7899 (N_7899,N_600,N_1770);
or U7900 (N_7900,N_1760,N_2976);
nand U7901 (N_7901,N_921,N_1412);
nand U7902 (N_7902,N_2760,N_1441);
nor U7903 (N_7903,N_306,N_3497);
or U7904 (N_7904,N_3247,N_1751);
nor U7905 (N_7905,N_672,N_2936);
and U7906 (N_7906,N_3311,N_2225);
and U7907 (N_7907,N_1959,N_2763);
and U7908 (N_7908,N_942,N_1546);
nand U7909 (N_7909,N_3570,N_386);
or U7910 (N_7910,N_2038,N_851);
nand U7911 (N_7911,N_1902,N_1168);
nand U7912 (N_7912,N_1245,N_3490);
and U7913 (N_7913,N_1298,N_2383);
nand U7914 (N_7914,N_933,N_794);
nor U7915 (N_7915,N_1980,N_3165);
xor U7916 (N_7916,N_3303,N_412);
and U7917 (N_7917,N_3487,N_3337);
nor U7918 (N_7918,N_912,N_1649);
and U7919 (N_7919,N_3893,N_3252);
or U7920 (N_7920,N_2888,N_2246);
or U7921 (N_7921,N_3457,N_1165);
and U7922 (N_7922,N_161,N_777);
nor U7923 (N_7923,N_441,N_2140);
and U7924 (N_7924,N_632,N_1601);
and U7925 (N_7925,N_1989,N_3613);
nor U7926 (N_7926,N_475,N_17);
or U7927 (N_7927,N_3598,N_534);
or U7928 (N_7928,N_3262,N_119);
nand U7929 (N_7929,N_3648,N_3019);
nand U7930 (N_7930,N_163,N_2754);
or U7931 (N_7931,N_2761,N_720);
nor U7932 (N_7932,N_2524,N_3847);
nor U7933 (N_7933,N_1154,N_1735);
and U7934 (N_7934,N_1138,N_1266);
or U7935 (N_7935,N_2804,N_1223);
nor U7936 (N_7936,N_113,N_3286);
nand U7937 (N_7937,N_62,N_783);
nor U7938 (N_7938,N_3697,N_1253);
and U7939 (N_7939,N_3421,N_3992);
or U7940 (N_7940,N_2040,N_1443);
and U7941 (N_7941,N_1076,N_3825);
nand U7942 (N_7942,N_3590,N_2806);
nand U7943 (N_7943,N_3985,N_1550);
nand U7944 (N_7944,N_2183,N_3957);
nor U7945 (N_7945,N_3850,N_3114);
nand U7946 (N_7946,N_3533,N_787);
or U7947 (N_7947,N_192,N_1758);
nor U7948 (N_7948,N_1777,N_1940);
nand U7949 (N_7949,N_2346,N_913);
nand U7950 (N_7950,N_828,N_2478);
or U7951 (N_7951,N_3457,N_2289);
nor U7952 (N_7952,N_536,N_1745);
xnor U7953 (N_7953,N_900,N_548);
nor U7954 (N_7954,N_2181,N_1614);
nor U7955 (N_7955,N_704,N_288);
nand U7956 (N_7956,N_1741,N_1719);
nand U7957 (N_7957,N_692,N_3604);
and U7958 (N_7958,N_3012,N_2276);
nand U7959 (N_7959,N_1245,N_73);
or U7960 (N_7960,N_3441,N_1081);
nor U7961 (N_7961,N_852,N_926);
nor U7962 (N_7962,N_1708,N_1072);
nor U7963 (N_7963,N_2765,N_1245);
nor U7964 (N_7964,N_3568,N_1761);
nand U7965 (N_7965,N_914,N_1686);
nand U7966 (N_7966,N_1367,N_460);
nor U7967 (N_7967,N_2955,N_1289);
nand U7968 (N_7968,N_2756,N_2933);
and U7969 (N_7969,N_2636,N_2012);
and U7970 (N_7970,N_3515,N_945);
or U7971 (N_7971,N_1853,N_3155);
and U7972 (N_7972,N_2498,N_259);
nor U7973 (N_7973,N_1564,N_1492);
or U7974 (N_7974,N_1269,N_3958);
nand U7975 (N_7975,N_3800,N_1378);
nor U7976 (N_7976,N_1957,N_160);
and U7977 (N_7977,N_1049,N_1402);
and U7978 (N_7978,N_739,N_803);
nor U7979 (N_7979,N_3859,N_2363);
nor U7980 (N_7980,N_1624,N_2453);
nand U7981 (N_7981,N_469,N_3717);
and U7982 (N_7982,N_535,N_2915);
or U7983 (N_7983,N_1066,N_910);
nor U7984 (N_7984,N_3356,N_3698);
or U7985 (N_7985,N_1528,N_463);
nand U7986 (N_7986,N_1833,N_2176);
nor U7987 (N_7987,N_1946,N_804);
or U7988 (N_7988,N_2045,N_2430);
or U7989 (N_7989,N_2476,N_2990);
or U7990 (N_7990,N_3868,N_3129);
nor U7991 (N_7991,N_2809,N_1752);
nor U7992 (N_7992,N_517,N_1862);
nor U7993 (N_7993,N_775,N_3663);
nand U7994 (N_7994,N_2797,N_2267);
and U7995 (N_7995,N_1139,N_1410);
and U7996 (N_7996,N_2085,N_324);
nand U7997 (N_7997,N_3037,N_3534);
nand U7998 (N_7998,N_436,N_2009);
nand U7999 (N_7999,N_730,N_1419);
and U8000 (N_8000,N_6860,N_7787);
and U8001 (N_8001,N_7904,N_5174);
nor U8002 (N_8002,N_4881,N_5649);
nand U8003 (N_8003,N_5757,N_4985);
or U8004 (N_8004,N_7750,N_6804);
or U8005 (N_8005,N_6831,N_5761);
nand U8006 (N_8006,N_4840,N_7994);
nand U8007 (N_8007,N_4649,N_6020);
nor U8008 (N_8008,N_7114,N_6569);
nor U8009 (N_8009,N_7394,N_7215);
and U8010 (N_8010,N_4213,N_4344);
nand U8011 (N_8011,N_4000,N_6941);
or U8012 (N_8012,N_5229,N_6885);
and U8013 (N_8013,N_7222,N_5596);
nor U8014 (N_8014,N_6062,N_5656);
or U8015 (N_8015,N_5218,N_6698);
or U8016 (N_8016,N_5186,N_6963);
or U8017 (N_8017,N_7213,N_7855);
or U8018 (N_8018,N_6735,N_7118);
or U8019 (N_8019,N_7637,N_5880);
and U8020 (N_8020,N_4694,N_5549);
or U8021 (N_8021,N_6081,N_7751);
and U8022 (N_8022,N_4369,N_5489);
or U8023 (N_8023,N_6503,N_5758);
nand U8024 (N_8024,N_6111,N_5230);
nor U8025 (N_8025,N_4681,N_4025);
or U8026 (N_8026,N_5414,N_7798);
nand U8027 (N_8027,N_7683,N_6093);
nand U8028 (N_8028,N_7032,N_6934);
and U8029 (N_8029,N_5665,N_4218);
or U8030 (N_8030,N_7916,N_7599);
nand U8031 (N_8031,N_5578,N_7077);
and U8032 (N_8032,N_7703,N_6590);
and U8033 (N_8033,N_6059,N_6468);
and U8034 (N_8034,N_4393,N_4342);
nand U8035 (N_8035,N_5553,N_4550);
or U8036 (N_8036,N_5144,N_6067);
nor U8037 (N_8037,N_7565,N_7176);
nand U8038 (N_8038,N_5477,N_6178);
nor U8039 (N_8039,N_4933,N_4440);
nor U8040 (N_8040,N_4276,N_4825);
nand U8041 (N_8041,N_7341,N_7296);
nor U8042 (N_8042,N_5251,N_7762);
or U8043 (N_8043,N_6460,N_7854);
or U8044 (N_8044,N_6207,N_5001);
nor U8045 (N_8045,N_5211,N_7616);
or U8046 (N_8046,N_6088,N_7698);
nand U8047 (N_8047,N_7123,N_6034);
nand U8048 (N_8048,N_6136,N_6216);
nand U8049 (N_8049,N_7397,N_7321);
and U8050 (N_8050,N_7194,N_5637);
nand U8051 (N_8051,N_6398,N_7314);
nor U8052 (N_8052,N_4786,N_6488);
and U8053 (N_8053,N_7808,N_7187);
nor U8054 (N_8054,N_4208,N_6624);
nor U8055 (N_8055,N_6445,N_7468);
nor U8056 (N_8056,N_6104,N_4051);
nand U8057 (N_8057,N_6800,N_6975);
and U8058 (N_8058,N_6637,N_6461);
nand U8059 (N_8059,N_6899,N_7426);
nand U8060 (N_8060,N_4711,N_4511);
and U8061 (N_8061,N_6415,N_4596);
and U8062 (N_8062,N_6879,N_7151);
nor U8063 (N_8063,N_5690,N_4905);
xnor U8064 (N_8064,N_6039,N_4376);
and U8065 (N_8065,N_5160,N_7046);
nand U8066 (N_8066,N_4091,N_5399);
and U8067 (N_8067,N_4613,N_5616);
nor U8068 (N_8068,N_6709,N_7582);
nand U8069 (N_8069,N_7066,N_5600);
nor U8070 (N_8070,N_6772,N_4003);
nand U8071 (N_8071,N_4193,N_7635);
or U8072 (N_8072,N_6725,N_5082);
nand U8073 (N_8073,N_5599,N_5155);
or U8074 (N_8074,N_7210,N_5954);
and U8075 (N_8075,N_4332,N_5793);
nor U8076 (N_8076,N_5413,N_5460);
nor U8077 (N_8077,N_5928,N_4124);
and U8078 (N_8078,N_6898,N_7303);
nand U8079 (N_8079,N_4976,N_6965);
nor U8080 (N_8080,N_6385,N_6563);
nand U8081 (N_8081,N_5106,N_4549);
or U8082 (N_8082,N_4456,N_7668);
nand U8083 (N_8083,N_4484,N_6537);
or U8084 (N_8084,N_7769,N_7116);
nand U8085 (N_8085,N_6937,N_6349);
and U8086 (N_8086,N_7970,N_6049);
nand U8087 (N_8087,N_4210,N_6674);
nor U8088 (N_8088,N_6376,N_6351);
and U8089 (N_8089,N_6274,N_5712);
and U8090 (N_8090,N_6163,N_7773);
nor U8091 (N_8091,N_6213,N_6528);
or U8092 (N_8092,N_4837,N_6949);
nor U8093 (N_8093,N_7083,N_4648);
nor U8094 (N_8094,N_5499,N_4771);
nor U8095 (N_8095,N_7090,N_6966);
nand U8096 (N_8096,N_4064,N_6433);
nor U8097 (N_8097,N_5012,N_7880);
and U8098 (N_8098,N_7913,N_6337);
or U8099 (N_8099,N_4716,N_4886);
and U8100 (N_8100,N_6521,N_7596);
nor U8101 (N_8101,N_7955,N_6515);
nor U8102 (N_8102,N_6310,N_7792);
or U8103 (N_8103,N_4253,N_4423);
nand U8104 (N_8104,N_6419,N_5925);
nand U8105 (N_8105,N_6620,N_4274);
nand U8106 (N_8106,N_7575,N_4975);
nand U8107 (N_8107,N_6649,N_7659);
or U8108 (N_8108,N_5114,N_5347);
nand U8109 (N_8109,N_5848,N_4250);
nand U8110 (N_8110,N_4008,N_4726);
nand U8111 (N_8111,N_5977,N_5785);
nor U8112 (N_8112,N_6380,N_5754);
nor U8113 (N_8113,N_4535,N_5492);
and U8114 (N_8114,N_5854,N_4782);
or U8115 (N_8115,N_4357,N_4979);
or U8116 (N_8116,N_6580,N_7950);
nor U8117 (N_8117,N_6648,N_4912);
nor U8118 (N_8118,N_6399,N_7841);
nand U8119 (N_8119,N_7137,N_5339);
and U8120 (N_8120,N_4058,N_7931);
nand U8121 (N_8121,N_4972,N_6016);
and U8122 (N_8122,N_4690,N_5225);
and U8123 (N_8123,N_5070,N_6742);
nor U8124 (N_8124,N_4134,N_6044);
nand U8125 (N_8125,N_7814,N_7153);
and U8126 (N_8126,N_4426,N_7908);
or U8127 (N_8127,N_5372,N_7622);
nand U8128 (N_8128,N_6317,N_4103);
nand U8129 (N_8129,N_7172,N_6440);
and U8130 (N_8130,N_6366,N_5691);
nor U8131 (N_8131,N_7856,N_6409);
nor U8132 (N_8132,N_4620,N_7593);
or U8133 (N_8133,N_5828,N_6189);
nor U8134 (N_8134,N_7337,N_5165);
or U8135 (N_8135,N_5159,N_6751);
and U8136 (N_8136,N_5940,N_6245);
nor U8137 (N_8137,N_7544,N_4927);
nand U8138 (N_8138,N_4278,N_6237);
nand U8139 (N_8139,N_4396,N_7483);
nor U8140 (N_8140,N_4849,N_7382);
and U8141 (N_8141,N_5411,N_6623);
nor U8142 (N_8142,N_5102,N_4759);
nor U8143 (N_8143,N_5836,N_6434);
xnor U8144 (N_8144,N_6268,N_4523);
nand U8145 (N_8145,N_4340,N_5993);
nand U8146 (N_8146,N_7155,N_7470);
and U8147 (N_8147,N_6630,N_5167);
nand U8148 (N_8148,N_6747,N_4778);
and U8149 (N_8149,N_6917,N_7467);
and U8150 (N_8150,N_6548,N_4071);
nor U8151 (N_8151,N_5926,N_4546);
and U8152 (N_8152,N_6066,N_6718);
nand U8153 (N_8153,N_6706,N_7237);
nor U8154 (N_8154,N_7371,N_7358);
and U8155 (N_8155,N_5528,N_7523);
and U8156 (N_8156,N_4413,N_6824);
nand U8157 (N_8157,N_7121,N_6991);
nand U8158 (N_8158,N_4223,N_5502);
or U8159 (N_8159,N_6462,N_7474);
nor U8160 (N_8160,N_6651,N_4528);
nand U8161 (N_8161,N_6631,N_4816);
nand U8162 (N_8162,N_5279,N_6668);
nand U8163 (N_8163,N_4202,N_7852);
and U8164 (N_8164,N_5272,N_7402);
nand U8165 (N_8165,N_7869,N_6484);
nor U8166 (N_8166,N_5356,N_5135);
or U8167 (N_8167,N_4035,N_7369);
and U8168 (N_8168,N_7064,N_7475);
or U8169 (N_8169,N_7966,N_4317);
nor U8170 (N_8170,N_4285,N_5000);
nor U8171 (N_8171,N_5980,N_4920);
nor U8172 (N_8172,N_4536,N_4473);
or U8173 (N_8173,N_4352,N_7859);
and U8174 (N_8174,N_7251,N_5516);
nor U8175 (N_8175,N_6865,N_5810);
or U8176 (N_8176,N_7407,N_6888);
or U8177 (N_8177,N_4329,N_7995);
or U8178 (N_8178,N_4339,N_4733);
and U8179 (N_8179,N_6615,N_6300);
nand U8180 (N_8180,N_5444,N_4204);
nor U8181 (N_8181,N_5935,N_4950);
or U8182 (N_8182,N_5254,N_7516);
nor U8183 (N_8183,N_5608,N_6307);
nand U8184 (N_8184,N_7150,N_7858);
nand U8185 (N_8185,N_5455,N_5929);
and U8186 (N_8186,N_7466,N_4039);
and U8187 (N_8187,N_7364,N_5800);
or U8188 (N_8188,N_6301,N_7221);
or U8189 (N_8189,N_5282,N_5551);
nand U8190 (N_8190,N_4921,N_4990);
xnor U8191 (N_8191,N_7811,N_5393);
and U8192 (N_8192,N_6056,N_6732);
nor U8193 (N_8193,N_5451,N_4491);
nor U8194 (N_8194,N_4954,N_5344);
nand U8195 (N_8195,N_4043,N_7202);
nor U8196 (N_8196,N_5873,N_7008);
or U8197 (N_8197,N_7310,N_7585);
and U8198 (N_8198,N_5735,N_6295);
nor U8199 (N_8199,N_4970,N_7343);
and U8200 (N_8200,N_7646,N_6203);
nor U8201 (N_8201,N_7249,N_7765);
nor U8202 (N_8202,N_4389,N_5002);
or U8203 (N_8203,N_5483,N_6959);
or U8204 (N_8204,N_6856,N_4459);
nand U8205 (N_8205,N_4320,N_7193);
nand U8206 (N_8206,N_4655,N_6903);
and U8207 (N_8207,N_5052,N_7777);
and U8208 (N_8208,N_6240,N_4662);
nand U8209 (N_8209,N_5999,N_5410);
and U8210 (N_8210,N_6555,N_7772);
nand U8211 (N_8211,N_7556,N_6578);
nand U8212 (N_8212,N_7721,N_5972);
nor U8213 (N_8213,N_4443,N_6810);
and U8214 (N_8214,N_4852,N_4241);
nand U8215 (N_8215,N_5907,N_6101);
and U8216 (N_8216,N_4330,N_6769);
nand U8217 (N_8217,N_4495,N_5952);
or U8218 (N_8218,N_5653,N_5258);
or U8219 (N_8219,N_6184,N_4448);
nor U8220 (N_8220,N_4643,N_6471);
nor U8221 (N_8221,N_5922,N_6633);
nand U8222 (N_8222,N_7224,N_4179);
nor U8223 (N_8223,N_7685,N_4358);
and U8224 (N_8224,N_7590,N_5369);
nand U8225 (N_8225,N_4020,N_6100);
and U8226 (N_8226,N_4909,N_6680);
and U8227 (N_8227,N_7619,N_5299);
nand U8228 (N_8228,N_4719,N_5732);
nor U8229 (N_8229,N_4573,N_6156);
or U8230 (N_8230,N_4299,N_7633);
or U8231 (N_8231,N_7051,N_4186);
nor U8232 (N_8232,N_6004,N_5721);
nand U8233 (N_8233,N_7356,N_5287);
and U8234 (N_8234,N_6738,N_5425);
or U8235 (N_8235,N_5090,N_6996);
nand U8236 (N_8236,N_5728,N_7020);
and U8237 (N_8237,N_6140,N_5522);
nor U8238 (N_8238,N_5775,N_6513);
and U8239 (N_8239,N_4854,N_4054);
nor U8240 (N_8240,N_7197,N_7133);
nand U8241 (N_8241,N_5659,N_7812);
nand U8242 (N_8242,N_7420,N_6935);
and U8243 (N_8243,N_6449,N_5564);
nor U8244 (N_8244,N_6343,N_5998);
nand U8245 (N_8245,N_6318,N_4458);
or U8246 (N_8246,N_4752,N_6597);
nor U8247 (N_8247,N_6873,N_4325);
nor U8248 (N_8248,N_4705,N_6582);
nor U8249 (N_8249,N_4031,N_7152);
and U8250 (N_8250,N_4034,N_7447);
nor U8251 (N_8251,N_5835,N_5724);
nand U8252 (N_8252,N_4296,N_5628);
nand U8253 (N_8253,N_6962,N_4206);
nand U8254 (N_8254,N_6008,N_4140);
and U8255 (N_8255,N_6608,N_5651);
and U8256 (N_8256,N_4216,N_6520);
nor U8257 (N_8257,N_7649,N_7952);
nor U8258 (N_8258,N_4085,N_6566);
nand U8259 (N_8259,N_4370,N_5910);
or U8260 (N_8260,N_4552,N_5196);
and U8261 (N_8261,N_4670,N_5898);
nand U8262 (N_8262,N_6906,N_4621);
and U8263 (N_8263,N_5717,N_5971);
xnor U8264 (N_8264,N_4373,N_6269);
nor U8265 (N_8265,N_4251,N_7824);
nor U8266 (N_8266,N_6667,N_7126);
and U8267 (N_8267,N_7177,N_5085);
nand U8268 (N_8268,N_5139,N_5981);
nand U8269 (N_8269,N_5037,N_7156);
and U8270 (N_8270,N_4505,N_7315);
or U8271 (N_8271,N_4326,N_5015);
or U8272 (N_8272,N_5213,N_7240);
and U8273 (N_8273,N_5725,N_6206);
and U8274 (N_8274,N_4539,N_5541);
xor U8275 (N_8275,N_7910,N_4403);
nor U8276 (N_8276,N_5358,N_5953);
nand U8277 (N_8277,N_4214,N_6276);
and U8278 (N_8278,N_4499,N_4823);
or U8279 (N_8279,N_4321,N_6666);
or U8280 (N_8280,N_5141,N_4334);
nand U8281 (N_8281,N_7429,N_5367);
nand U8282 (N_8282,N_4835,N_5113);
nor U8283 (N_8283,N_6129,N_4591);
and U8284 (N_8284,N_6767,N_7014);
and U8285 (N_8285,N_7306,N_5171);
nor U8286 (N_8286,N_4521,N_7398);
or U8287 (N_8287,N_4864,N_6086);
nand U8288 (N_8288,N_4319,N_5116);
nor U8289 (N_8289,N_4481,N_4520);
or U8290 (N_8290,N_5920,N_7778);
nor U8291 (N_8291,N_7862,N_5666);
nor U8292 (N_8292,N_6703,N_6985);
and U8293 (N_8293,N_7362,N_6181);
nand U8294 (N_8294,N_4745,N_5058);
nor U8295 (N_8295,N_4502,N_4693);
and U8296 (N_8296,N_4130,N_5812);
or U8297 (N_8297,N_6055,N_7530);
or U8298 (N_8298,N_4887,N_5603);
nor U8299 (N_8299,N_7641,N_7609);
or U8300 (N_8300,N_5719,N_5346);
nand U8301 (N_8301,N_7050,N_6371);
and U8302 (N_8302,N_5654,N_6726);
or U8303 (N_8303,N_7360,N_4347);
or U8304 (N_8304,N_5049,N_4906);
nor U8305 (N_8305,N_7879,N_4984);
nand U8306 (N_8306,N_5019,N_5901);
and U8307 (N_8307,N_5678,N_5267);
or U8308 (N_8308,N_5777,N_7361);
nor U8309 (N_8309,N_7623,N_7159);
nor U8310 (N_8310,N_6496,N_7891);
and U8311 (N_8311,N_6697,N_4534);
nor U8312 (N_8312,N_4245,N_7374);
nand U8313 (N_8313,N_6614,N_5166);
nor U8314 (N_8314,N_5945,N_7104);
or U8315 (N_8315,N_7431,N_5805);
and U8316 (N_8316,N_7553,N_7686);
and U8317 (N_8317,N_4683,N_6143);
nand U8318 (N_8318,N_5244,N_6524);
nor U8319 (N_8319,N_5066,N_4472);
or U8320 (N_8320,N_4100,N_4266);
and U8321 (N_8321,N_7632,N_6723);
nand U8322 (N_8322,N_5210,N_7250);
nand U8323 (N_8323,N_5479,N_7831);
nand U8324 (N_8324,N_5786,N_7018);
nor U8325 (N_8325,N_5547,N_7044);
and U8326 (N_8326,N_5905,N_6737);
and U8327 (N_8327,N_6481,N_5632);
and U8328 (N_8328,N_6822,N_4437);
nor U8329 (N_8329,N_4163,N_7849);
nand U8330 (N_8330,N_7330,N_6739);
nor U8331 (N_8331,N_6116,N_4496);
or U8332 (N_8332,N_4259,N_7112);
and U8333 (N_8333,N_6979,N_4112);
and U8334 (N_8334,N_7851,N_7333);
nor U8335 (N_8335,N_4601,N_5017);
and U8336 (N_8336,N_7318,N_6716);
or U8337 (N_8337,N_6227,N_4217);
and U8338 (N_8338,N_4780,N_4430);
xor U8339 (N_8339,N_5512,N_4879);
nor U8340 (N_8340,N_6131,N_6830);
nand U8341 (N_8341,N_7372,N_6685);
and U8342 (N_8342,N_7975,N_5041);
nor U8343 (N_8343,N_7456,N_5426);
or U8344 (N_8344,N_7500,N_6816);
and U8345 (N_8345,N_5673,N_7166);
nand U8346 (N_8346,N_7157,N_6015);
nor U8347 (N_8347,N_4850,N_4501);
or U8348 (N_8348,N_4736,N_4627);
nor U8349 (N_8349,N_4148,N_4857);
and U8350 (N_8350,N_7907,N_5860);
nand U8351 (N_8351,N_5055,N_7503);
or U8352 (N_8352,N_6893,N_6541);
nand U8353 (N_8353,N_4009,N_7411);
and U8354 (N_8354,N_4172,N_5310);
xor U8355 (N_8355,N_6426,N_4615);
nor U8356 (N_8356,N_5759,N_4853);
nor U8357 (N_8357,N_6525,N_7457);
nand U8358 (N_8358,N_6644,N_5028);
nor U8359 (N_8359,N_5449,N_5417);
and U8360 (N_8360,N_5474,N_6785);
xnor U8361 (N_8361,N_7232,N_4305);
nor U8362 (N_8362,N_5527,N_4399);
nand U8363 (N_8363,N_7746,N_6900);
and U8364 (N_8364,N_5996,N_7007);
and U8365 (N_8365,N_4754,N_6316);
or U8366 (N_8366,N_5190,N_7983);
and U8367 (N_8367,N_6846,N_6042);
or U8368 (N_8368,N_5014,N_6545);
nand U8369 (N_8369,N_6378,N_6479);
and U8370 (N_8370,N_6612,N_5223);
or U8371 (N_8371,N_7185,N_7980);
nor U8372 (N_8372,N_4303,N_4181);
and U8373 (N_8373,N_4311,N_4135);
nor U8374 (N_8374,N_5872,N_7233);
nor U8375 (N_8375,N_5164,N_5534);
and U8376 (N_8376,N_4384,N_7549);
nor U8377 (N_8377,N_5330,N_7900);
and U8378 (N_8378,N_7796,N_6263);
or U8379 (N_8379,N_5386,N_4557);
or U8380 (N_8380,N_7675,N_5079);
nor U8381 (N_8381,N_7996,N_6625);
or U8382 (N_8382,N_4519,N_7028);
nand U8383 (N_8383,N_7822,N_4318);
or U8384 (N_8384,N_4488,N_5312);
nor U8385 (N_8385,N_4758,N_5695);
nor U8386 (N_8386,N_7557,N_4232);
or U8387 (N_8387,N_4947,N_4783);
or U8388 (N_8388,N_7282,N_7508);
nand U8389 (N_8389,N_5882,N_5480);
nand U8390 (N_8390,N_6741,N_5365);
or U8391 (N_8391,N_4692,N_6601);
or U8392 (N_8392,N_6880,N_6549);
nand U8393 (N_8393,N_6872,N_7510);
nor U8394 (N_8394,N_5622,N_4556);
or U8395 (N_8395,N_7903,N_6094);
nor U8396 (N_8396,N_7894,N_4993);
or U8397 (N_8397,N_6466,N_7419);
and U8398 (N_8398,N_4848,N_4061);
nor U8399 (N_8399,N_4514,N_7347);
or U8400 (N_8400,N_6339,N_7267);
and U8401 (N_8401,N_5422,N_4587);
nor U8402 (N_8402,N_7953,N_6596);
and U8403 (N_8403,N_5948,N_7489);
nor U8404 (N_8404,N_6895,N_5539);
nor U8405 (N_8405,N_4688,N_7352);
or U8406 (N_8406,N_5032,N_4885);
or U8407 (N_8407,N_4616,N_7179);
nor U8408 (N_8408,N_4504,N_5518);
and U8409 (N_8409,N_5183,N_6807);
or U8410 (N_8410,N_7208,N_4657);
nor U8411 (N_8411,N_6095,N_7705);
nand U8412 (N_8412,N_7766,N_6878);
and U8413 (N_8413,N_6091,N_6740);
and U8414 (N_8414,N_7063,N_4784);
or U8415 (N_8415,N_4966,N_5217);
nand U8416 (N_8416,N_5380,N_7963);
and U8417 (N_8417,N_6050,N_7048);
or U8418 (N_8418,N_4343,N_4660);
or U8419 (N_8419,N_6491,N_4184);
nor U8420 (N_8420,N_4236,N_7482);
or U8421 (N_8421,N_4830,N_5611);
or U8422 (N_8422,N_4331,N_5189);
or U8423 (N_8423,N_4569,N_5962);
and U8424 (N_8424,N_7485,N_4199);
or U8425 (N_8425,N_5787,N_5069);
or U8426 (N_8426,N_6711,N_4027);
or U8427 (N_8427,N_5104,N_7513);
nor U8428 (N_8428,N_5441,N_7265);
and U8429 (N_8429,N_6406,N_6565);
nand U8430 (N_8430,N_4412,N_6286);
nor U8431 (N_8431,N_7477,N_4858);
or U8432 (N_8432,N_5080,N_4012);
or U8433 (N_8433,N_6818,N_7829);
and U8434 (N_8434,N_7459,N_7570);
or U8435 (N_8435,N_4076,N_6334);
or U8436 (N_8436,N_5643,N_6705);
nor U8437 (N_8437,N_6600,N_7514);
or U8438 (N_8438,N_6588,N_6388);
nand U8439 (N_8439,N_7386,N_5784);
and U8440 (N_8440,N_4165,N_4659);
or U8441 (N_8441,N_5874,N_6108);
nand U8442 (N_8442,N_5550,N_5222);
or U8443 (N_8443,N_6914,N_6944);
nand U8444 (N_8444,N_6238,N_6106);
or U8445 (N_8445,N_6744,N_7892);
and U8446 (N_8446,N_6704,N_7947);
nand U8447 (N_8447,N_5206,N_4903);
nor U8448 (N_8448,N_5525,N_6325);
nor U8449 (N_8449,N_4682,N_6423);
and U8450 (N_8450,N_5604,N_6876);
or U8451 (N_8451,N_6158,N_6657);
nor U8452 (N_8452,N_7257,N_6511);
nand U8453 (N_8453,N_7001,N_5228);
or U8454 (N_8454,N_6562,N_4518);
or U8455 (N_8455,N_5974,N_5313);
nor U8456 (N_8456,N_5892,N_6407);
nor U8457 (N_8457,N_5143,N_5679);
nand U8458 (N_8458,N_4701,N_6688);
nand U8459 (N_8459,N_6862,N_4777);
nor U8460 (N_8460,N_5542,N_4781);
nand U8461 (N_8461,N_4767,N_6877);
nand U8462 (N_8462,N_7587,N_7367);
and U8463 (N_8463,N_4271,N_7010);
nand U8464 (N_8464,N_4255,N_4605);
and U8465 (N_8465,N_7143,N_5245);
nand U8466 (N_8466,N_6646,N_4588);
nor U8467 (N_8467,N_5086,N_5884);
nor U8468 (N_8468,N_7785,N_4564);
and U8469 (N_8469,N_5877,N_5073);
or U8470 (N_8470,N_6841,N_6572);
and U8471 (N_8471,N_7899,N_6027);
and U8472 (N_8472,N_7478,N_5484);
and U8473 (N_8473,N_4364,N_7075);
nand U8474 (N_8474,N_6714,N_4871);
nor U8475 (N_8475,N_5598,N_7370);
nand U8476 (N_8476,N_7334,N_6721);
and U8477 (N_8477,N_6169,N_7793);
nor U8478 (N_8478,N_4914,N_5683);
nand U8479 (N_8479,N_5231,N_5033);
or U8480 (N_8480,N_4454,N_6743);
nand U8481 (N_8481,N_7375,N_4575);
and U8482 (N_8482,N_4590,N_4151);
or U8483 (N_8483,N_7989,N_6281);
or U8484 (N_8484,N_5689,N_5638);
and U8485 (N_8485,N_6874,N_7759);
nand U8486 (N_8486,N_5772,N_4592);
nand U8487 (N_8487,N_4227,N_4866);
and U8488 (N_8488,N_6950,N_4312);
nor U8489 (N_8489,N_7833,N_7231);
or U8490 (N_8490,N_6060,N_4467);
nor U8491 (N_8491,N_5519,N_5768);
and U8492 (N_8492,N_7928,N_4397);
nand U8493 (N_8493,N_6369,N_7325);
nor U8494 (N_8494,N_4589,N_7211);
nor U8495 (N_8495,N_6478,N_5341);
nand U8496 (N_8496,N_7624,N_5890);
nor U8497 (N_8497,N_4943,N_4308);
or U8498 (N_8498,N_6465,N_7584);
nor U8499 (N_8499,N_6282,N_5390);
nand U8500 (N_8500,N_5490,N_7640);
or U8501 (N_8501,N_7129,N_7427);
and U8502 (N_8502,N_7068,N_7089);
nor U8503 (N_8503,N_5389,N_6639);
or U8504 (N_8504,N_5606,N_6581);
nor U8505 (N_8505,N_6558,N_6535);
and U8506 (N_8506,N_6353,N_4964);
and U8507 (N_8507,N_7052,N_7284);
or U8508 (N_8508,N_7768,N_5852);
nor U8509 (N_8509,N_4656,N_4626);
nor U8510 (N_8510,N_7122,N_5841);
nor U8511 (N_8511,N_5685,N_6538);
or U8512 (N_8512,N_7422,N_6997);
and U8513 (N_8513,N_4333,N_7648);
or U8514 (N_8514,N_6375,N_5625);
and U8515 (N_8515,N_4558,N_7460);
or U8516 (N_8516,N_7758,N_5241);
or U8517 (N_8517,N_5428,N_7586);
and U8518 (N_8518,N_6137,N_4429);
nor U8519 (N_8519,N_5736,N_4961);
nor U8520 (N_8520,N_4439,N_6041);
or U8521 (N_8521,N_6075,N_4161);
nor U8522 (N_8522,N_6082,N_6319);
and U8523 (N_8523,N_6662,N_6686);
nand U8524 (N_8524,N_4597,N_5957);
nor U8525 (N_8525,N_4538,N_6180);
and U8526 (N_8526,N_7026,N_7340);
nand U8527 (N_8527,N_6995,N_5595);
nand U8528 (N_8528,N_6437,N_4102);
or U8529 (N_8529,N_6463,N_6218);
and U8530 (N_8530,N_6670,N_7102);
and U8531 (N_8531,N_6809,N_7543);
nand U8532 (N_8532,N_5081,N_5464);
and U8533 (N_8533,N_5232,N_7932);
and U8534 (N_8534,N_6724,N_7276);
nand U8535 (N_8535,N_7304,N_4740);
or U8536 (N_8536,N_5896,N_4060);
nand U8537 (N_8537,N_7368,N_5212);
nand U8538 (N_8538,N_6185,N_4045);
nor U8539 (N_8539,N_5983,N_4418);
nor U8540 (N_8540,N_7441,N_6892);
nand U8541 (N_8541,N_5684,N_5481);
nor U8542 (N_8542,N_4930,N_6146);
or U8543 (N_8543,N_5457,N_5302);
or U8544 (N_8544,N_6789,N_7711);
or U8545 (N_8545,N_5915,N_4883);
and U8546 (N_8546,N_7967,N_5126);
and U8547 (N_8547,N_4451,N_5989);
and U8548 (N_8548,N_5323,N_6064);
or U8549 (N_8549,N_7732,N_6190);
and U8550 (N_8550,N_5558,N_7079);
or U8551 (N_8551,N_4956,N_6540);
and U8552 (N_8552,N_5024,N_4992);
or U8553 (N_8553,N_5237,N_5048);
nand U8554 (N_8554,N_5388,N_5209);
nand U8555 (N_8555,N_7597,N_5994);
nand U8556 (N_8556,N_6978,N_7308);
and U8557 (N_8557,N_7699,N_7499);
or U8558 (N_8558,N_4667,N_4050);
nor U8559 (N_8559,N_7702,N_5091);
or U8560 (N_8560,N_6530,N_5292);
and U8561 (N_8561,N_6457,N_5508);
nand U8562 (N_8562,N_4028,N_4220);
nor U8563 (N_8563,N_4962,N_6354);
xor U8564 (N_8564,N_7610,N_6172);
and U8565 (N_8565,N_5491,N_6359);
or U8566 (N_8566,N_5511,N_5343);
nand U8567 (N_8567,N_4424,N_4194);
or U8568 (N_8568,N_4322,N_4324);
or U8569 (N_8569,N_6090,N_7918);
nand U8570 (N_8570,N_6261,N_7244);
nor U8571 (N_8571,N_6661,N_5587);
and U8572 (N_8572,N_4841,N_6840);
or U8573 (N_8573,N_7322,N_5939);
nor U8574 (N_8574,N_5566,N_4249);
nand U8575 (N_8575,N_6915,N_7815);
and U8576 (N_8576,N_5710,N_5010);
or U8577 (N_8577,N_7025,N_5875);
nand U8578 (N_8578,N_6473,N_4828);
nand U8579 (N_8579,N_5976,N_4428);
and U8580 (N_8580,N_7542,N_4486);
or U8581 (N_8581,N_7978,N_5722);
nand U8582 (N_8582,N_6539,N_6073);
nand U8583 (N_8583,N_7103,N_4554);
and U8584 (N_8584,N_5615,N_4047);
or U8585 (N_8585,N_6194,N_6749);
and U8586 (N_8586,N_6838,N_6547);
nand U8587 (N_8587,N_4599,N_5328);
and U8588 (N_8588,N_5593,N_4803);
nand U8589 (N_8589,N_7348,N_7909);
and U8590 (N_8590,N_5713,N_5973);
or U8591 (N_8591,N_4476,N_5133);
and U8592 (N_8592,N_6855,N_7830);
nor U8593 (N_8593,N_4863,N_6235);
and U8594 (N_8594,N_6654,N_7576);
and U8595 (N_8595,N_7607,N_7444);
nor U8596 (N_8596,N_4700,N_4444);
and U8597 (N_8597,N_4477,N_4177);
and U8598 (N_8598,N_7782,N_6322);
xor U8599 (N_8599,N_6208,N_6160);
nand U8600 (N_8600,N_6036,N_4049);
nand U8601 (N_8601,N_5715,N_7404);
or U8602 (N_8602,N_7943,N_6610);
and U8603 (N_8603,N_4182,N_6288);
nand U8604 (N_8604,N_7658,N_4658);
and U8605 (N_8605,N_7307,N_4545);
nand U8606 (N_8606,N_7455,N_4731);
nand U8607 (N_8607,N_6621,N_7412);
xnor U8608 (N_8608,N_4088,N_7248);
or U8609 (N_8609,N_4982,N_4704);
nor U8610 (N_8610,N_7449,N_6258);
nor U8611 (N_8611,N_6727,N_7689);
nand U8612 (N_8612,N_7255,N_7071);
or U8613 (N_8613,N_7438,N_5956);
nand U8614 (N_8614,N_4378,N_4260);
nor U8615 (N_8615,N_7573,N_7520);
or U8616 (N_8616,N_6664,N_6854);
and U8617 (N_8617,N_6438,N_4663);
nor U8618 (N_8618,N_5145,N_5657);
nand U8619 (N_8619,N_4080,N_6119);
nor U8620 (N_8620,N_7567,N_4918);
and U8621 (N_8621,N_6701,N_6604);
or U8622 (N_8622,N_6516,N_5377);
and U8623 (N_8623,N_7781,N_4619);
nor U8624 (N_8624,N_5261,N_4636);
nor U8625 (N_8625,N_7490,N_7784);
or U8626 (N_8626,N_5284,N_4191);
nor U8627 (N_8627,N_6598,N_6135);
nor U8628 (N_8628,N_4541,N_5937);
nor U8629 (N_8629,N_5439,N_5975);
nor U8630 (N_8630,N_7884,N_6068);
or U8631 (N_8631,N_7219,N_7998);
nand U8632 (N_8632,N_6886,N_6554);
or U8633 (N_8633,N_7806,N_5554);
nand U8634 (N_8634,N_7469,N_5631);
nand U8635 (N_8635,N_7350,N_5692);
nand U8636 (N_8636,N_4345,N_6498);
or U8637 (N_8637,N_5830,N_6321);
nand U8638 (N_8638,N_5582,N_4790);
nand U8639 (N_8639,N_4760,N_6902);
or U8640 (N_8640,N_7138,N_4288);
xnor U8641 (N_8641,N_6120,N_7682);
nor U8642 (N_8642,N_5569,N_5461);
or U8643 (N_8643,N_7132,N_6532);
nor U8644 (N_8644,N_5242,N_7788);
or U8645 (N_8645,N_6887,N_6593);
and U8646 (N_8646,N_4446,N_6866);
nand U8647 (N_8647,N_6992,N_4727);
nand U8648 (N_8648,N_5886,N_5556);
and U8649 (N_8649,N_7163,N_5808);
and U8650 (N_8650,N_4379,N_5409);
or U8651 (N_8651,N_4113,N_7606);
or U8652 (N_8652,N_7690,N_6571);
nand U8653 (N_8653,N_4968,N_7065);
and U8654 (N_8654,N_7629,N_7546);
or U8655 (N_8655,N_4046,N_7561);
nand U8656 (N_8656,N_6331,N_6788);
nor U8657 (N_8657,N_6294,N_5733);
and U8658 (N_8658,N_7301,N_5574);
or U8659 (N_8659,N_5644,N_5858);
nor U8660 (N_8660,N_5705,N_6863);
nand U8661 (N_8661,N_5112,N_4265);
or U8662 (N_8662,N_4106,N_4998);
and U8663 (N_8663,N_4017,N_5137);
or U8664 (N_8664,N_5291,N_4070);
and U8665 (N_8665,N_6010,N_7139);
nand U8666 (N_8666,N_6430,N_5333);
and U8667 (N_8667,N_6842,N_7381);
nand U8668 (N_8668,N_6138,N_4105);
and U8669 (N_8669,N_6332,N_4336);
and U8670 (N_8670,N_7687,N_6117);
nor U8671 (N_8671,N_7654,N_5008);
nand U8672 (N_8672,N_5463,N_6939);
and U8673 (N_8673,N_5089,N_4353);
or U8674 (N_8674,N_4785,N_5169);
and U8675 (N_8675,N_6609,N_6542);
nor U8676 (N_8676,N_5101,N_7644);
nand U8677 (N_8677,N_6656,N_6051);
nand U8678 (N_8678,N_7291,N_6533);
and U8679 (N_8679,N_5847,N_4512);
or U8680 (N_8680,N_5723,N_4044);
and U8681 (N_8681,N_7838,N_7959);
and U8682 (N_8682,N_7538,N_4603);
nand U8683 (N_8683,N_5194,N_7889);
or U8684 (N_8684,N_6710,N_7608);
nand U8685 (N_8685,N_4637,N_6556);
xnor U8686 (N_8686,N_4284,N_6947);
and U8687 (N_8687,N_6404,N_6089);
and U8688 (N_8688,N_6504,N_7186);
nor U8689 (N_8689,N_5744,N_6272);
or U8690 (N_8690,N_5170,N_4089);
and U8691 (N_8691,N_7605,N_5098);
or U8692 (N_8692,N_4416,N_4144);
and U8693 (N_8693,N_4793,N_7239);
nor U8694 (N_8694,N_4125,N_7521);
nor U8695 (N_8695,N_4809,N_5022);
or U8696 (N_8696,N_7663,N_4128);
nor U8697 (N_8697,N_6032,N_5340);
nor U8698 (N_8698,N_4264,N_7770);
nand U8699 (N_8699,N_5645,N_5075);
nand U8700 (N_8700,N_5969,N_7275);
and U8701 (N_8701,N_4360,N_4137);
and U8702 (N_8702,N_4122,N_6825);
nor U8703 (N_8703,N_7384,N_5130);
nor U8704 (N_8704,N_7515,N_7725);
and U8705 (N_8705,N_4773,N_4917);
or U8706 (N_8706,N_6115,N_7897);
nand U8707 (N_8707,N_5982,N_7704);
nor U8708 (N_8708,N_5111,N_5584);
nand U8709 (N_8709,N_7359,N_7938);
or U8710 (N_8710,N_6499,N_4057);
or U8711 (N_8711,N_5280,N_5609);
and U8712 (N_8712,N_7106,N_6982);
nor U8713 (N_8713,N_7024,N_6188);
or U8714 (N_8714,N_4238,N_7471);
or U8715 (N_8715,N_4974,N_6074);
nor U8716 (N_8716,N_7481,N_4666);
and U8717 (N_8717,N_4408,N_5577);
nor U8718 (N_8718,N_5958,N_4434);
and U8719 (N_8719,N_7262,N_4814);
or U8720 (N_8720,N_4800,N_5097);
or U8721 (N_8721,N_6925,N_5968);
nand U8722 (N_8722,N_7613,N_7578);
nor U8723 (N_8723,N_6713,N_7120);
and U8724 (N_8724,N_7652,N_7053);
and U8725 (N_8725,N_6635,N_7986);
and U8726 (N_8726,N_6765,N_6259);
nand U8727 (N_8727,N_7378,N_5176);
nor U8728 (N_8728,N_6489,N_5268);
nor U8729 (N_8729,N_5985,N_4703);
nor U8730 (N_8730,N_6271,N_4508);
nor U8731 (N_8731,N_4753,N_4720);
or U8732 (N_8732,N_4926,N_7035);
and U8733 (N_8733,N_5967,N_7512);
or U8734 (N_8734,N_6025,N_5315);
or U8735 (N_8735,N_7266,N_5855);
nor U8736 (N_8736,N_7192,N_5680);
or U8737 (N_8737,N_4233,N_4856);
or U8738 (N_8738,N_5942,N_6219);
nand U8739 (N_8739,N_6309,N_6356);
nand U8740 (N_8740,N_6311,N_7722);
nand U8741 (N_8741,N_7800,N_7254);
nand U8742 (N_8742,N_4689,N_5175);
nor U8743 (N_8743,N_6266,N_7294);
nor U8744 (N_8744,N_4517,N_4097);
and U8745 (N_8745,N_4107,N_6587);
and U8746 (N_8746,N_7774,N_5368);
and U8747 (N_8747,N_6183,N_5394);
nand U8748 (N_8748,N_6839,N_6071);
nand U8749 (N_8749,N_5497,N_5696);
nand U8750 (N_8750,N_6191,N_7272);
or U8751 (N_8751,N_4942,N_6217);
or U8752 (N_8752,N_4896,N_4638);
or U8753 (N_8753,N_4081,N_4141);
and U8754 (N_8754,N_5859,N_4445);
nand U8755 (N_8755,N_4832,N_4108);
or U8756 (N_8756,N_4170,N_6557);
and U8757 (N_8757,N_4944,N_5763);
and U8758 (N_8758,N_6759,N_7655);
xor U8759 (N_8759,N_6011,N_4390);
and U8760 (N_8760,N_6442,N_4374);
and U8761 (N_8761,N_7285,N_7757);
nand U8762 (N_8762,N_6676,N_7191);
or U8763 (N_8763,N_4686,N_5072);
nand U8764 (N_8764,N_6125,N_4297);
nand U8765 (N_8765,N_6501,N_7256);
nand U8766 (N_8766,N_6752,N_5308);
or U8767 (N_8767,N_7828,N_7188);
or U8768 (N_8768,N_7738,N_5370);
nor U8769 (N_8769,N_6340,N_6373);
nand U8770 (N_8770,N_4386,N_6342);
and U8771 (N_8771,N_5933,N_4684);
and U8772 (N_8772,N_4973,N_5867);
and U8773 (N_8773,N_4751,N_7988);
or U8774 (N_8774,N_5373,N_5158);
nor U8775 (N_8775,N_7408,N_6441);
or U8776 (N_8776,N_4169,N_4453);
nand U8777 (N_8777,N_7189,N_5557);
nand U8778 (N_8778,N_6352,N_6907);
nor U8779 (N_8779,N_6901,N_5324);
and U8780 (N_8780,N_4842,N_6092);
or U8781 (N_8781,N_5003,N_4366);
and U8782 (N_8782,N_4226,N_6647);
xnor U8783 (N_8783,N_7742,N_5845);
and U8784 (N_8784,N_4913,N_7005);
nand U8785 (N_8785,N_4729,N_7279);
and U8786 (N_8786,N_6076,N_5168);
or U8787 (N_8787,N_7351,N_7295);
nand U8788 (N_8788,N_7990,N_7958);
nor U8789 (N_8789,N_6605,N_4136);
and U8790 (N_8790,N_6779,N_6170);
and U8791 (N_8791,N_4544,N_5997);
or U8792 (N_8792,N_4053,N_4957);
nand U8793 (N_8793,N_4222,N_4433);
nand U8794 (N_8794,N_6750,N_4316);
and U8795 (N_8795,N_4515,N_4908);
and U8796 (N_8796,N_6330,N_6687);
or U8797 (N_8797,N_7115,N_6225);
nand U8798 (N_8798,N_6377,N_7708);
nand U8799 (N_8799,N_5687,N_7043);
xor U8800 (N_8800,N_7719,N_4411);
nor U8801 (N_8801,N_6882,N_5765);
nand U8802 (N_8802,N_6940,N_7817);
nor U8803 (N_8803,N_6447,N_7162);
nor U8804 (N_8804,N_7264,N_4059);
or U8805 (N_8805,N_7688,N_4270);
or U8806 (N_8806,N_4500,N_7826);
or U8807 (N_8807,N_7571,N_6796);
nor U8808 (N_8808,N_4506,N_6070);
nor U8809 (N_8809,N_7809,N_7409);
and U8810 (N_8810,N_5507,N_5263);
and U8811 (N_8811,N_7230,N_4668);
and U8812 (N_8812,N_5140,N_7921);
nand U8813 (N_8813,N_7207,N_5184);
nand U8814 (N_8814,N_7505,N_4310);
or U8815 (N_8815,N_6033,N_4899);
nand U8816 (N_8816,N_6396,N_6999);
or U8817 (N_8817,N_5397,N_5797);
xor U8818 (N_8818,N_6753,N_5927);
nor U8819 (N_8819,N_5791,N_7320);
and U8820 (N_8820,N_6162,N_7863);
and U8821 (N_8821,N_5862,N_6147);
nand U8822 (N_8822,N_5096,N_5259);
and U8823 (N_8823,N_4623,N_7925);
nand U8824 (N_8824,N_7425,N_6374);
nand U8825 (N_8825,N_6122,N_7807);
or U8826 (N_8826,N_6884,N_4404);
and U8827 (N_8827,N_4965,N_5662);
and U8828 (N_8828,N_5543,N_6561);
nor U8829 (N_8829,N_4665,N_6124);
or U8830 (N_8830,N_4651,N_7015);
and U8831 (N_8831,N_5742,N_5658);
nor U8832 (N_8832,N_6464,N_6355);
nor U8833 (N_8833,N_4652,N_5992);
nor U8834 (N_8834,N_7498,N_6381);
nand U8835 (N_8835,N_5573,N_4280);
nor U8836 (N_8836,N_5921,N_5851);
or U8837 (N_8837,N_7487,N_6429);
nand U8838 (N_8838,N_4622,N_5703);
nand U8839 (N_8839,N_4461,N_5514);
nor U8840 (N_8840,N_6798,N_5088);
nand U8841 (N_8841,N_6905,N_5142);
xor U8842 (N_8842,N_5594,N_6149);
and U8843 (N_8843,N_5908,N_6255);
or U8844 (N_8844,N_5342,N_7181);
nor U8845 (N_8845,N_4699,N_5866);
or U8846 (N_8846,N_5592,N_6243);
and U8847 (N_8847,N_6171,N_4197);
or U8848 (N_8848,N_6916,N_7748);
nor U8849 (N_8849,N_5051,N_5078);
or U8850 (N_8850,N_6401,N_4860);
nor U8851 (N_8851,N_6455,N_5509);
and U8852 (N_8852,N_4997,N_5911);
nand U8853 (N_8853,N_5699,N_5103);
and U8854 (N_8854,N_7860,N_5498);
nor U8855 (N_8855,N_7666,N_4811);
or U8856 (N_8856,N_5430,N_6383);
and U8857 (N_8857,N_6617,N_5693);
nand U8858 (N_8858,N_7754,N_6969);
and U8859 (N_8859,N_4873,N_5433);
nand U8860 (N_8860,N_4254,N_5729);
or U8861 (N_8861,N_5238,N_4388);
nor U8862 (N_8862,N_5843,N_6177);
or U8863 (N_8863,N_4457,N_5149);
nor U8864 (N_8864,N_7550,N_4160);
nand U8865 (N_8865,N_5163,N_6717);
nand U8866 (N_8866,N_7993,N_5006);
nand U8867 (N_8867,N_7676,N_4300);
and U8868 (N_8868,N_5249,N_5265);
nand U8869 (N_8869,N_7560,N_5661);
and U8870 (N_8870,N_5178,N_5005);
nand U8871 (N_8871,N_6833,N_5794);
or U8872 (N_8872,N_5320,N_6955);
nor U8873 (N_8873,N_6589,N_7302);
nor U8874 (N_8874,N_4629,N_4821);
nor U8875 (N_8875,N_5350,N_7896);
nand U8876 (N_8876,N_4859,N_5057);
and U8877 (N_8877,N_4279,N_7479);
and U8878 (N_8878,N_7552,N_5769);
or U8879 (N_8879,N_7670,N_4647);
nor U8880 (N_8880,N_5260,N_6835);
nor U8881 (N_8881,N_5620,N_6977);
and U8882 (N_8882,N_6372,N_7540);
nand U8883 (N_8883,N_6927,N_5630);
nand U8884 (N_8884,N_7280,N_7096);
nor U8885 (N_8885,N_7881,N_4844);
or U8886 (N_8886,N_4234,N_5750);
or U8887 (N_8887,N_6467,N_5361);
nand U8888 (N_8888,N_6205,N_7141);
nand U8889 (N_8889,N_7317,N_4774);
or U8890 (N_8890,N_7128,N_4354);
nor U8891 (N_8891,N_4565,N_7991);
or U8892 (N_8892,N_5737,N_7023);
nand U8893 (N_8893,N_6078,N_6803);
and U8894 (N_8894,N_5252,N_7242);
and U8895 (N_8895,N_5806,N_5401);
or U8896 (N_8896,N_4298,N_5918);
or U8897 (N_8897,N_4882,N_7864);
or U8898 (N_8898,N_5792,N_5182);
nor U8899 (N_8899,N_5154,N_5235);
nand U8900 (N_8900,N_7873,N_4907);
nor U8901 (N_8901,N_7541,N_5552);
or U8902 (N_8902,N_4738,N_4600);
or U8903 (N_8903,N_4375,N_6003);
and U8904 (N_8904,N_6256,N_6009);
or U8905 (N_8905,N_7270,N_6346);
or U8906 (N_8906,N_7464,N_4945);
nor U8907 (N_8907,N_5109,N_4846);
nand U8908 (N_8908,N_6506,N_5834);
nand U8909 (N_8909,N_6881,N_6929);
and U8910 (N_8910,N_4455,N_4561);
nor U8911 (N_8911,N_5607,N_4725);
or U8912 (N_8912,N_7519,N_5432);
or U8913 (N_8913,N_6942,N_4205);
and U8914 (N_8914,N_6784,N_6290);
nand U8915 (N_8915,N_7803,N_7982);
nor U8916 (N_8916,N_6970,N_5899);
and U8917 (N_8917,N_7009,N_6913);
and U8918 (N_8918,N_5469,N_5850);
and U8919 (N_8919,N_7577,N_7465);
nor U8920 (N_8920,N_6622,N_5275);
and U8921 (N_8921,N_7756,N_5187);
or U8922 (N_8922,N_6702,N_5788);
nand U8923 (N_8923,N_6980,N_5203);
nand U8924 (N_8924,N_4127,N_5730);
nor U8925 (N_8925,N_4287,N_7653);
and U8926 (N_8926,N_7865,N_4465);
nor U8927 (N_8927,N_4362,N_5462);
nand U8928 (N_8928,N_5567,N_6665);
nor U8929 (N_8929,N_6079,N_7218);
nor U8930 (N_8930,N_5153,N_4986);
nand U8931 (N_8931,N_6477,N_6320);
nand U8932 (N_8932,N_4586,N_5819);
nand U8933 (N_8933,N_6981,N_6226);
nor U8934 (N_8934,N_6144,N_5150);
nand U8935 (N_8935,N_4872,N_4555);
nor U8936 (N_8936,N_5276,N_4839);
and U8937 (N_8937,N_7395,N_7660);
or U8938 (N_8938,N_4797,N_5688);
or U8939 (N_8939,N_5290,N_5876);
and U8940 (N_8940,N_5076,N_7002);
nor U8941 (N_8941,N_5779,N_6014);
or U8942 (N_8942,N_4685,N_4024);
nand U8943 (N_8943,N_6517,N_5783);
nor U8944 (N_8944,N_7945,N_7127);
nor U8945 (N_8945,N_7526,N_7973);
nor U8946 (N_8946,N_5288,N_7396);
nand U8947 (N_8947,N_4104,N_7293);
or U8948 (N_8948,N_6629,N_4653);
nor U8949 (N_8949,N_5741,N_4410);
and U8950 (N_8950,N_7813,N_7446);
nor U8951 (N_8951,N_5586,N_6814);
nand U8952 (N_8952,N_7697,N_4563);
and U8953 (N_8953,N_7805,N_7042);
nor U8954 (N_8954,N_4818,N_7589);
or U8955 (N_8955,N_7810,N_7662);
or U8956 (N_8956,N_7558,N_5612);
nand U8957 (N_8957,N_5988,N_6040);
nand U8958 (N_8958,N_4916,N_6773);
nand U8959 (N_8959,N_5932,N_7309);
and U8960 (N_8960,N_6848,N_7964);
and U8961 (N_8961,N_6313,N_5674);
or U8962 (N_8962,N_4272,N_6199);
nand U8963 (N_8963,N_6476,N_5871);
nand U8964 (N_8964,N_5904,N_6422);
or U8965 (N_8965,N_5650,N_4614);
and U8966 (N_8966,N_4211,N_5047);
and U8967 (N_8967,N_4380,N_7645);
nor U8968 (N_8968,N_5256,N_6065);
and U8969 (N_8969,N_4946,N_4898);
nor U8970 (N_8970,N_7450,N_7491);
and U8971 (N_8971,N_6640,N_6948);
or U8972 (N_8972,N_6552,N_7868);
or U8973 (N_8973,N_7893,N_6712);
or U8974 (N_8974,N_5385,N_5357);
nand U8975 (N_8975,N_4677,N_7528);
and U8976 (N_8976,N_7021,N_5071);
or U8977 (N_8977,N_6708,N_5354);
nor U8978 (N_8978,N_6159,N_6118);
nand U8979 (N_8979,N_7729,N_5466);
nor U8980 (N_8980,N_6659,N_5513);
nand U8981 (N_8981,N_4676,N_4351);
nand U8982 (N_8982,N_7522,N_6022);
nor U8983 (N_8983,N_5415,N_6165);
nand U8984 (N_8984,N_7492,N_5039);
nor U8985 (N_8985,N_6432,N_5173);
nor U8986 (N_8986,N_6001,N_5585);
nor U8987 (N_8987,N_6870,N_7494);
or U8988 (N_8988,N_5488,N_6431);
or U8989 (N_8989,N_7283,N_7657);
nor U8990 (N_8990,N_5826,N_4018);
nand U8991 (N_8991,N_5436,N_4750);
nand U8992 (N_8992,N_5234,N_4507);
or U8993 (N_8993,N_7715,N_5327);
nand U8994 (N_8994,N_7843,N_4543);
nor U8995 (N_8995,N_5545,N_5161);
nand U8996 (N_8996,N_7486,N_6573);
and U8997 (N_8997,N_6500,N_4769);
and U8998 (N_8998,N_7673,N_5801);
or U8999 (N_8999,N_7363,N_6510);
nor U9000 (N_9000,N_7085,N_6019);
and U9001 (N_9001,N_7760,N_6602);
nor U9002 (N_9002,N_6692,N_5470);
and U9003 (N_9003,N_6946,N_5938);
nand U9004 (N_9004,N_4994,N_5930);
nand U9005 (N_9005,N_6922,N_7984);
and U9006 (N_9006,N_7037,N_4171);
and U9007 (N_9007,N_6968,N_4196);
nor U9008 (N_9008,N_7168,N_4119);
and U9009 (N_9009,N_6613,N_7452);
nand U9010 (N_9010,N_5694,N_6038);
nand U9011 (N_9011,N_5838,N_4129);
and U9012 (N_9012,N_4069,N_5568);
or U9013 (N_9013,N_5815,N_6257);
or U9014 (N_9014,N_7312,N_5063);
nor U9015 (N_9015,N_4256,N_6897);
or U9016 (N_9016,N_4067,N_4307);
and U9017 (N_9017,N_5362,N_7823);
nand U9018 (N_9018,N_5984,N_4640);
nand U9019 (N_9019,N_4493,N_6345);
and U9020 (N_9020,N_7154,N_5888);
nand U9021 (N_9021,N_4350,N_7518);
nand U9022 (N_9022,N_6584,N_5355);
or U9023 (N_9023,N_4513,N_7131);
nor U9024 (N_9024,N_6348,N_4902);
xor U9025 (N_9025,N_7246,N_4642);
nand U9026 (N_9026,N_6215,N_5059);
nand U9027 (N_9027,N_7941,N_5338);
nand U9028 (N_9028,N_7681,N_5046);
nand U9029 (N_9029,N_6790,N_4995);
and U9030 (N_9030,N_7563,N_6719);
nand U9031 (N_9031,N_4527,N_4855);
nor U9032 (N_9032,N_5640,N_5629);
or U9033 (N_9033,N_4407,N_5857);
and U9034 (N_9034,N_7171,N_5074);
nor U9035 (N_9035,N_6641,N_7878);
and U9036 (N_9036,N_4219,N_7278);
and U9037 (N_9037,N_4240,N_6273);
nor U9038 (N_9038,N_5883,N_6247);
and U9039 (N_9039,N_5523,N_6926);
and U9040 (N_9040,N_4611,N_5961);
nand U9041 (N_9041,N_6972,N_5042);
and U9042 (N_9042,N_4005,N_4040);
or U9043 (N_9043,N_4876,N_7373);
xnor U9044 (N_9044,N_5965,N_7488);
nand U9045 (N_9045,N_4207,N_6857);
or U9046 (N_9046,N_6952,N_5431);
nand U9047 (N_9047,N_4178,N_6397);
or U9048 (N_9048,N_4734,N_5709);
or U9049 (N_9049,N_5421,N_5960);
or U9050 (N_9050,N_4875,N_4796);
and U9051 (N_9051,N_7840,N_4432);
or U9052 (N_9052,N_5745,N_5832);
nor U9053 (N_9053,N_5192,N_7214);
nand U9054 (N_9054,N_4644,N_6575);
nor U9055 (N_9055,N_4804,N_4789);
and U9056 (N_9056,N_5822,N_7442);
and U9057 (N_9057,N_4478,N_5579);
or U9058 (N_9058,N_6096,N_4747);
and U9059 (N_9059,N_4829,N_5307);
nor U9060 (N_9060,N_5205,N_6298);
nor U9061 (N_9061,N_4158,N_7771);
nand U9062 (N_9062,N_4313,N_6599);
and U9063 (N_9063,N_7906,N_6891);
or U9064 (N_9064,N_4547,N_6861);
and U9065 (N_9065,N_5278,N_4062);
nand U9066 (N_9066,N_6161,N_6813);
or U9067 (N_9067,N_7614,N_7041);
and U9068 (N_9068,N_5289,N_6497);
nor U9069 (N_9069,N_4674,N_6911);
or U9070 (N_9070,N_7583,N_6123);
and U9071 (N_9071,N_4176,N_4768);
or U9072 (N_9072,N_5248,N_5198);
and U9073 (N_9073,N_7846,N_6270);
or U9074 (N_9074,N_6994,N_4087);
or U9075 (N_9075,N_4139,N_4155);
and U9076 (N_9076,N_5273,N_6350);
and U9077 (N_9077,N_5314,N_4891);
or U9078 (N_9078,N_7581,N_4540);
or U9079 (N_9079,N_6153,N_5127);
nand U9080 (N_9080,N_6234,N_4988);
nor U9081 (N_9081,N_6291,N_4395);
or U9082 (N_9082,N_6224,N_7136);
nand U9083 (N_9083,N_4980,N_6923);
and U9084 (N_9084,N_5803,N_7818);
nor U9085 (N_9085,N_7439,N_7125);
nor U9086 (N_9086,N_5949,N_4435);
or U9087 (N_9087,N_5068,N_4910);
nor U9088 (N_9088,N_6591,N_4138);
or U9089 (N_9089,N_6412,N_7885);
nor U9090 (N_9090,N_5152,N_6778);
or U9091 (N_9091,N_5084,N_7844);
or U9092 (N_9092,N_6658,N_6699);
nand U9093 (N_9093,N_6837,N_6277);
xor U9094 (N_9094,N_7413,N_7038);
nand U9095 (N_9095,N_4687,N_4805);
or U9096 (N_9096,N_4235,N_5243);
nor U9097 (N_9097,N_7049,N_7227);
and U9098 (N_9098,N_6828,N_5332);
and U9099 (N_9099,N_6675,N_6387);
xor U9100 (N_9100,N_5065,N_7626);
nor U9101 (N_9101,N_4743,N_6439);
and U9102 (N_9102,N_7055,N_7866);
nand U9103 (N_9103,N_7484,N_6035);
and U9104 (N_9104,N_7451,N_7327);
nor U9105 (N_9105,N_7795,N_6249);
or U9106 (N_9106,N_5303,N_6964);
nor U9107 (N_9107,N_6634,N_6628);
nand U9108 (N_9108,N_5914,N_7418);
and U9109 (N_9109,N_5591,N_7235);
and U9110 (N_9110,N_7776,N_6819);
or U9111 (N_9111,N_5146,N_5752);
or U9112 (N_9112,N_5789,N_6936);
nand U9113 (N_9113,N_4870,N_4450);
and U9114 (N_9114,N_6048,N_6919);
nand U9115 (N_9115,N_4359,N_4706);
nand U9116 (N_9116,N_5619,N_7461);
nor U9117 (N_9117,N_5427,N_7847);
and U9118 (N_9118,N_4417,N_7332);
nor U9119 (N_9119,N_7091,N_7473);
or U9120 (N_9120,N_4099,N_4709);
and U9121 (N_9121,N_5748,N_6720);
and U9122 (N_9122,N_6845,N_4522);
nor U9123 (N_9123,N_4937,N_5917);
and U9124 (N_9124,N_7839,N_4654);
nor U9125 (N_9125,N_6142,N_4290);
nor U9126 (N_9126,N_4082,N_7016);
and U9127 (N_9127,N_4661,N_7997);
and U9128 (N_9128,N_4277,N_6672);
nand U9129 (N_9129,N_5220,N_6000);
or U9130 (N_9130,N_5500,N_5077);
nand U9131 (N_9131,N_4094,N_7164);
nor U9132 (N_9132,N_4383,N_4892);
and U9133 (N_9133,N_4237,N_5583);
nand U9134 (N_9134,N_5107,N_7110);
or U9135 (N_9135,N_6486,N_4869);
and U9136 (N_9136,N_5642,N_4201);
and U9137 (N_9137,N_7600,N_5200);
nand U9138 (N_9138,N_4166,N_7707);
xnor U9139 (N_9139,N_4203,N_6053);
or U9140 (N_9140,N_7816,N_6998);
nor U9141 (N_9141,N_7954,N_6748);
and U9142 (N_9142,N_5524,N_7234);
nand U9143 (N_9143,N_5747,N_7263);
or U9144 (N_9144,N_7203,N_4548);
nand U9145 (N_9145,N_7400,N_5863);
or U9146 (N_9146,N_5156,N_6871);
or U9147 (N_9147,N_5995,N_7949);
or U9148 (N_9148,N_5799,N_5083);
nand U9149 (N_9149,N_7100,N_4578);
nand U9150 (N_9150,N_6166,N_6490);
and U9151 (N_9151,N_4365,N_7060);
or U9152 (N_9152,N_6774,N_4093);
nor U9153 (N_9153,N_5950,N_4819);
nor U9154 (N_9154,N_7743,N_7311);
or U9155 (N_9155,N_4822,N_7923);
nand U9156 (N_9156,N_5493,N_6389);
nand U9157 (N_9157,N_7316,N_5749);
and U9158 (N_9158,N_6777,N_5162);
or U9159 (N_9159,N_7525,N_4133);
and U9160 (N_9160,N_7393,N_5300);
nor U9161 (N_9161,N_6522,N_6007);
nand U9162 (N_9162,N_5418,N_7319);
or U9163 (N_9163,N_6890,N_5311);
nand U9164 (N_9164,N_7735,N_6006);
and U9165 (N_9165,N_6080,N_6794);
nand U9166 (N_9166,N_5559,N_4801);
or U9167 (N_9167,N_4077,N_4645);
nand U9168 (N_9168,N_6233,N_6921);
nand U9169 (N_9169,N_7642,N_5503);
nand U9170 (N_9170,N_4901,N_4862);
nor U9171 (N_9171,N_7730,N_7592);
nor U9172 (N_9172,N_7366,N_5216);
and U9173 (N_9173,N_6518,N_4867);
and U9174 (N_9174,N_7618,N_7930);
or U9175 (N_9175,N_4487,N_4581);
nand U9176 (N_9176,N_7097,N_6636);
or U9177 (N_9177,N_6771,N_6210);
nor U9178 (N_9178,N_6250,N_7252);
or U9179 (N_9179,N_6781,N_6454);
and U9180 (N_9180,N_5056,N_6768);
or U9181 (N_9181,N_4680,N_7365);
nor U9182 (N_9182,N_5562,N_5770);
nand U9183 (N_9183,N_4721,N_6148);
nor U9184 (N_9184,N_4749,N_4585);
or U9185 (N_9185,N_5478,N_6420);
and U9186 (N_9186,N_5405,N_6364);
nand U9187 (N_9187,N_6052,N_7497);
or U9188 (N_9188,N_7740,N_5944);
or U9189 (N_9189,N_5701,N_5027);
nand U9190 (N_9190,N_4485,N_6943);
and U9191 (N_9191,N_5445,N_4730);
nand U9192 (N_9192,N_7591,N_5636);
nand U9193 (N_9193,N_7380,N_7006);
or U9194 (N_9194,N_5467,N_5134);
nand U9195 (N_9195,N_4273,N_4221);
or U9196 (N_9196,N_6791,N_7634);
nand U9197 (N_9197,N_7269,N_6594);
nand U9198 (N_9198,N_7349,N_6595);
or U9199 (N_9199,N_5437,N_7999);
or U9200 (N_9200,N_6421,N_6326);
or U9201 (N_9201,N_4056,N_6783);
nand U9202 (N_9202,N_5094,N_4932);
and U9203 (N_9203,N_7387,N_6239);
nor U9204 (N_9204,N_6474,N_6262);
or U9205 (N_9205,N_6693,N_4791);
or U9206 (N_9206,N_6303,N_7509);
nand U9207 (N_9207,N_7598,N_6394);
or U9208 (N_9208,N_6909,N_4770);
and U9209 (N_9209,N_4953,N_4262);
nand U9210 (N_9210,N_4958,N_7679);
or U9211 (N_9211,N_4971,N_4335);
nor U9212 (N_9212,N_4900,N_5532);
or U9213 (N_9213,N_5283,N_4466);
nor U9214 (N_9214,N_6293,N_5776);
or U9215 (N_9215,N_7119,N_4808);
nor U9216 (N_9216,N_7842,N_5240);
nor U9217 (N_9217,N_4574,N_6512);
nor U9218 (N_9218,N_4671,N_7229);
or U9219 (N_9219,N_5322,N_5648);
and U9220 (N_9220,N_6904,N_7929);
or U9221 (N_9221,N_4696,N_7962);
and U9222 (N_9222,N_4503,N_7206);
and U9223 (N_9223,N_6408,N_6678);
nor U9224 (N_9224,N_6444,N_6924);
xnor U9225 (N_9225,N_7902,N_4635);
nor U9226 (N_9226,N_5570,N_6069);
and U9227 (N_9227,N_6694,N_5092);
or U9228 (N_9228,N_7047,N_7580);
and U9229 (N_9229,N_4618,N_6730);
or U9230 (N_9230,N_5364,N_6024);
nand U9231 (N_9231,N_6228,N_5286);
nand U9232 (N_9232,N_7535,N_7948);
or U9233 (N_9233,N_4772,N_5816);
and U9234 (N_9234,N_4029,N_6894);
and U9235 (N_9235,N_4919,N_6786);
or U9236 (N_9236,N_6176,N_7200);
nand U9237 (N_9237,N_7346,N_4086);
or U9238 (N_9238,N_7175,N_4022);
or U9239 (N_9239,N_5726,N_7111);
and U9240 (N_9240,N_4571,N_5751);
nand U9241 (N_9241,N_4229,N_7939);
and U9242 (N_9242,N_6418,N_4224);
or U9243 (N_9243,N_5912,N_5352);
nor U9244 (N_9244,N_4938,N_5007);
nor U9245 (N_9245,N_4646,N_4425);
nand U9246 (N_9246,N_4143,N_6386);
nor U9247 (N_9247,N_4987,N_7196);
and U9248 (N_9248,N_7946,N_7101);
and U9249 (N_9249,N_6690,N_6736);
nor U9250 (N_9250,N_7095,N_6017);
and U9251 (N_9251,N_6391,N_7779);
nand U9252 (N_9252,N_7819,N_7731);
and U9253 (N_9253,N_4895,N_7241);
and U9254 (N_9254,N_5538,N_5923);
and U9255 (N_9255,N_6797,N_5903);
nor U9256 (N_9256,N_6155,N_6850);
nor U9257 (N_9257,N_7615,N_6795);
nand U9258 (N_9258,N_6244,N_7108);
nor U9259 (N_9259,N_6023,N_7453);
nand U9260 (N_9260,N_6209,N_4372);
and U9261 (N_9261,N_4301,N_5515);
and U9262 (N_9262,N_7458,N_6204);
xor U9263 (N_9263,N_7184,N_6728);
nand U9264 (N_9264,N_4810,N_4959);
or U9265 (N_9265,N_6684,N_4714);
nor U9266 (N_9266,N_5271,N_5129);
nor U9267 (N_9267,N_6265,N_7837);
or U9268 (N_9268,N_5780,N_7872);
or U9269 (N_9269,N_4880,N_5202);
or U9270 (N_9270,N_7749,N_5520);
nor U9271 (N_9271,N_5698,N_7680);
nand U9272 (N_9272,N_5087,N_5536);
or U9273 (N_9273,N_5681,N_7965);
and U9274 (N_9274,N_6167,N_4787);
nand U9275 (N_9275,N_5325,N_6187);
nor U9276 (N_9276,N_7238,N_7299);
nand U9277 (N_9277,N_6956,N_5807);
nand U9278 (N_9278,N_5121,N_4960);
nor U9279 (N_9279,N_6695,N_5756);
nand U9280 (N_9280,N_5951,N_4115);
nand U9281 (N_9281,N_7148,N_5345);
nor U9282 (N_9282,N_4120,N_5708);
or U9283 (N_9283,N_4632,N_6043);
nand U9284 (N_9284,N_6212,N_5849);
or U9285 (N_9285,N_7480,N_7559);
nor U9286 (N_9286,N_6618,N_5823);
or U9287 (N_9287,N_4302,N_7124);
nor U9288 (N_9288,N_5239,N_6085);
and U9289 (N_9289,N_4559,N_5727);
and U9290 (N_9290,N_5204,N_6425);
or U9291 (N_9291,N_4669,N_5215);
and U9292 (N_9292,N_4792,N_7985);
or U9293 (N_9293,N_5576,N_4612);
and U9294 (N_9294,N_5660,N_6246);
nand U9295 (N_9295,N_6360,N_5614);
nand U9296 (N_9296,N_6336,N_7226);
or U9297 (N_9297,N_4079,N_4510);
nand U9298 (N_9298,N_6519,N_7274);
or U9299 (N_9299,N_7059,N_7149);
nor U9300 (N_9300,N_7752,N_6853);
or U9301 (N_9301,N_7495,N_6164);
nand U9302 (N_9302,N_6812,N_7882);
and U9303 (N_9303,N_5020,N_6834);
or U9304 (N_9304,N_4498,N_7638);
and U9305 (N_9305,N_6931,N_5045);
or U9306 (N_9306,N_5468,N_4114);
and U9307 (N_9307,N_6691,N_6058);
and U9308 (N_9308,N_7454,N_6883);
nor U9309 (N_9309,N_4756,N_4949);
or U9310 (N_9310,N_4083,N_7545);
nand U9311 (N_9311,N_4978,N_7391);
xor U9312 (N_9312,N_5214,N_7534);
or U9313 (N_9313,N_6175,N_7820);
and U9314 (N_9314,N_6308,N_7170);
nor U9315 (N_9315,N_5298,N_4269);
and U9316 (N_9316,N_5934,N_6761);
nor U9317 (N_9317,N_4824,N_6005);
nand U9318 (N_9318,N_7223,N_4014);
and U9319 (N_9319,N_5382,N_6312);
or U9320 (N_9320,N_5605,N_4951);
or U9321 (N_9321,N_4939,N_6746);
nand U9322 (N_9322,N_6560,N_7934);
nand U9323 (N_9323,N_6127,N_4717);
and U9324 (N_9324,N_7974,N_7287);
or U9325 (N_9325,N_6976,N_6182);
or U9326 (N_9326,N_7554,N_5309);
nand U9327 (N_9327,N_4185,N_4327);
nand U9328 (N_9328,N_6957,N_7667);
nor U9329 (N_9329,N_7924,N_6329);
nand U9330 (N_9330,N_4553,N_4431);
nand U9331 (N_9331,N_5669,N_7780);
or U9332 (N_9332,N_4935,N_4579);
nor U9333 (N_9333,N_7328,N_7709);
or U9334 (N_9334,N_6368,N_6832);
and U9335 (N_9335,N_7960,N_6221);
or U9336 (N_9336,N_6435,N_4452);
or U9337 (N_9337,N_4610,N_7228);
nand U9338 (N_9338,N_6475,N_7920);
or U9339 (N_9339,N_4363,N_4111);
nand U9340 (N_9340,N_6145,N_7448);
or U9341 (N_9341,N_5396,N_7339);
or U9342 (N_9342,N_4631,N_5269);
or U9343 (N_9343,N_5486,N_5304);
or U9344 (N_9344,N_5459,N_6054);
and U9345 (N_9345,N_4490,N_4006);
and U9346 (N_9346,N_5817,N_6103);
and U9347 (N_9347,N_4542,N_4074);
and U9348 (N_9348,N_4526,N_5760);
nand U9349 (N_9349,N_6097,N_6393);
or U9350 (N_9350,N_7887,N_6361);
nand U9351 (N_9351,N_4368,N_5105);
or U9352 (N_9352,N_4026,N_4582);
or U9353 (N_9353,N_6663,N_6984);
nand U9354 (N_9354,N_4168,N_6436);
nor U9355 (N_9355,N_6179,N_6762);
and U9356 (N_9356,N_6469,N_4724);
nor U9357 (N_9357,N_4595,N_5827);
nand U9358 (N_9358,N_4925,N_5406);
nand U9359 (N_9359,N_4402,N_5277);
nand U9360 (N_9360,N_5947,N_6037);
nand U9361 (N_9361,N_5771,N_4678);
nor U9362 (N_9362,N_5964,N_6113);
or U9363 (N_9363,N_4757,N_7298);
or U9364 (N_9364,N_6536,N_6174);
nor U9365 (N_9365,N_5247,N_7493);
nand U9366 (N_9366,N_5861,N_6990);
nand U9367 (N_9367,N_4673,N_4977);
and U9368 (N_9368,N_6817,N_6338);
and U9369 (N_9369,N_5119,N_6495);
nor U9370 (N_9370,N_4189,N_5434);
or U9371 (N_9371,N_7969,N_5293);
and U9372 (N_9372,N_7665,N_5179);
and U9373 (N_9373,N_4394,N_5646);
and U9374 (N_9374,N_5870,N_4560);
or U9375 (N_9375,N_6083,N_4242);
or U9376 (N_9376,N_7437,N_7300);
and U9377 (N_9377,N_4897,N_7936);
and U9378 (N_9378,N_4275,N_6974);
nor U9379 (N_9379,N_6729,N_5885);
and U9380 (N_9380,N_4475,N_7183);
or U9381 (N_9381,N_5030,N_5458);
or U9382 (N_9382,N_6787,N_7000);
and U9383 (N_9383,N_5506,N_6251);
and U9384 (N_9384,N_6395,N_7443);
and U9385 (N_9385,N_7603,N_4016);
or U9386 (N_9386,N_4246,N_4419);
and U9387 (N_9387,N_4494,N_4315);
or U9388 (N_9388,N_6586,N_6502);
or U9389 (N_9389,N_7564,N_6132);
and U9390 (N_9390,N_7684,N_6577);
or U9391 (N_9391,N_6299,N_7062);
and U9392 (N_9392,N_5371,N_6046);
nor U9393 (N_9393,N_5236,N_4532);
nand U9394 (N_9394,N_6232,N_6912);
and U9395 (N_9395,N_6403,N_6918);
nor U9396 (N_9396,N_7195,N_5936);
nor U9397 (N_9397,N_4030,N_7353);
and U9398 (N_9398,N_7956,N_6344);
or U9399 (N_9399,N_5128,N_6451);
nand U9400 (N_9400,N_6983,N_5376);
nor U9401 (N_9401,N_5025,N_6047);
and U9402 (N_9402,N_7620,N_5842);
nand U9403 (N_9403,N_4991,N_5575);
nand U9404 (N_9404,N_6868,N_7917);
nand U9405 (N_9405,N_4802,N_5766);
nor U9406 (N_9406,N_7113,N_7440);
nor U9407 (N_9407,N_6660,N_6619);
and U9408 (N_9408,N_4346,N_4367);
nor U9409 (N_9409,N_4723,N_4463);
or U9410 (N_9410,N_4698,N_7355);
nor U9411 (N_9411,N_7261,N_7117);
and U9412 (N_9412,N_4763,N_4697);
and U9413 (N_9413,N_5601,N_7260);
nand U9414 (N_9414,N_6775,N_6057);
nor U9415 (N_9415,N_4713,N_4248);
and U9416 (N_9416,N_6405,N_7045);
or U9417 (N_9417,N_7423,N_6681);
or U9418 (N_9418,N_7915,N_5704);
nand U9419 (N_9419,N_6279,N_6102);
nand U9420 (N_9420,N_7435,N_6328);
or U9421 (N_9421,N_6493,N_6358);
nor U9422 (N_9422,N_7022,N_5533);
nand U9423 (N_9423,N_5040,N_4737);
nor U9424 (N_9424,N_7212,N_7107);
nand U9425 (N_9425,N_6201,N_4464);
and U9426 (N_9426,N_4409,N_5351);
or U9427 (N_9427,N_7182,N_5359);
and U9428 (N_9428,N_5635,N_6570);
nand U9429 (N_9429,N_7694,N_5738);
xor U9430 (N_9430,N_6390,N_5755);
and U9431 (N_9431,N_5820,N_7678);
or U9432 (N_9432,N_5697,N_5897);
nor U9433 (N_9433,N_6202,N_7625);
xor U9434 (N_9434,N_7099,N_7871);
nor U9435 (N_9435,N_7421,N_5610);
nand U9436 (N_9436,N_7677,N_4314);
or U9437 (N_9437,N_7017,N_5824);
nand U9438 (N_9438,N_7292,N_4516);
nor U9439 (N_9439,N_6642,N_7714);
nor U9440 (N_9440,N_4608,N_6324);
nor U9441 (N_9441,N_7912,N_7802);
nor U9442 (N_9442,N_6627,N_4023);
nor U9443 (N_9443,N_4438,N_5906);
and U9444 (N_9444,N_6801,N_4295);
xor U9445 (N_9445,N_5301,N_4624);
and U9446 (N_9446,N_4258,N_4981);
nand U9447 (N_9447,N_4096,N_5318);
and U9448 (N_9448,N_7329,N_7243);
nand U9449 (N_9449,N_4762,N_7517);
nand U9450 (N_9450,N_4480,N_4382);
nand U9451 (N_9451,N_6150,N_4338);
and U9452 (N_9452,N_6304,N_5716);
and U9453 (N_9453,N_5837,N_5053);
or U9454 (N_9454,N_6114,N_7718);
and U9455 (N_9455,N_5714,N_5496);
or U9456 (N_9456,N_7672,N_6611);
and U9457 (N_9457,N_7639,N_4149);
nor U9458 (N_9458,N_5285,N_5442);
or U9459 (N_9459,N_6254,N_6836);
or U9460 (N_9460,N_4282,N_7647);
nor U9461 (N_9461,N_5597,N_4131);
or U9462 (N_9462,N_5197,N_7036);
nor U9463 (N_9463,N_5435,N_7019);
or U9464 (N_9464,N_5664,N_7057);
nand U9465 (N_9465,N_5224,N_6130);
nor U9466 (N_9466,N_4741,N_6689);
and U9467 (N_9467,N_7911,N_7376);
or U9468 (N_9468,N_5720,N_4004);
and U9469 (N_9469,N_6222,N_5811);
or U9470 (N_9470,N_4098,N_4530);
nor U9471 (N_9471,N_4156,N_5013);
or U9472 (N_9472,N_4650,N_6514);
nand U9473 (N_9473,N_7161,N_5540);
or U9474 (N_9474,N_7588,N_4068);
or U9475 (N_9475,N_5560,N_5639);
or U9476 (N_9476,N_5246,N_5924);
and U9477 (N_9477,N_5521,N_7527);
nand U9478 (N_9478,N_5360,N_4286);
and U9479 (N_9479,N_4524,N_7734);
nor U9480 (N_9480,N_7258,N_5487);
or U9481 (N_9481,N_4710,N_4019);
and U9482 (N_9482,N_6823,N_4798);
nor U9483 (N_9483,N_6564,N_5321);
nand U9484 (N_9484,N_5978,N_7504);
nor U9485 (N_9485,N_7354,N_7217);
xor U9486 (N_9486,N_7383,N_7726);
nand U9487 (N_9487,N_6196,N_7763);
or U9488 (N_9488,N_6987,N_5668);
and U9489 (N_9489,N_6151,N_6453);
nor U9490 (N_9490,N_4007,N_7942);
nand U9491 (N_9491,N_5633,N_7031);
and U9492 (N_9492,N_5667,N_7786);
nand U9493 (N_9493,N_4497,N_6236);
and U9494 (N_9494,N_6958,N_6715);
or U9495 (N_9495,N_7140,N_5110);
nor U9496 (N_9496,N_4209,N_6297);
nand U9497 (N_9497,N_6357,N_4922);
nand U9498 (N_9498,N_7030,N_6173);
and U9499 (N_9499,N_4983,N_6945);
or U9500 (N_9500,N_4999,N_6780);
or U9501 (N_9501,N_7403,N_7574);
nand U9502 (N_9502,N_6230,N_6574);
nor U9503 (N_9503,N_4292,N_6278);
or U9504 (N_9504,N_7845,N_4799);
or U9505 (N_9505,N_7146,N_4735);
nand U9506 (N_9506,N_6214,N_7336);
and U9507 (N_9507,N_6508,N_6030);
and U9508 (N_9508,N_6529,N_7981);
nand U9509 (N_9509,N_5123,N_7547);
nor U9510 (N_9510,N_4011,N_5329);
nor U9511 (N_9511,N_6315,N_7305);
nor U9512 (N_9512,N_6109,N_5093);
and U9513 (N_9513,N_7992,N_6400);
nand U9514 (N_9514,N_7012,N_6028);
and U9515 (N_9515,N_7080,N_7636);
and U9516 (N_9516,N_6526,N_7987);
or U9517 (N_9517,N_7602,N_5634);
nand U9518 (N_9518,N_6302,N_7039);
or U9519 (N_9519,N_7529,N_6653);
nor U9520 (N_9520,N_7167,N_4761);
nor U9521 (N_9521,N_7890,N_6063);
nor U9522 (N_9522,N_6960,N_7628);
or U9523 (N_9523,N_7084,N_4664);
nor U9524 (N_9524,N_5061,N_6284);
nand U9525 (N_9525,N_7531,N_4641);
or U9526 (N_9526,N_5840,N_7579);
nor U9527 (N_9527,N_7972,N_6195);
nor U9528 (N_9528,N_6673,N_5798);
and U9529 (N_9529,N_4630,N_7506);
nor U9530 (N_9530,N_5894,N_7783);
and U9531 (N_9531,N_7886,N_7612);
or U9532 (N_9532,N_5966,N_7072);
nand U9533 (N_9533,N_7253,N_6347);
nor U9534 (N_9534,N_6456,N_6731);
or U9535 (N_9535,N_6792,N_4847);
and U9536 (N_9536,N_5740,N_4826);
nor U9537 (N_9537,N_5856,N_7502);
or U9538 (N_9538,N_6843,N_7617);
or U9539 (N_9539,N_7790,N_6679);
or U9540 (N_9540,N_4150,N_5407);
and U9541 (N_9541,N_5677,N_6869);
and U9542 (N_9542,N_5818,N_4955);
and U9543 (N_9543,N_4355,N_7003);
and U9544 (N_9544,N_5349,N_5900);
nor U9545 (N_9545,N_4483,N_4154);
nor U9546 (N_9546,N_7651,N_4748);
nand U9547 (N_9547,N_5739,N_4948);
or U9548 (N_9548,N_4042,N_7476);
nand U9549 (N_9549,N_7775,N_5043);
or U9550 (N_9550,N_5809,N_5136);
nor U9551 (N_9551,N_7832,N_4533);
nor U9552 (N_9552,N_7357,N_7716);
and U9553 (N_9553,N_7004,N_4187);
and U9554 (N_9554,N_6072,N_6424);
and U9555 (N_9555,N_4562,N_5295);
nand U9556 (N_9556,N_4447,N_5023);
nand U9557 (N_9557,N_5453,N_4195);
nor U9558 (N_9558,N_7061,N_6875);
nor U9559 (N_9559,N_4145,N_7835);
nor U9560 (N_9560,N_4744,N_7643);
or U9561 (N_9561,N_6402,N_6951);
and U9562 (N_9562,N_5227,N_4252);
and U9563 (N_9563,N_5782,N_4441);
and U9564 (N_9564,N_7524,N_6820);
nand U9565 (N_9565,N_7710,N_4877);
nor U9566 (N_9566,N_7056,N_5495);
nor U9567 (N_9567,N_4092,N_7204);
and U9568 (N_9568,N_5009,N_4583);
or U9569 (N_9569,N_4063,N_6186);
nor U9570 (N_9570,N_5990,N_7825);
nor U9571 (N_9571,N_5450,N_5623);
and U9572 (N_9572,N_7827,N_6139);
nor U9573 (N_9573,N_5067,N_5831);
nand U9574 (N_9574,N_4525,N_7410);
or U9575 (N_9575,N_4609,N_5537);
nor U9576 (N_9576,N_4570,N_7331);
nor U9577 (N_9577,N_6553,N_7379);
and U9578 (N_9578,N_5257,N_7979);
and U9579 (N_9579,N_4594,N_6821);
or U9580 (N_9580,N_4118,N_4198);
nand U9581 (N_9581,N_4788,N_5676);
nand U9582 (N_9582,N_7073,N_4294);
nand U9583 (N_9583,N_4679,N_7271);
and U9584 (N_9584,N_6652,N_6722);
nand U9585 (N_9585,N_4146,N_6683);
or U9586 (N_9586,N_5336,N_7791);
or U9587 (N_9587,N_7245,N_5400);
nor U9588 (N_9588,N_6733,N_4479);
nor U9589 (N_9589,N_4923,N_5018);
nand U9590 (N_9590,N_6154,N_7836);
or U9591 (N_9591,N_6756,N_6306);
or U9592 (N_9592,N_5790,N_5580);
or U9593 (N_9593,N_6534,N_6029);
nor U9594 (N_9594,N_4090,N_4391);
or U9595 (N_9595,N_5115,N_4567);
nand U9596 (N_9596,N_7081,N_5700);
nand U9597 (N_9597,N_5531,N_7664);
or U9598 (N_9598,N_4794,N_4037);
and U9599 (N_9599,N_5108,N_7533);
and U9600 (N_9600,N_6953,N_4462);
or U9601 (N_9601,N_7789,N_4164);
and U9602 (N_9602,N_7428,N_7728);
nor U9603 (N_9603,N_6285,N_7147);
or U9604 (N_9604,N_4361,N_7135);
nor U9605 (N_9605,N_6805,N_6341);
or U9606 (N_9606,N_4414,N_6757);
nor U9607 (N_9607,N_5624,N_5471);
nand U9608 (N_9608,N_6241,N_7268);
nand U9609 (N_9609,N_4834,N_4392);
or U9610 (N_9610,N_5505,N_5865);
and U9611 (N_9611,N_4776,N_6099);
nor U9612 (N_9612,N_7436,N_6896);
and U9613 (N_9613,N_5374,N_4742);
nand U9614 (N_9614,N_6734,N_7723);
nand U9615 (N_9615,N_7671,N_7424);
or U9616 (N_9616,N_7568,N_5034);
nand U9617 (N_9617,N_5959,N_5151);
nand U9618 (N_9618,N_7551,N_5821);
nand U9619 (N_9619,N_5424,N_4101);
and U9620 (N_9620,N_4568,N_5099);
or U9621 (N_9621,N_6126,N_7737);
or U9622 (N_9622,N_4337,N_7385);
or U9623 (N_9623,N_6802,N_7532);
nand U9624 (N_9624,N_5762,N_7977);
nand U9625 (N_9625,N_4489,N_5652);
nand U9626 (N_9626,N_7712,N_7011);
nor U9627 (N_9627,N_5016,N_7741);
or U9628 (N_9628,N_5476,N_7092);
or U9629 (N_9629,N_6087,N_7968);
or U9630 (N_9630,N_4157,N_5029);
nand U9631 (N_9631,N_4833,N_7190);
nor U9632 (N_9632,N_6827,N_4888);
nand U9633 (N_9633,N_7390,N_6551);
or U9634 (N_9634,N_7313,N_4371);
and U9635 (N_9635,N_6410,N_6808);
or U9636 (N_9636,N_7445,N_4230);
or U9637 (N_9637,N_6021,N_4940);
nand U9638 (N_9638,N_7134,N_7937);
nor U9639 (N_9639,N_7717,N_7861);
or U9640 (N_9640,N_6287,N_4225);
nand U9641 (N_9641,N_6459,N_6428);
and U9642 (N_9642,N_5226,N_5408);
and U9643 (N_9643,N_7323,N_5913);
nor U9644 (N_9644,N_7236,N_7745);
or U9645 (N_9645,N_7536,N_6507);
or U9646 (N_9646,N_7604,N_5157);
nor U9647 (N_9647,N_6452,N_5118);
nand U9648 (N_9648,N_4911,N_6487);
nor U9649 (N_9649,N_6606,N_4420);
and U9650 (N_9650,N_5475,N_5813);
or U9651 (N_9651,N_4607,N_4936);
xor U9652 (N_9652,N_6248,N_6546);
or U9653 (N_9653,N_4531,N_6930);
nand U9654 (N_9654,N_7594,N_7630);
nor U9655 (N_9655,N_7867,N_7877);
and U9656 (N_9656,N_7919,N_7180);
and U9657 (N_9657,N_7848,N_7700);
nor U9658 (N_9658,N_5208,N_6755);
nand U9659 (N_9659,N_6782,N_4174);
nor U9660 (N_9660,N_4283,N_4718);
and U9661 (N_9661,N_5262,N_6002);
nand U9662 (N_9662,N_5526,N_6928);
or U9663 (N_9663,N_5895,N_5031);
nor U9664 (N_9664,N_6986,N_6932);
or U9665 (N_9665,N_4577,N_7627);
nor U9666 (N_9666,N_6567,N_5773);
nand U9667 (N_9667,N_6107,N_4868);
or U9668 (N_9668,N_5138,N_4072);
nand U9669 (N_9669,N_5963,N_7338);
nand U9670 (N_9670,N_6989,N_5572);
nor U9671 (N_9671,N_7971,N_4377);
nor U9672 (N_9672,N_5731,N_5255);
nand U9673 (N_9673,N_4739,N_4695);
and U9674 (N_9674,N_5844,N_6098);
nor U9675 (N_9675,N_4915,N_7794);
nor U9676 (N_9676,N_6505,N_7888);
nand U9677 (N_9677,N_5420,N_5191);
nor U9678 (N_9678,N_6677,N_6973);
nand U9679 (N_9679,N_5682,N_7074);
and U9680 (N_9680,N_7130,N_4291);
or U9681 (N_9681,N_6362,N_4470);
or U9682 (N_9682,N_4142,N_5281);
nand U9683 (N_9683,N_7692,N_5296);
nor U9684 (N_9684,N_7087,N_6961);
nor U9685 (N_9685,N_4231,N_6583);
and U9686 (N_9686,N_5120,N_7611);
or U9687 (N_9687,N_6411,N_5294);
nor U9688 (N_9688,N_6643,N_5887);
and U9689 (N_9689,N_6485,N_4183);
nor U9690 (N_9690,N_6867,N_4123);
nor U9691 (N_9691,N_5987,N_5909);
nand U9692 (N_9692,N_5563,N_7414);
nor U9693 (N_9693,N_4306,N_6527);
nand U9694 (N_9694,N_5004,N_5379);
nand U9695 (N_9695,N_6492,N_5879);
and U9696 (N_9696,N_7595,N_7406);
nor U9697 (N_9697,N_4551,N_6253);
nand U9698 (N_9698,N_5026,N_7566);
or U9699 (N_9699,N_7286,N_4349);
nor U9700 (N_9700,N_7082,N_6323);
nand U9701 (N_9701,N_5122,N_4878);
nor U9702 (N_9702,N_7548,N_6494);
and U9703 (N_9703,N_4634,N_5423);
nand U9704 (N_9704,N_7290,N_7883);
or U9705 (N_9705,N_7094,N_4827);
and U9706 (N_9706,N_6283,N_5561);
nand U9707 (N_9707,N_6134,N_7415);
or U9708 (N_9708,N_5814,N_4836);
nand U9709 (N_9709,N_6305,N_4732);
nand U9710 (N_9710,N_7069,N_7144);
nand U9711 (N_9711,N_7342,N_5456);
nor U9712 (N_9712,N_6446,N_7801);
or U9713 (N_9713,N_6267,N_7927);
or U9714 (N_9714,N_7821,N_7755);
nand U9715 (N_9715,N_5931,N_7713);
or U9716 (N_9716,N_5686,N_7661);
nand U9717 (N_9717,N_5743,N_6045);
nor U9718 (N_9718,N_5306,N_6509);
or U9719 (N_9719,N_5147,N_7922);
or U9720 (N_9720,N_6012,N_7744);
nor U9721 (N_9721,N_7753,N_4889);
nand U9722 (N_9722,N_5902,N_5718);
nor U9723 (N_9723,N_6242,N_7695);
nor U9724 (N_9724,N_7198,N_5363);
and U9725 (N_9725,N_7739,N_6482);
and U9726 (N_9726,N_7462,N_4247);
and U9727 (N_9727,N_6760,N_6543);
or U9728 (N_9728,N_6671,N_5270);
and U9729 (N_9729,N_7656,N_5391);
nor U9730 (N_9730,N_4261,N_5185);
and U9731 (N_9731,N_6157,N_5117);
and U9732 (N_9732,N_6252,N_5869);
and U9733 (N_9733,N_6152,N_5588);
and U9734 (N_9734,N_7701,N_6971);
nand U9735 (N_9735,N_5446,N_7165);
and U9736 (N_9736,N_6650,N_7399);
and U9737 (N_9737,N_5331,N_6592);
or U9738 (N_9738,N_5233,N_7281);
nor U9739 (N_9739,N_6121,N_4421);
nor U9740 (N_9740,N_4929,N_7463);
nand U9741 (N_9741,N_6745,N_7377);
nor U9742 (N_9742,N_4041,N_4764);
or U9743 (N_9743,N_6370,N_7501);
and U9744 (N_9744,N_4200,N_5250);
nand U9745 (N_9745,N_7898,N_4066);
nand U9746 (N_9746,N_7058,N_4639);
or U9747 (N_9747,N_6585,N_5535);
nor U9748 (N_9748,N_4537,N_6579);
nor U9749 (N_9749,N_5734,N_6920);
and U9750 (N_9750,N_7417,N_5317);
nand U9751 (N_9751,N_6084,N_4215);
or U9752 (N_9752,N_7142,N_5764);
nor U9753 (N_9753,N_4010,N_4293);
and U9754 (N_9754,N_7905,N_6707);
or U9755 (N_9755,N_5991,N_4584);
and U9756 (N_9756,N_4815,N_4775);
and U9757 (N_9757,N_7797,N_4633);
nor U9758 (N_9758,N_5617,N_5881);
nand U9759 (N_9759,N_5193,N_6275);
nor U9760 (N_9760,N_5011,N_7093);
nand U9761 (N_9761,N_6365,N_7401);
and U9762 (N_9762,N_6938,N_5555);
nand U9763 (N_9763,N_5348,N_6568);
or U9764 (N_9764,N_4013,N_7472);
and U9765 (N_9765,N_7199,N_5181);
nand U9766 (N_9766,N_6458,N_7901);
nand U9767 (N_9767,N_6559,N_6576);
or U9768 (N_9768,N_4468,N_4449);
or U9769 (N_9769,N_4385,N_5986);
nor U9770 (N_9770,N_4398,N_4173);
nand U9771 (N_9771,N_6450,N_5675);
and U9772 (N_9772,N_6413,N_6700);
and U9773 (N_9773,N_5448,N_5366);
and U9774 (N_9774,N_5465,N_4268);
nor U9775 (N_9775,N_5221,N_7105);
and U9776 (N_9776,N_6264,N_4904);
or U9777 (N_9777,N_6844,N_5188);
and U9778 (N_9778,N_6229,N_7178);
nand U9779 (N_9779,N_6211,N_7926);
nor U9780 (N_9780,N_7761,N_7572);
nand U9781 (N_9781,N_4482,N_4928);
nor U9782 (N_9782,N_6626,N_4289);
and U9783 (N_9783,N_5581,N_4566);
and U9784 (N_9784,N_7895,N_7696);
nand U9785 (N_9785,N_4593,N_5438);
and U9786 (N_9786,N_6655,N_7569);
or U9787 (N_9787,N_7976,N_4038);
and U9788 (N_9788,N_7078,N_6289);
nand U9789 (N_9789,N_4015,N_4167);
and U9790 (N_9790,N_6168,N_7961);
and U9791 (N_9791,N_6669,N_7174);
nor U9792 (N_9792,N_5671,N_4884);
or U9793 (N_9793,N_6112,N_4469);
nand U9794 (N_9794,N_7029,N_7631);
nand U9795 (N_9795,N_4055,N_4401);
nor U9796 (N_9796,N_4243,N_5443);
nor U9797 (N_9797,N_5946,N_4817);
nand U9798 (N_9798,N_6632,N_5753);
nand U9799 (N_9799,N_7562,N_4471);
nor U9800 (N_9800,N_7034,N_4065);
or U9801 (N_9801,N_4890,N_6110);
nand U9802 (N_9802,N_5565,N_4033);
nand U9803 (N_9803,N_7067,N_5504);
nor U9804 (N_9804,N_4812,N_7247);
and U9805 (N_9805,N_7724,N_5825);
and U9806 (N_9806,N_5180,N_4628);
nor U9807 (N_9807,N_5472,N_5839);
and U9808 (N_9808,N_4147,N_6799);
nor U9809 (N_9809,N_4002,N_4672);
or U9810 (N_9810,N_6993,N_5655);
or U9811 (N_9811,N_6480,N_6198);
nor U9812 (N_9812,N_5781,N_6763);
or U9813 (N_9813,N_4708,N_5916);
and U9814 (N_9814,N_5746,N_5979);
or U9815 (N_9815,N_7277,N_7289);
nand U9816 (N_9816,N_4117,N_4121);
and U9817 (N_9817,N_5353,N_4492);
or U9818 (N_9818,N_7389,N_6133);
or U9819 (N_9819,N_7691,N_4162);
nor U9820 (N_9820,N_4795,N_5613);
nor U9821 (N_9821,N_4722,N_7736);
nand U9822 (N_9822,N_4328,N_5060);
and U9823 (N_9823,N_5378,N_5767);
nor U9824 (N_9824,N_4831,N_5412);
or U9825 (N_9825,N_6314,N_5485);
nor U9826 (N_9826,N_5440,N_5627);
or U9827 (N_9827,N_4707,N_5419);
nand U9828 (N_9828,N_5672,N_4341);
xnor U9829 (N_9829,N_6531,N_5501);
nor U9830 (N_9830,N_6645,N_7070);
and U9831 (N_9831,N_5473,N_6696);
xnor U9832 (N_9832,N_5062,N_5778);
nor U9833 (N_9833,N_7507,N_4934);
nor U9834 (N_9834,N_6416,N_6806);
nor U9835 (N_9835,N_4602,N_6607);
nand U9836 (N_9836,N_7496,N_7259);
and U9837 (N_9837,N_5548,N_4021);
or U9838 (N_9838,N_4116,N_5530);
and U9839 (N_9839,N_6223,N_4598);
and U9840 (N_9840,N_6192,N_4348);
nor U9841 (N_9841,N_6220,N_4996);
xor U9842 (N_9842,N_4281,N_5482);
nand U9843 (N_9843,N_7086,N_5054);
nor U9844 (N_9844,N_6851,N_4422);
and U9845 (N_9845,N_6889,N_5095);
or U9846 (N_9846,N_6292,N_4267);
nor U9847 (N_9847,N_7335,N_5381);
and U9848 (N_9848,N_7220,N_5429);
nor U9849 (N_9849,N_6603,N_5050);
nand U9850 (N_9850,N_4001,N_6910);
or U9851 (N_9851,N_4323,N_7951);
or U9852 (N_9852,N_6849,N_5618);
nor U9853 (N_9853,N_4820,N_6231);
nor U9854 (N_9854,N_7434,N_4075);
nand U9855 (N_9855,N_4807,N_6858);
or U9856 (N_9856,N_4893,N_5864);
nand U9857 (N_9857,N_5707,N_7405);
nor U9858 (N_9858,N_4604,N_7433);
nand U9859 (N_9859,N_4084,N_7850);
and U9860 (N_9860,N_7555,N_6811);
nand U9861 (N_9861,N_5044,N_6379);
or U9862 (N_9862,N_4095,N_5833);
nand U9863 (N_9863,N_7933,N_7033);
and U9864 (N_9864,N_5326,N_6327);
nand U9865 (N_9865,N_6018,N_7326);
or U9866 (N_9866,N_4228,N_7225);
nand U9867 (N_9867,N_5955,N_4415);
or U9868 (N_9868,N_4109,N_6077);
nand U9869 (N_9869,N_6550,N_6280);
or U9870 (N_9870,N_4755,N_4073);
or U9871 (N_9871,N_4263,N_5941);
nor U9872 (N_9872,N_7804,N_7205);
nand U9873 (N_9873,N_5626,N_4110);
nand U9874 (N_9874,N_7537,N_5384);
nand U9875 (N_9875,N_5404,N_4576);
xor U9876 (N_9876,N_5131,N_6105);
nor U9877 (N_9877,N_6363,N_4436);
nor U9878 (N_9878,N_7145,N_4529);
nor U9879 (N_9879,N_6193,N_7539);
nor U9880 (N_9880,N_6335,N_7273);
nor U9881 (N_9881,N_5510,N_7216);
nor U9882 (N_9882,N_6754,N_4132);
and U9883 (N_9883,N_7733,N_4180);
and U9884 (N_9884,N_7076,N_7914);
and U9885 (N_9885,N_6367,N_4257);
nor U9886 (N_9886,N_4941,N_6766);
nor U9887 (N_9887,N_4851,N_4989);
nor U9888 (N_9888,N_6382,N_6443);
xnor U9889 (N_9889,N_5517,N_5264);
nand U9890 (N_9890,N_5546,N_5663);
nor U9891 (N_9891,N_4159,N_4078);
nand U9892 (N_9892,N_6031,N_5316);
and U9893 (N_9893,N_5878,N_7432);
nor U9894 (N_9894,N_5641,N_5774);
nor U9895 (N_9895,N_7767,N_6908);
nand U9896 (N_9896,N_4304,N_4728);
nand U9897 (N_9897,N_5846,N_5335);
and U9898 (N_9898,N_5195,N_6392);
xnor U9899 (N_9899,N_7706,N_5266);
nand U9900 (N_9900,N_5891,N_6414);
nor U9901 (N_9901,N_5207,N_5035);
nor U9902 (N_9902,N_4152,N_7054);
and U9903 (N_9903,N_6523,N_7875);
nor U9904 (N_9904,N_4779,N_6061);
nor U9905 (N_9905,N_5274,N_4838);
and U9906 (N_9906,N_5297,N_6829);
nor U9907 (N_9907,N_4861,N_7857);
or U9908 (N_9908,N_6764,N_7650);
nand U9909 (N_9909,N_4580,N_5132);
nand U9910 (N_9910,N_6483,N_7169);
and U9911 (N_9911,N_5387,N_4153);
nor U9912 (N_9912,N_5602,N_6448);
nand U9913 (N_9913,N_4212,N_7209);
or U9914 (N_9914,N_7764,N_4606);
nand U9915 (N_9915,N_5621,N_5124);
nor U9916 (N_9916,N_5172,N_7297);
nor U9917 (N_9917,N_5334,N_6544);
nand U9918 (N_9918,N_7799,N_6427);
or U9919 (N_9919,N_7834,N_4356);
and U9920 (N_9920,N_5375,N_6470);
nand U9921 (N_9921,N_5337,N_5253);
or U9922 (N_9922,N_6200,N_7669);
nor U9923 (N_9923,N_7344,N_4381);
nand U9924 (N_9924,N_7201,N_5064);
xnor U9925 (N_9925,N_5416,N_5219);
nand U9926 (N_9926,N_7727,N_6141);
nand U9927 (N_9927,N_4192,N_7511);
and U9928 (N_9928,N_5796,N_5494);
or U9929 (N_9929,N_7040,N_4712);
nor U9930 (N_9930,N_6758,N_5711);
and U9931 (N_9931,N_6472,N_5647);
or U9932 (N_9932,N_5201,N_7160);
or U9933 (N_9933,N_6638,N_4924);
or U9934 (N_9934,N_5452,N_4400);
or U9935 (N_9935,N_7693,N_4845);
nand U9936 (N_9936,N_6417,N_5305);
or U9937 (N_9937,N_4406,N_7173);
or U9938 (N_9938,N_5571,N_7621);
and U9939 (N_9939,N_5670,N_4032);
nor U9940 (N_9940,N_7158,N_7674);
nand U9941 (N_9941,N_4952,N_4746);
nand U9942 (N_9942,N_4405,N_5125);
nand U9943 (N_9943,N_4239,N_4474);
or U9944 (N_9944,N_5021,N_6826);
and U9945 (N_9945,N_5919,N_4036);
nor U9946 (N_9946,N_4387,N_5454);
nor U9947 (N_9947,N_6852,N_6128);
or U9948 (N_9948,N_5038,N_6384);
or U9949 (N_9949,N_7935,N_7088);
and U9950 (N_9950,N_4052,N_7853);
nor U9951 (N_9951,N_5319,N_5447);
or U9952 (N_9952,N_4617,N_7940);
nor U9953 (N_9953,N_7601,N_6815);
or U9954 (N_9954,N_7388,N_4894);
nor U9955 (N_9955,N_4969,N_7870);
nor U9956 (N_9956,N_4625,N_7392);
nand U9957 (N_9957,N_6954,N_4963);
nor U9958 (N_9958,N_7747,N_7430);
and U9959 (N_9959,N_5398,N_4967);
nor U9960 (N_9960,N_6933,N_7098);
nand U9961 (N_9961,N_4175,N_7957);
and U9962 (N_9962,N_6682,N_4766);
nand U9963 (N_9963,N_4702,N_7720);
or U9964 (N_9964,N_5829,N_4675);
and U9965 (N_9965,N_4442,N_5529);
nand U9966 (N_9966,N_4427,N_6296);
or U9967 (N_9967,N_6859,N_5395);
nor U9968 (N_9968,N_5177,N_4460);
nand U9969 (N_9969,N_5706,N_4806);
and U9970 (N_9970,N_5544,N_4813);
nand U9971 (N_9971,N_4188,N_6260);
nor U9972 (N_9972,N_7109,N_5943);
and U9973 (N_9973,N_5590,N_5589);
or U9974 (N_9974,N_4765,N_6988);
nor U9975 (N_9975,N_5868,N_6864);
nor U9976 (N_9976,N_5100,N_4309);
or U9977 (N_9977,N_4190,N_4126);
and U9978 (N_9978,N_7416,N_7013);
and U9979 (N_9979,N_4874,N_7027);
and U9980 (N_9980,N_4572,N_6333);
nor U9981 (N_9981,N_5148,N_6197);
and U9982 (N_9982,N_7944,N_6776);
and U9983 (N_9983,N_5403,N_5802);
nand U9984 (N_9984,N_5889,N_6967);
or U9985 (N_9985,N_6770,N_5383);
or U9986 (N_9986,N_6847,N_7288);
nand U9987 (N_9987,N_6793,N_7345);
nor U9988 (N_9988,N_4715,N_5795);
nor U9989 (N_9989,N_4048,N_7324);
nand U9990 (N_9990,N_5804,N_5036);
nand U9991 (N_9991,N_6013,N_5402);
nand U9992 (N_9992,N_5702,N_6616);
and U9993 (N_9993,N_5392,N_5853);
or U9994 (N_9994,N_5199,N_4843);
and U9995 (N_9995,N_4509,N_4244);
nand U9996 (N_9996,N_6026,N_4865);
nor U9997 (N_9997,N_4931,N_5970);
nor U9998 (N_9998,N_7876,N_4691);
nor U9999 (N_9999,N_5893,N_7874);
or U10000 (N_10000,N_5513,N_7156);
and U10001 (N_10001,N_6280,N_5572);
nor U10002 (N_10002,N_4409,N_4134);
or U10003 (N_10003,N_7564,N_5575);
or U10004 (N_10004,N_6533,N_5690);
nor U10005 (N_10005,N_7072,N_5191);
and U10006 (N_10006,N_5315,N_6766);
or U10007 (N_10007,N_6333,N_6134);
and U10008 (N_10008,N_4881,N_7366);
nand U10009 (N_10009,N_4091,N_5565);
and U10010 (N_10010,N_7782,N_5755);
nand U10011 (N_10011,N_5809,N_6735);
or U10012 (N_10012,N_7633,N_5127);
and U10013 (N_10013,N_5296,N_7991);
and U10014 (N_10014,N_4331,N_5475);
and U10015 (N_10015,N_5562,N_7782);
nand U10016 (N_10016,N_7044,N_4752);
or U10017 (N_10017,N_7680,N_7724);
and U10018 (N_10018,N_5475,N_5995);
nor U10019 (N_10019,N_7809,N_6812);
nor U10020 (N_10020,N_6555,N_4251);
nor U10021 (N_10021,N_6423,N_7122);
and U10022 (N_10022,N_5055,N_7994);
nor U10023 (N_10023,N_6814,N_5184);
nand U10024 (N_10024,N_7288,N_6235);
nor U10025 (N_10025,N_4831,N_4779);
nand U10026 (N_10026,N_5046,N_4147);
nor U10027 (N_10027,N_5014,N_7082);
nand U10028 (N_10028,N_5631,N_4469);
nor U10029 (N_10029,N_4463,N_5374);
nand U10030 (N_10030,N_5916,N_5466);
nand U10031 (N_10031,N_6051,N_6526);
or U10032 (N_10032,N_4318,N_7014);
nand U10033 (N_10033,N_5571,N_6335);
nand U10034 (N_10034,N_4990,N_6291);
and U10035 (N_10035,N_4610,N_7914);
or U10036 (N_10036,N_7644,N_7064);
nand U10037 (N_10037,N_5464,N_6766);
nor U10038 (N_10038,N_5929,N_7397);
or U10039 (N_10039,N_5646,N_5124);
and U10040 (N_10040,N_4327,N_7464);
nor U10041 (N_10041,N_5466,N_4708);
or U10042 (N_10042,N_6752,N_5274);
nand U10043 (N_10043,N_4079,N_6262);
nand U10044 (N_10044,N_6509,N_7019);
nand U10045 (N_10045,N_5388,N_6473);
nor U10046 (N_10046,N_5523,N_7034);
nor U10047 (N_10047,N_7446,N_5941);
and U10048 (N_10048,N_5780,N_7507);
and U10049 (N_10049,N_5905,N_5604);
or U10050 (N_10050,N_6129,N_7354);
nand U10051 (N_10051,N_4225,N_6558);
and U10052 (N_10052,N_5855,N_5498);
nor U10053 (N_10053,N_5368,N_6886);
nand U10054 (N_10054,N_6601,N_4503);
and U10055 (N_10055,N_4475,N_7244);
nand U10056 (N_10056,N_4859,N_4340);
nand U10057 (N_10057,N_5055,N_6887);
nand U10058 (N_10058,N_6345,N_6497);
or U10059 (N_10059,N_6162,N_6978);
nor U10060 (N_10060,N_7719,N_4740);
nor U10061 (N_10061,N_5078,N_4694);
nor U10062 (N_10062,N_5887,N_7635);
nor U10063 (N_10063,N_7640,N_6984);
nor U10064 (N_10064,N_7755,N_5750);
and U10065 (N_10065,N_5508,N_5311);
nor U10066 (N_10066,N_5376,N_6549);
and U10067 (N_10067,N_5134,N_7863);
nand U10068 (N_10068,N_5533,N_6433);
nor U10069 (N_10069,N_6144,N_5798);
and U10070 (N_10070,N_5036,N_4231);
nand U10071 (N_10071,N_7018,N_5629);
or U10072 (N_10072,N_7118,N_7629);
or U10073 (N_10073,N_6283,N_4666);
nand U10074 (N_10074,N_6804,N_7747);
or U10075 (N_10075,N_6684,N_4112);
and U10076 (N_10076,N_6003,N_7427);
and U10077 (N_10077,N_6219,N_7163);
and U10078 (N_10078,N_4767,N_6843);
or U10079 (N_10079,N_6847,N_5766);
nor U10080 (N_10080,N_7261,N_6065);
or U10081 (N_10081,N_4502,N_4931);
or U10082 (N_10082,N_4983,N_7103);
and U10083 (N_10083,N_4636,N_5269);
or U10084 (N_10084,N_5412,N_4524);
and U10085 (N_10085,N_7302,N_4660);
nand U10086 (N_10086,N_7167,N_4766);
or U10087 (N_10087,N_7069,N_4637);
or U10088 (N_10088,N_5021,N_5092);
nand U10089 (N_10089,N_5108,N_6924);
and U10090 (N_10090,N_6701,N_5961);
and U10091 (N_10091,N_5757,N_7272);
nand U10092 (N_10092,N_7878,N_6649);
or U10093 (N_10093,N_5967,N_5549);
nand U10094 (N_10094,N_4007,N_4516);
nand U10095 (N_10095,N_4489,N_4458);
and U10096 (N_10096,N_6059,N_4688);
nand U10097 (N_10097,N_7409,N_7797);
nand U10098 (N_10098,N_4005,N_5768);
nor U10099 (N_10099,N_5709,N_6626);
nor U10100 (N_10100,N_4479,N_5275);
nor U10101 (N_10101,N_5255,N_7316);
or U10102 (N_10102,N_5667,N_4156);
nand U10103 (N_10103,N_4452,N_5319);
or U10104 (N_10104,N_6751,N_5624);
nor U10105 (N_10105,N_6558,N_4776);
or U10106 (N_10106,N_5560,N_6624);
xnor U10107 (N_10107,N_7501,N_4129);
and U10108 (N_10108,N_6532,N_6495);
nor U10109 (N_10109,N_7925,N_7090);
and U10110 (N_10110,N_6768,N_5675);
or U10111 (N_10111,N_5829,N_4836);
or U10112 (N_10112,N_5605,N_5342);
and U10113 (N_10113,N_6706,N_5669);
nor U10114 (N_10114,N_5174,N_4590);
or U10115 (N_10115,N_6002,N_4647);
or U10116 (N_10116,N_5849,N_5934);
or U10117 (N_10117,N_7642,N_4446);
and U10118 (N_10118,N_4682,N_4307);
or U10119 (N_10119,N_4708,N_4214);
and U10120 (N_10120,N_4880,N_5769);
and U10121 (N_10121,N_5352,N_4130);
or U10122 (N_10122,N_5542,N_5412);
nand U10123 (N_10123,N_6883,N_5273);
and U10124 (N_10124,N_5256,N_7679);
nand U10125 (N_10125,N_6835,N_7517);
and U10126 (N_10126,N_5005,N_4322);
nor U10127 (N_10127,N_4927,N_7378);
and U10128 (N_10128,N_4850,N_6578);
and U10129 (N_10129,N_6864,N_5284);
or U10130 (N_10130,N_7094,N_6038);
nand U10131 (N_10131,N_5059,N_5211);
or U10132 (N_10132,N_4061,N_6185);
nand U10133 (N_10133,N_4197,N_7836);
and U10134 (N_10134,N_5316,N_4339);
nand U10135 (N_10135,N_4767,N_4581);
nor U10136 (N_10136,N_5255,N_5316);
nand U10137 (N_10137,N_6477,N_6014);
and U10138 (N_10138,N_6570,N_7073);
or U10139 (N_10139,N_6824,N_6261);
or U10140 (N_10140,N_6967,N_7773);
and U10141 (N_10141,N_5256,N_7082);
nand U10142 (N_10142,N_4438,N_5578);
and U10143 (N_10143,N_4397,N_4009);
or U10144 (N_10144,N_4040,N_4981);
and U10145 (N_10145,N_5230,N_4929);
nor U10146 (N_10146,N_7112,N_7232);
nor U10147 (N_10147,N_6881,N_5496);
nand U10148 (N_10148,N_7787,N_7857);
nor U10149 (N_10149,N_6557,N_7547);
and U10150 (N_10150,N_5216,N_7331);
and U10151 (N_10151,N_7610,N_6665);
or U10152 (N_10152,N_6028,N_6896);
nor U10153 (N_10153,N_4698,N_5367);
nor U10154 (N_10154,N_5209,N_4422);
and U10155 (N_10155,N_6470,N_4709);
or U10156 (N_10156,N_4561,N_5661);
and U10157 (N_10157,N_7535,N_5532);
and U10158 (N_10158,N_5656,N_6725);
nand U10159 (N_10159,N_7532,N_7600);
or U10160 (N_10160,N_4280,N_7896);
nand U10161 (N_10161,N_7751,N_7555);
nand U10162 (N_10162,N_7443,N_6756);
xor U10163 (N_10163,N_6970,N_7387);
or U10164 (N_10164,N_5568,N_7543);
nand U10165 (N_10165,N_7636,N_7207);
nor U10166 (N_10166,N_6339,N_4846);
or U10167 (N_10167,N_7320,N_4784);
nand U10168 (N_10168,N_5423,N_6610);
nor U10169 (N_10169,N_7301,N_4662);
nor U10170 (N_10170,N_7284,N_4919);
nand U10171 (N_10171,N_7521,N_6921);
nand U10172 (N_10172,N_5915,N_6365);
nand U10173 (N_10173,N_4839,N_6744);
and U10174 (N_10174,N_5773,N_6304);
and U10175 (N_10175,N_6681,N_4498);
xor U10176 (N_10176,N_5648,N_4979);
nor U10177 (N_10177,N_6323,N_4410);
and U10178 (N_10178,N_6818,N_5474);
nor U10179 (N_10179,N_4338,N_7309);
and U10180 (N_10180,N_5389,N_4943);
nand U10181 (N_10181,N_7812,N_6427);
and U10182 (N_10182,N_7278,N_6082);
nand U10183 (N_10183,N_4053,N_7204);
nor U10184 (N_10184,N_5489,N_5414);
or U10185 (N_10185,N_4242,N_7154);
and U10186 (N_10186,N_5404,N_6312);
or U10187 (N_10187,N_5997,N_5373);
nor U10188 (N_10188,N_5098,N_6353);
nor U10189 (N_10189,N_7131,N_7891);
and U10190 (N_10190,N_7158,N_7323);
or U10191 (N_10191,N_7225,N_4096);
nand U10192 (N_10192,N_7230,N_5420);
and U10193 (N_10193,N_4060,N_5997);
nand U10194 (N_10194,N_5111,N_5833);
nor U10195 (N_10195,N_6824,N_7468);
and U10196 (N_10196,N_4252,N_5254);
or U10197 (N_10197,N_4182,N_7650);
nor U10198 (N_10198,N_5236,N_5213);
nor U10199 (N_10199,N_6113,N_6578);
nor U10200 (N_10200,N_4402,N_4347);
nor U10201 (N_10201,N_6705,N_7216);
or U10202 (N_10202,N_7040,N_4964);
nor U10203 (N_10203,N_7083,N_6997);
or U10204 (N_10204,N_6984,N_4568);
nand U10205 (N_10205,N_4581,N_7240);
nor U10206 (N_10206,N_4209,N_6499);
nor U10207 (N_10207,N_4563,N_4130);
nand U10208 (N_10208,N_4427,N_7896);
xor U10209 (N_10209,N_7303,N_6123);
nand U10210 (N_10210,N_4323,N_4763);
nor U10211 (N_10211,N_5177,N_5943);
and U10212 (N_10212,N_6432,N_5193);
and U10213 (N_10213,N_5359,N_4037);
nor U10214 (N_10214,N_5141,N_5996);
nor U10215 (N_10215,N_6477,N_5818);
nand U10216 (N_10216,N_6270,N_6392);
and U10217 (N_10217,N_6540,N_6423);
nand U10218 (N_10218,N_5222,N_7912);
and U10219 (N_10219,N_6475,N_5337);
and U10220 (N_10220,N_4124,N_6098);
nand U10221 (N_10221,N_6689,N_4100);
or U10222 (N_10222,N_5248,N_6053);
nand U10223 (N_10223,N_6773,N_7658);
or U10224 (N_10224,N_7970,N_5653);
and U10225 (N_10225,N_7572,N_5456);
nor U10226 (N_10226,N_7782,N_4701);
and U10227 (N_10227,N_4407,N_5652);
and U10228 (N_10228,N_5617,N_7790);
nor U10229 (N_10229,N_4379,N_5158);
or U10230 (N_10230,N_6165,N_4128);
or U10231 (N_10231,N_7440,N_5137);
nand U10232 (N_10232,N_6839,N_5505);
or U10233 (N_10233,N_4088,N_6399);
and U10234 (N_10234,N_4068,N_6771);
nand U10235 (N_10235,N_6191,N_7324);
nand U10236 (N_10236,N_7826,N_7425);
nor U10237 (N_10237,N_7110,N_7687);
nand U10238 (N_10238,N_4287,N_5974);
or U10239 (N_10239,N_5017,N_7160);
and U10240 (N_10240,N_4439,N_6401);
or U10241 (N_10241,N_6459,N_4667);
nand U10242 (N_10242,N_4316,N_6161);
nand U10243 (N_10243,N_6422,N_7347);
nand U10244 (N_10244,N_4009,N_7613);
or U10245 (N_10245,N_7665,N_6758);
and U10246 (N_10246,N_7511,N_4318);
nand U10247 (N_10247,N_5563,N_6898);
or U10248 (N_10248,N_7340,N_7394);
nand U10249 (N_10249,N_5083,N_5765);
nand U10250 (N_10250,N_4840,N_7642);
or U10251 (N_10251,N_4258,N_5645);
nand U10252 (N_10252,N_5479,N_6784);
or U10253 (N_10253,N_5804,N_4450);
and U10254 (N_10254,N_5461,N_4112);
and U10255 (N_10255,N_4726,N_7826);
and U10256 (N_10256,N_4395,N_7144);
or U10257 (N_10257,N_5847,N_4609);
nor U10258 (N_10258,N_6259,N_5170);
and U10259 (N_10259,N_4744,N_4868);
nor U10260 (N_10260,N_4830,N_7764);
nor U10261 (N_10261,N_6743,N_5829);
nor U10262 (N_10262,N_7319,N_7419);
and U10263 (N_10263,N_6460,N_6217);
and U10264 (N_10264,N_7240,N_4664);
and U10265 (N_10265,N_7206,N_7389);
and U10266 (N_10266,N_5047,N_7463);
and U10267 (N_10267,N_6369,N_7786);
nand U10268 (N_10268,N_6150,N_6335);
nor U10269 (N_10269,N_7648,N_4186);
or U10270 (N_10270,N_5944,N_6440);
or U10271 (N_10271,N_5618,N_7538);
and U10272 (N_10272,N_6963,N_4381);
or U10273 (N_10273,N_7397,N_4570);
or U10274 (N_10274,N_5742,N_6950);
nand U10275 (N_10275,N_7014,N_7489);
or U10276 (N_10276,N_6552,N_5432);
or U10277 (N_10277,N_4080,N_7759);
nand U10278 (N_10278,N_5732,N_5773);
or U10279 (N_10279,N_7656,N_5211);
nor U10280 (N_10280,N_5726,N_6565);
nor U10281 (N_10281,N_5457,N_5088);
and U10282 (N_10282,N_4091,N_4642);
or U10283 (N_10283,N_5489,N_4811);
nor U10284 (N_10284,N_5804,N_4345);
nor U10285 (N_10285,N_7453,N_4701);
nand U10286 (N_10286,N_4497,N_7870);
nand U10287 (N_10287,N_4039,N_6289);
nand U10288 (N_10288,N_7899,N_6285);
xor U10289 (N_10289,N_4668,N_6329);
nand U10290 (N_10290,N_6333,N_6184);
nand U10291 (N_10291,N_4532,N_6004);
nand U10292 (N_10292,N_6900,N_4250);
and U10293 (N_10293,N_4677,N_4862);
nor U10294 (N_10294,N_5274,N_4047);
nor U10295 (N_10295,N_4300,N_5276);
or U10296 (N_10296,N_6008,N_5788);
or U10297 (N_10297,N_5321,N_7606);
or U10298 (N_10298,N_6082,N_6815);
nor U10299 (N_10299,N_6530,N_7399);
or U10300 (N_10300,N_4443,N_5501);
and U10301 (N_10301,N_7528,N_4681);
nor U10302 (N_10302,N_4008,N_6540);
and U10303 (N_10303,N_5280,N_7471);
nor U10304 (N_10304,N_6047,N_7733);
and U10305 (N_10305,N_7957,N_7766);
nand U10306 (N_10306,N_4049,N_4816);
or U10307 (N_10307,N_4085,N_6486);
and U10308 (N_10308,N_4201,N_7459);
or U10309 (N_10309,N_6587,N_7162);
or U10310 (N_10310,N_7860,N_4071);
or U10311 (N_10311,N_5344,N_7992);
nand U10312 (N_10312,N_4823,N_7870);
or U10313 (N_10313,N_6422,N_4389);
and U10314 (N_10314,N_4909,N_7607);
and U10315 (N_10315,N_6736,N_6281);
or U10316 (N_10316,N_4356,N_6933);
or U10317 (N_10317,N_5454,N_7641);
nand U10318 (N_10318,N_5454,N_5310);
and U10319 (N_10319,N_5889,N_4921);
and U10320 (N_10320,N_4357,N_6063);
nand U10321 (N_10321,N_6406,N_6719);
and U10322 (N_10322,N_4179,N_7337);
nand U10323 (N_10323,N_4286,N_6674);
and U10324 (N_10324,N_6675,N_6880);
or U10325 (N_10325,N_5495,N_5825);
nor U10326 (N_10326,N_4865,N_6967);
nor U10327 (N_10327,N_4139,N_4238);
or U10328 (N_10328,N_7102,N_4250);
and U10329 (N_10329,N_5669,N_7369);
nand U10330 (N_10330,N_6398,N_5966);
nand U10331 (N_10331,N_7227,N_6439);
or U10332 (N_10332,N_5532,N_7817);
nand U10333 (N_10333,N_6259,N_4475);
or U10334 (N_10334,N_5215,N_7043);
nor U10335 (N_10335,N_5687,N_6207);
nor U10336 (N_10336,N_6929,N_6781);
nor U10337 (N_10337,N_6346,N_4343);
nor U10338 (N_10338,N_6836,N_4334);
and U10339 (N_10339,N_6470,N_6266);
nor U10340 (N_10340,N_6418,N_6091);
nand U10341 (N_10341,N_7251,N_6736);
or U10342 (N_10342,N_5184,N_4959);
nor U10343 (N_10343,N_5369,N_4409);
nand U10344 (N_10344,N_5199,N_7819);
nand U10345 (N_10345,N_6843,N_6708);
nand U10346 (N_10346,N_4122,N_5365);
or U10347 (N_10347,N_6981,N_7136);
and U10348 (N_10348,N_6400,N_4696);
or U10349 (N_10349,N_4172,N_6965);
or U10350 (N_10350,N_5649,N_5486);
nand U10351 (N_10351,N_5112,N_5183);
and U10352 (N_10352,N_6462,N_5301);
or U10353 (N_10353,N_6950,N_6128);
nand U10354 (N_10354,N_5152,N_7650);
nand U10355 (N_10355,N_6700,N_6826);
nor U10356 (N_10356,N_6632,N_7874);
and U10357 (N_10357,N_6719,N_6620);
nand U10358 (N_10358,N_5649,N_4619);
or U10359 (N_10359,N_4157,N_7962);
nand U10360 (N_10360,N_6691,N_5044);
nor U10361 (N_10361,N_5237,N_4729);
nand U10362 (N_10362,N_4895,N_4085);
nand U10363 (N_10363,N_7312,N_6207);
and U10364 (N_10364,N_4131,N_7461);
nand U10365 (N_10365,N_7234,N_7466);
nand U10366 (N_10366,N_7560,N_5074);
nor U10367 (N_10367,N_6078,N_6537);
nand U10368 (N_10368,N_7504,N_7028);
nand U10369 (N_10369,N_4408,N_6610);
nand U10370 (N_10370,N_5390,N_5653);
nand U10371 (N_10371,N_7233,N_7080);
nor U10372 (N_10372,N_6472,N_5656);
nor U10373 (N_10373,N_4307,N_6522);
or U10374 (N_10374,N_7953,N_4199);
and U10375 (N_10375,N_4062,N_6139);
or U10376 (N_10376,N_6528,N_6601);
nand U10377 (N_10377,N_6527,N_7726);
nor U10378 (N_10378,N_5919,N_6531);
nand U10379 (N_10379,N_4790,N_7443);
or U10380 (N_10380,N_7578,N_6012);
nor U10381 (N_10381,N_7836,N_7960);
or U10382 (N_10382,N_5125,N_6749);
nor U10383 (N_10383,N_4819,N_7119);
nor U10384 (N_10384,N_5048,N_5726);
or U10385 (N_10385,N_5698,N_5187);
nand U10386 (N_10386,N_6889,N_5558);
nor U10387 (N_10387,N_7758,N_5170);
and U10388 (N_10388,N_7259,N_5243);
nor U10389 (N_10389,N_7680,N_7076);
and U10390 (N_10390,N_4032,N_6843);
and U10391 (N_10391,N_4226,N_4291);
or U10392 (N_10392,N_4587,N_4150);
or U10393 (N_10393,N_5986,N_6217);
nand U10394 (N_10394,N_4759,N_6305);
nor U10395 (N_10395,N_4927,N_5791);
nor U10396 (N_10396,N_7705,N_7607);
or U10397 (N_10397,N_5918,N_5368);
nor U10398 (N_10398,N_4094,N_7256);
or U10399 (N_10399,N_5008,N_6691);
nand U10400 (N_10400,N_7885,N_4619);
and U10401 (N_10401,N_7118,N_6005);
and U10402 (N_10402,N_4139,N_5409);
or U10403 (N_10403,N_7251,N_6688);
and U10404 (N_10404,N_4507,N_4509);
nand U10405 (N_10405,N_6289,N_7819);
or U10406 (N_10406,N_7374,N_6858);
and U10407 (N_10407,N_4251,N_6940);
nand U10408 (N_10408,N_7953,N_5455);
or U10409 (N_10409,N_4244,N_7335);
and U10410 (N_10410,N_7413,N_5588);
nor U10411 (N_10411,N_6837,N_5177);
or U10412 (N_10412,N_5883,N_5449);
nor U10413 (N_10413,N_7420,N_4628);
or U10414 (N_10414,N_4788,N_6879);
or U10415 (N_10415,N_5849,N_4760);
or U10416 (N_10416,N_7196,N_6232);
or U10417 (N_10417,N_5438,N_7294);
or U10418 (N_10418,N_7091,N_7020);
and U10419 (N_10419,N_7314,N_4957);
nand U10420 (N_10420,N_7085,N_4631);
nand U10421 (N_10421,N_4003,N_7330);
nor U10422 (N_10422,N_7853,N_4541);
nor U10423 (N_10423,N_4004,N_5885);
and U10424 (N_10424,N_5537,N_7646);
or U10425 (N_10425,N_6812,N_5073);
nand U10426 (N_10426,N_7402,N_5138);
nor U10427 (N_10427,N_7037,N_5052);
or U10428 (N_10428,N_5157,N_4149);
and U10429 (N_10429,N_5933,N_5014);
or U10430 (N_10430,N_6608,N_7928);
or U10431 (N_10431,N_6823,N_5045);
or U10432 (N_10432,N_4304,N_5998);
or U10433 (N_10433,N_4282,N_7698);
nor U10434 (N_10434,N_6724,N_4128);
xor U10435 (N_10435,N_7925,N_5268);
nand U10436 (N_10436,N_5533,N_6317);
and U10437 (N_10437,N_6926,N_7713);
or U10438 (N_10438,N_4828,N_5897);
nor U10439 (N_10439,N_7784,N_6511);
or U10440 (N_10440,N_6765,N_5656);
or U10441 (N_10441,N_7315,N_4586);
nand U10442 (N_10442,N_6510,N_7714);
nand U10443 (N_10443,N_7706,N_6936);
or U10444 (N_10444,N_4491,N_7290);
nor U10445 (N_10445,N_5173,N_6275);
nand U10446 (N_10446,N_7961,N_7067);
and U10447 (N_10447,N_7398,N_6777);
nor U10448 (N_10448,N_6582,N_6870);
nand U10449 (N_10449,N_7119,N_7953);
nor U10450 (N_10450,N_5272,N_4211);
nor U10451 (N_10451,N_4874,N_4388);
nor U10452 (N_10452,N_5877,N_5536);
xnor U10453 (N_10453,N_5697,N_4164);
or U10454 (N_10454,N_6997,N_4330);
or U10455 (N_10455,N_5323,N_5159);
nand U10456 (N_10456,N_6639,N_5805);
nand U10457 (N_10457,N_4282,N_6917);
or U10458 (N_10458,N_5579,N_5848);
nand U10459 (N_10459,N_4105,N_5670);
and U10460 (N_10460,N_6662,N_7492);
nand U10461 (N_10461,N_7933,N_6925);
and U10462 (N_10462,N_5084,N_4423);
and U10463 (N_10463,N_7022,N_6053);
or U10464 (N_10464,N_7607,N_7328);
nor U10465 (N_10465,N_5796,N_5359);
and U10466 (N_10466,N_5304,N_4600);
nand U10467 (N_10467,N_5296,N_7321);
or U10468 (N_10468,N_7878,N_4990);
nand U10469 (N_10469,N_7405,N_5459);
or U10470 (N_10470,N_5852,N_7053);
nor U10471 (N_10471,N_7283,N_6154);
and U10472 (N_10472,N_7925,N_5314);
nor U10473 (N_10473,N_6503,N_4514);
xor U10474 (N_10474,N_6623,N_4565);
nor U10475 (N_10475,N_7606,N_7275);
or U10476 (N_10476,N_6749,N_5457);
nor U10477 (N_10477,N_6028,N_6492);
xnor U10478 (N_10478,N_5858,N_6780);
or U10479 (N_10479,N_4733,N_7106);
or U10480 (N_10480,N_5228,N_4502);
nand U10481 (N_10481,N_4766,N_7302);
nand U10482 (N_10482,N_7853,N_4345);
and U10483 (N_10483,N_6704,N_7452);
and U10484 (N_10484,N_5858,N_7275);
and U10485 (N_10485,N_6609,N_4606);
nand U10486 (N_10486,N_6727,N_6825);
nor U10487 (N_10487,N_6765,N_4997);
nand U10488 (N_10488,N_5200,N_4523);
nor U10489 (N_10489,N_5437,N_7661);
or U10490 (N_10490,N_7103,N_5241);
nand U10491 (N_10491,N_7329,N_4592);
and U10492 (N_10492,N_7959,N_5446);
or U10493 (N_10493,N_7309,N_6804);
nand U10494 (N_10494,N_5247,N_5212);
nor U10495 (N_10495,N_4427,N_4862);
and U10496 (N_10496,N_4503,N_6695);
nand U10497 (N_10497,N_5567,N_4432);
xnor U10498 (N_10498,N_4251,N_5416);
nand U10499 (N_10499,N_6174,N_6859);
and U10500 (N_10500,N_4405,N_4770);
nor U10501 (N_10501,N_4090,N_5574);
nor U10502 (N_10502,N_5289,N_7042);
and U10503 (N_10503,N_7347,N_5577);
nor U10504 (N_10504,N_7542,N_6967);
and U10505 (N_10505,N_7647,N_6205);
and U10506 (N_10506,N_4534,N_7458);
xor U10507 (N_10507,N_6391,N_6840);
nand U10508 (N_10508,N_6153,N_4093);
or U10509 (N_10509,N_6804,N_6083);
and U10510 (N_10510,N_7662,N_6711);
and U10511 (N_10511,N_6467,N_7932);
or U10512 (N_10512,N_5573,N_6569);
nor U10513 (N_10513,N_6584,N_7310);
nand U10514 (N_10514,N_7135,N_7300);
nand U10515 (N_10515,N_5710,N_4584);
or U10516 (N_10516,N_5639,N_4986);
nand U10517 (N_10517,N_6311,N_5986);
or U10518 (N_10518,N_6245,N_5533);
nor U10519 (N_10519,N_5796,N_7896);
nand U10520 (N_10520,N_5888,N_5397);
and U10521 (N_10521,N_4066,N_6007);
and U10522 (N_10522,N_4303,N_4324);
nand U10523 (N_10523,N_6384,N_4272);
and U10524 (N_10524,N_7985,N_6489);
and U10525 (N_10525,N_7564,N_6587);
or U10526 (N_10526,N_5993,N_6135);
nand U10527 (N_10527,N_4089,N_6406);
nor U10528 (N_10528,N_4998,N_4861);
nand U10529 (N_10529,N_7703,N_6673);
or U10530 (N_10530,N_6225,N_5326);
or U10531 (N_10531,N_5859,N_6664);
nand U10532 (N_10532,N_6027,N_5309);
or U10533 (N_10533,N_6114,N_6765);
or U10534 (N_10534,N_5487,N_4519);
and U10535 (N_10535,N_7719,N_5875);
and U10536 (N_10536,N_6230,N_5174);
and U10537 (N_10537,N_6548,N_6809);
xnor U10538 (N_10538,N_7696,N_6539);
nor U10539 (N_10539,N_6777,N_4146);
nand U10540 (N_10540,N_4570,N_7439);
nor U10541 (N_10541,N_4366,N_6726);
nand U10542 (N_10542,N_5961,N_4177);
nand U10543 (N_10543,N_7553,N_5436);
nor U10544 (N_10544,N_6960,N_4559);
and U10545 (N_10545,N_5939,N_7769);
nand U10546 (N_10546,N_5878,N_4351);
nand U10547 (N_10547,N_6825,N_7599);
and U10548 (N_10548,N_4099,N_6009);
nor U10549 (N_10549,N_7029,N_5376);
or U10550 (N_10550,N_4879,N_6999);
or U10551 (N_10551,N_5191,N_6718);
nor U10552 (N_10552,N_5416,N_5381);
or U10553 (N_10553,N_4763,N_7747);
or U10554 (N_10554,N_4799,N_7224);
nor U10555 (N_10555,N_5985,N_7533);
or U10556 (N_10556,N_7831,N_4664);
or U10557 (N_10557,N_4731,N_6293);
or U10558 (N_10558,N_7882,N_6293);
or U10559 (N_10559,N_4113,N_5751);
or U10560 (N_10560,N_4132,N_5425);
nand U10561 (N_10561,N_4590,N_7354);
or U10562 (N_10562,N_5993,N_5305);
nor U10563 (N_10563,N_6366,N_6767);
nor U10564 (N_10564,N_4121,N_6534);
and U10565 (N_10565,N_5213,N_4510);
nor U10566 (N_10566,N_7816,N_5868);
nand U10567 (N_10567,N_7344,N_7661);
or U10568 (N_10568,N_5896,N_7973);
and U10569 (N_10569,N_6173,N_5890);
nor U10570 (N_10570,N_7714,N_4303);
nand U10571 (N_10571,N_5240,N_6170);
nor U10572 (N_10572,N_5230,N_5881);
and U10573 (N_10573,N_6377,N_5258);
and U10574 (N_10574,N_4057,N_6031);
or U10575 (N_10575,N_4720,N_6592);
nor U10576 (N_10576,N_5530,N_4851);
or U10577 (N_10577,N_7405,N_7748);
nor U10578 (N_10578,N_7376,N_7562);
nand U10579 (N_10579,N_5608,N_7581);
or U10580 (N_10580,N_5465,N_7753);
and U10581 (N_10581,N_5961,N_7849);
nor U10582 (N_10582,N_5129,N_4414);
or U10583 (N_10583,N_4987,N_7660);
nand U10584 (N_10584,N_5739,N_4086);
and U10585 (N_10585,N_6447,N_7948);
nand U10586 (N_10586,N_7258,N_6280);
nor U10587 (N_10587,N_4383,N_4133);
or U10588 (N_10588,N_4788,N_4216);
and U10589 (N_10589,N_7594,N_5052);
and U10590 (N_10590,N_5989,N_5082);
or U10591 (N_10591,N_7583,N_7257);
and U10592 (N_10592,N_5666,N_7729);
and U10593 (N_10593,N_6576,N_7817);
or U10594 (N_10594,N_4305,N_6248);
nor U10595 (N_10595,N_5455,N_6817);
nand U10596 (N_10596,N_5975,N_4930);
nand U10597 (N_10597,N_5897,N_4735);
and U10598 (N_10598,N_5567,N_5685);
or U10599 (N_10599,N_7840,N_4632);
nand U10600 (N_10600,N_5658,N_5703);
and U10601 (N_10601,N_4669,N_4269);
nor U10602 (N_10602,N_4478,N_6956);
or U10603 (N_10603,N_5734,N_4528);
or U10604 (N_10604,N_5599,N_4408);
or U10605 (N_10605,N_6719,N_6590);
nor U10606 (N_10606,N_4630,N_5449);
or U10607 (N_10607,N_4064,N_4882);
and U10608 (N_10608,N_4945,N_4322);
nand U10609 (N_10609,N_7399,N_7291);
nand U10610 (N_10610,N_7504,N_7885);
or U10611 (N_10611,N_5402,N_6548);
or U10612 (N_10612,N_7328,N_4189);
and U10613 (N_10613,N_7296,N_6658);
or U10614 (N_10614,N_5633,N_4333);
and U10615 (N_10615,N_6269,N_5569);
nand U10616 (N_10616,N_4586,N_7246);
nor U10617 (N_10617,N_4295,N_5174);
or U10618 (N_10618,N_6649,N_4730);
nor U10619 (N_10619,N_7044,N_4324);
or U10620 (N_10620,N_7390,N_7184);
nand U10621 (N_10621,N_7146,N_6933);
nor U10622 (N_10622,N_5613,N_7215);
and U10623 (N_10623,N_5760,N_7120);
nor U10624 (N_10624,N_4466,N_7907);
or U10625 (N_10625,N_5800,N_4202);
nor U10626 (N_10626,N_5673,N_5697);
and U10627 (N_10627,N_4063,N_5426);
nand U10628 (N_10628,N_7448,N_7844);
and U10629 (N_10629,N_7628,N_4022);
nand U10630 (N_10630,N_6110,N_7430);
and U10631 (N_10631,N_6204,N_7711);
nor U10632 (N_10632,N_6428,N_7620);
nor U10633 (N_10633,N_7499,N_5391);
nor U10634 (N_10634,N_6976,N_4823);
nand U10635 (N_10635,N_7198,N_7337);
and U10636 (N_10636,N_4120,N_6563);
or U10637 (N_10637,N_7996,N_4735);
or U10638 (N_10638,N_4716,N_6467);
nor U10639 (N_10639,N_7503,N_5008);
nor U10640 (N_10640,N_7120,N_5514);
or U10641 (N_10641,N_7246,N_4071);
nand U10642 (N_10642,N_7190,N_5539);
nand U10643 (N_10643,N_4275,N_5647);
nand U10644 (N_10644,N_4375,N_6201);
nand U10645 (N_10645,N_7384,N_4813);
and U10646 (N_10646,N_6778,N_6999);
or U10647 (N_10647,N_4168,N_5571);
or U10648 (N_10648,N_6501,N_6487);
nand U10649 (N_10649,N_6118,N_5035);
nor U10650 (N_10650,N_4802,N_5965);
and U10651 (N_10651,N_6050,N_4685);
and U10652 (N_10652,N_5750,N_7965);
nor U10653 (N_10653,N_7543,N_6338);
nand U10654 (N_10654,N_6870,N_4739);
nand U10655 (N_10655,N_7619,N_5508);
or U10656 (N_10656,N_4018,N_4957);
or U10657 (N_10657,N_4847,N_6535);
or U10658 (N_10658,N_4477,N_6315);
nor U10659 (N_10659,N_5935,N_4840);
nand U10660 (N_10660,N_7274,N_5728);
and U10661 (N_10661,N_5123,N_7788);
nand U10662 (N_10662,N_5767,N_5343);
nor U10663 (N_10663,N_5301,N_7457);
nor U10664 (N_10664,N_7049,N_5964);
nand U10665 (N_10665,N_5801,N_6107);
or U10666 (N_10666,N_6932,N_6346);
nor U10667 (N_10667,N_7967,N_6979);
or U10668 (N_10668,N_7819,N_7709);
and U10669 (N_10669,N_7459,N_5471);
and U10670 (N_10670,N_5494,N_6362);
nor U10671 (N_10671,N_6999,N_6220);
or U10672 (N_10672,N_6004,N_4403);
or U10673 (N_10673,N_6115,N_4255);
nor U10674 (N_10674,N_4470,N_6330);
nand U10675 (N_10675,N_6697,N_4811);
and U10676 (N_10676,N_5593,N_4812);
or U10677 (N_10677,N_4026,N_4776);
or U10678 (N_10678,N_6384,N_7081);
and U10679 (N_10679,N_4129,N_5488);
and U10680 (N_10680,N_4601,N_5938);
and U10681 (N_10681,N_5589,N_4240);
nor U10682 (N_10682,N_7150,N_5343);
or U10683 (N_10683,N_4743,N_4010);
and U10684 (N_10684,N_7175,N_4278);
and U10685 (N_10685,N_5934,N_5657);
nand U10686 (N_10686,N_7638,N_5244);
nand U10687 (N_10687,N_5477,N_4313);
nand U10688 (N_10688,N_6461,N_4993);
or U10689 (N_10689,N_5354,N_4592);
and U10690 (N_10690,N_5606,N_6319);
nor U10691 (N_10691,N_6115,N_5107);
and U10692 (N_10692,N_4093,N_6423);
and U10693 (N_10693,N_4460,N_4768);
nor U10694 (N_10694,N_5788,N_7580);
xnor U10695 (N_10695,N_7095,N_5691);
nor U10696 (N_10696,N_4549,N_4866);
nor U10697 (N_10697,N_6381,N_6122);
and U10698 (N_10698,N_6238,N_7153);
nand U10699 (N_10699,N_5406,N_6988);
and U10700 (N_10700,N_7199,N_5515);
nand U10701 (N_10701,N_5193,N_4108);
nand U10702 (N_10702,N_7996,N_5505);
or U10703 (N_10703,N_7717,N_6122);
nor U10704 (N_10704,N_6667,N_6233);
nor U10705 (N_10705,N_7738,N_5900);
or U10706 (N_10706,N_7190,N_6154);
and U10707 (N_10707,N_5118,N_5729);
or U10708 (N_10708,N_5724,N_6989);
or U10709 (N_10709,N_6839,N_6591);
or U10710 (N_10710,N_6883,N_6022);
nand U10711 (N_10711,N_7954,N_6072);
and U10712 (N_10712,N_7981,N_7623);
or U10713 (N_10713,N_6521,N_6569);
or U10714 (N_10714,N_4658,N_5681);
and U10715 (N_10715,N_5001,N_7030);
or U10716 (N_10716,N_4624,N_5853);
or U10717 (N_10717,N_7754,N_4077);
or U10718 (N_10718,N_4663,N_4707);
nand U10719 (N_10719,N_6949,N_7989);
or U10720 (N_10720,N_6097,N_7408);
or U10721 (N_10721,N_7338,N_5475);
or U10722 (N_10722,N_7535,N_4356);
or U10723 (N_10723,N_4900,N_7370);
nor U10724 (N_10724,N_5916,N_7046);
nand U10725 (N_10725,N_5140,N_7513);
or U10726 (N_10726,N_7052,N_7159);
xor U10727 (N_10727,N_4237,N_7024);
nand U10728 (N_10728,N_7304,N_4074);
and U10729 (N_10729,N_5359,N_6218);
or U10730 (N_10730,N_7302,N_4514);
nor U10731 (N_10731,N_4444,N_4668);
and U10732 (N_10732,N_6944,N_6211);
nor U10733 (N_10733,N_6831,N_5585);
nand U10734 (N_10734,N_7294,N_5138);
and U10735 (N_10735,N_6799,N_6282);
and U10736 (N_10736,N_5735,N_5796);
nor U10737 (N_10737,N_5351,N_7588);
or U10738 (N_10738,N_7495,N_5257);
nand U10739 (N_10739,N_4405,N_5688);
nand U10740 (N_10740,N_4467,N_6945);
and U10741 (N_10741,N_7255,N_7203);
and U10742 (N_10742,N_7475,N_7596);
or U10743 (N_10743,N_5790,N_4887);
nor U10744 (N_10744,N_5679,N_6191);
and U10745 (N_10745,N_5036,N_7489);
nand U10746 (N_10746,N_6485,N_4471);
nor U10747 (N_10747,N_4263,N_5785);
or U10748 (N_10748,N_4197,N_5804);
or U10749 (N_10749,N_4389,N_4762);
nor U10750 (N_10750,N_6131,N_7258);
and U10751 (N_10751,N_6285,N_7435);
nand U10752 (N_10752,N_7469,N_7957);
nor U10753 (N_10753,N_5513,N_6781);
or U10754 (N_10754,N_5988,N_7419);
or U10755 (N_10755,N_6861,N_5527);
or U10756 (N_10756,N_6233,N_4728);
nand U10757 (N_10757,N_4478,N_4090);
and U10758 (N_10758,N_5551,N_6834);
or U10759 (N_10759,N_7906,N_7836);
nand U10760 (N_10760,N_5663,N_5148);
and U10761 (N_10761,N_5222,N_4133);
and U10762 (N_10762,N_4548,N_4328);
and U10763 (N_10763,N_4175,N_7808);
nor U10764 (N_10764,N_4882,N_4420);
nand U10765 (N_10765,N_5848,N_6348);
or U10766 (N_10766,N_7722,N_5296);
nand U10767 (N_10767,N_6882,N_4132);
nor U10768 (N_10768,N_7846,N_4559);
or U10769 (N_10769,N_6331,N_6225);
and U10770 (N_10770,N_7888,N_5298);
nor U10771 (N_10771,N_5302,N_7849);
nor U10772 (N_10772,N_5203,N_6180);
or U10773 (N_10773,N_5452,N_6542);
or U10774 (N_10774,N_5414,N_7834);
and U10775 (N_10775,N_7005,N_5572);
nand U10776 (N_10776,N_4503,N_4440);
nor U10777 (N_10777,N_7618,N_6072);
xor U10778 (N_10778,N_4305,N_5913);
nand U10779 (N_10779,N_7898,N_5115);
or U10780 (N_10780,N_4396,N_6234);
or U10781 (N_10781,N_4579,N_4555);
and U10782 (N_10782,N_7424,N_6374);
nand U10783 (N_10783,N_6242,N_6792);
or U10784 (N_10784,N_7138,N_5308);
or U10785 (N_10785,N_4701,N_5677);
nand U10786 (N_10786,N_7546,N_4637);
and U10787 (N_10787,N_6734,N_4155);
or U10788 (N_10788,N_6958,N_7550);
and U10789 (N_10789,N_5669,N_7196);
and U10790 (N_10790,N_4195,N_5589);
nor U10791 (N_10791,N_6730,N_4400);
nand U10792 (N_10792,N_6332,N_4108);
and U10793 (N_10793,N_7636,N_5991);
or U10794 (N_10794,N_4032,N_4502);
nor U10795 (N_10795,N_5548,N_7669);
and U10796 (N_10796,N_7386,N_5953);
and U10797 (N_10797,N_7158,N_6999);
nand U10798 (N_10798,N_6584,N_4793);
nand U10799 (N_10799,N_4974,N_5195);
nor U10800 (N_10800,N_6028,N_4578);
nand U10801 (N_10801,N_5642,N_5420);
or U10802 (N_10802,N_7300,N_4893);
nand U10803 (N_10803,N_4837,N_6057);
nor U10804 (N_10804,N_6536,N_5835);
or U10805 (N_10805,N_6147,N_5347);
nand U10806 (N_10806,N_6128,N_5502);
or U10807 (N_10807,N_7426,N_6110);
and U10808 (N_10808,N_5972,N_6499);
and U10809 (N_10809,N_5013,N_7487);
or U10810 (N_10810,N_6215,N_4300);
and U10811 (N_10811,N_5312,N_6874);
nor U10812 (N_10812,N_4256,N_4518);
or U10813 (N_10813,N_6590,N_7916);
or U10814 (N_10814,N_5012,N_7269);
nor U10815 (N_10815,N_4750,N_5830);
nand U10816 (N_10816,N_7051,N_6665);
and U10817 (N_10817,N_4635,N_7051);
nand U10818 (N_10818,N_7919,N_6494);
nand U10819 (N_10819,N_7699,N_4378);
or U10820 (N_10820,N_5759,N_7752);
or U10821 (N_10821,N_5382,N_6068);
or U10822 (N_10822,N_7071,N_7759);
or U10823 (N_10823,N_4150,N_7480);
nand U10824 (N_10824,N_5619,N_4032);
nor U10825 (N_10825,N_6589,N_7842);
nor U10826 (N_10826,N_6112,N_6038);
nand U10827 (N_10827,N_4903,N_4127);
nor U10828 (N_10828,N_6158,N_6528);
and U10829 (N_10829,N_5062,N_4519);
nor U10830 (N_10830,N_5926,N_7421);
nor U10831 (N_10831,N_4602,N_6744);
or U10832 (N_10832,N_5666,N_6739);
or U10833 (N_10833,N_5316,N_7267);
and U10834 (N_10834,N_4110,N_6021);
or U10835 (N_10835,N_5692,N_5635);
and U10836 (N_10836,N_7451,N_5093);
nor U10837 (N_10837,N_7136,N_5269);
or U10838 (N_10838,N_7414,N_7354);
nor U10839 (N_10839,N_5646,N_7842);
nand U10840 (N_10840,N_4711,N_4118);
or U10841 (N_10841,N_7582,N_4313);
nor U10842 (N_10842,N_7181,N_6648);
or U10843 (N_10843,N_5813,N_6101);
nand U10844 (N_10844,N_6169,N_5892);
nand U10845 (N_10845,N_4747,N_7210);
nor U10846 (N_10846,N_7742,N_5339);
nor U10847 (N_10847,N_4277,N_5290);
or U10848 (N_10848,N_6886,N_7304);
and U10849 (N_10849,N_6980,N_4120);
and U10850 (N_10850,N_7185,N_4324);
or U10851 (N_10851,N_7820,N_4764);
or U10852 (N_10852,N_6257,N_7204);
or U10853 (N_10853,N_4488,N_6644);
and U10854 (N_10854,N_6460,N_6667);
nand U10855 (N_10855,N_6790,N_7950);
xor U10856 (N_10856,N_4209,N_5122);
or U10857 (N_10857,N_4258,N_7273);
nand U10858 (N_10858,N_5481,N_7923);
xnor U10859 (N_10859,N_6639,N_4806);
or U10860 (N_10860,N_6567,N_6868);
or U10861 (N_10861,N_4696,N_4464);
and U10862 (N_10862,N_6328,N_4773);
nor U10863 (N_10863,N_5566,N_7341);
or U10864 (N_10864,N_5049,N_6599);
nand U10865 (N_10865,N_5795,N_6497);
and U10866 (N_10866,N_6517,N_7119);
nor U10867 (N_10867,N_5341,N_5603);
nor U10868 (N_10868,N_4174,N_6329);
and U10869 (N_10869,N_6221,N_6643);
and U10870 (N_10870,N_5390,N_7575);
or U10871 (N_10871,N_7248,N_7877);
xor U10872 (N_10872,N_5286,N_6450);
or U10873 (N_10873,N_5495,N_4861);
and U10874 (N_10874,N_5363,N_6482);
nor U10875 (N_10875,N_7349,N_6688);
or U10876 (N_10876,N_4112,N_6919);
nand U10877 (N_10877,N_6447,N_6595);
and U10878 (N_10878,N_4921,N_6301);
nor U10879 (N_10879,N_7419,N_5843);
nor U10880 (N_10880,N_5453,N_6218);
nand U10881 (N_10881,N_7311,N_6735);
nor U10882 (N_10882,N_6714,N_7896);
and U10883 (N_10883,N_6452,N_5766);
and U10884 (N_10884,N_7682,N_4175);
and U10885 (N_10885,N_6618,N_5579);
and U10886 (N_10886,N_4778,N_6116);
or U10887 (N_10887,N_6818,N_6115);
nor U10888 (N_10888,N_5040,N_7994);
nand U10889 (N_10889,N_4353,N_6180);
or U10890 (N_10890,N_6562,N_7579);
nor U10891 (N_10891,N_6114,N_5697);
and U10892 (N_10892,N_7354,N_6107);
nand U10893 (N_10893,N_5438,N_5134);
nand U10894 (N_10894,N_5644,N_7039);
nor U10895 (N_10895,N_6870,N_7820);
nor U10896 (N_10896,N_7018,N_7009);
nor U10897 (N_10897,N_4567,N_6787);
nand U10898 (N_10898,N_5075,N_5288);
nor U10899 (N_10899,N_6563,N_7966);
nand U10900 (N_10900,N_4606,N_6025);
xor U10901 (N_10901,N_4195,N_5736);
or U10902 (N_10902,N_7629,N_6261);
nand U10903 (N_10903,N_7848,N_6743);
and U10904 (N_10904,N_7214,N_5835);
nand U10905 (N_10905,N_6666,N_4100);
nand U10906 (N_10906,N_6662,N_7776);
nand U10907 (N_10907,N_5215,N_6374);
nor U10908 (N_10908,N_5990,N_4139);
and U10909 (N_10909,N_5782,N_4524);
xnor U10910 (N_10910,N_7009,N_4903);
nand U10911 (N_10911,N_4837,N_4298);
nand U10912 (N_10912,N_7548,N_7832);
nor U10913 (N_10913,N_7563,N_7687);
xor U10914 (N_10914,N_4048,N_6385);
nor U10915 (N_10915,N_5943,N_4043);
nand U10916 (N_10916,N_5535,N_5489);
and U10917 (N_10917,N_6335,N_4171);
nand U10918 (N_10918,N_4821,N_7229);
nand U10919 (N_10919,N_5886,N_4013);
nor U10920 (N_10920,N_6791,N_4641);
and U10921 (N_10921,N_6403,N_5287);
nor U10922 (N_10922,N_5854,N_5959);
xnor U10923 (N_10923,N_4061,N_5315);
nand U10924 (N_10924,N_7902,N_4919);
or U10925 (N_10925,N_7797,N_7035);
nand U10926 (N_10926,N_4487,N_4601);
xor U10927 (N_10927,N_4152,N_6036);
and U10928 (N_10928,N_4405,N_4745);
nand U10929 (N_10929,N_6161,N_6964);
or U10930 (N_10930,N_7670,N_5589);
xor U10931 (N_10931,N_6717,N_4897);
nor U10932 (N_10932,N_4641,N_6786);
nor U10933 (N_10933,N_5054,N_6966);
and U10934 (N_10934,N_4365,N_6567);
or U10935 (N_10935,N_6742,N_6563);
or U10936 (N_10936,N_4216,N_4479);
nand U10937 (N_10937,N_5621,N_4727);
xnor U10938 (N_10938,N_6023,N_6866);
or U10939 (N_10939,N_6491,N_4046);
or U10940 (N_10940,N_7983,N_6734);
nand U10941 (N_10941,N_5276,N_5015);
nor U10942 (N_10942,N_6784,N_6983);
or U10943 (N_10943,N_5815,N_6011);
and U10944 (N_10944,N_5327,N_7905);
xor U10945 (N_10945,N_4230,N_7186);
nor U10946 (N_10946,N_5462,N_6769);
or U10947 (N_10947,N_5306,N_5018);
or U10948 (N_10948,N_5133,N_6848);
or U10949 (N_10949,N_5094,N_5482);
and U10950 (N_10950,N_5401,N_5646);
or U10951 (N_10951,N_5698,N_4294);
or U10952 (N_10952,N_7263,N_5380);
or U10953 (N_10953,N_7177,N_6643);
nand U10954 (N_10954,N_5391,N_5723);
nor U10955 (N_10955,N_6879,N_6000);
or U10956 (N_10956,N_7337,N_4473);
nor U10957 (N_10957,N_5928,N_5062);
and U10958 (N_10958,N_5584,N_5527);
nand U10959 (N_10959,N_6937,N_7463);
or U10960 (N_10960,N_6074,N_6964);
nand U10961 (N_10961,N_6637,N_6589);
or U10962 (N_10962,N_5779,N_4479);
and U10963 (N_10963,N_7919,N_5550);
or U10964 (N_10964,N_7436,N_5166);
nand U10965 (N_10965,N_5544,N_6954);
or U10966 (N_10966,N_4954,N_4961);
or U10967 (N_10967,N_6875,N_4099);
nor U10968 (N_10968,N_4158,N_5523);
nor U10969 (N_10969,N_4831,N_6139);
or U10970 (N_10970,N_7100,N_4419);
or U10971 (N_10971,N_6020,N_7115);
or U10972 (N_10972,N_7953,N_6368);
nor U10973 (N_10973,N_6623,N_6254);
nor U10974 (N_10974,N_6240,N_4051);
nor U10975 (N_10975,N_6652,N_4360);
nand U10976 (N_10976,N_5104,N_4634);
nand U10977 (N_10977,N_4887,N_5759);
or U10978 (N_10978,N_7420,N_5625);
and U10979 (N_10979,N_6228,N_7834);
nor U10980 (N_10980,N_4555,N_5943);
nor U10981 (N_10981,N_6902,N_6279);
or U10982 (N_10982,N_7947,N_7196);
nand U10983 (N_10983,N_5147,N_7933);
nand U10984 (N_10984,N_6532,N_7398);
and U10985 (N_10985,N_4411,N_5619);
nor U10986 (N_10986,N_6240,N_7017);
nor U10987 (N_10987,N_6567,N_5685);
and U10988 (N_10988,N_7221,N_4285);
nor U10989 (N_10989,N_5299,N_6284);
and U10990 (N_10990,N_6430,N_5545);
or U10991 (N_10991,N_7046,N_4509);
nor U10992 (N_10992,N_4197,N_5849);
or U10993 (N_10993,N_6183,N_6591);
and U10994 (N_10994,N_5002,N_7233);
and U10995 (N_10995,N_6794,N_4434);
or U10996 (N_10996,N_4843,N_7275);
nor U10997 (N_10997,N_4928,N_4839);
and U10998 (N_10998,N_4612,N_4924);
nand U10999 (N_10999,N_5768,N_6867);
and U11000 (N_11000,N_7354,N_6441);
and U11001 (N_11001,N_6594,N_4205);
or U11002 (N_11002,N_7649,N_7355);
or U11003 (N_11003,N_5075,N_7364);
or U11004 (N_11004,N_5859,N_4421);
nand U11005 (N_11005,N_5883,N_5867);
and U11006 (N_11006,N_7797,N_4156);
nand U11007 (N_11007,N_4253,N_5789);
nor U11008 (N_11008,N_6243,N_7383);
nand U11009 (N_11009,N_7476,N_7527);
nor U11010 (N_11010,N_6339,N_6007);
and U11011 (N_11011,N_5652,N_4282);
and U11012 (N_11012,N_6680,N_5626);
and U11013 (N_11013,N_6581,N_7022);
or U11014 (N_11014,N_7748,N_6349);
and U11015 (N_11015,N_4697,N_4066);
nor U11016 (N_11016,N_7424,N_4367);
or U11017 (N_11017,N_5024,N_4567);
nand U11018 (N_11018,N_5242,N_5269);
or U11019 (N_11019,N_5650,N_6607);
and U11020 (N_11020,N_6549,N_7383);
and U11021 (N_11021,N_7450,N_4547);
and U11022 (N_11022,N_5974,N_6851);
nor U11023 (N_11023,N_5997,N_4206);
nand U11024 (N_11024,N_6277,N_6198);
or U11025 (N_11025,N_6168,N_6187);
nand U11026 (N_11026,N_4772,N_5694);
and U11027 (N_11027,N_7029,N_5973);
nor U11028 (N_11028,N_4371,N_4099);
or U11029 (N_11029,N_6757,N_5770);
nor U11030 (N_11030,N_4128,N_6815);
nand U11031 (N_11031,N_6064,N_7803);
or U11032 (N_11032,N_4457,N_4176);
nand U11033 (N_11033,N_5116,N_6150);
and U11034 (N_11034,N_4628,N_4547);
nor U11035 (N_11035,N_5668,N_7532);
or U11036 (N_11036,N_5086,N_6938);
nand U11037 (N_11037,N_7469,N_4728);
nor U11038 (N_11038,N_7100,N_4535);
and U11039 (N_11039,N_4726,N_5247);
nor U11040 (N_11040,N_4820,N_5249);
and U11041 (N_11041,N_5589,N_6500);
nor U11042 (N_11042,N_7324,N_4741);
or U11043 (N_11043,N_7825,N_7016);
and U11044 (N_11044,N_4227,N_6558);
nor U11045 (N_11045,N_6637,N_4262);
and U11046 (N_11046,N_6981,N_6245);
nand U11047 (N_11047,N_4962,N_7142);
and U11048 (N_11048,N_6572,N_6634);
and U11049 (N_11049,N_4137,N_4446);
and U11050 (N_11050,N_5653,N_7985);
nor U11051 (N_11051,N_6432,N_4401);
and U11052 (N_11052,N_6818,N_6582);
and U11053 (N_11053,N_4462,N_7631);
nand U11054 (N_11054,N_5444,N_7789);
nand U11055 (N_11055,N_4788,N_6607);
or U11056 (N_11056,N_5722,N_6164);
nand U11057 (N_11057,N_6386,N_5170);
and U11058 (N_11058,N_7660,N_4998);
nor U11059 (N_11059,N_4728,N_5883);
or U11060 (N_11060,N_6181,N_7479);
and U11061 (N_11061,N_7773,N_6460);
nor U11062 (N_11062,N_6942,N_5984);
and U11063 (N_11063,N_7381,N_7637);
and U11064 (N_11064,N_6002,N_7519);
nor U11065 (N_11065,N_6494,N_7661);
or U11066 (N_11066,N_6222,N_7519);
and U11067 (N_11067,N_4488,N_5286);
nor U11068 (N_11068,N_4651,N_6950);
and U11069 (N_11069,N_6970,N_5331);
and U11070 (N_11070,N_7155,N_4520);
nand U11071 (N_11071,N_4214,N_4622);
and U11072 (N_11072,N_5411,N_6885);
nand U11073 (N_11073,N_7491,N_4343);
or U11074 (N_11074,N_6328,N_6025);
or U11075 (N_11075,N_7053,N_7428);
nor U11076 (N_11076,N_4443,N_6511);
nor U11077 (N_11077,N_7218,N_4099);
nand U11078 (N_11078,N_7157,N_6108);
and U11079 (N_11079,N_5944,N_6546);
nand U11080 (N_11080,N_6422,N_4502);
nor U11081 (N_11081,N_6752,N_6329);
or U11082 (N_11082,N_6979,N_4975);
nor U11083 (N_11083,N_7405,N_4869);
nand U11084 (N_11084,N_4434,N_4044);
nor U11085 (N_11085,N_7531,N_7066);
nor U11086 (N_11086,N_6554,N_5454);
nor U11087 (N_11087,N_7154,N_7400);
or U11088 (N_11088,N_6841,N_5896);
nor U11089 (N_11089,N_6637,N_6330);
nor U11090 (N_11090,N_4936,N_4110);
or U11091 (N_11091,N_5472,N_7893);
nor U11092 (N_11092,N_5305,N_6608);
or U11093 (N_11093,N_6244,N_7643);
and U11094 (N_11094,N_6006,N_6253);
or U11095 (N_11095,N_4478,N_7220);
nand U11096 (N_11096,N_5362,N_5558);
nand U11097 (N_11097,N_4184,N_7228);
nor U11098 (N_11098,N_7262,N_6131);
nor U11099 (N_11099,N_7975,N_7974);
and U11100 (N_11100,N_4983,N_4024);
and U11101 (N_11101,N_5357,N_7369);
nor U11102 (N_11102,N_5015,N_4925);
and U11103 (N_11103,N_5079,N_4860);
or U11104 (N_11104,N_6842,N_6313);
nand U11105 (N_11105,N_5212,N_7169);
or U11106 (N_11106,N_5580,N_7411);
and U11107 (N_11107,N_6719,N_5247);
and U11108 (N_11108,N_6674,N_7685);
or U11109 (N_11109,N_4549,N_6115);
nor U11110 (N_11110,N_6176,N_6687);
and U11111 (N_11111,N_5856,N_4590);
or U11112 (N_11112,N_5632,N_6200);
and U11113 (N_11113,N_7970,N_5519);
nand U11114 (N_11114,N_4482,N_7243);
and U11115 (N_11115,N_7751,N_7259);
nand U11116 (N_11116,N_5173,N_7821);
nor U11117 (N_11117,N_7486,N_5378);
and U11118 (N_11118,N_7936,N_6915);
or U11119 (N_11119,N_4673,N_5070);
nor U11120 (N_11120,N_7261,N_4145);
nand U11121 (N_11121,N_7833,N_4476);
nor U11122 (N_11122,N_7367,N_7043);
nor U11123 (N_11123,N_5191,N_7390);
nor U11124 (N_11124,N_7775,N_5260);
and U11125 (N_11125,N_5935,N_5145);
or U11126 (N_11126,N_7463,N_4328);
and U11127 (N_11127,N_5445,N_5987);
and U11128 (N_11128,N_6615,N_5429);
and U11129 (N_11129,N_7349,N_7301);
and U11130 (N_11130,N_5962,N_5763);
nor U11131 (N_11131,N_5828,N_4992);
nand U11132 (N_11132,N_7328,N_4151);
or U11133 (N_11133,N_6226,N_5300);
nor U11134 (N_11134,N_4130,N_6982);
or U11135 (N_11135,N_5346,N_7245);
or U11136 (N_11136,N_7021,N_5896);
nand U11137 (N_11137,N_6985,N_4178);
and U11138 (N_11138,N_5115,N_6162);
or U11139 (N_11139,N_7662,N_6002);
and U11140 (N_11140,N_4512,N_6987);
and U11141 (N_11141,N_6005,N_4335);
nand U11142 (N_11142,N_5683,N_7210);
or U11143 (N_11143,N_6935,N_7818);
nor U11144 (N_11144,N_6445,N_4750);
nand U11145 (N_11145,N_4535,N_6138);
nand U11146 (N_11146,N_7220,N_7540);
or U11147 (N_11147,N_7773,N_7436);
nand U11148 (N_11148,N_4437,N_6301);
nor U11149 (N_11149,N_5899,N_6346);
nand U11150 (N_11150,N_5497,N_5799);
and U11151 (N_11151,N_6291,N_6146);
and U11152 (N_11152,N_5153,N_7551);
and U11153 (N_11153,N_4521,N_5605);
nor U11154 (N_11154,N_6848,N_5246);
nand U11155 (N_11155,N_7360,N_7009);
nor U11156 (N_11156,N_4774,N_4036);
nor U11157 (N_11157,N_6497,N_6343);
nor U11158 (N_11158,N_7542,N_7149);
and U11159 (N_11159,N_7840,N_6575);
nor U11160 (N_11160,N_5588,N_7226);
and U11161 (N_11161,N_7680,N_4186);
nand U11162 (N_11162,N_4955,N_7831);
nor U11163 (N_11163,N_6468,N_5750);
nor U11164 (N_11164,N_6860,N_5812);
and U11165 (N_11165,N_7116,N_6629);
and U11166 (N_11166,N_5719,N_7215);
nand U11167 (N_11167,N_5621,N_4188);
nor U11168 (N_11168,N_6888,N_5466);
nand U11169 (N_11169,N_6266,N_4051);
nor U11170 (N_11170,N_4177,N_4264);
nor U11171 (N_11171,N_7165,N_7404);
nor U11172 (N_11172,N_5608,N_4611);
nand U11173 (N_11173,N_6543,N_4953);
nand U11174 (N_11174,N_5540,N_4086);
nor U11175 (N_11175,N_7740,N_6308);
or U11176 (N_11176,N_4568,N_4508);
and U11177 (N_11177,N_5648,N_7012);
xnor U11178 (N_11178,N_4195,N_5652);
nor U11179 (N_11179,N_6515,N_4029);
nor U11180 (N_11180,N_6756,N_5322);
nor U11181 (N_11181,N_7468,N_6232);
nor U11182 (N_11182,N_5542,N_4851);
nor U11183 (N_11183,N_6290,N_6318);
and U11184 (N_11184,N_7040,N_5903);
or U11185 (N_11185,N_6418,N_4839);
or U11186 (N_11186,N_7271,N_4502);
and U11187 (N_11187,N_4816,N_6905);
nor U11188 (N_11188,N_7563,N_4866);
or U11189 (N_11189,N_6038,N_4601);
and U11190 (N_11190,N_4519,N_4701);
or U11191 (N_11191,N_7710,N_6747);
or U11192 (N_11192,N_4730,N_6109);
nand U11193 (N_11193,N_6092,N_5923);
or U11194 (N_11194,N_6122,N_5133);
and U11195 (N_11195,N_6112,N_5670);
nor U11196 (N_11196,N_5234,N_5757);
nor U11197 (N_11197,N_7417,N_6962);
xnor U11198 (N_11198,N_4959,N_4021);
nand U11199 (N_11199,N_7408,N_7321);
or U11200 (N_11200,N_4614,N_4742);
nor U11201 (N_11201,N_7863,N_6417);
and U11202 (N_11202,N_5842,N_5028);
nor U11203 (N_11203,N_6273,N_4191);
and U11204 (N_11204,N_5833,N_5136);
or U11205 (N_11205,N_5078,N_7241);
or U11206 (N_11206,N_7376,N_6234);
or U11207 (N_11207,N_5452,N_4033);
or U11208 (N_11208,N_7029,N_7692);
nor U11209 (N_11209,N_7564,N_4895);
nor U11210 (N_11210,N_7678,N_6739);
xnor U11211 (N_11211,N_6942,N_6322);
or U11212 (N_11212,N_6185,N_4711);
and U11213 (N_11213,N_5153,N_4120);
xnor U11214 (N_11214,N_5087,N_6224);
or U11215 (N_11215,N_7869,N_4821);
nand U11216 (N_11216,N_4518,N_4760);
or U11217 (N_11217,N_7325,N_5529);
and U11218 (N_11218,N_6110,N_5501);
or U11219 (N_11219,N_4930,N_4133);
and U11220 (N_11220,N_7879,N_7782);
and U11221 (N_11221,N_6106,N_7704);
nor U11222 (N_11222,N_5399,N_5583);
nand U11223 (N_11223,N_7624,N_6440);
nor U11224 (N_11224,N_6525,N_4533);
nor U11225 (N_11225,N_4568,N_5499);
nor U11226 (N_11226,N_6763,N_7435);
nand U11227 (N_11227,N_4204,N_7155);
nor U11228 (N_11228,N_5413,N_4959);
nand U11229 (N_11229,N_4867,N_7916);
nand U11230 (N_11230,N_6718,N_7317);
nand U11231 (N_11231,N_6257,N_4596);
and U11232 (N_11232,N_4012,N_6133);
and U11233 (N_11233,N_6004,N_5958);
and U11234 (N_11234,N_5701,N_5419);
and U11235 (N_11235,N_5361,N_4379);
and U11236 (N_11236,N_5634,N_4085);
nor U11237 (N_11237,N_7248,N_4351);
nand U11238 (N_11238,N_6482,N_4313);
nor U11239 (N_11239,N_5403,N_7304);
and U11240 (N_11240,N_7909,N_7181);
or U11241 (N_11241,N_5114,N_4986);
or U11242 (N_11242,N_4985,N_7626);
nor U11243 (N_11243,N_4225,N_4731);
and U11244 (N_11244,N_6067,N_6494);
nand U11245 (N_11245,N_6332,N_4914);
nor U11246 (N_11246,N_7143,N_6053);
nor U11247 (N_11247,N_6743,N_6226);
nor U11248 (N_11248,N_4108,N_5018);
and U11249 (N_11249,N_7699,N_6631);
nor U11250 (N_11250,N_5526,N_5426);
and U11251 (N_11251,N_6797,N_5284);
or U11252 (N_11252,N_5595,N_6516);
or U11253 (N_11253,N_7379,N_5747);
nand U11254 (N_11254,N_7615,N_7542);
nor U11255 (N_11255,N_7326,N_7806);
or U11256 (N_11256,N_5106,N_6440);
nor U11257 (N_11257,N_7609,N_6861);
nand U11258 (N_11258,N_5999,N_5623);
and U11259 (N_11259,N_5660,N_5722);
nand U11260 (N_11260,N_5575,N_5651);
nand U11261 (N_11261,N_7646,N_4355);
nand U11262 (N_11262,N_6601,N_4286);
and U11263 (N_11263,N_7939,N_4765);
nor U11264 (N_11264,N_5582,N_4826);
nor U11265 (N_11265,N_5867,N_6721);
and U11266 (N_11266,N_7566,N_5270);
or U11267 (N_11267,N_4974,N_4522);
xnor U11268 (N_11268,N_5387,N_7722);
and U11269 (N_11269,N_7919,N_5920);
nand U11270 (N_11270,N_7820,N_6689);
and U11271 (N_11271,N_4907,N_5858);
nand U11272 (N_11272,N_7770,N_5453);
or U11273 (N_11273,N_7524,N_5096);
nor U11274 (N_11274,N_6992,N_5156);
or U11275 (N_11275,N_7908,N_7202);
or U11276 (N_11276,N_6392,N_5550);
or U11277 (N_11277,N_4447,N_5132);
and U11278 (N_11278,N_4340,N_4845);
nor U11279 (N_11279,N_4214,N_4308);
or U11280 (N_11280,N_4943,N_5334);
or U11281 (N_11281,N_7014,N_6115);
nand U11282 (N_11282,N_5961,N_6525);
nand U11283 (N_11283,N_5846,N_6333);
nand U11284 (N_11284,N_6292,N_4890);
nor U11285 (N_11285,N_5801,N_5641);
nor U11286 (N_11286,N_7710,N_7417);
nor U11287 (N_11287,N_7535,N_4504);
and U11288 (N_11288,N_7552,N_7100);
or U11289 (N_11289,N_4527,N_4699);
and U11290 (N_11290,N_5056,N_4691);
and U11291 (N_11291,N_5672,N_7549);
nor U11292 (N_11292,N_7292,N_6731);
or U11293 (N_11293,N_7861,N_6933);
and U11294 (N_11294,N_5400,N_6255);
and U11295 (N_11295,N_6706,N_7922);
nor U11296 (N_11296,N_5664,N_5174);
and U11297 (N_11297,N_5338,N_5181);
and U11298 (N_11298,N_7496,N_7530);
nor U11299 (N_11299,N_4133,N_5689);
or U11300 (N_11300,N_5871,N_6995);
and U11301 (N_11301,N_7629,N_6592);
nor U11302 (N_11302,N_5181,N_5722);
and U11303 (N_11303,N_4876,N_5973);
and U11304 (N_11304,N_6590,N_7911);
or U11305 (N_11305,N_6880,N_4675);
or U11306 (N_11306,N_7658,N_4442);
or U11307 (N_11307,N_7958,N_4394);
nor U11308 (N_11308,N_4528,N_5156);
nand U11309 (N_11309,N_7289,N_6431);
nor U11310 (N_11310,N_6267,N_5845);
nand U11311 (N_11311,N_7951,N_4228);
and U11312 (N_11312,N_7492,N_6446);
nor U11313 (N_11313,N_5339,N_5469);
nand U11314 (N_11314,N_7877,N_4012);
nand U11315 (N_11315,N_4167,N_4316);
nor U11316 (N_11316,N_5327,N_7355);
nand U11317 (N_11317,N_4844,N_7328);
xor U11318 (N_11318,N_6700,N_7100);
nand U11319 (N_11319,N_5877,N_6626);
nor U11320 (N_11320,N_4426,N_6051);
nand U11321 (N_11321,N_4275,N_4332);
xor U11322 (N_11322,N_6388,N_7539);
nor U11323 (N_11323,N_4156,N_5970);
nand U11324 (N_11324,N_5751,N_6803);
nor U11325 (N_11325,N_5689,N_7133);
nor U11326 (N_11326,N_4124,N_5823);
or U11327 (N_11327,N_5637,N_5568);
or U11328 (N_11328,N_5490,N_6287);
nor U11329 (N_11329,N_7648,N_4045);
or U11330 (N_11330,N_4673,N_6643);
nand U11331 (N_11331,N_7259,N_4378);
nor U11332 (N_11332,N_6012,N_6117);
nor U11333 (N_11333,N_7896,N_6117);
nor U11334 (N_11334,N_6704,N_4487);
and U11335 (N_11335,N_4698,N_5094);
or U11336 (N_11336,N_5299,N_6432);
or U11337 (N_11337,N_4840,N_4172);
nor U11338 (N_11338,N_5498,N_6922);
or U11339 (N_11339,N_6605,N_6104);
and U11340 (N_11340,N_5130,N_4854);
and U11341 (N_11341,N_4672,N_4136);
xnor U11342 (N_11342,N_7268,N_5385);
nand U11343 (N_11343,N_6320,N_5371);
or U11344 (N_11344,N_4192,N_5132);
or U11345 (N_11345,N_4932,N_6377);
nand U11346 (N_11346,N_5057,N_7827);
nand U11347 (N_11347,N_4406,N_4891);
or U11348 (N_11348,N_6863,N_7274);
or U11349 (N_11349,N_4529,N_7840);
nor U11350 (N_11350,N_6462,N_6596);
nor U11351 (N_11351,N_7743,N_4125);
xor U11352 (N_11352,N_7722,N_7149);
nand U11353 (N_11353,N_5974,N_7851);
nand U11354 (N_11354,N_5516,N_7593);
or U11355 (N_11355,N_4001,N_7875);
nor U11356 (N_11356,N_7815,N_7863);
and U11357 (N_11357,N_5716,N_5775);
or U11358 (N_11358,N_7579,N_4319);
or U11359 (N_11359,N_4757,N_6776);
nand U11360 (N_11360,N_6923,N_6383);
or U11361 (N_11361,N_7953,N_7079);
nor U11362 (N_11362,N_7135,N_6062);
or U11363 (N_11363,N_6324,N_6762);
nand U11364 (N_11364,N_4291,N_4417);
or U11365 (N_11365,N_6620,N_6642);
or U11366 (N_11366,N_6694,N_4919);
nor U11367 (N_11367,N_5972,N_5904);
and U11368 (N_11368,N_6606,N_4697);
or U11369 (N_11369,N_6124,N_7937);
or U11370 (N_11370,N_5175,N_5720);
nand U11371 (N_11371,N_6109,N_5818);
nor U11372 (N_11372,N_6412,N_5287);
nor U11373 (N_11373,N_4646,N_4801);
nor U11374 (N_11374,N_6964,N_7992);
or U11375 (N_11375,N_5080,N_4093);
or U11376 (N_11376,N_7010,N_7989);
nor U11377 (N_11377,N_6316,N_5313);
nor U11378 (N_11378,N_7652,N_6268);
nand U11379 (N_11379,N_4050,N_6820);
and U11380 (N_11380,N_7180,N_6355);
and U11381 (N_11381,N_6970,N_4883);
or U11382 (N_11382,N_6910,N_4555);
and U11383 (N_11383,N_4163,N_7082);
nor U11384 (N_11384,N_5748,N_4844);
nor U11385 (N_11385,N_7781,N_6827);
nand U11386 (N_11386,N_7542,N_6270);
and U11387 (N_11387,N_7371,N_4032);
and U11388 (N_11388,N_5882,N_6001);
or U11389 (N_11389,N_7693,N_5888);
nor U11390 (N_11390,N_4612,N_5069);
nor U11391 (N_11391,N_6769,N_7772);
nand U11392 (N_11392,N_7795,N_4325);
nand U11393 (N_11393,N_6981,N_7906);
nor U11394 (N_11394,N_5095,N_4669);
nand U11395 (N_11395,N_4196,N_6176);
and U11396 (N_11396,N_6647,N_6122);
or U11397 (N_11397,N_7174,N_4302);
or U11398 (N_11398,N_4644,N_4010);
nor U11399 (N_11399,N_7304,N_5654);
or U11400 (N_11400,N_4874,N_4048);
nand U11401 (N_11401,N_7518,N_7352);
nor U11402 (N_11402,N_4684,N_7086);
or U11403 (N_11403,N_5334,N_7663);
and U11404 (N_11404,N_6557,N_4492);
or U11405 (N_11405,N_4074,N_4597);
nor U11406 (N_11406,N_6401,N_7541);
nor U11407 (N_11407,N_4757,N_4626);
and U11408 (N_11408,N_7450,N_4267);
nor U11409 (N_11409,N_7695,N_4217);
nor U11410 (N_11410,N_4646,N_5190);
and U11411 (N_11411,N_7611,N_4960);
nor U11412 (N_11412,N_7187,N_7525);
or U11413 (N_11413,N_6695,N_5886);
and U11414 (N_11414,N_6129,N_7016);
nor U11415 (N_11415,N_4124,N_5727);
and U11416 (N_11416,N_4113,N_5228);
nand U11417 (N_11417,N_5307,N_4766);
nand U11418 (N_11418,N_6298,N_5538);
nor U11419 (N_11419,N_6399,N_4108);
nand U11420 (N_11420,N_4779,N_7019);
or U11421 (N_11421,N_5840,N_6862);
nor U11422 (N_11422,N_5908,N_6858);
or U11423 (N_11423,N_5280,N_7967);
or U11424 (N_11424,N_7998,N_6504);
nand U11425 (N_11425,N_5889,N_6714);
nand U11426 (N_11426,N_4937,N_7970);
or U11427 (N_11427,N_4631,N_4672);
nor U11428 (N_11428,N_6111,N_6607);
or U11429 (N_11429,N_5526,N_6766);
and U11430 (N_11430,N_5391,N_7075);
nand U11431 (N_11431,N_5777,N_5741);
nor U11432 (N_11432,N_5973,N_5305);
nor U11433 (N_11433,N_5455,N_7906);
and U11434 (N_11434,N_5812,N_5318);
or U11435 (N_11435,N_7157,N_5001);
or U11436 (N_11436,N_7015,N_7125);
nor U11437 (N_11437,N_5456,N_5258);
or U11438 (N_11438,N_6281,N_5484);
nor U11439 (N_11439,N_4783,N_6913);
and U11440 (N_11440,N_5707,N_7861);
or U11441 (N_11441,N_5406,N_6981);
and U11442 (N_11442,N_6469,N_5743);
or U11443 (N_11443,N_6205,N_4905);
or U11444 (N_11444,N_7358,N_7593);
or U11445 (N_11445,N_6434,N_4806);
nand U11446 (N_11446,N_6244,N_6332);
and U11447 (N_11447,N_4163,N_6967);
and U11448 (N_11448,N_4213,N_7943);
nand U11449 (N_11449,N_6535,N_7837);
and U11450 (N_11450,N_4585,N_7969);
xnor U11451 (N_11451,N_4294,N_4877);
and U11452 (N_11452,N_4362,N_5113);
or U11453 (N_11453,N_7242,N_5827);
nand U11454 (N_11454,N_6736,N_7165);
and U11455 (N_11455,N_4872,N_7913);
or U11456 (N_11456,N_5115,N_6031);
nor U11457 (N_11457,N_5047,N_4926);
nor U11458 (N_11458,N_6756,N_6140);
and U11459 (N_11459,N_7701,N_4561);
or U11460 (N_11460,N_7449,N_7447);
or U11461 (N_11461,N_5317,N_6455);
nand U11462 (N_11462,N_5078,N_4045);
or U11463 (N_11463,N_4838,N_7704);
nor U11464 (N_11464,N_6880,N_7476);
and U11465 (N_11465,N_7569,N_5880);
and U11466 (N_11466,N_6650,N_6143);
nand U11467 (N_11467,N_7184,N_4382);
nand U11468 (N_11468,N_4978,N_4083);
or U11469 (N_11469,N_4471,N_4580);
and U11470 (N_11470,N_5428,N_4970);
nand U11471 (N_11471,N_4460,N_6353);
and U11472 (N_11472,N_6573,N_7700);
nor U11473 (N_11473,N_5764,N_5833);
or U11474 (N_11474,N_6207,N_6379);
nor U11475 (N_11475,N_6279,N_7039);
and U11476 (N_11476,N_5117,N_6913);
and U11477 (N_11477,N_7398,N_7190);
nand U11478 (N_11478,N_5359,N_5575);
nand U11479 (N_11479,N_5122,N_7290);
or U11480 (N_11480,N_5344,N_5815);
or U11481 (N_11481,N_5890,N_5963);
nand U11482 (N_11482,N_6925,N_5351);
or U11483 (N_11483,N_4183,N_7197);
and U11484 (N_11484,N_7497,N_7906);
and U11485 (N_11485,N_4521,N_7346);
and U11486 (N_11486,N_6947,N_6491);
nor U11487 (N_11487,N_4286,N_6741);
nand U11488 (N_11488,N_4202,N_4406);
and U11489 (N_11489,N_5362,N_6263);
or U11490 (N_11490,N_4015,N_6484);
or U11491 (N_11491,N_7004,N_4592);
and U11492 (N_11492,N_5381,N_4620);
nor U11493 (N_11493,N_4263,N_7302);
nand U11494 (N_11494,N_4575,N_4597);
or U11495 (N_11495,N_5540,N_6761);
and U11496 (N_11496,N_5441,N_5584);
nand U11497 (N_11497,N_4353,N_4835);
or U11498 (N_11498,N_7011,N_6030);
nor U11499 (N_11499,N_6823,N_5880);
xor U11500 (N_11500,N_5724,N_5214);
nor U11501 (N_11501,N_7907,N_5982);
or U11502 (N_11502,N_5402,N_7624);
and U11503 (N_11503,N_5036,N_6245);
or U11504 (N_11504,N_5283,N_4707);
nor U11505 (N_11505,N_7047,N_4738);
or U11506 (N_11506,N_5551,N_6361);
or U11507 (N_11507,N_4809,N_6507);
nor U11508 (N_11508,N_6965,N_6036);
nor U11509 (N_11509,N_6781,N_7218);
or U11510 (N_11510,N_7301,N_7498);
or U11511 (N_11511,N_7952,N_6639);
nor U11512 (N_11512,N_6451,N_4943);
nor U11513 (N_11513,N_6066,N_6775);
nor U11514 (N_11514,N_5217,N_6614);
nor U11515 (N_11515,N_7989,N_6224);
nor U11516 (N_11516,N_5905,N_7735);
nor U11517 (N_11517,N_7241,N_4959);
nor U11518 (N_11518,N_6030,N_6145);
or U11519 (N_11519,N_6856,N_4535);
nand U11520 (N_11520,N_4700,N_5955);
nand U11521 (N_11521,N_4422,N_6877);
and U11522 (N_11522,N_6251,N_7110);
nor U11523 (N_11523,N_6902,N_5941);
or U11524 (N_11524,N_4640,N_6755);
or U11525 (N_11525,N_4734,N_4501);
and U11526 (N_11526,N_7408,N_6125);
nor U11527 (N_11527,N_5132,N_5662);
or U11528 (N_11528,N_5952,N_5387);
xnor U11529 (N_11529,N_7470,N_5589);
nand U11530 (N_11530,N_4719,N_7607);
and U11531 (N_11531,N_7313,N_6140);
and U11532 (N_11532,N_7147,N_6202);
nor U11533 (N_11533,N_5623,N_6436);
or U11534 (N_11534,N_7533,N_6460);
nand U11535 (N_11535,N_6719,N_7774);
nand U11536 (N_11536,N_4698,N_5135);
and U11537 (N_11537,N_5785,N_4446);
and U11538 (N_11538,N_5142,N_6623);
and U11539 (N_11539,N_6243,N_6832);
and U11540 (N_11540,N_4323,N_4729);
or U11541 (N_11541,N_4270,N_5578);
and U11542 (N_11542,N_7765,N_7658);
nor U11543 (N_11543,N_6818,N_6316);
nor U11544 (N_11544,N_6591,N_6820);
and U11545 (N_11545,N_4042,N_7442);
nor U11546 (N_11546,N_6419,N_4736);
and U11547 (N_11547,N_6874,N_4110);
nand U11548 (N_11548,N_5826,N_4328);
or U11549 (N_11549,N_6552,N_4976);
xor U11550 (N_11550,N_5046,N_7344);
nand U11551 (N_11551,N_6710,N_7702);
or U11552 (N_11552,N_4812,N_4978);
or U11553 (N_11553,N_6111,N_7359);
nand U11554 (N_11554,N_7525,N_5377);
and U11555 (N_11555,N_6737,N_7501);
nand U11556 (N_11556,N_4623,N_4689);
nor U11557 (N_11557,N_7095,N_6221);
nand U11558 (N_11558,N_7405,N_7209);
nor U11559 (N_11559,N_4193,N_5198);
or U11560 (N_11560,N_5995,N_7926);
or U11561 (N_11561,N_7296,N_5768);
or U11562 (N_11562,N_4170,N_7375);
nor U11563 (N_11563,N_4129,N_6250);
or U11564 (N_11564,N_7278,N_4331);
nand U11565 (N_11565,N_7375,N_7481);
and U11566 (N_11566,N_6291,N_6914);
nor U11567 (N_11567,N_7094,N_4251);
or U11568 (N_11568,N_6478,N_7848);
nand U11569 (N_11569,N_4618,N_5009);
and U11570 (N_11570,N_5983,N_5525);
nand U11571 (N_11571,N_7454,N_7471);
nand U11572 (N_11572,N_4813,N_5673);
nor U11573 (N_11573,N_4764,N_7940);
nand U11574 (N_11574,N_4358,N_6717);
or U11575 (N_11575,N_6810,N_4408);
nor U11576 (N_11576,N_6122,N_7890);
nand U11577 (N_11577,N_7992,N_4813);
nand U11578 (N_11578,N_4802,N_5773);
or U11579 (N_11579,N_5597,N_5569);
nor U11580 (N_11580,N_4346,N_5542);
nor U11581 (N_11581,N_5025,N_4813);
nand U11582 (N_11582,N_4726,N_4956);
or U11583 (N_11583,N_7426,N_7148);
nand U11584 (N_11584,N_6122,N_6391);
or U11585 (N_11585,N_4163,N_6907);
nor U11586 (N_11586,N_4369,N_6145);
and U11587 (N_11587,N_6116,N_4114);
or U11588 (N_11588,N_4006,N_5351);
nor U11589 (N_11589,N_6638,N_5283);
or U11590 (N_11590,N_4566,N_6968);
nor U11591 (N_11591,N_7653,N_7648);
nor U11592 (N_11592,N_6766,N_4823);
and U11593 (N_11593,N_4003,N_4016);
nor U11594 (N_11594,N_6014,N_7103);
or U11595 (N_11595,N_4804,N_6768);
nand U11596 (N_11596,N_5148,N_4823);
nor U11597 (N_11597,N_5127,N_4503);
nor U11598 (N_11598,N_6360,N_7084);
or U11599 (N_11599,N_7315,N_7485);
or U11600 (N_11600,N_5309,N_5957);
nand U11601 (N_11601,N_7447,N_6069);
and U11602 (N_11602,N_4822,N_7960);
nand U11603 (N_11603,N_4193,N_5500);
and U11604 (N_11604,N_7684,N_7267);
nor U11605 (N_11605,N_4893,N_4497);
or U11606 (N_11606,N_6762,N_5667);
or U11607 (N_11607,N_5626,N_4087);
or U11608 (N_11608,N_7790,N_5853);
or U11609 (N_11609,N_5380,N_5510);
nand U11610 (N_11610,N_6339,N_7426);
or U11611 (N_11611,N_4799,N_5099);
and U11612 (N_11612,N_7070,N_4887);
or U11613 (N_11613,N_6656,N_5330);
or U11614 (N_11614,N_4195,N_6707);
or U11615 (N_11615,N_5722,N_5705);
or U11616 (N_11616,N_5817,N_4789);
and U11617 (N_11617,N_5215,N_4841);
and U11618 (N_11618,N_6980,N_4033);
nand U11619 (N_11619,N_6688,N_6080);
and U11620 (N_11620,N_7660,N_4101);
and U11621 (N_11621,N_5131,N_7967);
and U11622 (N_11622,N_5417,N_5240);
nor U11623 (N_11623,N_4742,N_5905);
and U11624 (N_11624,N_6199,N_7309);
or U11625 (N_11625,N_7351,N_6833);
nand U11626 (N_11626,N_4172,N_6573);
nand U11627 (N_11627,N_4974,N_4709);
or U11628 (N_11628,N_5404,N_4159);
or U11629 (N_11629,N_6146,N_7108);
and U11630 (N_11630,N_6945,N_7672);
or U11631 (N_11631,N_6002,N_6627);
or U11632 (N_11632,N_4983,N_6571);
or U11633 (N_11633,N_4750,N_7110);
and U11634 (N_11634,N_5909,N_4001);
and U11635 (N_11635,N_5516,N_7365);
or U11636 (N_11636,N_4174,N_5014);
nand U11637 (N_11637,N_5571,N_5985);
nand U11638 (N_11638,N_7697,N_7810);
nor U11639 (N_11639,N_6649,N_6983);
nand U11640 (N_11640,N_5424,N_6749);
or U11641 (N_11641,N_7515,N_7808);
nand U11642 (N_11642,N_5439,N_4086);
or U11643 (N_11643,N_7274,N_7150);
nand U11644 (N_11644,N_4425,N_6789);
nor U11645 (N_11645,N_4920,N_5462);
or U11646 (N_11646,N_6508,N_5368);
and U11647 (N_11647,N_6473,N_7317);
nand U11648 (N_11648,N_5585,N_4103);
and U11649 (N_11649,N_4720,N_6580);
nor U11650 (N_11650,N_5998,N_5454);
and U11651 (N_11651,N_5499,N_7884);
or U11652 (N_11652,N_4449,N_7790);
and U11653 (N_11653,N_6649,N_4780);
and U11654 (N_11654,N_5462,N_4986);
nand U11655 (N_11655,N_6768,N_4068);
nand U11656 (N_11656,N_4440,N_4537);
nand U11657 (N_11657,N_4679,N_4147);
and U11658 (N_11658,N_4200,N_4009);
and U11659 (N_11659,N_5347,N_4766);
or U11660 (N_11660,N_6530,N_7224);
or U11661 (N_11661,N_4710,N_4958);
nand U11662 (N_11662,N_4782,N_5747);
or U11663 (N_11663,N_4948,N_4543);
nand U11664 (N_11664,N_6110,N_5875);
and U11665 (N_11665,N_4040,N_4619);
and U11666 (N_11666,N_6368,N_6825);
nand U11667 (N_11667,N_4156,N_7364);
and U11668 (N_11668,N_4131,N_6130);
and U11669 (N_11669,N_5638,N_5042);
or U11670 (N_11670,N_7816,N_6099);
and U11671 (N_11671,N_5471,N_4584);
and U11672 (N_11672,N_6835,N_4385);
nand U11673 (N_11673,N_5066,N_6760);
or U11674 (N_11674,N_4670,N_7770);
nand U11675 (N_11675,N_6482,N_7662);
nand U11676 (N_11676,N_5069,N_5580);
nor U11677 (N_11677,N_5049,N_6863);
or U11678 (N_11678,N_4117,N_6173);
and U11679 (N_11679,N_7827,N_5857);
and U11680 (N_11680,N_5958,N_5471);
or U11681 (N_11681,N_4960,N_6385);
or U11682 (N_11682,N_7019,N_5650);
xor U11683 (N_11683,N_5867,N_7687);
and U11684 (N_11684,N_5345,N_4550);
nand U11685 (N_11685,N_7046,N_4654);
and U11686 (N_11686,N_4784,N_6531);
nand U11687 (N_11687,N_4528,N_5328);
nand U11688 (N_11688,N_6003,N_6970);
nor U11689 (N_11689,N_4352,N_4956);
and U11690 (N_11690,N_4223,N_5666);
nand U11691 (N_11691,N_4901,N_4681);
and U11692 (N_11692,N_4787,N_4216);
nand U11693 (N_11693,N_5321,N_4966);
nor U11694 (N_11694,N_6211,N_5356);
nor U11695 (N_11695,N_6590,N_6958);
nor U11696 (N_11696,N_4588,N_5894);
nor U11697 (N_11697,N_6045,N_5599);
or U11698 (N_11698,N_4094,N_5523);
and U11699 (N_11699,N_4234,N_5984);
nor U11700 (N_11700,N_4552,N_7098);
and U11701 (N_11701,N_6884,N_7757);
nand U11702 (N_11702,N_4500,N_7715);
or U11703 (N_11703,N_6900,N_7299);
nand U11704 (N_11704,N_6392,N_6495);
or U11705 (N_11705,N_5014,N_4946);
nor U11706 (N_11706,N_5515,N_5835);
nor U11707 (N_11707,N_5899,N_5071);
and U11708 (N_11708,N_6515,N_6145);
nand U11709 (N_11709,N_6545,N_4522);
nand U11710 (N_11710,N_6981,N_6489);
or U11711 (N_11711,N_4553,N_7325);
or U11712 (N_11712,N_6985,N_7774);
nor U11713 (N_11713,N_6461,N_7082);
xor U11714 (N_11714,N_4490,N_4658);
or U11715 (N_11715,N_6994,N_7905);
nor U11716 (N_11716,N_4030,N_6579);
or U11717 (N_11717,N_6040,N_7375);
and U11718 (N_11718,N_6803,N_4271);
nor U11719 (N_11719,N_5790,N_7268);
or U11720 (N_11720,N_4235,N_6352);
nand U11721 (N_11721,N_5636,N_6648);
and U11722 (N_11722,N_6593,N_5510);
or U11723 (N_11723,N_7470,N_4483);
nor U11724 (N_11724,N_7202,N_6664);
or U11725 (N_11725,N_4034,N_6749);
and U11726 (N_11726,N_5362,N_7304);
nand U11727 (N_11727,N_5054,N_7707);
or U11728 (N_11728,N_4044,N_4068);
nand U11729 (N_11729,N_6100,N_7920);
nand U11730 (N_11730,N_5587,N_6385);
nor U11731 (N_11731,N_6073,N_6945);
nor U11732 (N_11732,N_6480,N_5820);
and U11733 (N_11733,N_6108,N_4971);
nand U11734 (N_11734,N_6205,N_7097);
nand U11735 (N_11735,N_6921,N_6395);
nor U11736 (N_11736,N_4526,N_4395);
nand U11737 (N_11737,N_6487,N_7744);
nor U11738 (N_11738,N_6215,N_4944);
or U11739 (N_11739,N_4899,N_4976);
nand U11740 (N_11740,N_7360,N_5689);
nor U11741 (N_11741,N_6412,N_6186);
and U11742 (N_11742,N_4989,N_5640);
nand U11743 (N_11743,N_6519,N_4717);
or U11744 (N_11744,N_6385,N_7053);
nand U11745 (N_11745,N_6179,N_6720);
nor U11746 (N_11746,N_4591,N_7820);
and U11747 (N_11747,N_7622,N_6239);
nand U11748 (N_11748,N_5819,N_4272);
or U11749 (N_11749,N_5764,N_5042);
or U11750 (N_11750,N_6197,N_4373);
nand U11751 (N_11751,N_4103,N_7299);
and U11752 (N_11752,N_6921,N_7839);
nor U11753 (N_11753,N_6598,N_6158);
and U11754 (N_11754,N_5823,N_6534);
and U11755 (N_11755,N_5772,N_5799);
and U11756 (N_11756,N_7606,N_6561);
or U11757 (N_11757,N_7158,N_6263);
nand U11758 (N_11758,N_5789,N_5231);
or U11759 (N_11759,N_7534,N_4881);
nor U11760 (N_11760,N_5258,N_4498);
nor U11761 (N_11761,N_5056,N_7603);
nand U11762 (N_11762,N_5123,N_6289);
nand U11763 (N_11763,N_7707,N_4874);
or U11764 (N_11764,N_4275,N_7254);
nand U11765 (N_11765,N_4740,N_5376);
nand U11766 (N_11766,N_6224,N_7490);
and U11767 (N_11767,N_6012,N_7371);
nand U11768 (N_11768,N_7634,N_5447);
and U11769 (N_11769,N_4018,N_5508);
or U11770 (N_11770,N_6272,N_7955);
nand U11771 (N_11771,N_4060,N_7642);
and U11772 (N_11772,N_5558,N_6638);
nand U11773 (N_11773,N_5742,N_7025);
and U11774 (N_11774,N_6849,N_6013);
and U11775 (N_11775,N_6976,N_7858);
and U11776 (N_11776,N_4781,N_4912);
and U11777 (N_11777,N_4316,N_6241);
or U11778 (N_11778,N_6618,N_6290);
and U11779 (N_11779,N_7047,N_4909);
or U11780 (N_11780,N_7729,N_5800);
or U11781 (N_11781,N_7756,N_6471);
nor U11782 (N_11782,N_7982,N_7591);
and U11783 (N_11783,N_4484,N_5306);
or U11784 (N_11784,N_7608,N_4832);
or U11785 (N_11785,N_5057,N_5405);
and U11786 (N_11786,N_5683,N_6290);
nor U11787 (N_11787,N_4167,N_5567);
nand U11788 (N_11788,N_4345,N_6627);
or U11789 (N_11789,N_4406,N_7073);
nand U11790 (N_11790,N_7846,N_7581);
or U11791 (N_11791,N_6631,N_6159);
xnor U11792 (N_11792,N_6798,N_4638);
and U11793 (N_11793,N_5295,N_6429);
nand U11794 (N_11794,N_6478,N_4648);
nor U11795 (N_11795,N_4210,N_5603);
nor U11796 (N_11796,N_6031,N_5740);
nor U11797 (N_11797,N_4167,N_7254);
and U11798 (N_11798,N_5930,N_4545);
nand U11799 (N_11799,N_4360,N_7862);
and U11800 (N_11800,N_6082,N_4437);
and U11801 (N_11801,N_7708,N_4087);
nand U11802 (N_11802,N_4429,N_7593);
or U11803 (N_11803,N_4625,N_4433);
and U11804 (N_11804,N_5646,N_7042);
and U11805 (N_11805,N_5912,N_4157);
nand U11806 (N_11806,N_4003,N_5715);
nor U11807 (N_11807,N_4051,N_5510);
and U11808 (N_11808,N_7576,N_6792);
and U11809 (N_11809,N_7012,N_6740);
nand U11810 (N_11810,N_7198,N_7299);
nor U11811 (N_11811,N_4949,N_7132);
nor U11812 (N_11812,N_5391,N_7350);
xnor U11813 (N_11813,N_7485,N_6955);
nand U11814 (N_11814,N_4440,N_7032);
nor U11815 (N_11815,N_5600,N_4474);
nor U11816 (N_11816,N_4737,N_5288);
or U11817 (N_11817,N_7810,N_5216);
nor U11818 (N_11818,N_5669,N_4994);
nor U11819 (N_11819,N_6839,N_7232);
and U11820 (N_11820,N_4140,N_7403);
and U11821 (N_11821,N_7074,N_7652);
nor U11822 (N_11822,N_4511,N_6343);
or U11823 (N_11823,N_7966,N_7490);
nand U11824 (N_11824,N_4050,N_7451);
and U11825 (N_11825,N_4597,N_7824);
or U11826 (N_11826,N_6076,N_7903);
and U11827 (N_11827,N_6559,N_6161);
and U11828 (N_11828,N_4698,N_7089);
nand U11829 (N_11829,N_5510,N_5934);
nand U11830 (N_11830,N_6379,N_6513);
nor U11831 (N_11831,N_6334,N_6933);
nor U11832 (N_11832,N_5483,N_7695);
or U11833 (N_11833,N_4894,N_5653);
xnor U11834 (N_11834,N_5868,N_4154);
nor U11835 (N_11835,N_7948,N_6807);
or U11836 (N_11836,N_4528,N_4595);
and U11837 (N_11837,N_5619,N_7072);
and U11838 (N_11838,N_5333,N_6765);
and U11839 (N_11839,N_4207,N_4500);
or U11840 (N_11840,N_4209,N_6212);
nor U11841 (N_11841,N_4248,N_4254);
or U11842 (N_11842,N_5156,N_6225);
and U11843 (N_11843,N_7849,N_7434);
nor U11844 (N_11844,N_6207,N_4458);
nor U11845 (N_11845,N_4080,N_4819);
or U11846 (N_11846,N_7505,N_4485);
and U11847 (N_11847,N_6972,N_7818);
nand U11848 (N_11848,N_6355,N_5682);
or U11849 (N_11849,N_4433,N_4117);
or U11850 (N_11850,N_5634,N_6736);
nand U11851 (N_11851,N_7709,N_4944);
and U11852 (N_11852,N_5156,N_7666);
nor U11853 (N_11853,N_5065,N_7638);
nand U11854 (N_11854,N_6850,N_6982);
and U11855 (N_11855,N_6535,N_4519);
nor U11856 (N_11856,N_7031,N_4984);
nand U11857 (N_11857,N_4658,N_7820);
or U11858 (N_11858,N_7288,N_7891);
and U11859 (N_11859,N_6482,N_7636);
nand U11860 (N_11860,N_5580,N_6051);
and U11861 (N_11861,N_7577,N_7227);
or U11862 (N_11862,N_4220,N_7785);
and U11863 (N_11863,N_6053,N_7469);
and U11864 (N_11864,N_5166,N_7503);
and U11865 (N_11865,N_5157,N_5190);
and U11866 (N_11866,N_7933,N_6268);
or U11867 (N_11867,N_7899,N_7079);
nor U11868 (N_11868,N_7830,N_4884);
or U11869 (N_11869,N_4494,N_4145);
nand U11870 (N_11870,N_4019,N_6365);
and U11871 (N_11871,N_6002,N_7246);
and U11872 (N_11872,N_4344,N_5578);
and U11873 (N_11873,N_6063,N_7476);
or U11874 (N_11874,N_5385,N_5946);
and U11875 (N_11875,N_5458,N_5105);
and U11876 (N_11876,N_7126,N_6811);
nand U11877 (N_11877,N_7016,N_7200);
or U11878 (N_11878,N_6893,N_7918);
nand U11879 (N_11879,N_5216,N_6377);
and U11880 (N_11880,N_5929,N_5377);
or U11881 (N_11881,N_4190,N_7426);
or U11882 (N_11882,N_6215,N_6978);
and U11883 (N_11883,N_6701,N_4122);
and U11884 (N_11884,N_4832,N_6494);
nand U11885 (N_11885,N_5056,N_5926);
nand U11886 (N_11886,N_7528,N_7072);
and U11887 (N_11887,N_4252,N_4088);
nand U11888 (N_11888,N_6628,N_4632);
nor U11889 (N_11889,N_6973,N_5640);
nor U11890 (N_11890,N_5858,N_7596);
and U11891 (N_11891,N_5324,N_7821);
nand U11892 (N_11892,N_6338,N_4483);
and U11893 (N_11893,N_7091,N_6130);
nor U11894 (N_11894,N_7659,N_4645);
and U11895 (N_11895,N_6213,N_4286);
nand U11896 (N_11896,N_5999,N_6284);
nand U11897 (N_11897,N_6639,N_7278);
or U11898 (N_11898,N_4151,N_4916);
nor U11899 (N_11899,N_5147,N_6086);
xor U11900 (N_11900,N_7408,N_7601);
or U11901 (N_11901,N_4073,N_7294);
nor U11902 (N_11902,N_6380,N_5014);
nor U11903 (N_11903,N_6277,N_6493);
and U11904 (N_11904,N_4848,N_6775);
and U11905 (N_11905,N_4057,N_7969);
or U11906 (N_11906,N_7903,N_6338);
and U11907 (N_11907,N_4647,N_7566);
nand U11908 (N_11908,N_4711,N_4321);
nor U11909 (N_11909,N_6756,N_7319);
or U11910 (N_11910,N_4393,N_4000);
or U11911 (N_11911,N_5127,N_4020);
or U11912 (N_11912,N_7133,N_7799);
or U11913 (N_11913,N_5501,N_5753);
or U11914 (N_11914,N_4738,N_5126);
or U11915 (N_11915,N_5856,N_4089);
and U11916 (N_11916,N_7341,N_7508);
nor U11917 (N_11917,N_6670,N_5104);
or U11918 (N_11918,N_7193,N_6019);
nand U11919 (N_11919,N_4706,N_4654);
nor U11920 (N_11920,N_5121,N_4912);
nand U11921 (N_11921,N_5257,N_4529);
or U11922 (N_11922,N_4738,N_6196);
nand U11923 (N_11923,N_6883,N_7649);
and U11924 (N_11924,N_7506,N_6926);
or U11925 (N_11925,N_6177,N_7737);
or U11926 (N_11926,N_6395,N_5903);
and U11927 (N_11927,N_4034,N_5132);
nand U11928 (N_11928,N_7979,N_6862);
nor U11929 (N_11929,N_6095,N_6145);
and U11930 (N_11930,N_6953,N_4545);
and U11931 (N_11931,N_4706,N_6016);
nand U11932 (N_11932,N_4181,N_4740);
and U11933 (N_11933,N_6002,N_4624);
nand U11934 (N_11934,N_6471,N_4039);
nor U11935 (N_11935,N_5884,N_6986);
or U11936 (N_11936,N_4463,N_6219);
and U11937 (N_11937,N_6185,N_7908);
and U11938 (N_11938,N_6190,N_5572);
or U11939 (N_11939,N_6588,N_6725);
nor U11940 (N_11940,N_5114,N_7167);
nand U11941 (N_11941,N_6462,N_5425);
nand U11942 (N_11942,N_7723,N_7380);
and U11943 (N_11943,N_5005,N_7060);
nor U11944 (N_11944,N_5486,N_6775);
and U11945 (N_11945,N_7261,N_5190);
nor U11946 (N_11946,N_7697,N_6125);
nor U11947 (N_11947,N_7360,N_6627);
or U11948 (N_11948,N_4210,N_5046);
nor U11949 (N_11949,N_7395,N_6671);
nor U11950 (N_11950,N_5667,N_5048);
and U11951 (N_11951,N_4248,N_5856);
nor U11952 (N_11952,N_4991,N_6439);
nor U11953 (N_11953,N_6430,N_4351);
and U11954 (N_11954,N_6476,N_7667);
nand U11955 (N_11955,N_4276,N_6294);
nor U11956 (N_11956,N_4120,N_5735);
and U11957 (N_11957,N_5994,N_4008);
nand U11958 (N_11958,N_5603,N_6157);
and U11959 (N_11959,N_4794,N_5157);
or U11960 (N_11960,N_4090,N_5637);
nor U11961 (N_11961,N_6114,N_4603);
or U11962 (N_11962,N_4469,N_5926);
and U11963 (N_11963,N_7940,N_6823);
and U11964 (N_11964,N_6620,N_6059);
or U11965 (N_11965,N_7758,N_5563);
or U11966 (N_11966,N_5078,N_6147);
nor U11967 (N_11967,N_4129,N_5943);
and U11968 (N_11968,N_5584,N_5346);
nor U11969 (N_11969,N_5588,N_7563);
and U11970 (N_11970,N_7640,N_5242);
nand U11971 (N_11971,N_7020,N_4917);
nand U11972 (N_11972,N_7547,N_5637);
nor U11973 (N_11973,N_7188,N_4156);
and U11974 (N_11974,N_7812,N_5615);
and U11975 (N_11975,N_6664,N_6793);
nand U11976 (N_11976,N_4473,N_7580);
nor U11977 (N_11977,N_6643,N_5946);
nor U11978 (N_11978,N_7117,N_7240);
nand U11979 (N_11979,N_6139,N_4412);
or U11980 (N_11980,N_5984,N_4306);
xor U11981 (N_11981,N_7689,N_7527);
or U11982 (N_11982,N_4027,N_4160);
nand U11983 (N_11983,N_7477,N_4099);
nand U11984 (N_11984,N_6991,N_5960);
or U11985 (N_11985,N_4332,N_5341);
nor U11986 (N_11986,N_4375,N_4586);
nand U11987 (N_11987,N_7943,N_4827);
and U11988 (N_11988,N_6287,N_5718);
or U11989 (N_11989,N_5745,N_5730);
and U11990 (N_11990,N_4896,N_7250);
nor U11991 (N_11991,N_7751,N_4905);
nand U11992 (N_11992,N_6203,N_6877);
nand U11993 (N_11993,N_4226,N_6097);
or U11994 (N_11994,N_6202,N_6894);
nand U11995 (N_11995,N_5917,N_4221);
nor U11996 (N_11996,N_5357,N_4859);
or U11997 (N_11997,N_7880,N_4624);
and U11998 (N_11998,N_5087,N_5965);
nor U11999 (N_11999,N_6870,N_7875);
and U12000 (N_12000,N_11342,N_10084);
nor U12001 (N_12001,N_11595,N_11509);
and U12002 (N_12002,N_10278,N_8012);
nand U12003 (N_12003,N_8680,N_9268);
and U12004 (N_12004,N_11117,N_9676);
nand U12005 (N_12005,N_8470,N_8142);
xor U12006 (N_12006,N_10486,N_11851);
and U12007 (N_12007,N_8460,N_10822);
or U12008 (N_12008,N_8160,N_11877);
and U12009 (N_12009,N_10636,N_11217);
nand U12010 (N_12010,N_10770,N_9538);
or U12011 (N_12011,N_11749,N_9009);
or U12012 (N_12012,N_8639,N_10623);
nand U12013 (N_12013,N_9472,N_11312);
and U12014 (N_12014,N_10480,N_11896);
nor U12015 (N_12015,N_10938,N_11604);
nand U12016 (N_12016,N_9111,N_10397);
and U12017 (N_12017,N_11937,N_10026);
nor U12018 (N_12018,N_8951,N_10362);
or U12019 (N_12019,N_9267,N_10483);
nor U12020 (N_12020,N_8032,N_10400);
nor U12021 (N_12021,N_8857,N_8945);
and U12022 (N_12022,N_10191,N_9673);
xnor U12023 (N_12023,N_8802,N_9156);
and U12024 (N_12024,N_8300,N_11576);
nand U12025 (N_12025,N_8441,N_8363);
nand U12026 (N_12026,N_8276,N_10305);
and U12027 (N_12027,N_11722,N_10217);
and U12028 (N_12028,N_10686,N_11285);
and U12029 (N_12029,N_8906,N_10898);
nand U12030 (N_12030,N_9315,N_11613);
and U12031 (N_12031,N_11485,N_8289);
nand U12032 (N_12032,N_10885,N_9912);
nor U12033 (N_12033,N_9557,N_8166);
and U12034 (N_12034,N_10440,N_10621);
nand U12035 (N_12035,N_8941,N_8590);
or U12036 (N_12036,N_8874,N_8294);
nor U12037 (N_12037,N_10341,N_11904);
nand U12038 (N_12038,N_9048,N_8255);
and U12039 (N_12039,N_8690,N_9917);
and U12040 (N_12040,N_8675,N_11003);
nand U12041 (N_12041,N_9715,N_10069);
and U12042 (N_12042,N_11524,N_10167);
or U12043 (N_12043,N_9858,N_11736);
nor U12044 (N_12044,N_10658,N_11548);
nor U12045 (N_12045,N_8402,N_10399);
and U12046 (N_12046,N_9145,N_9155);
and U12047 (N_12047,N_9840,N_8340);
nor U12048 (N_12048,N_9570,N_11328);
or U12049 (N_12049,N_8625,N_8665);
and U12050 (N_12050,N_10860,N_11711);
nand U12051 (N_12051,N_10116,N_10450);
nor U12052 (N_12052,N_10939,N_9940);
nand U12053 (N_12053,N_8650,N_8643);
nand U12054 (N_12054,N_10465,N_11667);
and U12055 (N_12055,N_10025,N_11290);
nor U12056 (N_12056,N_9656,N_11822);
nand U12057 (N_12057,N_10408,N_10209);
and U12058 (N_12058,N_8637,N_11570);
nand U12059 (N_12059,N_11743,N_9028);
nor U12060 (N_12060,N_11377,N_10169);
nand U12061 (N_12061,N_11925,N_10716);
nor U12062 (N_12062,N_8522,N_8054);
nand U12063 (N_12063,N_8751,N_9446);
or U12064 (N_12064,N_9195,N_11383);
nor U12065 (N_12065,N_10256,N_10171);
nand U12066 (N_12066,N_9835,N_9959);
nor U12067 (N_12067,N_9704,N_8345);
nor U12068 (N_12068,N_10604,N_8278);
nor U12069 (N_12069,N_9292,N_8664);
nor U12070 (N_12070,N_8275,N_11910);
and U12071 (N_12071,N_8956,N_11634);
or U12072 (N_12072,N_9851,N_8656);
or U12073 (N_12073,N_11766,N_11958);
nand U12074 (N_12074,N_9432,N_11070);
nand U12075 (N_12075,N_9277,N_8872);
nand U12076 (N_12076,N_10456,N_8417);
nor U12077 (N_12077,N_9168,N_10033);
or U12078 (N_12078,N_11337,N_10335);
nor U12079 (N_12079,N_9493,N_9394);
or U12080 (N_12080,N_8888,N_11861);
nand U12081 (N_12081,N_10331,N_8057);
nor U12082 (N_12082,N_8817,N_11039);
nand U12083 (N_12083,N_8626,N_10005);
or U12084 (N_12084,N_9924,N_9342);
nand U12085 (N_12085,N_10911,N_10142);
nand U12086 (N_12086,N_10926,N_9494);
and U12087 (N_12087,N_10760,N_9757);
and U12088 (N_12088,N_11410,N_11187);
and U12089 (N_12089,N_10119,N_9211);
and U12090 (N_12090,N_8086,N_9030);
or U12091 (N_12091,N_10462,N_9122);
nor U12092 (N_12092,N_11515,N_10637);
nand U12093 (N_12093,N_11374,N_8673);
or U12094 (N_12094,N_10539,N_11905);
and U12095 (N_12095,N_9084,N_9995);
nor U12096 (N_12096,N_10192,N_9659);
nor U12097 (N_12097,N_10311,N_9876);
nor U12098 (N_12098,N_11840,N_9371);
xnor U12099 (N_12099,N_9541,N_8954);
and U12100 (N_12100,N_9126,N_9958);
nand U12101 (N_12101,N_11565,N_8394);
and U12102 (N_12102,N_10837,N_11615);
nand U12103 (N_12103,N_8213,N_10366);
nand U12104 (N_12104,N_11335,N_10742);
or U12105 (N_12105,N_11409,N_9230);
xor U12106 (N_12106,N_8988,N_8467);
or U12107 (N_12107,N_8575,N_9583);
nand U12108 (N_12108,N_11894,N_11735);
and U12109 (N_12109,N_8715,N_10394);
nand U12110 (N_12110,N_11493,N_11418);
or U12111 (N_12111,N_9669,N_11620);
nand U12112 (N_12112,N_10106,N_10523);
and U12113 (N_12113,N_9117,N_10502);
or U12114 (N_12114,N_9784,N_10086);
and U12115 (N_12115,N_10055,N_9745);
nand U12116 (N_12116,N_11541,N_10471);
nand U12117 (N_12117,N_11519,N_9564);
or U12118 (N_12118,N_10600,N_10920);
and U12119 (N_12119,N_8725,N_9161);
or U12120 (N_12120,N_11975,N_8567);
nor U12121 (N_12121,N_9593,N_8783);
and U12122 (N_12122,N_11994,N_10891);
and U12123 (N_12123,N_10886,N_10390);
and U12124 (N_12124,N_10349,N_11372);
or U12125 (N_12125,N_9590,N_9597);
nand U12126 (N_12126,N_11564,N_10093);
or U12127 (N_12127,N_11303,N_11249);
and U12128 (N_12128,N_11927,N_8246);
nor U12129 (N_12129,N_11072,N_9154);
nor U12130 (N_12130,N_9044,N_9439);
or U12131 (N_12131,N_10029,N_9334);
and U12132 (N_12132,N_9772,N_9120);
nand U12133 (N_12133,N_10384,N_11890);
nor U12134 (N_12134,N_9068,N_10446);
nor U12135 (N_12135,N_10546,N_8514);
or U12136 (N_12136,N_9610,N_9857);
xnor U12137 (N_12137,N_9611,N_11288);
or U12138 (N_12138,N_9531,N_8288);
nand U12139 (N_12139,N_8759,N_10620);
or U12140 (N_12140,N_9584,N_8488);
nand U12141 (N_12141,N_11608,N_11734);
nor U12142 (N_12142,N_11996,N_10152);
or U12143 (N_12143,N_11833,N_11776);
or U12144 (N_12144,N_9470,N_9206);
nor U12145 (N_12145,N_11394,N_9183);
and U12146 (N_12146,N_11148,N_10490);
nand U12147 (N_12147,N_9534,N_11528);
nor U12148 (N_12148,N_11049,N_9299);
nor U12149 (N_12149,N_9499,N_9992);
nor U12150 (N_12150,N_10754,N_10518);
xor U12151 (N_12151,N_10238,N_9109);
and U12152 (N_12152,N_10099,N_10975);
or U12153 (N_12153,N_8842,N_9916);
nor U12154 (N_12154,N_10965,N_9599);
nand U12155 (N_12155,N_10160,N_8471);
and U12156 (N_12156,N_8104,N_9215);
and U12157 (N_12157,N_10771,N_8846);
and U12158 (N_12158,N_8138,N_9083);
and U12159 (N_12159,N_9838,N_9407);
nand U12160 (N_12160,N_10221,N_11078);
and U12161 (N_12161,N_11081,N_10113);
nor U12162 (N_12162,N_11431,N_9633);
nand U12163 (N_12163,N_9485,N_10285);
nand U12164 (N_12164,N_8611,N_9424);
or U12165 (N_12165,N_8122,N_10413);
nor U12166 (N_12166,N_8862,N_11046);
or U12167 (N_12167,N_10818,N_11286);
nand U12168 (N_12168,N_10847,N_11522);
nand U12169 (N_12169,N_9953,N_11345);
nand U12170 (N_12170,N_11508,N_10946);
and U12171 (N_12171,N_10892,N_8020);
nand U12172 (N_12172,N_8808,N_8531);
nor U12173 (N_12173,N_8425,N_9212);
and U12174 (N_12174,N_8434,N_11464);
or U12175 (N_12175,N_8666,N_9535);
or U12176 (N_12176,N_9519,N_9073);
nor U12177 (N_12177,N_9790,N_10650);
nor U12178 (N_12178,N_9164,N_11650);
and U12179 (N_12179,N_9910,N_9844);
or U12180 (N_12180,N_8899,N_10125);
and U12181 (N_12181,N_9635,N_8310);
or U12182 (N_12182,N_11683,N_11741);
nor U12183 (N_12183,N_8173,N_8458);
or U12184 (N_12184,N_10003,N_11820);
nand U12185 (N_12185,N_10286,N_8655);
and U12186 (N_12186,N_8962,N_11752);
and U12187 (N_12187,N_9771,N_11916);
or U12188 (N_12188,N_8169,N_8306);
or U12189 (N_12189,N_10109,N_8062);
or U12190 (N_12190,N_8612,N_11503);
or U12191 (N_12191,N_10201,N_10448);
or U12192 (N_12192,N_11102,N_8630);
nor U12193 (N_12193,N_10479,N_11566);
nand U12194 (N_12194,N_9678,N_9140);
nand U12195 (N_12195,N_8823,N_10075);
nor U12196 (N_12196,N_8309,N_11255);
and U12197 (N_12197,N_9850,N_10706);
or U12198 (N_12198,N_10810,N_9675);
or U12199 (N_12199,N_11992,N_11662);
nor U12200 (N_12200,N_10163,N_11582);
nor U12201 (N_12201,N_9974,N_9730);
and U12202 (N_12202,N_9779,N_11853);
and U12203 (N_12203,N_9809,N_9276);
nand U12204 (N_12204,N_11474,N_9588);
nor U12205 (N_12205,N_10629,N_10264);
or U12206 (N_12206,N_11154,N_9795);
and U12207 (N_12207,N_9194,N_10309);
nor U12208 (N_12208,N_11147,N_11484);
nand U12209 (N_12209,N_11583,N_8800);
and U12210 (N_12210,N_8125,N_9740);
nor U12211 (N_12211,N_9888,N_11980);
nor U12212 (N_12212,N_8192,N_8555);
nor U12213 (N_12213,N_10387,N_8442);
nand U12214 (N_12214,N_8421,N_11118);
or U12215 (N_12215,N_8430,N_11309);
and U12216 (N_12216,N_11351,N_8787);
and U12217 (N_12217,N_9454,N_9889);
nand U12218 (N_12218,N_11450,N_8498);
and U12219 (N_12219,N_8006,N_8815);
nand U12220 (N_12220,N_8068,N_10582);
nor U12221 (N_12221,N_9294,N_9280);
and U12222 (N_12222,N_9142,N_10591);
and U12223 (N_12223,N_9387,N_9725);
nor U12224 (N_12224,N_9688,N_8709);
or U12225 (N_12225,N_8948,N_9563);
or U12226 (N_12226,N_9124,N_9138);
nand U12227 (N_12227,N_8557,N_10333);
and U12228 (N_12228,N_10615,N_8033);
or U12229 (N_12229,N_11126,N_9748);
nand U12230 (N_12230,N_9020,N_9004);
or U12231 (N_12231,N_9094,N_9556);
nand U12232 (N_12232,N_10094,N_11499);
nor U12233 (N_12233,N_11220,N_10098);
or U12234 (N_12234,N_11965,N_11647);
nand U12235 (N_12235,N_11557,N_11703);
or U12236 (N_12236,N_11966,N_10469);
or U12237 (N_12237,N_9349,N_9234);
or U12238 (N_12238,N_11918,N_8970);
or U12239 (N_12239,N_11543,N_11844);
or U12240 (N_12240,N_10897,N_10375);
and U12241 (N_12241,N_10510,N_9753);
and U12242 (N_12242,N_11325,N_10701);
or U12243 (N_12243,N_8355,N_9104);
and U12244 (N_12244,N_10261,N_11502);
nand U12245 (N_12245,N_11691,N_10454);
or U12246 (N_12246,N_10583,N_8745);
nor U12247 (N_12247,N_11350,N_11511);
or U12248 (N_12248,N_10673,N_11213);
and U12249 (N_12249,N_11706,N_9674);
nand U12250 (N_12250,N_10964,N_9525);
nor U12251 (N_12251,N_8215,N_8359);
and U12252 (N_12252,N_9340,N_8194);
and U12253 (N_12253,N_8913,N_9724);
nand U12254 (N_12254,N_10932,N_8283);
and U12255 (N_12255,N_9150,N_10419);
nor U12256 (N_12256,N_11056,N_10787);
or U12257 (N_12257,N_10412,N_11322);
nand U12258 (N_12258,N_10213,N_10695);
nor U12259 (N_12259,N_8279,N_8238);
and U12260 (N_12260,N_11069,N_9899);
or U12261 (N_12261,N_9067,N_10208);
nor U12262 (N_12262,N_11804,N_11439);
or U12263 (N_12263,N_10095,N_11516);
and U12264 (N_12264,N_11919,N_9710);
nor U12265 (N_12265,N_9905,N_10194);
nand U12266 (N_12266,N_11641,N_11007);
or U12267 (N_12267,N_10269,N_10713);
nand U12268 (N_12268,N_9957,N_8143);
nor U12269 (N_12269,N_8195,N_8902);
or U12270 (N_12270,N_9241,N_9722);
nor U12271 (N_12271,N_11159,N_11600);
nor U12272 (N_12272,N_11184,N_11610);
nor U12273 (N_12273,N_8245,N_8632);
nand U12274 (N_12274,N_10628,N_8833);
nor U12275 (N_12275,N_9575,N_8649);
nor U12276 (N_12276,N_11866,N_10326);
or U12277 (N_12277,N_10157,N_11315);
nor U12278 (N_12278,N_8504,N_8876);
and U12279 (N_12279,N_10914,N_11441);
and U12280 (N_12280,N_9312,N_9655);
nor U12281 (N_12281,N_9062,N_10108);
or U12282 (N_12282,N_10193,N_10402);
xnor U12283 (N_12283,N_8079,N_8546);
or U12284 (N_12284,N_11035,N_11211);
and U12285 (N_12285,N_9647,N_8510);
and U12286 (N_12286,N_10556,N_10605);
nor U12287 (N_12287,N_10903,N_8569);
nor U12288 (N_12288,N_9650,N_11061);
and U12289 (N_12289,N_8181,N_11795);
and U12290 (N_12290,N_9727,N_8391);
and U12291 (N_12291,N_10291,N_9765);
and U12292 (N_12292,N_8197,N_9482);
nor U12293 (N_12293,N_11120,N_10571);
nor U12294 (N_12294,N_11505,N_10078);
or U12295 (N_12295,N_8864,N_9964);
nand U12296 (N_12296,N_8766,N_9359);
and U12297 (N_12297,N_11801,N_9598);
nand U12298 (N_12298,N_10350,N_8542);
or U12299 (N_12299,N_9479,N_9434);
or U12300 (N_12300,N_9954,N_9946);
nand U12301 (N_12301,N_10232,N_10536);
or U12302 (N_12302,N_9318,N_11589);
and U12303 (N_12303,N_9540,N_10596);
or U12304 (N_12304,N_10014,N_11802);
or U12305 (N_12305,N_11214,N_9732);
nand U12306 (N_12306,N_10352,N_9311);
and U12307 (N_12307,N_11205,N_11057);
nor U12308 (N_12308,N_11402,N_9481);
nor U12309 (N_12309,N_10149,N_9460);
nand U12310 (N_12310,N_10044,N_10246);
nor U12311 (N_12311,N_9660,N_9459);
or U12312 (N_12312,N_11097,N_8552);
nor U12313 (N_12313,N_10888,N_9198);
nor U12314 (N_12314,N_11770,N_9148);
and U12315 (N_12315,N_9592,N_8982);
or U12316 (N_12316,N_10519,N_11623);
and U12317 (N_12317,N_10534,N_11984);
xor U12318 (N_12318,N_11429,N_10184);
and U12319 (N_12319,N_11584,N_8834);
and U12320 (N_12320,N_9993,N_9372);
nand U12321 (N_12321,N_8399,N_9239);
or U12322 (N_12322,N_9613,N_9224);
and U12323 (N_12323,N_10531,N_11514);
or U12324 (N_12324,N_10659,N_10521);
nor U12325 (N_12325,N_11892,N_9373);
nand U12326 (N_12326,N_9928,N_10312);
nand U12327 (N_12327,N_10737,N_10243);
nor U12328 (N_12328,N_8856,N_11104);
and U12329 (N_12329,N_9783,N_8211);
and U12330 (N_12330,N_10477,N_10916);
and U12331 (N_12331,N_10931,N_8588);
or U12332 (N_12332,N_9248,N_11912);
or U12333 (N_12333,N_11852,N_10940);
nand U12334 (N_12334,N_9892,N_8485);
nor U12335 (N_12335,N_11614,N_10239);
or U12336 (N_12336,N_10494,N_8327);
or U12337 (N_12337,N_8495,N_9865);
or U12338 (N_12338,N_10685,N_10316);
nand U12339 (N_12339,N_10786,N_11875);
nand U12340 (N_12340,N_9622,N_11181);
nor U12341 (N_12341,N_11763,N_9400);
or U12342 (N_12342,N_10606,N_11863);
nand U12343 (N_12343,N_11062,N_10665);
nand U12344 (N_12344,N_11942,N_8468);
and U12345 (N_12345,N_10386,N_9685);
or U12346 (N_12346,N_9418,N_10730);
nand U12347 (N_12347,N_10065,N_10879);
nand U12348 (N_12348,N_10010,N_10838);
nand U12349 (N_12349,N_9602,N_11789);
and U12350 (N_12350,N_8087,N_10070);
or U12351 (N_12351,N_10758,N_10207);
and U12352 (N_12352,N_11920,N_10361);
nand U12353 (N_12353,N_8339,N_11730);
nor U12354 (N_12354,N_9329,N_9392);
and U12355 (N_12355,N_8227,N_11172);
and U12356 (N_12356,N_8868,N_10547);
and U12357 (N_12357,N_10773,N_10498);
and U12358 (N_12358,N_8628,N_10551);
and U12359 (N_12359,N_8593,N_8404);
nor U12360 (N_12360,N_11386,N_10991);
nand U12361 (N_12361,N_11272,N_9214);
nor U12362 (N_12362,N_9511,N_11532);
and U12363 (N_12363,N_9476,N_11228);
nor U12364 (N_12364,N_10042,N_8298);
or U12365 (N_12365,N_11999,N_9934);
nor U12366 (N_12366,N_9034,N_10175);
and U12367 (N_12367,N_9813,N_9537);
nand U12368 (N_12368,N_10865,N_11810);
nor U12369 (N_12369,N_11141,N_9546);
and U12370 (N_12370,N_8521,N_11713);
and U12371 (N_12371,N_8174,N_11670);
and U12372 (N_12372,N_8741,N_11343);
and U12373 (N_12373,N_9000,N_10420);
nor U12374 (N_12374,N_8040,N_9770);
nor U12375 (N_12375,N_9501,N_10962);
nand U12376 (N_12376,N_11066,N_10423);
nand U12377 (N_12377,N_8131,N_8882);
or U12378 (N_12378,N_8285,N_9877);
nor U12379 (N_12379,N_8570,N_9759);
nor U12380 (N_12380,N_9014,N_11242);
nand U12381 (N_12381,N_10218,N_9990);
or U12382 (N_12382,N_9042,N_8199);
or U12383 (N_12383,N_9384,N_11082);
or U12384 (N_12384,N_8201,N_8343);
or U12385 (N_12385,N_10712,N_9343);
and U12386 (N_12386,N_10196,N_10151);
nand U12387 (N_12387,N_11116,N_9799);
nor U12388 (N_12388,N_11478,N_11448);
nor U12389 (N_12389,N_9947,N_10825);
xnor U12390 (N_12390,N_10287,N_9587);
or U12391 (N_12391,N_8381,N_8223);
nor U12392 (N_12392,N_11948,N_10688);
or U12393 (N_12393,N_10128,N_11581);
nand U12394 (N_12394,N_10241,N_9792);
nor U12395 (N_12395,N_10705,N_8983);
and U12396 (N_12396,N_9997,N_10577);
or U12397 (N_12397,N_11700,N_11936);
and U12398 (N_12398,N_9011,N_10200);
nand U12399 (N_12399,N_9475,N_9064);
nand U12400 (N_12400,N_11024,N_11191);
nand U12401 (N_12401,N_9487,N_10907);
or U12402 (N_12402,N_8216,N_11512);
nor U12403 (N_12403,N_10781,N_10012);
nand U12404 (N_12404,N_9167,N_11510);
nor U12405 (N_12405,N_8676,N_11067);
nand U12406 (N_12406,N_8036,N_9843);
nand U12407 (N_12407,N_11127,N_11353);
xor U12408 (N_12408,N_10321,N_9737);
or U12409 (N_12409,N_11950,N_10899);
nand U12410 (N_12410,N_10460,N_8247);
nand U12411 (N_12411,N_11972,N_10908);
or U12412 (N_12412,N_8317,N_9093);
and U12413 (N_12413,N_8387,N_8738);
or U12414 (N_12414,N_10276,N_11000);
nor U12415 (N_12415,N_9679,N_11107);
nor U12416 (N_12416,N_9060,N_8648);
nand U12417 (N_12417,N_8536,N_8607);
nor U12418 (N_12418,N_11321,N_10757);
or U12419 (N_12419,N_9108,N_11696);
nor U12420 (N_12420,N_8616,N_9023);
or U12421 (N_12421,N_9015,N_8583);
nor U12422 (N_12422,N_9883,N_11277);
and U12423 (N_12423,N_9604,N_10631);
and U12424 (N_12424,N_10726,N_10370);
nand U12425 (N_12425,N_11777,N_10764);
nand U12426 (N_12426,N_11358,N_9290);
nor U12427 (N_12427,N_8384,N_11949);
or U12428 (N_12428,N_11506,N_11204);
nand U12429 (N_12429,N_11675,N_8221);
and U12430 (N_12430,N_8670,N_10247);
and U12431 (N_12431,N_10994,N_8809);
nor U12432 (N_12432,N_10953,N_9483);
and U12433 (N_12433,N_8953,N_11336);
and U12434 (N_12434,N_8157,N_11628);
or U12435 (N_12435,N_10784,N_10266);
or U12436 (N_12436,N_10874,N_9965);
nor U12437 (N_12437,N_10796,N_11563);
or U12438 (N_12438,N_9272,N_8475);
nor U12439 (N_12439,N_9542,N_9718);
nand U12440 (N_12440,N_11029,N_8700);
and U12441 (N_12441,N_9555,N_8537);
or U12442 (N_12442,N_9265,N_11855);
nand U12443 (N_12443,N_10776,N_8204);
and U12444 (N_12444,N_9202,N_8870);
nand U12445 (N_12445,N_11196,N_10626);
nand U12446 (N_12446,N_10210,N_11869);
and U12447 (N_12447,N_9505,N_10942);
and U12448 (N_12448,N_11079,N_10297);
nand U12449 (N_12449,N_8155,N_11481);
xnor U12450 (N_12450,N_11207,N_9119);
or U12451 (N_12451,N_8263,N_8291);
or U12452 (N_12452,N_10056,N_8580);
or U12453 (N_12453,N_11674,N_11324);
and U12454 (N_12454,N_11655,N_10609);
and U12455 (N_12455,N_10259,N_8248);
nand U12456 (N_12456,N_9890,N_10429);
or U12457 (N_12457,N_11546,N_11986);
nor U12458 (N_12458,N_10330,N_8711);
nor U12459 (N_12459,N_9869,N_11917);
nor U12460 (N_12460,N_11451,N_10585);
nor U12461 (N_12461,N_9378,N_8353);
and U12462 (N_12462,N_10587,N_10640);
and U12463 (N_12463,N_11001,N_11593);
nand U12464 (N_12464,N_10870,N_11672);
nor U12465 (N_12465,N_8739,N_11969);
nor U12466 (N_12466,N_9433,N_8513);
xor U12467 (N_12467,N_8875,N_10242);
or U12468 (N_12468,N_8686,N_8452);
nand U12469 (N_12469,N_10393,N_10206);
and U12470 (N_12470,N_9035,N_8017);
xor U12471 (N_12471,N_9099,N_8048);
or U12472 (N_12472,N_9072,N_8177);
or U12473 (N_12473,N_10348,N_8334);
and U12474 (N_12474,N_11824,N_8069);
nand U12475 (N_12475,N_9780,N_11629);
nand U12476 (N_12476,N_9352,N_10385);
or U12477 (N_12477,N_11656,N_9812);
and U12478 (N_12478,N_9262,N_11329);
and U12479 (N_12479,N_8074,N_10775);
xnor U12480 (N_12480,N_11605,N_8241);
nand U12481 (N_12481,N_10910,N_9750);
nand U12482 (N_12482,N_10154,N_9152);
nor U12483 (N_12483,N_9766,N_8010);
nor U12484 (N_12484,N_8968,N_9581);
nor U12485 (N_12485,N_9082,N_10048);
nor U12486 (N_12486,N_11018,N_9648);
or U12487 (N_12487,N_11279,N_11831);
xnor U12488 (N_12488,N_10622,N_11729);
nand U12489 (N_12489,N_8435,N_9733);
nor U12490 (N_12490,N_9654,N_9667);
xnor U12491 (N_12491,N_9381,N_9526);
and U12492 (N_12492,N_8478,N_10308);
nand U12493 (N_12493,N_8184,N_10988);
nand U12494 (N_12494,N_11292,N_10553);
nand U12495 (N_12495,N_10441,N_10590);
nand U12496 (N_12496,N_9188,N_9642);
or U12497 (N_12497,N_11426,N_11334);
and U12498 (N_12498,N_9039,N_11501);
nand U12499 (N_12499,N_8743,N_10057);
nor U12500 (N_12500,N_11415,N_10199);
nor U12501 (N_12501,N_9565,N_8149);
nor U12502 (N_12502,N_10129,N_9474);
nand U12503 (N_12503,N_11050,N_10438);
and U12504 (N_12504,N_11778,N_8971);
and U12505 (N_12505,N_10832,N_9741);
nor U12506 (N_12506,N_11470,N_8920);
and U12507 (N_12507,N_10873,N_10145);
nor U12508 (N_12508,N_11771,N_11253);
or U12509 (N_12509,N_8893,N_8146);
and U12510 (N_12510,N_10476,N_8507);
or U12511 (N_12511,N_11542,N_10105);
and U12512 (N_12512,N_8663,N_9951);
nor U12513 (N_12513,N_11371,N_9661);
nand U12514 (N_12514,N_10538,N_11883);
nor U12515 (N_12515,N_10262,N_11265);
and U12516 (N_12516,N_8793,N_9322);
or U12517 (N_12517,N_11862,N_9001);
or U12518 (N_12518,N_10499,N_10520);
and U12519 (N_12519,N_10294,N_11480);
and U12520 (N_12520,N_11122,N_9553);
nand U12521 (N_12521,N_11712,N_8919);
nand U12522 (N_12522,N_8813,N_10731);
nor U12523 (N_12523,N_8424,N_8183);
nor U12524 (N_12524,N_8440,N_10922);
and U12525 (N_12525,N_11412,N_8065);
or U12526 (N_12526,N_8796,N_11819);
and U12527 (N_12527,N_8329,N_10500);
nand U12528 (N_12528,N_8852,N_10651);
nor U12529 (N_12529,N_11168,N_9046);
or U12530 (N_12530,N_11437,N_8024);
nand U12531 (N_12531,N_10222,N_10833);
nand U12532 (N_12532,N_11128,N_10166);
or U12533 (N_12533,N_11176,N_8323);
nor U12534 (N_12534,N_8691,N_8679);
nand U12535 (N_12535,N_11622,N_11302);
nor U12536 (N_12536,N_10819,N_11268);
or U12537 (N_12537,N_10566,N_11270);
and U12538 (N_12538,N_8973,N_10054);
nand U12539 (N_12539,N_8096,N_11174);
and U12540 (N_12540,N_8820,N_10506);
and U12541 (N_12541,N_8763,N_10844);
and U12542 (N_12542,N_10180,N_10445);
nor U12543 (N_12543,N_10114,N_9457);
xnor U12544 (N_12544,N_11455,N_10662);
or U12545 (N_12545,N_10972,N_10182);
xnor U12546 (N_12546,N_11230,N_8810);
or U12547 (N_12547,N_9693,N_9856);
nor U12548 (N_12548,N_9217,N_11550);
nand U12549 (N_12549,N_10474,N_10027);
and U12550 (N_12550,N_8088,N_8185);
nand U12551 (N_12551,N_11161,N_11945);
nor U12552 (N_12552,N_8845,N_11707);
nand U12553 (N_12553,N_8118,N_10258);
nand U12554 (N_12554,N_10458,N_9275);
and U12555 (N_12555,N_11715,N_8647);
and U12556 (N_12556,N_11538,N_9477);
nand U12557 (N_12557,N_10852,N_9132);
or U12558 (N_12558,N_8747,N_9429);
or U12559 (N_12559,N_10608,N_8210);
and U12560 (N_12560,N_9353,N_10329);
nand U12561 (N_12561,N_9480,N_9716);
nor U12562 (N_12562,N_11682,N_10409);
nand U12563 (N_12563,N_9837,N_9269);
nand U12564 (N_12564,N_11224,N_10415);
or U12565 (N_12565,N_8449,N_9832);
and U12566 (N_12566,N_8943,N_8901);
xor U12567 (N_12567,N_11422,N_9517);
or U12568 (N_12568,N_10593,N_11616);
nand U12569 (N_12569,N_10744,N_8224);
nand U12570 (N_12570,N_11143,N_8547);
and U12571 (N_12571,N_8801,N_11596);
nand U12572 (N_12572,N_11076,N_11673);
or U12573 (N_12573,N_9904,N_10568);
nand U12574 (N_12574,N_11816,N_8009);
nor U12575 (N_12575,N_10364,N_8635);
nor U12576 (N_12576,N_9503,N_11644);
nand U12577 (N_12577,N_9668,N_11330);
and U12578 (N_12578,N_8392,N_11311);
nor U12579 (N_12579,N_8703,N_8117);
nor U12580 (N_12580,N_11850,N_11212);
or U12581 (N_12581,N_9266,N_9281);
nand U12582 (N_12582,N_11243,N_8073);
or U12583 (N_12583,N_11577,N_11040);
nand U12584 (N_12584,N_10550,N_10282);
or U12585 (N_12585,N_11721,N_8287);
nand U12586 (N_12586,N_11215,N_8301);
nand U12587 (N_12587,N_11836,N_10130);
nor U12588 (N_12588,N_11828,N_8346);
nor U12589 (N_12589,N_8313,N_9747);
and U12590 (N_12590,N_11814,N_11065);
or U12591 (N_12591,N_11258,N_8462);
nand U12592 (N_12592,N_11149,N_8307);
and U12593 (N_12593,N_11155,N_11014);
and U12594 (N_12594,N_11103,N_11637);
or U12595 (N_12595,N_8749,N_10342);
nand U12596 (N_12596,N_9348,N_8367);
or U12597 (N_12597,N_11702,N_9834);
nor U12598 (N_12598,N_10955,N_9225);
or U12599 (N_12599,N_9894,N_9708);
or U12600 (N_12600,N_8877,N_10422);
nand U12601 (N_12601,N_11864,N_10868);
nand U12602 (N_12602,N_9335,N_9929);
or U12603 (N_12603,N_9141,N_11256);
nand U12604 (N_12604,N_9742,N_11033);
and U12605 (N_12605,N_10883,N_10648);
or U12606 (N_12606,N_9366,N_8419);
and U12607 (N_12607,N_9121,N_8900);
nand U12608 (N_12608,N_11843,N_11504);
nor U12609 (N_12609,N_11135,N_11839);
and U12610 (N_12610,N_11739,N_9881);
nand U12611 (N_12611,N_8113,N_11880);
nor U12612 (N_12612,N_11299,N_9802);
nor U12613 (N_12613,N_10993,N_9607);
nor U12614 (N_12614,N_8832,N_8252);
and U12615 (N_12615,N_10655,N_9797);
nand U12616 (N_12616,N_11893,N_11888);
nor U12617 (N_12617,N_8556,N_11421);
and U12618 (N_12618,N_11240,N_9186);
and U12619 (N_12619,N_11408,N_10143);
nor U12620 (N_12620,N_8942,N_10353);
nand U12621 (N_12621,N_8697,N_10992);
nor U12622 (N_12622,N_9231,N_11575);
or U12623 (N_12623,N_8476,N_10064);
or U12624 (N_12624,N_10089,N_9736);
or U12625 (N_12625,N_8744,N_8258);
and U12626 (N_12626,N_8105,N_11071);
and U12627 (N_12627,N_10540,N_11578);
nand U12628 (N_12628,N_10624,N_11817);
nand U12629 (N_12629,N_9734,N_8944);
nor U12630 (N_12630,N_8847,N_11047);
nor U12631 (N_12631,N_11601,N_8539);
nor U12632 (N_12632,N_11206,N_11401);
and U12633 (N_12633,N_11976,N_10969);
nand U12634 (N_12634,N_8758,N_11643);
nor U12635 (N_12635,N_8375,N_9402);
and U12636 (N_12636,N_10733,N_10777);
or U12637 (N_12637,N_8844,N_9087);
or U12638 (N_12638,N_10525,N_9723);
nand U12639 (N_12639,N_9226,N_9440);
or U12640 (N_12640,N_8383,N_10317);
nor U12641 (N_12641,N_11473,N_9096);
and U12642 (N_12642,N_11027,N_11599);
and U12643 (N_12643,N_9819,N_8443);
and U12644 (N_12644,N_10816,N_11555);
and U12645 (N_12645,N_11640,N_11178);
or U12646 (N_12646,N_10467,N_11301);
or U12647 (N_12647,N_8447,N_10411);
and U12648 (N_12648,N_8964,N_8865);
and U12649 (N_12649,N_9692,N_8829);
nand U12650 (N_12650,N_8914,N_9764);
and U12651 (N_12651,N_9278,N_11015);
and U12652 (N_12652,N_9775,N_8677);
and U12653 (N_12653,N_9841,N_9356);
or U12654 (N_12654,N_10850,N_9339);
nor U12655 (N_12655,N_8066,N_9829);
nand U12656 (N_12656,N_11758,N_8786);
nand U12657 (N_12657,N_11060,N_10367);
and U12658 (N_12658,N_8162,N_10447);
nand U12659 (N_12659,N_9902,N_9102);
nand U12660 (N_12660,N_10672,N_11544);
nand U12661 (N_12661,N_9443,N_11826);
nor U12662 (N_12662,N_10449,N_10530);
and U12663 (N_12663,N_11276,N_10389);
and U12664 (N_12664,N_9252,N_11140);
or U12665 (N_12665,N_8894,N_8388);
nor U12666 (N_12666,N_10378,N_8141);
nor U12667 (N_12667,N_11395,N_9497);
or U12668 (N_12668,N_11167,N_9444);
nand U12669 (N_12669,N_11086,N_8529);
nand U12670 (N_12670,N_9413,N_9054);
and U12671 (N_12671,N_10170,N_11813);
nand U12672 (N_12672,N_10514,N_11423);
or U12673 (N_12673,N_8814,N_10388);
nor U12674 (N_12674,N_9097,N_9071);
nand U12675 (N_12675,N_8072,N_10036);
nand U12676 (N_12676,N_8179,N_10782);
nand U12677 (N_12677,N_8070,N_11746);
and U12678 (N_12678,N_11034,N_11585);
or U12679 (N_12679,N_8060,N_8008);
nand U12680 (N_12680,N_9939,N_8240);
nor U12681 (N_12681,N_9363,N_8734);
nand U12682 (N_12682,N_9107,N_10373);
nor U12683 (N_12683,N_9749,N_11940);
and U12684 (N_12684,N_9815,N_8273);
or U12685 (N_12685,N_8129,N_9706);
nand U12686 (N_12686,N_11931,N_9776);
nand U12687 (N_12687,N_8361,N_9326);
nor U12688 (N_12688,N_10489,N_11287);
nand U12689 (N_12689,N_8338,N_8761);
nand U12690 (N_12690,N_8463,N_10322);
and U12691 (N_12691,N_9077,N_8170);
nand U12692 (N_12692,N_9682,N_10987);
or U12693 (N_12693,N_11961,N_11051);
or U12694 (N_12694,N_8684,N_9702);
nor U12695 (N_12695,N_10008,N_11882);
nor U12696 (N_12696,N_11259,N_11792);
nor U12697 (N_12697,N_9976,N_8541);
nor U12698 (N_12698,N_11317,N_8947);
or U12699 (N_12699,N_11115,N_9833);
and U12700 (N_12700,N_8851,N_9041);
and U12701 (N_12701,N_8867,N_8979);
or U12702 (N_12702,N_10821,N_9360);
nand U12703 (N_12703,N_10324,N_11856);
nor U12704 (N_12704,N_8360,N_10410);
nor U12705 (N_12705,N_9728,N_8871);
and U12706 (N_12706,N_11109,N_10328);
or U12707 (N_12707,N_11044,N_11327);
nor U12708 (N_12708,N_11815,N_10711);
nor U12709 (N_12709,N_10343,N_9296);
and U12710 (N_12710,N_9337,N_8782);
or U12711 (N_12711,N_10371,N_10038);
or U12712 (N_12712,N_9498,N_8114);
nor U12713 (N_12713,N_9756,N_9190);
nand U12714 (N_12714,N_10225,N_9293);
or U12715 (N_12715,N_8389,N_9448);
and U12716 (N_12716,N_9625,N_10696);
and U12717 (N_12717,N_10976,N_11129);
nor U12718 (N_12718,N_9336,N_11179);
nand U12719 (N_12719,N_8621,N_9263);
and U12720 (N_12720,N_9382,N_8497);
nor U12721 (N_12721,N_8256,N_8806);
or U12722 (N_12722,N_8422,N_9118);
and U12723 (N_12723,N_10884,N_8642);
nor U12724 (N_12724,N_9738,N_8083);
xor U12725 (N_12725,N_9242,N_10800);
or U12726 (N_12726,N_11762,N_9462);
nor U12727 (N_12727,N_11513,N_9786);
or U12728 (N_12728,N_9798,N_10882);
nor U12729 (N_12729,N_9385,N_10789);
nor U12730 (N_12730,N_11002,N_9621);
nor U12731 (N_12731,N_10267,N_10657);
or U12732 (N_12732,N_11955,N_8411);
nand U12733 (N_12733,N_8589,N_9170);
nand U12734 (N_12734,N_11536,N_11274);
or U12735 (N_12735,N_9410,N_8318);
nor U12736 (N_12736,N_8581,N_11121);
and U12737 (N_12737,N_10303,N_9341);
nand U12738 (N_12738,N_11340,N_8661);
nor U12739 (N_12739,N_9486,N_8050);
nand U12740 (N_12740,N_8041,N_9510);
nand U12741 (N_12741,N_8853,N_10491);
nor U12742 (N_12742,N_10481,N_10022);
nor U12743 (N_12743,N_10377,N_9056);
or U12744 (N_12744,N_11346,N_8658);
and U12745 (N_12745,N_8601,N_8726);
nand U12746 (N_12746,N_9403,N_11988);
xor U12747 (N_12747,N_10594,N_10947);
and U12748 (N_12748,N_11093,N_10215);
and U12749 (N_12749,N_10338,N_10846);
and U12750 (N_12750,N_8879,N_9411);
xor U12751 (N_12751,N_11177,N_9762);
nand U12752 (N_12752,N_9984,N_9447);
or U12753 (N_12753,N_8727,N_11624);
nor U12754 (N_12754,N_8311,N_9092);
or U12755 (N_12755,N_8502,N_9091);
nor U12756 (N_12756,N_10150,N_8641);
nor U12757 (N_12757,N_8631,N_10866);
or U12758 (N_12758,N_10096,N_11125);
nor U12759 (N_12759,N_8490,N_11554);
nand U12760 (N_12760,N_11338,N_11239);
or U12761 (N_12761,N_8472,N_10292);
nand U12762 (N_12762,N_9003,N_11390);
or U12763 (N_12763,N_9512,N_9058);
nand U12764 (N_12764,N_8506,N_8895);
nor U12765 (N_12765,N_11708,N_11545);
or U12766 (N_12766,N_10619,N_11089);
nor U12767 (N_12767,N_11225,N_8769);
nor U12768 (N_12768,N_8206,N_8144);
nor U12769 (N_12769,N_11716,N_10998);
nor U12770 (N_12770,N_8826,N_8023);
nand U12771 (N_12771,N_8516,N_11957);
nand U12772 (N_12772,N_10061,N_10788);
nor U12773 (N_12773,N_11084,N_8534);
and U12774 (N_12774,N_9379,N_9273);
and U12775 (N_12775,N_8265,N_10951);
and U12776 (N_12776,N_8707,N_9197);
nor U12777 (N_12777,N_9128,N_11222);
or U12778 (N_12778,N_9136,N_10958);
or U12779 (N_12779,N_8843,N_10255);
nand U12780 (N_12780,N_9919,N_8564);
or U12781 (N_12781,N_10532,N_8825);
or U12782 (N_12782,N_8390,N_10382);
nand U12783 (N_12783,N_9711,N_9769);
nand U12784 (N_12784,N_8921,N_9358);
or U12785 (N_12785,N_10552,N_8757);
nand U12786 (N_12786,N_11947,N_8304);
xor U12787 (N_12787,N_9651,N_10793);
nor U12788 (N_12788,N_9074,N_9287);
and U12789 (N_12789,N_11316,N_9567);
nand U12790 (N_12790,N_11251,N_8595);
or U12791 (N_12791,N_8249,N_8325);
nor U12792 (N_12792,N_8908,N_11430);
xor U12793 (N_12793,N_10216,N_10251);
nor U12794 (N_12794,N_8651,N_11435);
nand U12795 (N_12795,N_10558,N_11921);
and U12796 (N_12796,N_9681,N_9697);
and U12797 (N_12797,N_9047,N_11989);
and U12798 (N_12798,N_10252,N_10007);
and U12799 (N_12799,N_9867,N_10318);
or U12800 (N_12800,N_8981,N_11806);
and U12801 (N_12801,N_8321,N_9925);
or U12802 (N_12802,N_8619,N_10727);
and U12803 (N_12803,N_9395,N_8451);
nand U12804 (N_12804,N_9895,N_10376);
xor U12805 (N_12805,N_10613,N_8175);
or U12806 (N_12806,N_10859,N_8214);
nand U12807 (N_12807,N_8558,N_9589);
nand U12808 (N_12808,N_11970,N_8623);
xnor U12809 (N_12809,N_9886,N_11389);
nor U12810 (N_12810,N_8406,N_9615);
nand U12811 (N_12811,N_9991,N_8494);
or U12812 (N_12812,N_9491,N_11419);
nand U12813 (N_12813,N_8171,N_11232);
nor U12814 (N_12814,N_8268,N_11818);
nand U12815 (N_12815,N_10740,N_8401);
nor U12816 (N_12816,N_11262,N_10000);
nor U12817 (N_12817,N_10060,N_9430);
nand U12818 (N_12818,N_11192,N_10178);
nor U12819 (N_12819,N_8858,N_10340);
nor U12820 (N_12820,N_8044,N_11194);
nor U12821 (N_12821,N_10302,N_9853);
or U12822 (N_12822,N_9825,N_9636);
and U12823 (N_12823,N_11490,N_10709);
or U12824 (N_12824,N_8455,N_11573);
or U12825 (N_12825,N_8620,N_8492);
nand U12826 (N_12826,N_9078,N_9911);
nand U12827 (N_12827,N_10652,N_9049);
nand U12828 (N_12828,N_10876,N_9609);
or U12829 (N_12829,N_11489,N_9222);
nand U12830 (N_12830,N_9467,N_11110);
nand U12831 (N_12831,N_10526,N_8076);
nor U12832 (N_12832,N_8898,N_10501);
nand U12833 (N_12833,N_9406,N_11540);
nand U12834 (N_12834,N_9842,N_9376);
nor U12835 (N_12835,N_8597,N_11879);
nand U12836 (N_12836,N_9007,N_9735);
nor U12837 (N_12837,N_10656,N_9513);
nor U12838 (N_12838,N_10890,N_11373);
nor U12839 (N_12839,N_9146,N_11923);
or U12840 (N_12840,N_11720,N_10802);
nand U12841 (N_12841,N_8115,N_11361);
nor U12842 (N_12842,N_10049,N_10398);
nand U12843 (N_12843,N_11261,N_11150);
and U12844 (N_12844,N_11203,N_11105);
nor U12845 (N_12845,N_11870,N_10183);
or U12846 (N_12846,N_9703,N_8508);
nand U12847 (N_12847,N_9090,N_9139);
or U12848 (N_12848,N_11619,N_10037);
and U12849 (N_12849,N_8849,N_8746);
and U12850 (N_12850,N_8234,N_10563);
and U12851 (N_12851,N_8337,N_8167);
nor U12852 (N_12852,N_10612,N_8187);
or U12853 (N_12853,N_8461,N_10901);
and U12854 (N_12854,N_9861,N_8958);
nand U12855 (N_12855,N_8152,N_9305);
nand U12856 (N_12856,N_9388,N_8609);
or U12857 (N_12857,N_11393,N_8332);
nand U12858 (N_12858,N_10719,N_8159);
or U12859 (N_12859,N_9973,N_8374);
or U12860 (N_12860,N_8614,N_10186);
or U12861 (N_12861,N_11132,N_11635);
and U12862 (N_12862,N_8189,N_8038);
nor U12863 (N_12863,N_10134,N_11901);
nor U12864 (N_12864,N_10561,N_11688);
or U12865 (N_12865,N_8752,N_11355);
nand U12866 (N_12866,N_11413,N_10396);
nand U12867 (N_12867,N_8230,N_8604);
and U12868 (N_12868,N_8840,N_10772);
nand U12869 (N_12869,N_10881,N_10301);
and U12870 (N_12870,N_8000,N_8770);
and U12871 (N_12871,N_10346,N_10974);
nor U12872 (N_12872,N_9684,N_9628);
nor U12873 (N_12873,N_10919,N_9308);
nand U12874 (N_12874,N_9309,N_10374);
and U12875 (N_12875,N_10195,N_9595);
and U12876 (N_12876,N_10081,N_10016);
or U12877 (N_12877,N_10750,N_10799);
nor U12878 (N_12878,N_9966,N_10843);
nand U12879 (N_12879,N_11663,N_9302);
and U12880 (N_12880,N_11250,N_8615);
or U12881 (N_12881,N_9431,N_8127);
or U12882 (N_12882,N_11341,N_10808);
and U12883 (N_12883,N_8924,N_9804);
nand U12884 (N_12884,N_11123,N_10714);
nand U12885 (N_12885,N_10365,N_10933);
nor U12886 (N_12886,N_8866,N_10104);
or U12887 (N_12887,N_11556,N_11446);
or U12888 (N_12888,N_8491,N_10945);
nor U12889 (N_12889,N_10405,N_9032);
or U12890 (N_12890,N_10952,N_8634);
and U12891 (N_12891,N_10692,N_10189);
and U12892 (N_12892,N_9839,N_10960);
nand U12893 (N_12893,N_11981,N_10040);
nor U12894 (N_12894,N_8721,N_8154);
or U12895 (N_12895,N_8828,N_8640);
or U12896 (N_12896,N_8487,N_10080);
and U12897 (N_12897,N_10485,N_8835);
or U12898 (N_12898,N_9773,N_9282);
and U12899 (N_12899,N_8937,N_11952);
and U12900 (N_12900,N_8295,N_9948);
or U12901 (N_12901,N_9805,N_10136);
nand U12902 (N_12902,N_9791,N_11830);
or U12903 (N_12903,N_10774,N_11924);
and U12904 (N_12904,N_8016,N_8963);
and U12905 (N_12905,N_10981,N_8103);
and U12906 (N_12906,N_11694,N_10812);
nor U12907 (N_12907,N_10724,N_10878);
or U12908 (N_12908,N_10140,N_9871);
nor U12909 (N_12909,N_11227,N_9181);
or U12910 (N_12910,N_11209,N_11621);
nor U12911 (N_12911,N_10747,N_9549);
nand U12912 (N_12912,N_8188,N_10580);
or U12913 (N_12913,N_11829,N_9380);
or U12914 (N_12914,N_8095,N_9821);
and U12915 (N_12915,N_8133,N_9110);
or U12916 (N_12916,N_10334,N_11930);
nand U12917 (N_12917,N_9696,N_10107);
nand U12918 (N_12918,N_8091,N_10032);
nand U12919 (N_12919,N_10841,N_8290);
nand U12920 (N_12920,N_11681,N_11075);
and U12921 (N_12921,N_10190,N_9666);
nor U12922 (N_12922,N_8453,N_8785);
nand U12923 (N_12923,N_11530,N_11461);
nand U12924 (N_12924,N_9778,N_10660);
or U12925 (N_12925,N_8511,N_10263);
and U12926 (N_12926,N_10720,N_8830);
nand U12927 (N_12927,N_9401,N_9002);
or U12928 (N_12928,N_11973,N_11453);
nand U12929 (N_12929,N_9324,N_8955);
or U12930 (N_12930,N_10047,N_8582);
nand U12931 (N_12931,N_10339,N_9488);
nor U12932 (N_12932,N_11756,N_8678);
and U12933 (N_12933,N_8191,N_10248);
nand U12934 (N_12934,N_11726,N_11897);
and U12935 (N_12935,N_9787,N_11699);
and U12936 (N_12936,N_8203,N_11171);
nor U12937 (N_12937,N_10795,N_11760);
nand U12938 (N_12938,N_9412,N_8022);
nor U12939 (N_12939,N_11260,N_11041);
or U12940 (N_12940,N_10589,N_10050);
or U12941 (N_12941,N_11684,N_9080);
and U12942 (N_12942,N_9350,N_10139);
xnor U12943 (N_12943,N_9279,N_8836);
nor U12944 (N_12944,N_9427,N_11360);
nor U12945 (N_12945,N_10272,N_11567);
nand U12946 (N_12946,N_11909,N_10427);
and U12947 (N_12947,N_10856,N_9166);
nand U12948 (N_12948,N_10572,N_10451);
nand U12949 (N_12949,N_10146,N_10355);
nor U12950 (N_12950,N_11010,N_10574);
nand U12951 (N_12951,N_11382,N_8135);
nor U12952 (N_12952,N_11359,N_10970);
and U12953 (N_12953,N_9820,N_10478);
nand U12954 (N_12954,N_10369,N_9134);
and U12955 (N_12955,N_11380,N_8515);
and U12956 (N_12956,N_10893,N_10565);
or U12957 (N_12957,N_9192,N_9291);
and U12958 (N_12958,N_9926,N_9405);
or U12959 (N_12959,N_8123,N_9731);
and U12960 (N_12960,N_8551,N_8314);
nor U12961 (N_12961,N_11226,N_10562);
nor U12962 (N_12962,N_8819,N_8014);
or U12963 (N_12963,N_8667,N_11438);
or U12964 (N_12964,N_10127,N_8544);
or U12965 (N_12965,N_8420,N_11747);
nor U12966 (N_12966,N_9514,N_11469);
nand U12967 (N_12967,N_8055,N_8218);
nand U12968 (N_12968,N_9036,N_11693);
nand U12969 (N_12969,N_8775,N_11821);
nand U12970 (N_12970,N_8357,N_9085);
and U12971 (N_12971,N_8994,N_11825);
nand U12972 (N_12972,N_11399,N_8107);
and U12973 (N_12973,N_8890,N_11305);
and U12974 (N_12974,N_11891,N_10851);
nand U12975 (N_12975,N_11551,N_11114);
nor U12976 (N_12976,N_10896,N_11951);
nor U12977 (N_12977,N_9527,N_10442);
nor U12978 (N_12978,N_8423,N_8863);
nor U12979 (N_12979,N_8168,N_10978);
nor U12980 (N_12980,N_9763,N_8816);
nand U12981 (N_12981,N_10588,N_9670);
nand U12982 (N_12982,N_10584,N_9199);
and U12983 (N_12983,N_11718,N_8768);
and U12984 (N_12984,N_9619,N_10240);
nor U12985 (N_12985,N_8755,N_9752);
nand U12986 (N_12986,N_11476,N_8771);
nor U12987 (N_12987,N_11296,N_9903);
nand U12988 (N_12988,N_10840,N_9456);
nor U12989 (N_12989,N_11872,N_8912);
or U12990 (N_12990,N_11602,N_8124);
and U12991 (N_12991,N_11420,N_10807);
nand U12992 (N_12992,N_8884,N_11934);
nor U12993 (N_12993,N_8489,N_10363);
and U12994 (N_12994,N_8960,N_9461);
or U12995 (N_12995,N_9969,N_10118);
and U12996 (N_12996,N_11185,N_9235);
and U12997 (N_12997,N_10237,N_9826);
or U12998 (N_12998,N_9551,N_11709);
nor U12999 (N_12999,N_10780,N_8097);
and U13000 (N_13000,N_11823,N_11848);
or U13001 (N_13001,N_8106,N_8997);
nor U13002 (N_13002,N_11195,N_10529);
nor U13003 (N_13003,N_10058,N_11648);
nand U13004 (N_13004,N_8733,N_11751);
or U13005 (N_13005,N_10559,N_10573);
or U13006 (N_13006,N_8474,N_10835);
nand U13007 (N_13007,N_8274,N_11182);
nand U13008 (N_13008,N_8685,N_10681);
or U13009 (N_13009,N_8235,N_10595);
nor U13010 (N_13010,N_8121,N_11724);
or U13011 (N_13011,N_8998,N_11424);
and U13012 (N_13012,N_9422,N_10906);
nand U13013 (N_13013,N_11004,N_9782);
and U13014 (N_13014,N_11349,N_11639);
or U13015 (N_13015,N_10404,N_10666);
nand U13016 (N_13016,N_9163,N_8969);
or U13017 (N_13017,N_9532,N_10414);
and U13018 (N_13018,N_11064,N_9923);
and U13019 (N_13019,N_9568,N_10827);
or U13020 (N_13020,N_10283,N_8450);
and U13021 (N_13021,N_8262,N_9368);
and U13022 (N_13022,N_10172,N_11138);
nor U13023 (N_13023,N_9515,N_11037);
and U13024 (N_13024,N_11865,N_9717);
nand U13025 (N_13025,N_9789,N_11748);
or U13026 (N_13026,N_9803,N_8322);
nand U13027 (N_13027,N_10416,N_8229);
or U13028 (N_13028,N_9489,N_9351);
nor U13029 (N_13029,N_8928,N_8439);
nand U13030 (N_13030,N_9125,N_10284);
and U13031 (N_13031,N_9558,N_10576);
or U13032 (N_13032,N_8056,N_9375);
nand U13033 (N_13033,N_10433,N_9601);
nand U13034 (N_13034,N_10344,N_10543);
and U13035 (N_13035,N_10135,N_10265);
nand U13036 (N_13036,N_8961,N_10187);
and U13037 (N_13037,N_9863,N_8457);
or U13038 (N_13038,N_8244,N_8519);
nand U13039 (N_13039,N_10074,N_10765);
nand U13040 (N_13040,N_11521,N_10887);
nand U13041 (N_13041,N_11008,N_11320);
and U13042 (N_13042,N_11348,N_8119);
and U13043 (N_13043,N_11974,N_10088);
or U13044 (N_13044,N_10020,N_11045);
nor U13045 (N_13045,N_8165,N_11773);
and U13046 (N_13046,N_11788,N_8730);
nor U13047 (N_13047,N_8377,N_9933);
nand U13048 (N_13048,N_8403,N_10845);
and U13049 (N_13049,N_11200,N_10202);
and U13050 (N_13050,N_8779,N_10679);
and U13051 (N_13051,N_8579,N_10395);
or U13052 (N_13052,N_11124,N_11827);
or U13053 (N_13053,N_9130,N_9203);
nand U13054 (N_13054,N_11052,N_8444);
and U13055 (N_13055,N_8600,N_11811);
and U13056 (N_13056,N_10725,N_9051);
and U13057 (N_13057,N_10031,N_10229);
nand U13058 (N_13058,N_9817,N_9317);
or U13059 (N_13059,N_8633,N_11314);
or U13060 (N_13060,N_9026,N_11561);
nor U13061 (N_13061,N_10368,N_10664);
nor U13062 (N_13062,N_11796,N_8728);
and U13063 (N_13063,N_8645,N_8077);
nand U13064 (N_13064,N_11692,N_8043);
nand U13065 (N_13065,N_11685,N_8015);
nor U13066 (N_13066,N_11356,N_11352);
and U13067 (N_13067,N_10638,N_9458);
and U13068 (N_13068,N_11190,N_10299);
or U13069 (N_13069,N_9055,N_9369);
and U13070 (N_13070,N_9261,N_11175);
nand U13071 (N_13071,N_11680,N_8158);
and U13072 (N_13072,N_9288,N_11434);
or U13073 (N_13073,N_11494,N_11058);
nand U13074 (N_13074,N_11636,N_11594);
or U13075 (N_13075,N_8584,N_10912);
nor U13076 (N_13076,N_10877,N_8704);
nor U13077 (N_13077,N_8266,N_9683);
nor U13078 (N_13078,N_8344,N_11953);
and U13079 (N_13079,N_8469,N_9577);
nand U13080 (N_13080,N_10071,N_11719);
and U13081 (N_13081,N_9414,N_10314);
nor U13082 (N_13082,N_9389,N_9463);
nand U13083 (N_13083,N_8482,N_11248);
and U13084 (N_13084,N_8446,N_11471);
and U13085 (N_13085,N_11590,N_11885);
nand U13086 (N_13086,N_8713,N_10300);
and U13087 (N_13087,N_10249,N_8722);
nor U13088 (N_13088,N_9013,N_11193);
nand U13089 (N_13089,N_10274,N_11452);
nor U13090 (N_13090,N_11876,N_8085);
nor U13091 (N_13091,N_11799,N_11289);
or U13092 (N_13092,N_9149,N_9386);
and U13093 (N_13093,N_10700,N_9981);
or U13094 (N_13094,N_9264,N_10792);
and U13095 (N_13095,N_9284,N_10245);
nor U13096 (N_13096,N_10909,N_11092);
nand U13097 (N_13097,N_9596,N_11889);
or U13098 (N_13098,N_9680,N_11664);
or U13099 (N_13099,N_10513,N_10668);
or U13100 (N_13100,N_8205,N_8978);
nand U13101 (N_13101,N_10682,N_8681);
nand U13102 (N_13102,N_11467,N_11907);
or U13103 (N_13103,N_10554,N_11580);
nor U13104 (N_13104,N_8172,N_9932);
nor U13105 (N_13105,N_10707,N_8596);
nand U13106 (N_13106,N_9390,N_8075);
and U13107 (N_13107,N_10250,N_11219);
nor U13108 (N_13108,N_8257,N_11367);
nand U13109 (N_13109,N_11130,N_8376);
nand U13110 (N_13110,N_8046,N_9112);
or U13111 (N_13111,N_11985,N_10277);
nor U13112 (N_13112,N_8538,N_9768);
nand U13113 (N_13113,N_9658,N_8549);
or U13114 (N_13114,N_8002,N_8407);
nor U13115 (N_13115,N_9744,N_11657);
or U13116 (N_13116,N_8305,N_9690);
and U13117 (N_13117,N_11186,N_11745);
xor U13118 (N_13118,N_11032,N_9788);
and U13119 (N_13119,N_8499,N_8250);
and U13120 (N_13120,N_10895,N_10434);
nand U13121 (N_13121,N_10633,N_11944);
and U13122 (N_13122,N_8412,N_9608);
and U13123 (N_13123,N_11618,N_9151);
and U13124 (N_13124,N_8788,N_11456);
nor U13125 (N_13125,N_11791,N_11444);
nand U13126 (N_13126,N_10137,N_9038);
and U13127 (N_13127,N_8315,N_9182);
nor U13128 (N_13128,N_9506,N_11432);
and U13129 (N_13129,N_9627,N_9533);
and U13130 (N_13130,N_9618,N_8225);
and U13131 (N_13131,N_9975,N_9915);
or U13132 (N_13132,N_9415,N_8350);
nand U13133 (N_13133,N_11404,N_11088);
or U13134 (N_13134,N_9938,N_10634);
nand U13135 (N_13135,N_11291,N_9113);
and U13136 (N_13136,N_11871,N_10505);
nor U13137 (N_13137,N_8860,N_9689);
nand U13138 (N_13138,N_8693,N_10824);
nand U13139 (N_13139,N_10281,N_8780);
nor U13140 (N_13140,N_10457,N_8153);
and U13141 (N_13141,N_8342,N_8991);
nor U13142 (N_13142,N_8878,N_10924);
nand U13143 (N_13143,N_11362,N_11267);
nor U13144 (N_13144,N_10011,N_8861);
or U13145 (N_13145,N_8957,N_8548);
and U13146 (N_13146,N_10708,N_8120);
nor U13147 (N_13147,N_10670,N_9550);
and U13148 (N_13148,N_10678,N_8694);
and U13149 (N_13149,N_11873,N_11835);
and U13150 (N_13150,N_10610,N_11928);
nand U13151 (N_13151,N_10732,N_9438);
or U13152 (N_13152,N_10858,N_8731);
or U13153 (N_13153,N_10004,N_10699);
or U13154 (N_13154,N_11364,N_11854);
nand U13155 (N_13155,N_11964,N_10372);
nand U13156 (N_13156,N_8984,N_8413);
or U13157 (N_13157,N_11495,N_8373);
and U13158 (N_13158,N_11632,N_10603);
and U13159 (N_13159,N_10430,N_9632);
and U13160 (N_13160,N_9174,N_8108);
or U13161 (N_13161,N_8989,N_8603);
nand U13162 (N_13162,N_8139,N_10185);
and U13163 (N_13163,N_8571,N_11113);
nand U13164 (N_13164,N_8051,N_10767);
nand U13165 (N_13165,N_11378,N_10954);
nand U13166 (N_13166,N_9900,N_11765);
or U13167 (N_13167,N_9253,N_9365);
and U13168 (N_13168,N_10537,N_11902);
and U13169 (N_13169,N_9758,N_11612);
and U13170 (N_13170,N_10028,N_10019);
or U13171 (N_13171,N_8550,N_10468);
or U13172 (N_13172,N_9393,N_9362);
or U13173 (N_13173,N_8891,N_11468);
nand U13174 (N_13174,N_9852,N_8705);
nand U13175 (N_13175,N_8668,N_10062);
or U13176 (N_13176,N_11568,N_11939);
nand U13177 (N_13177,N_11649,N_10354);
nor U13178 (N_13178,N_11202,N_10517);
nand U13179 (N_13179,N_9921,N_11458);
nor U13180 (N_13180,N_9306,N_11308);
nand U13181 (N_13181,N_9409,N_9228);
nor U13182 (N_13182,N_10722,N_10418);
nand U13183 (N_13183,N_9423,N_10956);
nand U13184 (N_13184,N_11727,N_11486);
nor U13185 (N_13185,N_10470,N_11642);
nor U13186 (N_13186,N_9025,N_11666);
and U13187 (N_13187,N_8965,N_8824);
and U13188 (N_13188,N_10046,N_9614);
or U13189 (N_13189,N_8518,N_10642);
or U13190 (N_13190,N_10889,N_10581);
nor U13191 (N_13191,N_10830,N_9310);
or U13192 (N_13192,N_10813,N_11677);
or U13193 (N_13193,N_9045,N_9831);
or U13194 (N_13194,N_11617,N_10966);
nor U13195 (N_13195,N_8735,N_11096);
and U13196 (N_13196,N_8636,N_11055);
or U13197 (N_13197,N_9536,N_8818);
nor U13198 (N_13198,N_10904,N_11460);
and U13199 (N_13199,N_10228,N_11357);
nand U13200 (N_13200,N_11053,N_10271);
or U13201 (N_13201,N_10524,N_9053);
or U13202 (N_13202,N_10473,N_8975);
or U13203 (N_13203,N_9712,N_11021);
nand U13204 (N_13204,N_10968,N_11160);
or U13205 (N_13205,N_10100,N_9254);
nor U13206 (N_13206,N_11943,N_8532);
nand U13207 (N_13207,N_8799,N_11300);
and U13208 (N_13208,N_9657,N_9955);
or U13209 (N_13209,N_8163,N_9767);
nor U13210 (N_13210,N_9629,N_9987);
nand U13211 (N_13211,N_10455,N_9859);
nand U13212 (N_13212,N_9059,N_10244);
and U13213 (N_13213,N_9464,N_11978);
nor U13214 (N_13214,N_8929,N_11646);
nand U13215 (N_13215,N_10971,N_8760);
or U13216 (N_13216,N_11183,N_9466);
or U13217 (N_13217,N_8525,N_8917);
nor U13218 (N_13218,N_9884,N_10880);
nand U13219 (N_13219,N_10203,N_10944);
nor U13220 (N_13220,N_9223,N_8737);
nand U13221 (N_13221,N_9066,N_10295);
nor U13222 (N_13222,N_9970,N_8911);
and U13223 (N_13223,N_10601,N_11714);
nand U13224 (N_13224,N_9022,N_11954);
and U13225 (N_13225,N_9258,N_8503);
and U13226 (N_13226,N_8299,N_11764);
or U13227 (N_13227,N_10013,N_11941);
xor U13228 (N_13228,N_10024,N_11725);
or U13229 (N_13229,N_10751,N_8887);
and U13230 (N_13230,N_11333,N_9316);
or U13231 (N_13231,N_10683,N_8484);
nor U13232 (N_13232,N_10159,N_11233);
nor U13233 (N_13233,N_8486,N_9116);
and U13234 (N_13234,N_11874,N_8896);
nor U13235 (N_13235,N_10503,N_9918);
nand U13236 (N_13236,N_11645,N_10849);
or U13237 (N_13237,N_8931,N_8145);
or U13238 (N_13238,N_10834,N_8527);
nand U13239 (N_13239,N_9634,N_8627);
or U13240 (N_13240,N_9398,N_8772);
xor U13241 (N_13241,N_8505,N_11750);
or U13242 (N_13242,N_8092,N_10541);
nand U13243 (N_13243,N_9304,N_8841);
nor U13244 (N_13244,N_11099,N_8101);
nor U13245 (N_13245,N_11679,N_9626);
nand U13246 (N_13246,N_8710,N_10212);
or U13247 (N_13247,N_11331,N_8764);
and U13248 (N_13248,N_8618,N_11073);
nand U13249 (N_13249,N_11652,N_10327);
nand U13250 (N_13250,N_10957,N_9147);
or U13251 (N_13251,N_8067,N_9095);
nand U13252 (N_13252,N_8638,N_8242);
nand U13253 (N_13253,N_9377,N_11520);
or U13254 (N_13254,N_8512,N_10989);
nor U13255 (N_13255,N_8395,N_8972);
nor U13256 (N_13256,N_9162,N_10823);
and U13257 (N_13257,N_9344,N_10820);
and U13258 (N_13258,N_11660,N_11009);
and U13259 (N_13259,N_11932,N_9236);
nor U13260 (N_13260,N_10304,N_10809);
nor U13261 (N_13261,N_10153,N_10986);
nor U13262 (N_13262,N_10855,N_9713);
nand U13263 (N_13263,N_9008,N_11507);
nand U13264 (N_13264,N_11534,N_11678);
nand U13265 (N_13265,N_11158,N_11990);
nor U13266 (N_13266,N_8939,N_8013);
and U13267 (N_13267,N_11633,N_10905);
or U13268 (N_13268,N_11218,N_9201);
nand U13269 (N_13269,N_10579,N_9814);
nand U13270 (N_13270,N_8672,N_11198);
nand U13271 (N_13271,N_9913,N_11769);
and U13272 (N_13272,N_9616,N_11733);
or U13273 (N_13273,N_10693,N_10406);
and U13274 (N_13274,N_11790,N_10401);
nor U13275 (N_13275,N_8178,N_8202);
nand U13276 (N_13276,N_8480,N_8566);
nand U13277 (N_13277,N_10144,N_9936);
or U13278 (N_13278,N_11216,N_8021);
nor U13279 (N_13279,N_9935,N_9952);
nor U13280 (N_13280,N_8193,N_8354);
and U13281 (N_13281,N_11326,N_11411);
and U13282 (N_13282,N_9133,N_11588);
nor U13283 (N_13283,N_10495,N_9972);
nor U13284 (N_13284,N_8669,N_10697);
nand U13285 (N_13285,N_9301,N_9332);
nor U13286 (N_13286,N_8025,N_9887);
and U13287 (N_13287,N_8251,N_11368);
nand U13288 (N_13288,N_10533,N_10360);
and U13289 (N_13289,N_8393,N_10997);
nand U13290 (N_13290,N_8729,N_11858);
and U13291 (N_13291,N_9793,N_9891);
and U13292 (N_13292,N_10351,N_10677);
and U13293 (N_13293,N_11914,N_10484);
nor U13294 (N_13294,N_10996,N_11868);
or U13295 (N_13295,N_10564,N_9492);
nor U13296 (N_13296,N_11080,N_8212);
nand U13297 (N_13297,N_9171,N_11414);
and U13298 (N_13298,N_9319,N_10738);
and U13299 (N_13299,N_11244,N_11100);
or U13300 (N_13300,N_9465,N_8112);
or U13301 (N_13301,N_10985,N_8903);
nor U13302 (N_13302,N_10425,N_9208);
nand U13303 (N_13303,N_11755,N_11388);
or U13304 (N_13304,N_8719,N_11732);
or U13305 (N_13305,N_11366,N_10743);
or U13306 (N_13306,N_9624,N_9846);
and U13307 (N_13307,N_11139,N_8341);
and U13308 (N_13308,N_10669,N_8368);
and U13309 (N_13309,N_10051,N_11111);
nor U13310 (N_13310,N_9901,N_10869);
and U13311 (N_13311,N_9229,N_9165);
and U13312 (N_13312,N_11163,N_10995);
nor U13313 (N_13313,N_8030,N_11134);
and U13314 (N_13314,N_9726,N_8372);
or U13315 (N_13315,N_11571,N_9739);
and U13316 (N_13316,N_8617,N_10625);
or U13317 (N_13317,N_9106,N_10336);
or U13318 (N_13318,N_10721,N_11459);
or U13319 (N_13319,N_9298,N_9695);
nor U13320 (N_13320,N_9435,N_11443);
nand U13321 (N_13321,N_11022,N_11723);
nor U13322 (N_13322,N_11381,N_11598);
nand U13323 (N_13323,N_8545,N_9760);
or U13324 (N_13324,N_9408,N_11959);
nand U13325 (N_13325,N_11526,N_11433);
nor U13326 (N_13326,N_11273,N_8176);
or U13327 (N_13327,N_11899,N_10936);
or U13328 (N_13328,N_9637,N_9518);
nand U13329 (N_13329,N_9754,N_11995);
or U13330 (N_13330,N_10437,N_8535);
nor U13331 (N_13331,N_11157,N_9455);
nor U13332 (N_13332,N_10875,N_11492);
and U13333 (N_13333,N_10436,N_8578);
nand U13334 (N_13334,N_10803,N_8599);
nand U13335 (N_13335,N_9196,N_8750);
or U13336 (N_13336,N_8662,N_10734);
nand U13337 (N_13337,N_10982,N_11319);
or U13338 (N_13338,N_10627,N_9286);
nand U13339 (N_13339,N_8333,N_8233);
and U13340 (N_13340,N_11173,N_9204);
or U13341 (N_13341,N_10611,N_8003);
or U13342 (N_13342,N_10233,N_11162);
and U13343 (N_13343,N_9232,N_9100);
nand U13344 (N_13344,N_8692,N_9325);
and U13345 (N_13345,N_8369,N_11137);
or U13346 (N_13346,N_11737,N_8236);
or U13347 (N_13347,N_10488,N_11533);
or U13348 (N_13348,N_8910,N_9283);
and U13349 (N_13349,N_9848,N_9950);
and U13350 (N_13350,N_11591,N_8456);
or U13351 (N_13351,N_8587,N_11235);
and U13352 (N_13352,N_9469,N_11572);
and U13353 (N_13353,N_9985,N_8272);
or U13354 (N_13354,N_11479,N_11059);
nor U13355 (N_13355,N_9024,N_11857);
and U13356 (N_13356,N_10544,N_10236);
or U13357 (N_13357,N_10894,N_10021);
or U13358 (N_13358,N_11794,N_10694);
nand U13359 (N_13359,N_11180,N_8585);
xnor U13360 (N_13360,N_8099,N_11396);
nor U13361 (N_13361,N_11271,N_9870);
and U13362 (N_13362,N_10805,N_10804);
or U13363 (N_13363,N_11370,N_8094);
nand U13364 (N_13364,N_11935,N_10015);
nand U13365 (N_13365,N_9671,N_8805);
nor U13366 (N_13366,N_10597,N_8437);
and U13367 (N_13367,N_8687,N_11282);
nand U13368 (N_13368,N_11631,N_9006);
nand U13369 (N_13369,N_9516,N_10948);
nand U13370 (N_13370,N_9478,N_10512);
nand U13371 (N_13371,N_8416,N_8732);
or U13372 (N_13372,N_10359,N_10205);
and U13373 (N_13373,N_8286,N_11237);
nand U13374 (N_13374,N_9983,N_9345);
and U13375 (N_13375,N_10929,N_8398);
and U13376 (N_13376,N_9963,N_11011);
or U13377 (N_13377,N_9639,N_9191);
or U13378 (N_13378,N_10923,N_8859);
or U13379 (N_13379,N_10522,N_11252);
nand U13380 (N_13380,N_9213,N_9496);
nor U13381 (N_13381,N_11475,N_10290);
nand U13382 (N_13382,N_10967,N_9643);
nand U13383 (N_13383,N_10817,N_9652);
nor U13384 (N_13384,N_10115,N_9885);
nor U13385 (N_13385,N_11144,N_9729);
or U13386 (N_13386,N_10674,N_11238);
nand U13387 (N_13387,N_8992,N_10198);
or U13388 (N_13388,N_9893,N_8431);
nor U13389 (N_13389,N_11809,N_10231);
and U13390 (N_13390,N_10663,N_10085);
nand U13391 (N_13391,N_9522,N_8267);
nand U13392 (N_13392,N_9827,N_10928);
and U13393 (N_13393,N_10332,N_8530);
or U13394 (N_13394,N_8208,N_11845);
and U13395 (N_13395,N_8509,N_9574);
nor U13396 (N_13396,N_8111,N_11405);
and U13397 (N_13397,N_11783,N_11659);
nand U13398 (N_13398,N_8880,N_10509);
and U13399 (N_13399,N_11294,N_8454);
nand U13400 (N_13400,N_9257,N_11687);
xor U13401 (N_13401,N_11846,N_9873);
and U13402 (N_13402,N_9127,N_11152);
nand U13403 (N_13403,N_11903,N_9677);
or U13404 (N_13404,N_8935,N_9370);
nor U13405 (N_13405,N_10842,N_11025);
nand U13406 (N_13406,N_10431,N_11442);
nand U13407 (N_13407,N_8302,N_8232);
or U13408 (N_13408,N_8716,N_10079);
nor U13409 (N_13409,N_8493,N_9956);
nor U13410 (N_13410,N_11023,N_8269);
and U13411 (N_13411,N_9785,N_10035);
xor U13412 (N_13412,N_8659,N_8280);
nor U13413 (N_13413,N_11449,N_10785);
nand U13414 (N_13414,N_10268,N_9638);
nand U13415 (N_13415,N_9061,N_9131);
nor U13416 (N_13416,N_8222,N_10279);
nand U13417 (N_13417,N_9205,N_10293);
nor U13418 (N_13418,N_10273,N_8848);
nand U13419 (N_13419,N_9828,N_10435);
nor U13420 (N_13420,N_11603,N_11587);
nor U13421 (N_13421,N_10288,N_9566);
nand U13422 (N_13422,N_10690,N_11403);
or U13423 (N_13423,N_10176,N_8563);
nor U13424 (N_13424,N_11753,N_9300);
and U13425 (N_13425,N_8093,N_8949);
and U13426 (N_13426,N_8946,N_9451);
nor U13427 (N_13427,N_8116,N_8427);
nand U13428 (N_13428,N_8885,N_8110);
nor U13429 (N_13429,N_9453,N_11189);
nand U13430 (N_13430,N_11483,N_8980);
nand U13431 (N_13431,N_10131,N_9364);
or U13432 (N_13432,N_9781,N_8807);
nand U13433 (N_13433,N_10432,N_9033);
nor U13434 (N_13434,N_8922,N_11030);
nor U13435 (N_13435,N_9806,N_8573);
nor U13436 (N_13436,N_10616,N_8320);
nand U13437 (N_13437,N_11607,N_10704);
or U13438 (N_13438,N_11223,N_11387);
nor U13439 (N_13439,N_8996,N_10296);
nand U13440 (N_13440,N_9207,N_11169);
nor U13441 (N_13441,N_10101,N_9437);
or U13442 (N_13442,N_9037,N_11087);
and U13443 (N_13443,N_10959,N_8622);
nor U13444 (N_13444,N_11210,N_11654);
and U13445 (N_13445,N_8259,N_8740);
and U13446 (N_13446,N_9404,N_11054);
nand U13447 (N_13447,N_10687,N_10121);
nor U13448 (N_13448,N_8109,N_8909);
nand U13449 (N_13449,N_11407,N_10310);
or U13450 (N_13450,N_11264,N_10507);
or U13451 (N_13451,N_11938,N_8804);
or U13452 (N_13452,N_9663,N_11586);
or U13453 (N_13453,N_9017,N_11658);
nand U13454 (N_13454,N_10766,N_11531);
or U13455 (N_13455,N_9591,N_10126);
or U13456 (N_13456,N_11529,N_11676);
or U13457 (N_13457,N_10617,N_11803);
or U13458 (N_13458,N_10979,N_8562);
nand U13459 (N_13459,N_8577,N_11993);
or U13460 (N_13460,N_9707,N_8045);
nor U13461 (N_13461,N_10569,N_8610);
nor U13462 (N_13462,N_8543,N_10689);
nor U13463 (N_13463,N_11539,N_10508);
nand U13464 (N_13464,N_10421,N_11012);
nand U13465 (N_13465,N_8608,N_10214);
nor U13466 (N_13466,N_8459,N_10197);
or U13467 (N_13467,N_11068,N_10745);
nand U13468 (N_13468,N_10320,N_8466);
and U13469 (N_13469,N_9441,N_11201);
or U13470 (N_13470,N_11946,N_9544);
nand U13471 (N_13471,N_9698,N_9179);
and U13472 (N_13472,N_10739,N_10289);
or U13473 (N_13473,N_8089,N_9019);
and U13474 (N_13474,N_10257,N_8281);
nor U13475 (N_13475,N_8881,N_10545);
nor U13476 (N_13476,N_8052,N_8078);
and U13477 (N_13477,N_11497,N_8130);
nand U13478 (N_13478,N_11787,N_11095);
nand U13479 (N_13479,N_8565,N_11295);
and U13480 (N_13480,N_8330,N_10459);
nand U13481 (N_13481,N_10124,N_9612);
or U13482 (N_13482,N_9807,N_10983);
and U13483 (N_13483,N_8781,N_10347);
nand U13484 (N_13484,N_9507,N_9751);
or U13485 (N_13485,N_11669,N_9079);
nor U13486 (N_13486,N_11754,N_11318);
and U13487 (N_13487,N_11231,N_10407);
nand U13488 (N_13488,N_9605,N_9855);
and U13489 (N_13489,N_10528,N_8410);
nor U13490 (N_13490,N_11781,N_8148);
nor U13491 (N_13491,N_9256,N_11560);
nand U13492 (N_13492,N_9314,N_8473);
or U13493 (N_13493,N_9578,N_11911);
and U13494 (N_13494,N_10018,N_10598);
nor U13495 (N_13495,N_11690,N_8366);
nor U13496 (N_13496,N_10599,N_9307);
nand U13497 (N_13497,N_11915,N_9509);
nor U13498 (N_13498,N_10950,N_10173);
or U13499 (N_13499,N_10864,N_10755);
nand U13500 (N_13500,N_10110,N_8987);
and U13501 (N_13501,N_11780,N_11275);
nand U13502 (N_13502,N_10748,N_9323);
and U13503 (N_13503,N_8352,N_10391);
nand U13504 (N_13504,N_9691,N_11805);
nor U13505 (N_13505,N_9559,N_8776);
or U13506 (N_13506,N_8967,N_11440);
nor U13507 (N_13507,N_8260,N_8324);
nand U13508 (N_13508,N_8397,N_8699);
nor U13509 (N_13509,N_10090,N_11638);
or U13510 (N_13510,N_10260,N_8049);
nor U13511 (N_13511,N_8652,N_8136);
or U13512 (N_13512,N_9259,N_9328);
or U13513 (N_13513,N_11457,N_8297);
and U13514 (N_13514,N_8219,N_9052);
or U13515 (N_13515,N_9818,N_9620);
or U13516 (N_13516,N_11517,N_9057);
nand U13517 (N_13517,N_10963,N_8312);
or U13518 (N_13518,N_8237,N_9701);
nand U13519 (N_13519,N_8754,N_10828);
or U13520 (N_13520,N_11344,N_8586);
nor U13521 (N_13521,N_10607,N_9854);
nor U13522 (N_13522,N_11425,N_9687);
or U13523 (N_13523,N_10718,N_11347);
nand U13524 (N_13524,N_8100,N_11842);
or U13525 (N_13525,N_8999,N_8380);
or U13526 (N_13526,N_11728,N_11523);
nor U13527 (N_13527,N_11761,N_8465);
and U13528 (N_13528,N_10806,N_8533);
and U13529 (N_13529,N_9135,N_9160);
and U13530 (N_13530,N_8990,N_9989);
nand U13531 (N_13531,N_8058,N_8501);
and U13532 (N_13532,N_10527,N_10602);
and U13533 (N_13533,N_9552,N_8239);
or U13534 (N_13534,N_8660,N_11254);
and U13535 (N_13535,N_10174,N_10443);
nor U13536 (N_13536,N_8822,N_8811);
and U13537 (N_13537,N_10155,N_9221);
nor U13538 (N_13538,N_9103,N_10068);
nor U13539 (N_13539,N_8035,N_10383);
or U13540 (N_13540,N_9586,N_8479);
or U13541 (N_13541,N_11962,N_9303);
or U13542 (N_13542,N_11376,N_11164);
nor U13543 (N_13543,N_8904,N_10270);
or U13544 (N_13544,N_9962,N_9686);
and U13545 (N_13545,N_9101,N_9338);
or U13546 (N_13546,N_10030,N_10063);
and U13547 (N_13547,N_9811,N_10235);
or U13548 (N_13548,N_11090,N_11929);
nor U13549 (N_13549,N_11569,N_8496);
and U13550 (N_13550,N_9665,N_10298);
and U13551 (N_13551,N_11166,N_8231);
nor U13552 (N_13552,N_11269,N_9027);
or U13553 (N_13553,N_9906,N_10211);
nand U13554 (N_13554,N_9200,N_11284);
or U13555 (N_13555,N_10729,N_9978);
or U13556 (N_13556,N_9606,N_9114);
or U13557 (N_13557,N_8748,N_10854);
or U13558 (N_13558,N_9860,N_11101);
or U13559 (N_13559,N_9297,N_9502);
or U13560 (N_13560,N_10990,N_8568);
nor U13561 (N_13561,N_11496,N_11742);
or U13562 (N_13562,N_8028,N_10204);
and U13563 (N_13563,N_8316,N_8688);
or U13564 (N_13564,N_9449,N_11759);
and U13565 (N_13565,N_10927,N_9209);
or U13566 (N_13566,N_9445,N_11417);
nor U13567 (N_13567,N_8850,N_10848);
or U13568 (N_13568,N_8606,N_10630);
and U13569 (N_13569,N_9777,N_11017);
nor U13570 (N_13570,N_8080,N_8714);
nand U13571 (N_13571,N_8164,N_10756);
nor U13572 (N_13572,N_10902,N_10570);
nor U13573 (N_13573,N_11363,N_8004);
and U13574 (N_13574,N_11906,N_9428);
nand U13575 (N_13575,N_10980,N_11020);
and U13576 (N_13576,N_9238,N_9600);
and U13577 (N_13577,N_9562,N_9018);
and U13578 (N_13578,N_10097,N_9193);
or U13579 (N_13579,N_10937,N_11454);
or U13580 (N_13580,N_9255,N_11379);
or U13581 (N_13581,N_10358,N_11744);
nor U13582 (N_13582,N_8695,N_9823);
nand U13583 (N_13583,N_9694,N_8385);
nor U13584 (N_13584,N_10504,N_9623);
or U13585 (N_13585,N_8974,N_9672);
and U13586 (N_13586,N_8277,N_10083);
xor U13587 (N_13587,N_9115,N_8671);
nand U13588 (N_13588,N_10337,N_11898);
nand U13589 (N_13589,N_9774,N_11445);
and U13590 (N_13590,N_10698,N_11983);
nor U13591 (N_13591,N_9243,N_9572);
or U13592 (N_13592,N_11208,N_11339);
nor U13593 (N_13593,N_11668,N_9979);
nand U13594 (N_13594,N_8063,N_9866);
nor U13595 (N_13595,N_11717,N_9031);
nand U13596 (N_13596,N_11369,N_10123);
nand U13597 (N_13597,N_10158,N_9571);
nor U13598 (N_13598,N_9646,N_10223);
or U13599 (N_13599,N_8147,N_10735);
nor U13600 (N_13600,N_9520,N_10578);
nand U13601 (N_13601,N_9630,N_10515);
and U13602 (N_13602,N_10671,N_11247);
nor U13603 (N_13603,N_11847,N_9271);
and U13604 (N_13604,N_10826,N_10077);
nor U13605 (N_13605,N_11146,N_9189);
nand U13606 (N_13606,N_8985,N_11661);
and U13607 (N_13607,N_11757,N_9878);
nor U13608 (N_13608,N_10043,N_11782);
or U13609 (N_13609,N_8190,N_10768);
nand U13610 (N_13610,N_8348,N_8892);
and U13611 (N_13611,N_8477,N_9012);
or U13612 (N_13612,N_9274,N_11043);
nand U13613 (N_13613,N_8001,N_10392);
or U13614 (N_13614,N_8653,N_9705);
or U13615 (N_13615,N_11391,N_8952);
nor U13616 (N_13616,N_10039,N_9246);
and U13617 (N_13617,N_11462,N_11332);
and U13618 (N_13618,N_10466,N_10177);
or U13619 (N_13619,N_8464,N_11042);
nand U13620 (N_13620,N_8084,N_8328);
nand U13621 (N_13621,N_8196,N_9523);
nor U13622 (N_13622,N_8784,N_8925);
nand U13623 (N_13623,N_10453,N_9347);
nor U13624 (N_13624,N_8356,N_9830);
or U13625 (N_13625,N_10164,N_10227);
nand U13626 (N_13626,N_10917,N_10675);
or U13627 (N_13627,N_8198,N_9244);
and U13628 (N_13628,N_11119,N_11527);
xnor U13629 (N_13629,N_10082,N_11436);
and U13630 (N_13630,N_9699,N_8426);
and U13631 (N_13631,N_11775,N_11834);
and U13632 (N_13632,N_11427,N_8702);
nor U13633 (N_13633,N_9585,N_10921);
and U13634 (N_13634,N_9346,N_11705);
nand U13635 (N_13635,N_9484,N_8150);
nand U13636 (N_13636,N_8228,N_8071);
nand U13637 (N_13637,N_11307,N_9425);
nor U13638 (N_13638,N_9524,N_9361);
and U13639 (N_13639,N_9050,N_8500);
nor U13640 (N_13640,N_9945,N_9529);
nand U13641 (N_13641,N_10148,N_11397);
nor U13642 (N_13642,N_10357,N_8682);
and U13643 (N_13643,N_10759,N_11786);
nand U13644 (N_13644,N_10111,N_10790);
and U13645 (N_13645,N_10034,N_11136);
and U13646 (N_13646,N_10023,N_8156);
nor U13647 (N_13647,N_9076,N_8396);
nor U13648 (N_13648,N_8837,N_8098);
nand U13649 (N_13649,N_10836,N_8064);
nand U13650 (N_13650,N_8950,N_10542);
and U13651 (N_13651,N_11807,N_10356);
or U13652 (N_13652,N_11922,N_11278);
or U13653 (N_13653,N_9980,N_9420);
nor U13654 (N_13654,N_10220,N_9530);
nand U13655 (N_13655,N_8576,N_11236);
nand U13656 (N_13656,N_11465,N_8371);
nand U13657 (N_13657,N_11313,N_10549);
nor U13658 (N_13658,N_10791,N_8243);
or U13659 (N_13659,N_10814,N_10133);
and U13660 (N_13660,N_8708,N_11701);
or U13661 (N_13661,N_8778,N_9836);
nor U13662 (N_13662,N_10872,N_9927);
nor U13663 (N_13663,N_8061,N_11028);
and U13664 (N_13664,N_10472,N_11298);
nand U13665 (N_13665,N_9755,N_11887);
nand U13666 (N_13666,N_9810,N_11686);
nor U13667 (N_13667,N_9986,N_10122);
nor U13668 (N_13668,N_9490,N_11477);
or U13669 (N_13669,N_9468,N_9399);
or U13670 (N_13670,N_9548,N_9021);
or U13671 (N_13671,N_8026,N_8927);
nand U13672 (N_13672,N_9065,N_11019);
nor U13673 (N_13673,N_8409,N_8432);
or U13674 (N_13674,N_9709,N_11579);
nor U13675 (N_13675,N_9721,N_10592);
nor U13676 (N_13676,N_8292,N_9937);
and U13677 (N_13677,N_10017,N_8382);
or U13678 (N_13678,N_8448,N_10560);
and U13679 (N_13679,N_10092,N_11900);
nand U13680 (N_13680,N_11537,N_8540);
nor U13681 (N_13681,N_11266,N_9442);
nand U13682 (N_13682,N_10839,N_8605);
nand U13683 (N_13683,N_8319,N_9631);
nor U13684 (N_13684,N_8915,N_11354);
nand U13685 (N_13685,N_9176,N_11558);
nor U13686 (N_13686,N_8646,N_8790);
or U13687 (N_13687,N_11229,N_10984);
or U13688 (N_13688,N_8264,N_11131);
and U13689 (N_13689,N_11257,N_9943);
or U13690 (N_13690,N_10426,N_9941);
nand U13691 (N_13691,N_8090,N_8559);
or U13692 (N_13692,N_8698,N_10915);
or U13693 (N_13693,N_11297,N_10752);
nor U13694 (N_13694,N_9641,N_11406);
nand U13695 (N_13695,N_9996,N_11785);
nand U13696 (N_13696,N_10710,N_8706);
or U13697 (N_13697,N_8261,N_11525);
or U13698 (N_13698,N_11574,N_8839);
nand U13699 (N_13699,N_8792,N_8400);
nor U13700 (N_13700,N_10045,N_8794);
nand U13701 (N_13701,N_8907,N_9988);
nor U13702 (N_13702,N_11293,N_10753);
nor U13703 (N_13703,N_11016,N_11881);
and U13704 (N_13704,N_11606,N_11998);
nand U13705 (N_13705,N_8415,N_8082);
and U13706 (N_13706,N_8717,N_9971);
or U13707 (N_13707,N_8007,N_9879);
or U13708 (N_13708,N_8572,N_11982);
nor U13709 (N_13709,N_11651,N_11812);
nor U13710 (N_13710,N_11145,N_8777);
xnor U13711 (N_13711,N_9105,N_9504);
and U13712 (N_13712,N_8528,N_9419);
nor U13713 (N_13713,N_8200,N_8855);
and U13714 (N_13714,N_10661,N_10794);
nand U13715 (N_13715,N_9295,N_11036);
or U13716 (N_13716,N_10112,N_9397);
nor U13717 (N_13717,N_8414,N_10424);
nand U13718 (N_13718,N_10862,N_10002);
nor U13719 (N_13719,N_9153,N_8995);
nand U13720 (N_13720,N_10487,N_8803);
nand U13721 (N_13721,N_10315,N_10702);
nor U13722 (N_13722,N_9069,N_8936);
xor U13723 (N_13723,N_10871,N_11860);
nor U13724 (N_13724,N_10941,N_11500);
or U13725 (N_13725,N_11153,N_10475);
or U13726 (N_13726,N_9086,N_8831);
nor U13727 (N_13727,N_9719,N_8827);
nand U13728 (N_13728,N_9251,N_10769);
and U13729 (N_13729,N_9158,N_11867);
and U13730 (N_13730,N_11283,N_11263);
xnor U13731 (N_13731,N_11710,N_9880);
nand U13732 (N_13732,N_10439,N_9005);
nor U13733 (N_13733,N_9089,N_9998);
or U13734 (N_13734,N_10763,N_9968);
or U13735 (N_13735,N_10120,N_9808);
nand U13736 (N_13736,N_11977,N_10811);
nand U13737 (N_13737,N_10345,N_9383);
nor U13738 (N_13738,N_11832,N_8923);
nand U13739 (N_13739,N_9355,N_9582);
and U13740 (N_13740,N_11671,N_11798);
nand U13741 (N_13741,N_8594,N_8303);
nor U13742 (N_13742,N_8905,N_11549);
and U13743 (N_13743,N_8436,N_8034);
nand U13744 (N_13744,N_8182,N_11026);
or U13745 (N_13745,N_10087,N_10275);
or U13746 (N_13746,N_10452,N_10815);
and U13747 (N_13747,N_10179,N_9862);
nor U13748 (N_13748,N_10417,N_11838);
or U13749 (N_13749,N_10313,N_9175);
nor U13750 (N_13750,N_8812,N_9868);
nor U13751 (N_13751,N_9098,N_9897);
or U13752 (N_13752,N_11837,N_9594);
and U13753 (N_13753,N_8657,N_8712);
nand U13754 (N_13754,N_8254,N_9949);
nand U13755 (N_13755,N_8128,N_11005);
nor U13756 (N_13756,N_11704,N_8378);
or U13757 (N_13757,N_8271,N_8773);
xor U13758 (N_13758,N_10380,N_8102);
nand U13759 (N_13759,N_8059,N_11597);
nand U13760 (N_13760,N_11304,N_10319);
nand U13761 (N_13761,N_9794,N_9450);
nand U13762 (N_13762,N_9543,N_10749);
or U13763 (N_13763,N_9922,N_10162);
or U13764 (N_13764,N_10586,N_8011);
nand U13765 (N_13765,N_11774,N_9187);
or U13766 (N_13766,N_11562,N_10761);
nor U13767 (N_13767,N_8358,N_11738);
nor U13768 (N_13768,N_10829,N_8591);
and U13769 (N_13769,N_11665,N_8408);
or U13770 (N_13770,N_11800,N_11895);
nand U13771 (N_13771,N_11626,N_10801);
and U13772 (N_13772,N_9088,N_8047);
or U13773 (N_13773,N_9961,N_9743);
or U13774 (N_13774,N_9994,N_8151);
nor U13775 (N_13775,N_8654,N_9357);
and U13776 (N_13776,N_8854,N_11106);
nand U13777 (N_13777,N_8966,N_9845);
nor U13778 (N_13778,N_11967,N_10949);
or U13779 (N_13779,N_11535,N_9999);
nor U13780 (N_13780,N_8938,N_11908);
or U13781 (N_13781,N_10913,N_9070);
or U13782 (N_13782,N_10961,N_9173);
nor U13783 (N_13783,N_9579,N_8296);
nand U13784 (N_13784,N_11365,N_9796);
nor U13785 (N_13785,N_8042,N_8613);
nand U13786 (N_13786,N_11491,N_9720);
nor U13787 (N_13787,N_10224,N_10783);
nor U13788 (N_13788,N_11108,N_8561);
or U13789 (N_13789,N_11689,N_11553);
nand U13790 (N_13790,N_8134,N_11797);
or U13791 (N_13791,N_9908,N_9545);
nand U13792 (N_13792,N_9875,N_10428);
nor U13793 (N_13793,N_10117,N_8933);
nor U13794 (N_13794,N_11310,N_9327);
nand U13795 (N_13795,N_10831,N_10059);
and U13796 (N_13796,N_8554,N_10323);
nand U13797 (N_13797,N_9547,N_11466);
nand U13798 (N_13798,N_10925,N_8934);
and U13799 (N_13799,N_8031,N_11197);
or U13800 (N_13800,N_11472,N_11968);
or U13801 (N_13801,N_9218,N_8977);
and U13802 (N_13802,N_9849,N_8027);
and U13803 (N_13803,N_8674,N_8293);
and U13804 (N_13804,N_9391,N_9313);
or U13805 (N_13805,N_10091,N_11487);
and U13806 (N_13806,N_11306,N_10168);
and U13807 (N_13807,N_10516,N_9573);
nor U13808 (N_13808,N_9270,N_11246);
and U13809 (N_13809,N_10691,N_11398);
nand U13810 (N_13810,N_10935,N_9640);
or U13811 (N_13811,N_8701,N_9043);
and U13812 (N_13812,N_8889,N_9942);
nand U13813 (N_13813,N_10548,N_11559);
and U13814 (N_13814,N_8517,N_11498);
nand U13815 (N_13815,N_9824,N_10555);
nor U13816 (N_13816,N_10379,N_8696);
nor U13817 (N_13817,N_10230,N_10618);
or U13818 (N_13818,N_8916,N_9075);
and U13819 (N_13819,N_11400,N_10736);
or U13820 (N_13820,N_9289,N_11085);
and U13821 (N_13821,N_8362,N_9245);
or U13822 (N_13822,N_10646,N_10717);
and U13823 (N_13823,N_10798,N_10797);
or U13824 (N_13824,N_8883,N_11142);
and U13825 (N_13825,N_9882,N_8993);
and U13826 (N_13826,N_8207,N_9560);
nand U13827 (N_13827,N_8005,N_9662);
or U13828 (N_13828,N_8724,N_8284);
nand U13829 (N_13829,N_8574,N_10676);
nand U13830 (N_13830,N_8753,N_10973);
and U13831 (N_13831,N_9210,N_11987);
and U13832 (N_13832,N_10867,N_8886);
or U13833 (N_13833,N_10723,N_10496);
nor U13834 (N_13834,N_9320,N_9143);
nor U13835 (N_13835,N_8723,N_10306);
nor U13836 (N_13836,N_9521,N_8140);
nor U13837 (N_13837,N_10226,N_10779);
or U13838 (N_13838,N_10463,N_8335);
nor U13839 (N_13839,N_9178,N_9649);
and U13840 (N_13840,N_9421,N_9473);
nor U13841 (N_13841,N_11772,N_8762);
and U13842 (N_13842,N_9816,N_11767);
and U13843 (N_13843,N_10641,N_9137);
or U13844 (N_13844,N_8873,N_9129);
and U13845 (N_13845,N_10900,N_8897);
or U13846 (N_13846,N_8226,N_9746);
and U13847 (N_13847,N_11112,N_11048);
nand U13848 (N_13848,N_9081,N_8331);
xor U13849 (N_13849,N_9237,N_11063);
or U13850 (N_13850,N_8282,N_9216);
nor U13851 (N_13851,N_10403,N_8351);
and U13852 (N_13852,N_11156,N_10667);
and U13853 (N_13853,N_11031,N_9874);
nand U13854 (N_13854,N_9645,N_8039);
nor U13855 (N_13855,N_11653,N_8932);
or U13856 (N_13856,N_10762,N_8349);
nor U13857 (N_13857,N_11960,N_11447);
xor U13858 (N_13858,N_8253,N_10535);
nand U13859 (N_13859,N_8789,N_11698);
nand U13860 (N_13860,N_11784,N_10645);
or U13861 (N_13861,N_9330,N_8736);
or U13862 (N_13862,N_9367,N_9396);
nor U13863 (N_13863,N_11731,N_8053);
or U13864 (N_13864,N_10461,N_8438);
and U13865 (N_13865,N_11151,N_8126);
nor U13866 (N_13866,N_9333,N_10703);
nor U13867 (N_13867,N_11416,N_10102);
or U13868 (N_13868,N_8869,N_8644);
and U13869 (N_13869,N_9169,N_10643);
and U13870 (N_13870,N_9508,N_11094);
and U13871 (N_13871,N_8326,N_10741);
nor U13872 (N_13872,N_9426,N_8918);
or U13873 (N_13873,N_11793,N_11245);
or U13874 (N_13874,N_11841,N_9653);
nor U13875 (N_13875,N_8428,N_8347);
or U13876 (N_13876,N_11038,N_8526);
nor U13877 (N_13877,N_9010,N_9896);
nor U13878 (N_13878,N_11697,N_11933);
nor U13879 (N_13879,N_11281,N_10482);
or U13880 (N_13880,N_10492,N_11547);
xnor U13881 (N_13881,N_10684,N_11091);
and U13882 (N_13882,N_8186,N_8217);
nor U13883 (N_13883,N_11077,N_8180);
and U13884 (N_13884,N_9644,N_9172);
nand U13885 (N_13885,N_10943,N_8797);
nor U13886 (N_13886,N_10654,N_10325);
nand U13887 (N_13887,N_9907,N_11779);
nand U13888 (N_13888,N_9416,N_11221);
nand U13889 (N_13889,N_11241,N_8209);
nor U13890 (N_13890,N_8742,N_8336);
nor U13891 (N_13891,N_9240,N_11098);
or U13892 (N_13892,N_9822,N_9500);
nand U13893 (N_13893,N_9321,N_11768);
and U13894 (N_13894,N_8270,N_8370);
nor U13895 (N_13895,N_9227,N_8308);
nor U13896 (N_13896,N_8523,N_10234);
or U13897 (N_13897,N_11695,N_9580);
or U13898 (N_13898,N_11518,N_9177);
or U13899 (N_13899,N_8520,N_10715);
and U13900 (N_13900,N_9180,N_9452);
or U13901 (N_13901,N_11609,N_11013);
nor U13902 (N_13902,N_11385,N_8037);
or U13903 (N_13903,N_8592,N_10497);
or U13904 (N_13904,N_9436,N_9864);
and U13905 (N_13905,N_10575,N_8553);
and U13906 (N_13906,N_9471,N_11625);
nor U13907 (N_13907,N_10930,N_8795);
nor U13908 (N_13908,N_8986,N_10653);
nor U13909 (N_13909,N_9040,N_10066);
or U13910 (N_13910,N_9285,N_9354);
nand U13911 (N_13911,N_8379,N_9603);
nand U13912 (N_13912,N_8838,N_9931);
or U13913 (N_13913,N_9247,N_11997);
or U13914 (N_13914,N_10076,N_11884);
nand U13915 (N_13915,N_8386,N_10861);
nand U13916 (N_13916,N_10253,N_11199);
or U13917 (N_13917,N_10132,N_10381);
nor U13918 (N_13918,N_9800,N_11375);
and U13919 (N_13919,N_10067,N_9219);
nand U13920 (N_13920,N_8137,N_11083);
nand U13921 (N_13921,N_9920,N_11552);
nor U13922 (N_13922,N_9417,N_11592);
and U13923 (N_13923,N_11926,N_10161);
and U13924 (N_13924,N_8774,N_10444);
nand U13925 (N_13925,N_9960,N_9967);
nand U13926 (N_13926,N_9700,N_10680);
and U13927 (N_13927,N_10728,N_9331);
nor U13928 (N_13928,N_9185,N_9374);
and U13929 (N_13929,N_9914,N_10647);
nand U13930 (N_13930,N_9220,N_11165);
or U13931 (N_13931,N_10188,N_8689);
or U13932 (N_13932,N_11234,N_9617);
nand U13933 (N_13933,N_8132,N_9714);
nor U13934 (N_13934,N_11170,N_10557);
nand U13935 (N_13935,N_10778,N_11627);
or U13936 (N_13936,N_11428,N_11991);
or U13937 (N_13937,N_8718,N_8976);
or U13938 (N_13938,N_9250,N_9260);
or U13939 (N_13939,N_10746,N_10147);
and U13940 (N_13940,N_10103,N_8624);
nand U13941 (N_13941,N_8940,N_9157);
and U13942 (N_13942,N_8365,N_8798);
nand U13943 (N_13943,N_10254,N_9539);
nand U13944 (N_13944,N_8029,N_9016);
and U13945 (N_13945,N_9977,N_8019);
or U13946 (N_13946,N_9029,N_11611);
nor U13947 (N_13947,N_10165,N_8429);
or U13948 (N_13948,N_10567,N_11849);
or U13949 (N_13949,N_8433,N_11384);
or U13950 (N_13950,N_8598,N_10635);
nand U13951 (N_13951,N_8926,N_10073);
xor U13952 (N_13952,N_8756,N_11740);
nor U13953 (N_13953,N_8483,N_11971);
or U13954 (N_13954,N_11280,N_10857);
nor U13955 (N_13955,N_9159,N_10977);
nand U13956 (N_13956,N_10493,N_10181);
nor U13957 (N_13957,N_9495,N_10511);
or U13958 (N_13958,N_11886,N_10138);
or U13959 (N_13959,N_8018,N_8445);
and U13960 (N_13960,N_8161,N_8418);
and U13961 (N_13961,N_10280,N_9801);
or U13962 (N_13962,N_11463,N_10853);
nor U13963 (N_13963,N_9528,N_8821);
xor U13964 (N_13964,N_10464,N_10639);
and U13965 (N_13965,N_11913,N_9554);
and U13966 (N_13966,N_11133,N_11323);
nand U13967 (N_13967,N_10632,N_8791);
and U13968 (N_13968,N_8765,N_10614);
and U13969 (N_13969,N_9909,N_8524);
nand U13970 (N_13970,N_11963,N_8767);
and U13971 (N_13971,N_9847,N_8560);
nor U13972 (N_13972,N_10072,N_10156);
and U13973 (N_13973,N_8220,N_9233);
nand U13974 (N_13974,N_8364,N_10052);
and U13975 (N_13975,N_11006,N_8481);
or U13976 (N_13976,N_11188,N_9930);
nor U13977 (N_13977,N_8405,N_8602);
nor U13978 (N_13978,N_9944,N_10219);
or U13979 (N_13979,N_10006,N_9569);
and U13980 (N_13980,N_11956,N_11482);
and U13981 (N_13981,N_10934,N_11630);
and U13982 (N_13982,N_9982,N_10307);
or U13983 (N_13983,N_10649,N_8081);
and U13984 (N_13984,N_10041,N_9761);
and U13985 (N_13985,N_9576,N_9184);
nand U13986 (N_13986,N_9898,N_9249);
or U13987 (N_13987,N_10053,N_9664);
nor U13988 (N_13988,N_11488,N_10644);
nor U13989 (N_13989,N_10009,N_10001);
and U13990 (N_13990,N_10999,N_8720);
or U13991 (N_13991,N_9123,N_9144);
nor U13992 (N_13992,N_11979,N_8930);
and U13993 (N_13993,N_11808,N_8629);
and U13994 (N_13994,N_11392,N_10141);
and U13995 (N_13995,N_11859,N_10863);
nand U13996 (N_13996,N_11074,N_9872);
or U13997 (N_13997,N_9063,N_8959);
or U13998 (N_13998,N_9561,N_10918);
nand U13999 (N_13999,N_11878,N_8683);
nand U14000 (N_14000,N_9655,N_9559);
and U14001 (N_14001,N_10174,N_10623);
or U14002 (N_14002,N_8332,N_11729);
or U14003 (N_14003,N_11480,N_8110);
nor U14004 (N_14004,N_10531,N_10797);
and U14005 (N_14005,N_9066,N_8698);
and U14006 (N_14006,N_11929,N_8147);
nand U14007 (N_14007,N_11648,N_10849);
xnor U14008 (N_14008,N_11057,N_11323);
or U14009 (N_14009,N_9607,N_11222);
and U14010 (N_14010,N_10679,N_9837);
nor U14011 (N_14011,N_8608,N_8009);
nand U14012 (N_14012,N_9692,N_10933);
or U14013 (N_14013,N_11369,N_11631);
and U14014 (N_14014,N_9926,N_9249);
or U14015 (N_14015,N_10875,N_10967);
nand U14016 (N_14016,N_11614,N_9860);
and U14017 (N_14017,N_9611,N_11958);
nand U14018 (N_14018,N_8071,N_11662);
nor U14019 (N_14019,N_11213,N_8638);
nor U14020 (N_14020,N_10279,N_11278);
and U14021 (N_14021,N_11914,N_9140);
or U14022 (N_14022,N_10384,N_8845);
and U14023 (N_14023,N_10552,N_9089);
nand U14024 (N_14024,N_11620,N_9448);
nor U14025 (N_14025,N_9590,N_9883);
nand U14026 (N_14026,N_10635,N_10541);
and U14027 (N_14027,N_8208,N_9508);
nand U14028 (N_14028,N_9580,N_9768);
and U14029 (N_14029,N_8044,N_11823);
nor U14030 (N_14030,N_10699,N_11495);
nor U14031 (N_14031,N_9119,N_11987);
and U14032 (N_14032,N_10251,N_10490);
nand U14033 (N_14033,N_11750,N_11557);
nor U14034 (N_14034,N_8184,N_11732);
and U14035 (N_14035,N_11373,N_11478);
or U14036 (N_14036,N_8941,N_11251);
or U14037 (N_14037,N_10189,N_9457);
nor U14038 (N_14038,N_9404,N_11093);
nand U14039 (N_14039,N_9908,N_9609);
and U14040 (N_14040,N_11653,N_8754);
nor U14041 (N_14041,N_11035,N_11581);
nor U14042 (N_14042,N_9208,N_11990);
or U14043 (N_14043,N_11682,N_11925);
or U14044 (N_14044,N_11500,N_11727);
nand U14045 (N_14045,N_8152,N_8041);
and U14046 (N_14046,N_11053,N_10992);
nand U14047 (N_14047,N_8321,N_10820);
nor U14048 (N_14048,N_10053,N_8829);
and U14049 (N_14049,N_10185,N_11844);
or U14050 (N_14050,N_8426,N_8889);
or U14051 (N_14051,N_10263,N_9743);
nor U14052 (N_14052,N_10149,N_11387);
or U14053 (N_14053,N_11725,N_9759);
nand U14054 (N_14054,N_8081,N_10180);
and U14055 (N_14055,N_10293,N_9100);
or U14056 (N_14056,N_11817,N_10496);
nor U14057 (N_14057,N_9109,N_10809);
nand U14058 (N_14058,N_9865,N_9303);
nor U14059 (N_14059,N_8254,N_11252);
or U14060 (N_14060,N_8849,N_11499);
nand U14061 (N_14061,N_11258,N_10376);
nor U14062 (N_14062,N_8249,N_10081);
nand U14063 (N_14063,N_9566,N_8968);
and U14064 (N_14064,N_8658,N_9912);
and U14065 (N_14065,N_9340,N_10533);
and U14066 (N_14066,N_10217,N_9815);
nand U14067 (N_14067,N_9248,N_10421);
nand U14068 (N_14068,N_11521,N_9900);
and U14069 (N_14069,N_9064,N_8049);
nor U14070 (N_14070,N_10286,N_9458);
and U14071 (N_14071,N_9789,N_10165);
or U14072 (N_14072,N_8394,N_11286);
nor U14073 (N_14073,N_11118,N_9330);
nor U14074 (N_14074,N_11598,N_9395);
nor U14075 (N_14075,N_10207,N_11350);
or U14076 (N_14076,N_9692,N_9452);
and U14077 (N_14077,N_8984,N_11091);
or U14078 (N_14078,N_9993,N_11489);
or U14079 (N_14079,N_10381,N_11947);
nor U14080 (N_14080,N_8008,N_8245);
nand U14081 (N_14081,N_8221,N_10918);
nor U14082 (N_14082,N_10339,N_11022);
nor U14083 (N_14083,N_10168,N_10480);
nand U14084 (N_14084,N_10953,N_10015);
nor U14085 (N_14085,N_11828,N_9041);
or U14086 (N_14086,N_9890,N_8846);
nand U14087 (N_14087,N_11217,N_9114);
nand U14088 (N_14088,N_11106,N_9979);
nand U14089 (N_14089,N_10049,N_8529);
nor U14090 (N_14090,N_9418,N_10824);
nand U14091 (N_14091,N_11630,N_10358);
nand U14092 (N_14092,N_11389,N_8784);
nor U14093 (N_14093,N_9025,N_8454);
or U14094 (N_14094,N_9694,N_11751);
and U14095 (N_14095,N_8294,N_10664);
and U14096 (N_14096,N_9221,N_11492);
and U14097 (N_14097,N_8603,N_8261);
and U14098 (N_14098,N_10546,N_11280);
or U14099 (N_14099,N_11393,N_8582);
nor U14100 (N_14100,N_8979,N_9276);
or U14101 (N_14101,N_11054,N_9005);
or U14102 (N_14102,N_11293,N_9338);
nand U14103 (N_14103,N_10212,N_8070);
or U14104 (N_14104,N_10899,N_9526);
nand U14105 (N_14105,N_11772,N_9083);
nand U14106 (N_14106,N_11468,N_9730);
and U14107 (N_14107,N_10821,N_8841);
or U14108 (N_14108,N_10401,N_8567);
or U14109 (N_14109,N_11522,N_8937);
and U14110 (N_14110,N_11127,N_9288);
nand U14111 (N_14111,N_10058,N_9836);
nor U14112 (N_14112,N_11453,N_11572);
nor U14113 (N_14113,N_11629,N_9631);
and U14114 (N_14114,N_9522,N_11525);
nand U14115 (N_14115,N_9355,N_9947);
and U14116 (N_14116,N_10811,N_10127);
or U14117 (N_14117,N_11605,N_8235);
nand U14118 (N_14118,N_11938,N_10034);
nor U14119 (N_14119,N_9214,N_11312);
and U14120 (N_14120,N_11256,N_9395);
and U14121 (N_14121,N_9656,N_11794);
and U14122 (N_14122,N_8236,N_10280);
or U14123 (N_14123,N_9659,N_9488);
or U14124 (N_14124,N_9831,N_11767);
nor U14125 (N_14125,N_9329,N_8809);
nor U14126 (N_14126,N_9144,N_11995);
nor U14127 (N_14127,N_9174,N_10224);
and U14128 (N_14128,N_9105,N_8603);
or U14129 (N_14129,N_11702,N_8174);
nand U14130 (N_14130,N_11835,N_10287);
and U14131 (N_14131,N_11617,N_8282);
nor U14132 (N_14132,N_8805,N_10724);
nand U14133 (N_14133,N_8024,N_8300);
and U14134 (N_14134,N_10142,N_9998);
and U14135 (N_14135,N_8158,N_9266);
nand U14136 (N_14136,N_11495,N_8999);
nand U14137 (N_14137,N_11174,N_8235);
or U14138 (N_14138,N_9484,N_8946);
nor U14139 (N_14139,N_11674,N_8732);
nor U14140 (N_14140,N_11475,N_11159);
or U14141 (N_14141,N_10012,N_11614);
nor U14142 (N_14142,N_9867,N_8099);
or U14143 (N_14143,N_11746,N_9703);
xor U14144 (N_14144,N_11070,N_8449);
and U14145 (N_14145,N_8442,N_10707);
nand U14146 (N_14146,N_9295,N_8167);
or U14147 (N_14147,N_11738,N_8269);
or U14148 (N_14148,N_8836,N_8432);
nand U14149 (N_14149,N_10531,N_11563);
or U14150 (N_14150,N_11545,N_8138);
nor U14151 (N_14151,N_11897,N_9079);
nor U14152 (N_14152,N_11346,N_8706);
nand U14153 (N_14153,N_8905,N_10131);
and U14154 (N_14154,N_11995,N_11667);
nor U14155 (N_14155,N_10244,N_9665);
nor U14156 (N_14156,N_10566,N_8417);
nand U14157 (N_14157,N_9101,N_11596);
nand U14158 (N_14158,N_9571,N_9434);
nand U14159 (N_14159,N_8778,N_9029);
and U14160 (N_14160,N_10064,N_11851);
and U14161 (N_14161,N_10748,N_11509);
and U14162 (N_14162,N_9276,N_8197);
or U14163 (N_14163,N_11813,N_9044);
or U14164 (N_14164,N_10727,N_8496);
nor U14165 (N_14165,N_8980,N_8405);
and U14166 (N_14166,N_10844,N_11190);
nor U14167 (N_14167,N_11392,N_9810);
nand U14168 (N_14168,N_10518,N_11433);
nand U14169 (N_14169,N_10421,N_8050);
nor U14170 (N_14170,N_11908,N_9155);
or U14171 (N_14171,N_8412,N_8226);
and U14172 (N_14172,N_11949,N_10590);
or U14173 (N_14173,N_11962,N_11852);
and U14174 (N_14174,N_9561,N_9484);
nor U14175 (N_14175,N_10915,N_8502);
nand U14176 (N_14176,N_11591,N_10346);
nor U14177 (N_14177,N_8919,N_9927);
or U14178 (N_14178,N_11342,N_10916);
nor U14179 (N_14179,N_10917,N_11863);
nor U14180 (N_14180,N_10399,N_9772);
or U14181 (N_14181,N_9689,N_9147);
and U14182 (N_14182,N_10694,N_8387);
or U14183 (N_14183,N_8040,N_10428);
nand U14184 (N_14184,N_8617,N_10491);
nor U14185 (N_14185,N_8318,N_11952);
and U14186 (N_14186,N_8291,N_9759);
or U14187 (N_14187,N_8753,N_11531);
and U14188 (N_14188,N_10952,N_10672);
nor U14189 (N_14189,N_11239,N_8479);
nor U14190 (N_14190,N_9378,N_8334);
nor U14191 (N_14191,N_11131,N_8723);
and U14192 (N_14192,N_9483,N_8150);
nor U14193 (N_14193,N_9713,N_11670);
or U14194 (N_14194,N_8392,N_8298);
nand U14195 (N_14195,N_9150,N_10673);
or U14196 (N_14196,N_11141,N_9174);
nand U14197 (N_14197,N_9719,N_11981);
or U14198 (N_14198,N_9920,N_10923);
nor U14199 (N_14199,N_10038,N_9800);
or U14200 (N_14200,N_9837,N_9301);
or U14201 (N_14201,N_9558,N_11908);
nand U14202 (N_14202,N_8995,N_9814);
and U14203 (N_14203,N_8891,N_10422);
nor U14204 (N_14204,N_8766,N_9890);
and U14205 (N_14205,N_10797,N_8428);
or U14206 (N_14206,N_10997,N_10283);
nor U14207 (N_14207,N_8175,N_8879);
and U14208 (N_14208,N_9017,N_9766);
nor U14209 (N_14209,N_8529,N_8698);
nand U14210 (N_14210,N_8911,N_11412);
nand U14211 (N_14211,N_10437,N_11578);
nor U14212 (N_14212,N_8087,N_8159);
nor U14213 (N_14213,N_9648,N_9278);
nand U14214 (N_14214,N_9714,N_9101);
nand U14215 (N_14215,N_10013,N_8261);
and U14216 (N_14216,N_11670,N_11295);
or U14217 (N_14217,N_11774,N_11255);
nand U14218 (N_14218,N_8645,N_10020);
nor U14219 (N_14219,N_9380,N_8941);
or U14220 (N_14220,N_10877,N_10109);
and U14221 (N_14221,N_9252,N_10793);
or U14222 (N_14222,N_11995,N_8308);
or U14223 (N_14223,N_10948,N_8728);
nand U14224 (N_14224,N_10713,N_9258);
nor U14225 (N_14225,N_10006,N_10557);
nand U14226 (N_14226,N_8512,N_9348);
nand U14227 (N_14227,N_8650,N_8958);
and U14228 (N_14228,N_8783,N_9243);
nand U14229 (N_14229,N_9952,N_10168);
nand U14230 (N_14230,N_8744,N_8706);
nand U14231 (N_14231,N_10937,N_8285);
nor U14232 (N_14232,N_8258,N_11128);
nor U14233 (N_14233,N_11080,N_8642);
and U14234 (N_14234,N_9964,N_10715);
nor U14235 (N_14235,N_11124,N_11685);
nor U14236 (N_14236,N_11661,N_10681);
and U14237 (N_14237,N_10602,N_10710);
or U14238 (N_14238,N_9512,N_11949);
nor U14239 (N_14239,N_11425,N_11558);
nor U14240 (N_14240,N_11292,N_8399);
nor U14241 (N_14241,N_8832,N_8117);
and U14242 (N_14242,N_11685,N_8145);
nand U14243 (N_14243,N_9770,N_9693);
and U14244 (N_14244,N_9572,N_8109);
and U14245 (N_14245,N_10532,N_9992);
and U14246 (N_14246,N_11536,N_11654);
nor U14247 (N_14247,N_8992,N_11494);
or U14248 (N_14248,N_8778,N_9863);
and U14249 (N_14249,N_9201,N_10942);
nand U14250 (N_14250,N_11147,N_9407);
or U14251 (N_14251,N_8213,N_9577);
nor U14252 (N_14252,N_8828,N_11735);
nand U14253 (N_14253,N_11806,N_10422);
and U14254 (N_14254,N_9552,N_10368);
or U14255 (N_14255,N_8072,N_8350);
and U14256 (N_14256,N_11042,N_11643);
nor U14257 (N_14257,N_8674,N_11115);
nand U14258 (N_14258,N_10577,N_11014);
nand U14259 (N_14259,N_11059,N_9809);
or U14260 (N_14260,N_11788,N_10721);
nor U14261 (N_14261,N_11581,N_9646);
nand U14262 (N_14262,N_8370,N_9006);
nor U14263 (N_14263,N_8832,N_9142);
or U14264 (N_14264,N_10252,N_10636);
and U14265 (N_14265,N_11218,N_8323);
and U14266 (N_14266,N_8667,N_11401);
and U14267 (N_14267,N_8483,N_8308);
and U14268 (N_14268,N_11848,N_9412);
nor U14269 (N_14269,N_11511,N_9799);
or U14270 (N_14270,N_9999,N_10430);
or U14271 (N_14271,N_8888,N_10835);
nand U14272 (N_14272,N_11555,N_8582);
nor U14273 (N_14273,N_9835,N_9886);
or U14274 (N_14274,N_9663,N_11871);
or U14275 (N_14275,N_8486,N_9615);
nor U14276 (N_14276,N_9377,N_9091);
xor U14277 (N_14277,N_11911,N_8877);
or U14278 (N_14278,N_11127,N_8162);
or U14279 (N_14279,N_9123,N_10164);
nor U14280 (N_14280,N_11739,N_8983);
or U14281 (N_14281,N_8357,N_10395);
and U14282 (N_14282,N_9021,N_9726);
nor U14283 (N_14283,N_11805,N_9347);
and U14284 (N_14284,N_10035,N_11798);
or U14285 (N_14285,N_11237,N_11837);
and U14286 (N_14286,N_8904,N_10877);
nand U14287 (N_14287,N_11324,N_8623);
or U14288 (N_14288,N_8141,N_9945);
or U14289 (N_14289,N_10771,N_10625);
nand U14290 (N_14290,N_8427,N_11688);
xnor U14291 (N_14291,N_8699,N_10932);
and U14292 (N_14292,N_10228,N_8780);
nor U14293 (N_14293,N_11870,N_9280);
and U14294 (N_14294,N_11934,N_11763);
nand U14295 (N_14295,N_8525,N_11839);
and U14296 (N_14296,N_8648,N_11424);
nand U14297 (N_14297,N_11430,N_10753);
nand U14298 (N_14298,N_10241,N_10625);
nand U14299 (N_14299,N_10477,N_11451);
or U14300 (N_14300,N_10437,N_9732);
or U14301 (N_14301,N_8643,N_11015);
and U14302 (N_14302,N_9433,N_8179);
or U14303 (N_14303,N_8301,N_9827);
nand U14304 (N_14304,N_8344,N_8282);
nor U14305 (N_14305,N_9614,N_9424);
or U14306 (N_14306,N_10859,N_10958);
or U14307 (N_14307,N_8337,N_9989);
or U14308 (N_14308,N_9804,N_10438);
nand U14309 (N_14309,N_9026,N_11687);
nand U14310 (N_14310,N_10236,N_9916);
or U14311 (N_14311,N_10322,N_10557);
or U14312 (N_14312,N_11514,N_10488);
nand U14313 (N_14313,N_11075,N_9511);
nor U14314 (N_14314,N_9001,N_11820);
and U14315 (N_14315,N_9365,N_10614);
and U14316 (N_14316,N_10616,N_8705);
and U14317 (N_14317,N_10818,N_10875);
nand U14318 (N_14318,N_8421,N_10393);
nand U14319 (N_14319,N_8992,N_11962);
nand U14320 (N_14320,N_8182,N_8054);
nor U14321 (N_14321,N_10772,N_8453);
or U14322 (N_14322,N_8357,N_11583);
nand U14323 (N_14323,N_8949,N_11914);
nand U14324 (N_14324,N_11812,N_10448);
nor U14325 (N_14325,N_10288,N_9824);
and U14326 (N_14326,N_10246,N_11131);
nor U14327 (N_14327,N_9715,N_8509);
and U14328 (N_14328,N_10982,N_8711);
and U14329 (N_14329,N_10177,N_10484);
or U14330 (N_14330,N_9178,N_9800);
and U14331 (N_14331,N_11536,N_10813);
or U14332 (N_14332,N_9592,N_9790);
or U14333 (N_14333,N_8829,N_11190);
nand U14334 (N_14334,N_11410,N_11619);
nand U14335 (N_14335,N_11777,N_10437);
or U14336 (N_14336,N_11155,N_10308);
nor U14337 (N_14337,N_10066,N_10070);
and U14338 (N_14338,N_8009,N_8866);
nor U14339 (N_14339,N_9044,N_8714);
nor U14340 (N_14340,N_9185,N_10042);
or U14341 (N_14341,N_9752,N_11067);
and U14342 (N_14342,N_11977,N_10196);
nor U14343 (N_14343,N_9968,N_10599);
or U14344 (N_14344,N_11039,N_8862);
nand U14345 (N_14345,N_11823,N_8384);
or U14346 (N_14346,N_9638,N_8634);
and U14347 (N_14347,N_10697,N_8819);
nor U14348 (N_14348,N_8246,N_10387);
nor U14349 (N_14349,N_9080,N_8221);
or U14350 (N_14350,N_9229,N_8001);
nor U14351 (N_14351,N_8352,N_9476);
nand U14352 (N_14352,N_9691,N_10715);
nor U14353 (N_14353,N_10627,N_11656);
or U14354 (N_14354,N_8103,N_8001);
or U14355 (N_14355,N_8135,N_11160);
and U14356 (N_14356,N_8189,N_10252);
or U14357 (N_14357,N_9623,N_11988);
nor U14358 (N_14358,N_9113,N_10125);
or U14359 (N_14359,N_10764,N_8449);
or U14360 (N_14360,N_9371,N_9507);
nand U14361 (N_14361,N_9454,N_10656);
nor U14362 (N_14362,N_9174,N_11035);
or U14363 (N_14363,N_11039,N_11023);
nand U14364 (N_14364,N_11342,N_8254);
or U14365 (N_14365,N_10000,N_10592);
nand U14366 (N_14366,N_10026,N_11045);
nor U14367 (N_14367,N_10423,N_9382);
or U14368 (N_14368,N_8036,N_10902);
or U14369 (N_14369,N_8642,N_10642);
nor U14370 (N_14370,N_11944,N_9673);
and U14371 (N_14371,N_9217,N_10220);
or U14372 (N_14372,N_9849,N_9036);
or U14373 (N_14373,N_9470,N_10217);
nor U14374 (N_14374,N_11897,N_9419);
or U14375 (N_14375,N_8924,N_9677);
and U14376 (N_14376,N_11927,N_8543);
or U14377 (N_14377,N_8633,N_11016);
or U14378 (N_14378,N_10277,N_8564);
or U14379 (N_14379,N_8443,N_9269);
nand U14380 (N_14380,N_9325,N_8137);
nor U14381 (N_14381,N_9284,N_10776);
and U14382 (N_14382,N_9610,N_10815);
nor U14383 (N_14383,N_8642,N_11623);
nand U14384 (N_14384,N_11637,N_8844);
nand U14385 (N_14385,N_8681,N_9415);
or U14386 (N_14386,N_9153,N_11113);
and U14387 (N_14387,N_11043,N_10872);
xor U14388 (N_14388,N_9710,N_11119);
nor U14389 (N_14389,N_9192,N_11204);
and U14390 (N_14390,N_11114,N_11186);
or U14391 (N_14391,N_10582,N_9236);
or U14392 (N_14392,N_10887,N_8433);
nand U14393 (N_14393,N_9148,N_8155);
nand U14394 (N_14394,N_10137,N_10469);
nand U14395 (N_14395,N_9114,N_11028);
and U14396 (N_14396,N_11851,N_10698);
nand U14397 (N_14397,N_9261,N_10046);
nor U14398 (N_14398,N_8654,N_10530);
and U14399 (N_14399,N_10802,N_10025);
nand U14400 (N_14400,N_11846,N_10387);
nand U14401 (N_14401,N_11814,N_9722);
or U14402 (N_14402,N_8734,N_9314);
or U14403 (N_14403,N_11311,N_10435);
or U14404 (N_14404,N_9853,N_8686);
or U14405 (N_14405,N_10678,N_10233);
nor U14406 (N_14406,N_9295,N_10148);
xnor U14407 (N_14407,N_8834,N_8306);
nand U14408 (N_14408,N_10444,N_10505);
nor U14409 (N_14409,N_8290,N_8795);
and U14410 (N_14410,N_9317,N_10112);
or U14411 (N_14411,N_11000,N_8416);
nand U14412 (N_14412,N_9402,N_8678);
nand U14413 (N_14413,N_8327,N_9536);
nor U14414 (N_14414,N_8591,N_9461);
and U14415 (N_14415,N_11206,N_8132);
nand U14416 (N_14416,N_9283,N_9102);
and U14417 (N_14417,N_8023,N_11247);
or U14418 (N_14418,N_11210,N_10527);
nand U14419 (N_14419,N_8157,N_11843);
nor U14420 (N_14420,N_9434,N_9903);
and U14421 (N_14421,N_9106,N_11094);
and U14422 (N_14422,N_9116,N_11783);
or U14423 (N_14423,N_10127,N_9726);
and U14424 (N_14424,N_11687,N_9324);
and U14425 (N_14425,N_10032,N_8782);
and U14426 (N_14426,N_8533,N_10019);
nor U14427 (N_14427,N_9804,N_9448);
or U14428 (N_14428,N_11758,N_11296);
nand U14429 (N_14429,N_9081,N_8985);
or U14430 (N_14430,N_8528,N_9028);
and U14431 (N_14431,N_9520,N_10232);
or U14432 (N_14432,N_8422,N_10718);
and U14433 (N_14433,N_11079,N_10659);
and U14434 (N_14434,N_9505,N_11774);
nand U14435 (N_14435,N_11042,N_10078);
and U14436 (N_14436,N_10828,N_10238);
nor U14437 (N_14437,N_8645,N_9373);
nor U14438 (N_14438,N_10904,N_9798);
nor U14439 (N_14439,N_8429,N_9025);
nand U14440 (N_14440,N_11189,N_11334);
nor U14441 (N_14441,N_11759,N_9136);
nor U14442 (N_14442,N_11393,N_9725);
nor U14443 (N_14443,N_11602,N_10890);
and U14444 (N_14444,N_9754,N_8280);
or U14445 (N_14445,N_10291,N_11880);
nor U14446 (N_14446,N_9235,N_10097);
or U14447 (N_14447,N_8692,N_8404);
or U14448 (N_14448,N_11003,N_11243);
or U14449 (N_14449,N_8298,N_9778);
nand U14450 (N_14450,N_10328,N_11021);
and U14451 (N_14451,N_9845,N_9940);
nor U14452 (N_14452,N_8087,N_8980);
nor U14453 (N_14453,N_11203,N_11037);
nor U14454 (N_14454,N_10170,N_11045);
nor U14455 (N_14455,N_9205,N_10931);
or U14456 (N_14456,N_9799,N_11109);
and U14457 (N_14457,N_9688,N_11820);
nand U14458 (N_14458,N_9473,N_8691);
nand U14459 (N_14459,N_8846,N_8483);
and U14460 (N_14460,N_11661,N_11712);
and U14461 (N_14461,N_11249,N_11134);
nand U14462 (N_14462,N_9091,N_8720);
and U14463 (N_14463,N_8356,N_10989);
nor U14464 (N_14464,N_11591,N_11244);
and U14465 (N_14465,N_8638,N_11973);
and U14466 (N_14466,N_9296,N_10548);
nand U14467 (N_14467,N_11157,N_10407);
and U14468 (N_14468,N_10104,N_9674);
nand U14469 (N_14469,N_9670,N_11379);
and U14470 (N_14470,N_10628,N_11150);
and U14471 (N_14471,N_9135,N_8899);
and U14472 (N_14472,N_9654,N_11530);
nand U14473 (N_14473,N_9483,N_10971);
or U14474 (N_14474,N_11479,N_9709);
and U14475 (N_14475,N_9744,N_9697);
and U14476 (N_14476,N_10125,N_11233);
nand U14477 (N_14477,N_11254,N_8259);
nor U14478 (N_14478,N_11094,N_9242);
nor U14479 (N_14479,N_10564,N_8362);
or U14480 (N_14480,N_8132,N_11003);
and U14481 (N_14481,N_8303,N_10549);
or U14482 (N_14482,N_10685,N_11520);
or U14483 (N_14483,N_10669,N_8608);
nor U14484 (N_14484,N_8769,N_10406);
and U14485 (N_14485,N_8435,N_10729);
nor U14486 (N_14486,N_10162,N_10091);
or U14487 (N_14487,N_11842,N_9281);
nor U14488 (N_14488,N_11673,N_10907);
or U14489 (N_14489,N_9800,N_9382);
nor U14490 (N_14490,N_11027,N_11512);
nor U14491 (N_14491,N_11845,N_11682);
nor U14492 (N_14492,N_9913,N_9178);
or U14493 (N_14493,N_9028,N_11283);
and U14494 (N_14494,N_9236,N_9761);
nor U14495 (N_14495,N_10254,N_10987);
or U14496 (N_14496,N_8955,N_9397);
nor U14497 (N_14497,N_8324,N_8198);
nand U14498 (N_14498,N_9019,N_9057);
nand U14499 (N_14499,N_11759,N_11994);
nand U14500 (N_14500,N_8169,N_10956);
or U14501 (N_14501,N_11614,N_8811);
nor U14502 (N_14502,N_10574,N_10069);
nor U14503 (N_14503,N_9845,N_9062);
nand U14504 (N_14504,N_9999,N_10240);
or U14505 (N_14505,N_8535,N_9918);
and U14506 (N_14506,N_11667,N_10438);
nand U14507 (N_14507,N_9540,N_11799);
and U14508 (N_14508,N_8195,N_10469);
nand U14509 (N_14509,N_11947,N_11996);
nand U14510 (N_14510,N_11691,N_11475);
nand U14511 (N_14511,N_9752,N_8303);
nand U14512 (N_14512,N_9737,N_10665);
and U14513 (N_14513,N_9601,N_10160);
or U14514 (N_14514,N_11366,N_11374);
and U14515 (N_14515,N_10439,N_9866);
and U14516 (N_14516,N_9101,N_8772);
nor U14517 (N_14517,N_11815,N_8239);
nand U14518 (N_14518,N_10158,N_8629);
and U14519 (N_14519,N_11894,N_8360);
nor U14520 (N_14520,N_8781,N_11810);
nand U14521 (N_14521,N_8094,N_10798);
nor U14522 (N_14522,N_8978,N_10498);
and U14523 (N_14523,N_8881,N_8465);
and U14524 (N_14524,N_10845,N_10494);
or U14525 (N_14525,N_11288,N_9338);
nand U14526 (N_14526,N_8834,N_11909);
nand U14527 (N_14527,N_8106,N_11122);
and U14528 (N_14528,N_11375,N_8994);
or U14529 (N_14529,N_8906,N_8507);
nand U14530 (N_14530,N_11459,N_8618);
nor U14531 (N_14531,N_10276,N_10251);
and U14532 (N_14532,N_8805,N_9924);
nor U14533 (N_14533,N_8951,N_9653);
nand U14534 (N_14534,N_8485,N_9937);
nor U14535 (N_14535,N_9179,N_8175);
and U14536 (N_14536,N_8550,N_9875);
or U14537 (N_14537,N_11597,N_11147);
nor U14538 (N_14538,N_9482,N_9408);
nor U14539 (N_14539,N_11746,N_9028);
nor U14540 (N_14540,N_8918,N_11785);
or U14541 (N_14541,N_8609,N_10963);
and U14542 (N_14542,N_11759,N_8309);
and U14543 (N_14543,N_8091,N_9840);
and U14544 (N_14544,N_8686,N_9741);
nand U14545 (N_14545,N_11649,N_9937);
nand U14546 (N_14546,N_11327,N_9620);
nand U14547 (N_14547,N_9748,N_8121);
nor U14548 (N_14548,N_8607,N_10495);
or U14549 (N_14549,N_10419,N_11989);
and U14550 (N_14550,N_11533,N_11452);
nand U14551 (N_14551,N_11548,N_11333);
and U14552 (N_14552,N_8435,N_8481);
or U14553 (N_14553,N_10434,N_11830);
or U14554 (N_14554,N_11801,N_8696);
nor U14555 (N_14555,N_11579,N_10781);
and U14556 (N_14556,N_10121,N_11718);
and U14557 (N_14557,N_8197,N_11194);
nor U14558 (N_14558,N_11791,N_10634);
or U14559 (N_14559,N_9960,N_8023);
nor U14560 (N_14560,N_8586,N_8932);
nand U14561 (N_14561,N_8663,N_10906);
nand U14562 (N_14562,N_8057,N_9358);
or U14563 (N_14563,N_8890,N_9257);
and U14564 (N_14564,N_10261,N_9107);
and U14565 (N_14565,N_10085,N_8136);
and U14566 (N_14566,N_11524,N_10604);
nor U14567 (N_14567,N_10761,N_9875);
and U14568 (N_14568,N_11729,N_10818);
nor U14569 (N_14569,N_10141,N_9678);
and U14570 (N_14570,N_10316,N_8669);
or U14571 (N_14571,N_11274,N_10241);
nor U14572 (N_14572,N_9183,N_9114);
nor U14573 (N_14573,N_10583,N_10898);
or U14574 (N_14574,N_9058,N_8257);
and U14575 (N_14575,N_8716,N_8601);
nand U14576 (N_14576,N_9873,N_10320);
nor U14577 (N_14577,N_11123,N_8083);
nor U14578 (N_14578,N_10490,N_8094);
and U14579 (N_14579,N_8602,N_10273);
nand U14580 (N_14580,N_8377,N_10260);
or U14581 (N_14581,N_8818,N_8645);
nor U14582 (N_14582,N_10908,N_8888);
or U14583 (N_14583,N_9639,N_8453);
nand U14584 (N_14584,N_11867,N_8967);
or U14585 (N_14585,N_10280,N_9921);
nand U14586 (N_14586,N_9861,N_8196);
or U14587 (N_14587,N_10707,N_10349);
and U14588 (N_14588,N_8369,N_8472);
or U14589 (N_14589,N_9459,N_10906);
and U14590 (N_14590,N_8071,N_8448);
nor U14591 (N_14591,N_8913,N_10818);
nor U14592 (N_14592,N_11881,N_9310);
and U14593 (N_14593,N_11317,N_9326);
and U14594 (N_14594,N_11528,N_10977);
nand U14595 (N_14595,N_11315,N_10138);
nor U14596 (N_14596,N_11851,N_10451);
nor U14597 (N_14597,N_11153,N_9235);
and U14598 (N_14598,N_10033,N_8496);
or U14599 (N_14599,N_8135,N_10865);
and U14600 (N_14600,N_10700,N_10854);
or U14601 (N_14601,N_11886,N_10470);
nand U14602 (N_14602,N_8731,N_8830);
or U14603 (N_14603,N_8231,N_10533);
nand U14604 (N_14604,N_9528,N_9571);
and U14605 (N_14605,N_9978,N_8366);
or U14606 (N_14606,N_9199,N_11504);
nand U14607 (N_14607,N_9072,N_10128);
nor U14608 (N_14608,N_10465,N_11939);
nor U14609 (N_14609,N_10998,N_10395);
nor U14610 (N_14610,N_8970,N_11479);
or U14611 (N_14611,N_11116,N_9230);
or U14612 (N_14612,N_8017,N_9285);
nor U14613 (N_14613,N_8918,N_8367);
or U14614 (N_14614,N_8533,N_8230);
nor U14615 (N_14615,N_11029,N_10968);
and U14616 (N_14616,N_10617,N_9681);
nand U14617 (N_14617,N_11550,N_10957);
nor U14618 (N_14618,N_9206,N_8057);
or U14619 (N_14619,N_9936,N_11320);
and U14620 (N_14620,N_8256,N_10032);
and U14621 (N_14621,N_11642,N_9203);
nor U14622 (N_14622,N_8194,N_10400);
nand U14623 (N_14623,N_11745,N_8430);
or U14624 (N_14624,N_11981,N_8673);
or U14625 (N_14625,N_9791,N_10933);
nand U14626 (N_14626,N_11814,N_9796);
nor U14627 (N_14627,N_8982,N_10030);
nand U14628 (N_14628,N_11252,N_8345);
nor U14629 (N_14629,N_10795,N_8029);
or U14630 (N_14630,N_9239,N_11052);
nor U14631 (N_14631,N_8284,N_8145);
nand U14632 (N_14632,N_11484,N_11462);
and U14633 (N_14633,N_10948,N_8098);
or U14634 (N_14634,N_11365,N_8001);
and U14635 (N_14635,N_10277,N_9192);
and U14636 (N_14636,N_10148,N_11912);
nor U14637 (N_14637,N_10039,N_10141);
and U14638 (N_14638,N_9889,N_10224);
or U14639 (N_14639,N_10512,N_11868);
or U14640 (N_14640,N_9466,N_9524);
nand U14641 (N_14641,N_11745,N_10099);
nand U14642 (N_14642,N_11815,N_8405);
nand U14643 (N_14643,N_11803,N_8407);
and U14644 (N_14644,N_11890,N_11117);
and U14645 (N_14645,N_10951,N_10911);
nand U14646 (N_14646,N_8942,N_10039);
and U14647 (N_14647,N_11612,N_9665);
or U14648 (N_14648,N_8916,N_9090);
and U14649 (N_14649,N_9113,N_10987);
nand U14650 (N_14650,N_8898,N_8022);
or U14651 (N_14651,N_11238,N_9370);
and U14652 (N_14652,N_8901,N_10892);
nor U14653 (N_14653,N_11552,N_11754);
or U14654 (N_14654,N_8295,N_9951);
and U14655 (N_14655,N_9858,N_11388);
and U14656 (N_14656,N_8139,N_10878);
and U14657 (N_14657,N_10622,N_11542);
nor U14658 (N_14658,N_11130,N_10133);
nand U14659 (N_14659,N_11467,N_10715);
and U14660 (N_14660,N_11831,N_8889);
or U14661 (N_14661,N_11581,N_8032);
and U14662 (N_14662,N_11033,N_11218);
and U14663 (N_14663,N_11980,N_10882);
nand U14664 (N_14664,N_9711,N_9991);
and U14665 (N_14665,N_10382,N_9835);
or U14666 (N_14666,N_8129,N_11126);
or U14667 (N_14667,N_9000,N_8558);
or U14668 (N_14668,N_8635,N_8687);
or U14669 (N_14669,N_11990,N_9175);
nor U14670 (N_14670,N_8560,N_11604);
and U14671 (N_14671,N_11585,N_11590);
or U14672 (N_14672,N_8852,N_10230);
or U14673 (N_14673,N_9121,N_9844);
nor U14674 (N_14674,N_11465,N_9208);
or U14675 (N_14675,N_9437,N_11700);
and U14676 (N_14676,N_9103,N_11287);
nand U14677 (N_14677,N_11972,N_8440);
or U14678 (N_14678,N_9836,N_9839);
or U14679 (N_14679,N_9298,N_11328);
and U14680 (N_14680,N_9202,N_10980);
or U14681 (N_14681,N_11185,N_9939);
and U14682 (N_14682,N_10327,N_11159);
or U14683 (N_14683,N_9116,N_9465);
nand U14684 (N_14684,N_11521,N_8028);
nor U14685 (N_14685,N_8043,N_8958);
nor U14686 (N_14686,N_11269,N_11102);
nand U14687 (N_14687,N_11642,N_9610);
and U14688 (N_14688,N_10506,N_8833);
nor U14689 (N_14689,N_8821,N_8645);
and U14690 (N_14690,N_10530,N_8986);
nor U14691 (N_14691,N_8003,N_9818);
or U14692 (N_14692,N_9671,N_8368);
or U14693 (N_14693,N_11319,N_11984);
or U14694 (N_14694,N_9159,N_9728);
and U14695 (N_14695,N_10496,N_11531);
or U14696 (N_14696,N_10673,N_10359);
and U14697 (N_14697,N_8938,N_10252);
nor U14698 (N_14698,N_8319,N_11227);
and U14699 (N_14699,N_9477,N_10874);
xnor U14700 (N_14700,N_11346,N_8164);
nor U14701 (N_14701,N_8189,N_10349);
and U14702 (N_14702,N_11785,N_9301);
nand U14703 (N_14703,N_8283,N_9307);
nand U14704 (N_14704,N_9801,N_9391);
nor U14705 (N_14705,N_11530,N_10872);
and U14706 (N_14706,N_10203,N_11465);
nor U14707 (N_14707,N_11247,N_10449);
nor U14708 (N_14708,N_9861,N_10068);
nand U14709 (N_14709,N_11076,N_9863);
or U14710 (N_14710,N_9635,N_8965);
nand U14711 (N_14711,N_8539,N_10295);
or U14712 (N_14712,N_11777,N_8896);
nand U14713 (N_14713,N_8371,N_8068);
and U14714 (N_14714,N_10435,N_8696);
nor U14715 (N_14715,N_9849,N_8175);
nand U14716 (N_14716,N_10794,N_10433);
nor U14717 (N_14717,N_9069,N_8056);
or U14718 (N_14718,N_9840,N_10638);
and U14719 (N_14719,N_10480,N_10601);
nand U14720 (N_14720,N_8046,N_8263);
and U14721 (N_14721,N_9887,N_10817);
or U14722 (N_14722,N_8576,N_9018);
nand U14723 (N_14723,N_11998,N_8713);
nand U14724 (N_14724,N_9663,N_8404);
nor U14725 (N_14725,N_11548,N_9684);
or U14726 (N_14726,N_8232,N_8660);
or U14727 (N_14727,N_8514,N_10679);
and U14728 (N_14728,N_9732,N_9394);
or U14729 (N_14729,N_11178,N_9844);
or U14730 (N_14730,N_11075,N_9371);
or U14731 (N_14731,N_9203,N_11312);
or U14732 (N_14732,N_9973,N_11873);
nor U14733 (N_14733,N_9696,N_10907);
or U14734 (N_14734,N_9136,N_8357);
and U14735 (N_14735,N_9629,N_11327);
nand U14736 (N_14736,N_11245,N_8137);
and U14737 (N_14737,N_9665,N_11547);
and U14738 (N_14738,N_11612,N_11390);
nor U14739 (N_14739,N_10580,N_11334);
nor U14740 (N_14740,N_11426,N_9638);
nand U14741 (N_14741,N_10835,N_8309);
and U14742 (N_14742,N_9237,N_9195);
or U14743 (N_14743,N_10732,N_8913);
nand U14744 (N_14744,N_8173,N_8612);
nand U14745 (N_14745,N_11607,N_9646);
nand U14746 (N_14746,N_9942,N_11268);
nand U14747 (N_14747,N_8427,N_10433);
nand U14748 (N_14748,N_10129,N_8215);
and U14749 (N_14749,N_11960,N_10659);
and U14750 (N_14750,N_11289,N_11111);
or U14751 (N_14751,N_8948,N_9347);
and U14752 (N_14752,N_8610,N_9554);
nor U14753 (N_14753,N_8114,N_8847);
nand U14754 (N_14754,N_10667,N_8038);
and U14755 (N_14755,N_10592,N_8502);
or U14756 (N_14756,N_11349,N_11235);
or U14757 (N_14757,N_10878,N_8390);
nor U14758 (N_14758,N_11519,N_11059);
nand U14759 (N_14759,N_8506,N_11219);
or U14760 (N_14760,N_8693,N_8167);
nand U14761 (N_14761,N_8998,N_8733);
nand U14762 (N_14762,N_8635,N_8624);
nand U14763 (N_14763,N_9121,N_9830);
and U14764 (N_14764,N_11070,N_8435);
nor U14765 (N_14765,N_8998,N_9600);
or U14766 (N_14766,N_11905,N_11162);
and U14767 (N_14767,N_11829,N_11511);
nand U14768 (N_14768,N_11951,N_9151);
and U14769 (N_14769,N_11536,N_9379);
or U14770 (N_14770,N_9768,N_10720);
and U14771 (N_14771,N_11559,N_9083);
or U14772 (N_14772,N_8334,N_11467);
or U14773 (N_14773,N_11744,N_10786);
and U14774 (N_14774,N_9989,N_11131);
or U14775 (N_14775,N_8593,N_11459);
nor U14776 (N_14776,N_9359,N_8210);
and U14777 (N_14777,N_11890,N_11239);
and U14778 (N_14778,N_10475,N_10196);
nand U14779 (N_14779,N_9180,N_8485);
nand U14780 (N_14780,N_10749,N_10972);
nor U14781 (N_14781,N_11897,N_8242);
or U14782 (N_14782,N_10020,N_8330);
and U14783 (N_14783,N_11380,N_9640);
and U14784 (N_14784,N_10575,N_10246);
or U14785 (N_14785,N_9904,N_11103);
nor U14786 (N_14786,N_11965,N_10727);
and U14787 (N_14787,N_11649,N_9695);
nand U14788 (N_14788,N_8254,N_9036);
nand U14789 (N_14789,N_10854,N_9087);
nand U14790 (N_14790,N_9176,N_10806);
xor U14791 (N_14791,N_11044,N_11254);
and U14792 (N_14792,N_11303,N_8483);
or U14793 (N_14793,N_9883,N_8711);
and U14794 (N_14794,N_11595,N_8056);
nor U14795 (N_14795,N_11672,N_9438);
or U14796 (N_14796,N_9846,N_10492);
or U14797 (N_14797,N_8560,N_11482);
or U14798 (N_14798,N_10656,N_9026);
nand U14799 (N_14799,N_11134,N_11866);
and U14800 (N_14800,N_11461,N_11144);
nor U14801 (N_14801,N_9428,N_11873);
nand U14802 (N_14802,N_8277,N_11240);
or U14803 (N_14803,N_9469,N_11441);
or U14804 (N_14804,N_9518,N_8927);
or U14805 (N_14805,N_8297,N_11145);
nor U14806 (N_14806,N_11759,N_8682);
or U14807 (N_14807,N_11664,N_8602);
nand U14808 (N_14808,N_9543,N_11164);
nor U14809 (N_14809,N_10757,N_9927);
nor U14810 (N_14810,N_8454,N_11210);
and U14811 (N_14811,N_8493,N_8034);
nand U14812 (N_14812,N_10929,N_10142);
nand U14813 (N_14813,N_11591,N_10079);
nor U14814 (N_14814,N_9414,N_9161);
and U14815 (N_14815,N_10337,N_9658);
and U14816 (N_14816,N_9450,N_11309);
nand U14817 (N_14817,N_10776,N_10357);
nor U14818 (N_14818,N_9812,N_11173);
or U14819 (N_14819,N_10850,N_9467);
nand U14820 (N_14820,N_11040,N_8916);
or U14821 (N_14821,N_10281,N_11675);
nand U14822 (N_14822,N_11949,N_9277);
nor U14823 (N_14823,N_8664,N_10525);
or U14824 (N_14824,N_9471,N_11020);
or U14825 (N_14825,N_8545,N_10819);
nand U14826 (N_14826,N_11015,N_8694);
nand U14827 (N_14827,N_9929,N_10922);
or U14828 (N_14828,N_8047,N_11720);
or U14829 (N_14829,N_10836,N_9286);
or U14830 (N_14830,N_11018,N_10411);
and U14831 (N_14831,N_11133,N_10091);
nand U14832 (N_14832,N_9129,N_8199);
nand U14833 (N_14833,N_11451,N_8458);
and U14834 (N_14834,N_9544,N_8676);
or U14835 (N_14835,N_10298,N_8971);
and U14836 (N_14836,N_9032,N_11207);
or U14837 (N_14837,N_9786,N_11248);
or U14838 (N_14838,N_11917,N_11498);
nand U14839 (N_14839,N_11458,N_8322);
nand U14840 (N_14840,N_9643,N_9003);
and U14841 (N_14841,N_11357,N_10203);
or U14842 (N_14842,N_11598,N_11460);
nor U14843 (N_14843,N_9332,N_10734);
and U14844 (N_14844,N_11137,N_11957);
or U14845 (N_14845,N_9746,N_8874);
and U14846 (N_14846,N_9823,N_10988);
and U14847 (N_14847,N_9861,N_9184);
nand U14848 (N_14848,N_9541,N_8714);
nor U14849 (N_14849,N_8272,N_10274);
nor U14850 (N_14850,N_8151,N_8871);
nor U14851 (N_14851,N_10409,N_8077);
nand U14852 (N_14852,N_10661,N_11849);
or U14853 (N_14853,N_10144,N_11262);
or U14854 (N_14854,N_11588,N_10937);
nor U14855 (N_14855,N_8865,N_11896);
nand U14856 (N_14856,N_10088,N_9741);
and U14857 (N_14857,N_8790,N_10575);
nand U14858 (N_14858,N_10464,N_10331);
nor U14859 (N_14859,N_8365,N_11368);
and U14860 (N_14860,N_10664,N_10787);
or U14861 (N_14861,N_8445,N_8986);
nor U14862 (N_14862,N_9987,N_8491);
nor U14863 (N_14863,N_8964,N_11504);
or U14864 (N_14864,N_8479,N_8725);
or U14865 (N_14865,N_9517,N_11384);
and U14866 (N_14866,N_8385,N_9981);
and U14867 (N_14867,N_10426,N_11091);
nand U14868 (N_14868,N_10954,N_11590);
nor U14869 (N_14869,N_10611,N_9807);
nand U14870 (N_14870,N_11768,N_8549);
or U14871 (N_14871,N_10783,N_11125);
or U14872 (N_14872,N_9392,N_9306);
nand U14873 (N_14873,N_11244,N_10365);
nand U14874 (N_14874,N_11346,N_8500);
and U14875 (N_14875,N_11211,N_10396);
nor U14876 (N_14876,N_9992,N_10632);
or U14877 (N_14877,N_9135,N_8981);
nor U14878 (N_14878,N_11581,N_11117);
nand U14879 (N_14879,N_10705,N_9164);
nor U14880 (N_14880,N_10218,N_8255);
and U14881 (N_14881,N_10386,N_11637);
or U14882 (N_14882,N_11313,N_11658);
or U14883 (N_14883,N_9207,N_11676);
or U14884 (N_14884,N_8043,N_9055);
and U14885 (N_14885,N_10391,N_9693);
nand U14886 (N_14886,N_8650,N_8801);
or U14887 (N_14887,N_10590,N_8622);
and U14888 (N_14888,N_11148,N_9170);
and U14889 (N_14889,N_11812,N_10086);
nor U14890 (N_14890,N_11633,N_11786);
and U14891 (N_14891,N_8852,N_9156);
nor U14892 (N_14892,N_9809,N_11998);
nand U14893 (N_14893,N_10642,N_9736);
nor U14894 (N_14894,N_9411,N_11519);
or U14895 (N_14895,N_10251,N_10019);
or U14896 (N_14896,N_10974,N_11216);
and U14897 (N_14897,N_10677,N_10512);
nand U14898 (N_14898,N_8360,N_9287);
nor U14899 (N_14899,N_10397,N_8297);
nor U14900 (N_14900,N_11461,N_10164);
and U14901 (N_14901,N_9841,N_11886);
nor U14902 (N_14902,N_8617,N_9091);
nand U14903 (N_14903,N_8590,N_9348);
and U14904 (N_14904,N_9840,N_9108);
or U14905 (N_14905,N_9253,N_8562);
or U14906 (N_14906,N_8223,N_9849);
nand U14907 (N_14907,N_11736,N_9998);
nor U14908 (N_14908,N_8395,N_10772);
nor U14909 (N_14909,N_8289,N_11616);
or U14910 (N_14910,N_11775,N_10105);
nand U14911 (N_14911,N_8142,N_11847);
nand U14912 (N_14912,N_8500,N_10399);
or U14913 (N_14913,N_9773,N_8382);
nor U14914 (N_14914,N_11186,N_10023);
or U14915 (N_14915,N_9275,N_10922);
nor U14916 (N_14916,N_9546,N_9210);
nor U14917 (N_14917,N_9733,N_9880);
nand U14918 (N_14918,N_11479,N_10058);
or U14919 (N_14919,N_10838,N_11088);
and U14920 (N_14920,N_8450,N_11820);
and U14921 (N_14921,N_9916,N_8118);
and U14922 (N_14922,N_11364,N_10018);
nand U14923 (N_14923,N_11276,N_9016);
nand U14924 (N_14924,N_10743,N_9658);
nor U14925 (N_14925,N_9543,N_11196);
and U14926 (N_14926,N_8492,N_11189);
and U14927 (N_14927,N_9846,N_8985);
or U14928 (N_14928,N_8803,N_10132);
and U14929 (N_14929,N_8382,N_10495);
nor U14930 (N_14930,N_9066,N_10661);
or U14931 (N_14931,N_9313,N_9502);
nand U14932 (N_14932,N_9511,N_8616);
nand U14933 (N_14933,N_9552,N_10511);
nor U14934 (N_14934,N_8359,N_11937);
or U14935 (N_14935,N_9882,N_8839);
nand U14936 (N_14936,N_10024,N_9936);
nand U14937 (N_14937,N_9957,N_10144);
nor U14938 (N_14938,N_10737,N_10639);
and U14939 (N_14939,N_8774,N_10458);
and U14940 (N_14940,N_10915,N_11441);
nor U14941 (N_14941,N_9947,N_10517);
or U14942 (N_14942,N_9226,N_11771);
nand U14943 (N_14943,N_10044,N_10825);
nand U14944 (N_14944,N_8218,N_8910);
nor U14945 (N_14945,N_11720,N_8730);
or U14946 (N_14946,N_11227,N_9350);
and U14947 (N_14947,N_10775,N_11381);
and U14948 (N_14948,N_11463,N_9073);
nor U14949 (N_14949,N_11307,N_10163);
nor U14950 (N_14950,N_10543,N_10231);
and U14951 (N_14951,N_11299,N_11025);
nand U14952 (N_14952,N_9301,N_8284);
and U14953 (N_14953,N_11551,N_9137);
or U14954 (N_14954,N_8681,N_9798);
nand U14955 (N_14955,N_9020,N_10141);
nor U14956 (N_14956,N_8165,N_10124);
or U14957 (N_14957,N_11480,N_8249);
and U14958 (N_14958,N_11205,N_8530);
nand U14959 (N_14959,N_8800,N_10936);
nand U14960 (N_14960,N_10540,N_8126);
and U14961 (N_14961,N_8024,N_11560);
nor U14962 (N_14962,N_11323,N_10990);
nor U14963 (N_14963,N_11464,N_8930);
and U14964 (N_14964,N_11126,N_11508);
or U14965 (N_14965,N_10346,N_10665);
and U14966 (N_14966,N_10206,N_9572);
or U14967 (N_14967,N_9165,N_10733);
or U14968 (N_14968,N_8582,N_11618);
nand U14969 (N_14969,N_11841,N_8299);
nand U14970 (N_14970,N_8532,N_8591);
and U14971 (N_14971,N_10016,N_9821);
nand U14972 (N_14972,N_9448,N_8908);
nor U14973 (N_14973,N_10294,N_8106);
and U14974 (N_14974,N_11303,N_10709);
nand U14975 (N_14975,N_10410,N_8504);
nor U14976 (N_14976,N_9834,N_9747);
and U14977 (N_14977,N_11454,N_8098);
nor U14978 (N_14978,N_10546,N_10303);
nor U14979 (N_14979,N_8161,N_8834);
nand U14980 (N_14980,N_9392,N_9057);
or U14981 (N_14981,N_8169,N_9070);
nor U14982 (N_14982,N_11519,N_9741);
or U14983 (N_14983,N_11686,N_10376);
nor U14984 (N_14984,N_10154,N_9248);
and U14985 (N_14985,N_9334,N_8678);
nand U14986 (N_14986,N_11973,N_8546);
xnor U14987 (N_14987,N_10768,N_10198);
nor U14988 (N_14988,N_9329,N_10458);
nand U14989 (N_14989,N_8161,N_11291);
or U14990 (N_14990,N_8194,N_9102);
nor U14991 (N_14991,N_9037,N_9383);
or U14992 (N_14992,N_10333,N_8703);
or U14993 (N_14993,N_8693,N_10777);
nand U14994 (N_14994,N_9860,N_11403);
and U14995 (N_14995,N_9239,N_11091);
or U14996 (N_14996,N_8989,N_11327);
nand U14997 (N_14997,N_10609,N_10718);
and U14998 (N_14998,N_8724,N_8009);
nand U14999 (N_14999,N_11540,N_10761);
nand U15000 (N_15000,N_10440,N_8670);
and U15001 (N_15001,N_11086,N_11429);
or U15002 (N_15002,N_8972,N_8945);
nand U15003 (N_15003,N_8591,N_8608);
or U15004 (N_15004,N_10724,N_9664);
nor U15005 (N_15005,N_11859,N_10598);
and U15006 (N_15006,N_9633,N_9626);
nor U15007 (N_15007,N_8384,N_9611);
or U15008 (N_15008,N_9007,N_9382);
or U15009 (N_15009,N_11009,N_8570);
nand U15010 (N_15010,N_8898,N_10106);
nand U15011 (N_15011,N_9900,N_8122);
nand U15012 (N_15012,N_11202,N_8557);
and U15013 (N_15013,N_11900,N_8601);
nor U15014 (N_15014,N_10687,N_11359);
or U15015 (N_15015,N_9123,N_11873);
nor U15016 (N_15016,N_9529,N_9803);
nand U15017 (N_15017,N_9008,N_11138);
or U15018 (N_15018,N_8536,N_9357);
nor U15019 (N_15019,N_11754,N_9393);
nand U15020 (N_15020,N_11855,N_8804);
and U15021 (N_15021,N_10373,N_9054);
nor U15022 (N_15022,N_10987,N_10765);
or U15023 (N_15023,N_8063,N_10306);
and U15024 (N_15024,N_11118,N_10102);
or U15025 (N_15025,N_8161,N_9093);
nor U15026 (N_15026,N_9446,N_11576);
nand U15027 (N_15027,N_9444,N_8584);
nand U15028 (N_15028,N_11778,N_9239);
nand U15029 (N_15029,N_10817,N_8563);
or U15030 (N_15030,N_11129,N_11421);
and U15031 (N_15031,N_10062,N_11056);
or U15032 (N_15032,N_9903,N_9955);
and U15033 (N_15033,N_11994,N_11927);
or U15034 (N_15034,N_11832,N_10547);
and U15035 (N_15035,N_11411,N_8552);
nor U15036 (N_15036,N_9543,N_8427);
xnor U15037 (N_15037,N_11796,N_11726);
and U15038 (N_15038,N_11874,N_10457);
nor U15039 (N_15039,N_8506,N_8010);
nor U15040 (N_15040,N_11907,N_8824);
and U15041 (N_15041,N_8926,N_8549);
nor U15042 (N_15042,N_9834,N_11230);
or U15043 (N_15043,N_10443,N_8842);
nand U15044 (N_15044,N_8134,N_9079);
nand U15045 (N_15045,N_8573,N_11855);
nor U15046 (N_15046,N_9023,N_11688);
nor U15047 (N_15047,N_10147,N_8181);
nor U15048 (N_15048,N_9518,N_8900);
and U15049 (N_15049,N_8876,N_8161);
and U15050 (N_15050,N_11572,N_9876);
and U15051 (N_15051,N_9837,N_11376);
or U15052 (N_15052,N_10871,N_10344);
and U15053 (N_15053,N_8938,N_9966);
nor U15054 (N_15054,N_11120,N_9455);
nand U15055 (N_15055,N_8179,N_9370);
and U15056 (N_15056,N_10172,N_11976);
and U15057 (N_15057,N_9303,N_10701);
or U15058 (N_15058,N_8221,N_9207);
or U15059 (N_15059,N_11780,N_8563);
or U15060 (N_15060,N_9584,N_9631);
or U15061 (N_15061,N_9749,N_11176);
and U15062 (N_15062,N_9927,N_11531);
and U15063 (N_15063,N_8326,N_9161);
and U15064 (N_15064,N_9447,N_8824);
nand U15065 (N_15065,N_10947,N_9257);
and U15066 (N_15066,N_10831,N_11263);
and U15067 (N_15067,N_9689,N_9294);
or U15068 (N_15068,N_11747,N_8932);
nand U15069 (N_15069,N_9908,N_10508);
and U15070 (N_15070,N_10833,N_9462);
and U15071 (N_15071,N_10287,N_11259);
and U15072 (N_15072,N_10873,N_9521);
nor U15073 (N_15073,N_8614,N_10149);
and U15074 (N_15074,N_9247,N_10133);
and U15075 (N_15075,N_10076,N_8190);
nand U15076 (N_15076,N_8555,N_9203);
nand U15077 (N_15077,N_10931,N_9863);
nor U15078 (N_15078,N_8491,N_11833);
or U15079 (N_15079,N_9932,N_11941);
or U15080 (N_15080,N_9516,N_8689);
nor U15081 (N_15081,N_11828,N_9976);
and U15082 (N_15082,N_9441,N_10985);
and U15083 (N_15083,N_10117,N_9619);
nor U15084 (N_15084,N_9531,N_10215);
and U15085 (N_15085,N_11499,N_8067);
and U15086 (N_15086,N_11685,N_11803);
or U15087 (N_15087,N_11957,N_10606);
nor U15088 (N_15088,N_11862,N_9622);
and U15089 (N_15089,N_11545,N_11567);
and U15090 (N_15090,N_8931,N_9431);
nand U15091 (N_15091,N_8956,N_11378);
nand U15092 (N_15092,N_8405,N_9610);
nor U15093 (N_15093,N_8116,N_10515);
and U15094 (N_15094,N_9706,N_8731);
or U15095 (N_15095,N_8084,N_11986);
and U15096 (N_15096,N_11746,N_11144);
nand U15097 (N_15097,N_8810,N_8581);
nand U15098 (N_15098,N_9895,N_10931);
and U15099 (N_15099,N_9841,N_9928);
nand U15100 (N_15100,N_10234,N_10088);
nor U15101 (N_15101,N_11519,N_9651);
or U15102 (N_15102,N_8465,N_11822);
and U15103 (N_15103,N_8871,N_9936);
or U15104 (N_15104,N_10754,N_9525);
or U15105 (N_15105,N_10355,N_8621);
and U15106 (N_15106,N_10085,N_10746);
or U15107 (N_15107,N_8230,N_10923);
nand U15108 (N_15108,N_8662,N_11715);
nand U15109 (N_15109,N_9099,N_9865);
and U15110 (N_15110,N_11992,N_11249);
or U15111 (N_15111,N_11029,N_11558);
or U15112 (N_15112,N_10877,N_9741);
and U15113 (N_15113,N_8569,N_10606);
or U15114 (N_15114,N_11383,N_9502);
nand U15115 (N_15115,N_9218,N_11439);
nor U15116 (N_15116,N_8219,N_11327);
nor U15117 (N_15117,N_8270,N_8987);
nand U15118 (N_15118,N_9283,N_10329);
nand U15119 (N_15119,N_10579,N_11051);
nand U15120 (N_15120,N_9423,N_10182);
nor U15121 (N_15121,N_9645,N_9178);
and U15122 (N_15122,N_8420,N_9514);
or U15123 (N_15123,N_9716,N_9001);
and U15124 (N_15124,N_10541,N_11859);
or U15125 (N_15125,N_8994,N_11274);
nor U15126 (N_15126,N_11355,N_9438);
nor U15127 (N_15127,N_10777,N_10083);
or U15128 (N_15128,N_8739,N_8770);
nand U15129 (N_15129,N_8309,N_10636);
nand U15130 (N_15130,N_9267,N_10010);
nand U15131 (N_15131,N_11866,N_9651);
or U15132 (N_15132,N_8922,N_11273);
and U15133 (N_15133,N_9445,N_9760);
nor U15134 (N_15134,N_11466,N_8950);
or U15135 (N_15135,N_10147,N_8676);
nor U15136 (N_15136,N_11784,N_11684);
or U15137 (N_15137,N_9174,N_11054);
and U15138 (N_15138,N_10336,N_9835);
nand U15139 (N_15139,N_9756,N_11791);
nor U15140 (N_15140,N_10414,N_10585);
nand U15141 (N_15141,N_9548,N_11843);
nand U15142 (N_15142,N_10170,N_11036);
nor U15143 (N_15143,N_8452,N_8042);
or U15144 (N_15144,N_8992,N_11616);
and U15145 (N_15145,N_9216,N_8743);
nor U15146 (N_15146,N_10806,N_11526);
nor U15147 (N_15147,N_10529,N_9283);
and U15148 (N_15148,N_10330,N_11672);
nand U15149 (N_15149,N_11110,N_11953);
or U15150 (N_15150,N_8394,N_9107);
nand U15151 (N_15151,N_9126,N_10773);
or U15152 (N_15152,N_9048,N_10865);
nand U15153 (N_15153,N_9884,N_11056);
nand U15154 (N_15154,N_10076,N_8232);
nor U15155 (N_15155,N_10919,N_8446);
or U15156 (N_15156,N_9573,N_10570);
nor U15157 (N_15157,N_11971,N_10723);
or U15158 (N_15158,N_11428,N_8084);
nor U15159 (N_15159,N_10964,N_11080);
or U15160 (N_15160,N_9526,N_9185);
and U15161 (N_15161,N_8972,N_11075);
or U15162 (N_15162,N_11034,N_11309);
nor U15163 (N_15163,N_9994,N_9192);
nor U15164 (N_15164,N_11774,N_11034);
or U15165 (N_15165,N_11533,N_9027);
or U15166 (N_15166,N_9416,N_11629);
or U15167 (N_15167,N_9800,N_8554);
or U15168 (N_15168,N_11765,N_11543);
nor U15169 (N_15169,N_11433,N_10668);
or U15170 (N_15170,N_8220,N_8312);
nand U15171 (N_15171,N_9081,N_9011);
and U15172 (N_15172,N_9139,N_9061);
nor U15173 (N_15173,N_10754,N_10567);
and U15174 (N_15174,N_9060,N_8794);
nand U15175 (N_15175,N_8863,N_10750);
or U15176 (N_15176,N_8175,N_9325);
nand U15177 (N_15177,N_9251,N_11395);
or U15178 (N_15178,N_8030,N_8071);
nor U15179 (N_15179,N_10153,N_10555);
nand U15180 (N_15180,N_10654,N_11131);
and U15181 (N_15181,N_8737,N_8266);
nand U15182 (N_15182,N_9759,N_10508);
or U15183 (N_15183,N_10496,N_9075);
nand U15184 (N_15184,N_10623,N_11976);
and U15185 (N_15185,N_10647,N_9958);
nor U15186 (N_15186,N_10384,N_11191);
nor U15187 (N_15187,N_11373,N_10281);
or U15188 (N_15188,N_10536,N_9415);
or U15189 (N_15189,N_11055,N_8555);
nor U15190 (N_15190,N_11360,N_11187);
nor U15191 (N_15191,N_11852,N_9924);
nand U15192 (N_15192,N_10007,N_9494);
nand U15193 (N_15193,N_8588,N_9072);
nand U15194 (N_15194,N_11198,N_9059);
or U15195 (N_15195,N_10555,N_11527);
and U15196 (N_15196,N_10478,N_8639);
or U15197 (N_15197,N_8930,N_8714);
nor U15198 (N_15198,N_11666,N_8615);
and U15199 (N_15199,N_9088,N_8736);
nand U15200 (N_15200,N_10394,N_10514);
nor U15201 (N_15201,N_9126,N_11972);
nor U15202 (N_15202,N_8738,N_9784);
nand U15203 (N_15203,N_9828,N_9139);
or U15204 (N_15204,N_11310,N_8805);
or U15205 (N_15205,N_10162,N_11652);
and U15206 (N_15206,N_8710,N_9702);
or U15207 (N_15207,N_9465,N_10209);
nand U15208 (N_15208,N_10295,N_9478);
and U15209 (N_15209,N_11576,N_10783);
nor U15210 (N_15210,N_10534,N_10560);
or U15211 (N_15211,N_8895,N_11939);
or U15212 (N_15212,N_11400,N_11372);
and U15213 (N_15213,N_11415,N_8107);
or U15214 (N_15214,N_8027,N_10945);
or U15215 (N_15215,N_9059,N_10904);
nor U15216 (N_15216,N_9206,N_10586);
or U15217 (N_15217,N_11706,N_11785);
or U15218 (N_15218,N_11558,N_11526);
and U15219 (N_15219,N_10211,N_8812);
and U15220 (N_15220,N_8395,N_9527);
nand U15221 (N_15221,N_8985,N_9185);
nor U15222 (N_15222,N_11590,N_10953);
nand U15223 (N_15223,N_11792,N_10983);
nand U15224 (N_15224,N_8730,N_10055);
nor U15225 (N_15225,N_8802,N_11198);
nor U15226 (N_15226,N_10527,N_11971);
nor U15227 (N_15227,N_10962,N_11882);
and U15228 (N_15228,N_9084,N_11327);
nand U15229 (N_15229,N_10142,N_8651);
and U15230 (N_15230,N_9488,N_8405);
nor U15231 (N_15231,N_10962,N_10410);
nor U15232 (N_15232,N_9764,N_10865);
nor U15233 (N_15233,N_10115,N_9247);
or U15234 (N_15234,N_8430,N_11109);
nand U15235 (N_15235,N_10922,N_11833);
nor U15236 (N_15236,N_8628,N_11608);
and U15237 (N_15237,N_8981,N_8787);
or U15238 (N_15238,N_10502,N_10672);
nor U15239 (N_15239,N_10120,N_11211);
and U15240 (N_15240,N_8507,N_10397);
or U15241 (N_15241,N_10776,N_8328);
and U15242 (N_15242,N_11891,N_9932);
and U15243 (N_15243,N_8985,N_9405);
nand U15244 (N_15244,N_9475,N_11045);
nand U15245 (N_15245,N_11843,N_9142);
nand U15246 (N_15246,N_9788,N_8357);
and U15247 (N_15247,N_11355,N_11040);
nor U15248 (N_15248,N_10136,N_11617);
nand U15249 (N_15249,N_10148,N_9469);
and U15250 (N_15250,N_10888,N_11070);
or U15251 (N_15251,N_11945,N_10449);
nand U15252 (N_15252,N_11766,N_10034);
nor U15253 (N_15253,N_11550,N_8441);
nor U15254 (N_15254,N_8977,N_9267);
and U15255 (N_15255,N_11948,N_11596);
nand U15256 (N_15256,N_11997,N_8009);
or U15257 (N_15257,N_10671,N_11161);
or U15258 (N_15258,N_11612,N_11881);
nor U15259 (N_15259,N_10224,N_10574);
nor U15260 (N_15260,N_8292,N_10731);
or U15261 (N_15261,N_10722,N_10277);
nand U15262 (N_15262,N_8080,N_10815);
nand U15263 (N_15263,N_9843,N_11032);
nand U15264 (N_15264,N_11209,N_11112);
nand U15265 (N_15265,N_11260,N_11113);
nor U15266 (N_15266,N_8154,N_8858);
nand U15267 (N_15267,N_10416,N_10524);
and U15268 (N_15268,N_8209,N_8803);
and U15269 (N_15269,N_10720,N_9375);
and U15270 (N_15270,N_8357,N_9546);
or U15271 (N_15271,N_11360,N_11564);
nand U15272 (N_15272,N_8417,N_10127);
nor U15273 (N_15273,N_8461,N_11377);
nor U15274 (N_15274,N_8262,N_9129);
and U15275 (N_15275,N_10128,N_9951);
and U15276 (N_15276,N_11769,N_11984);
or U15277 (N_15277,N_11443,N_9744);
or U15278 (N_15278,N_11568,N_8347);
nor U15279 (N_15279,N_11297,N_9402);
or U15280 (N_15280,N_8385,N_9159);
and U15281 (N_15281,N_8505,N_10961);
nor U15282 (N_15282,N_9688,N_9741);
or U15283 (N_15283,N_10714,N_11594);
and U15284 (N_15284,N_11447,N_9290);
or U15285 (N_15285,N_9390,N_9113);
or U15286 (N_15286,N_9468,N_8917);
nand U15287 (N_15287,N_8671,N_11685);
and U15288 (N_15288,N_9011,N_10078);
nor U15289 (N_15289,N_10811,N_10132);
or U15290 (N_15290,N_11711,N_10533);
nand U15291 (N_15291,N_10245,N_10850);
nand U15292 (N_15292,N_9860,N_11717);
and U15293 (N_15293,N_11233,N_9195);
or U15294 (N_15294,N_8452,N_8075);
and U15295 (N_15295,N_9796,N_9022);
nor U15296 (N_15296,N_11258,N_10269);
or U15297 (N_15297,N_9322,N_9792);
nand U15298 (N_15298,N_8050,N_9654);
nor U15299 (N_15299,N_8303,N_11487);
or U15300 (N_15300,N_10690,N_11312);
or U15301 (N_15301,N_9847,N_11599);
or U15302 (N_15302,N_10226,N_10438);
xnor U15303 (N_15303,N_8732,N_8030);
nand U15304 (N_15304,N_9972,N_9712);
and U15305 (N_15305,N_8980,N_11934);
nor U15306 (N_15306,N_11238,N_9169);
nor U15307 (N_15307,N_11175,N_9067);
nor U15308 (N_15308,N_9013,N_8109);
nor U15309 (N_15309,N_9920,N_11144);
nand U15310 (N_15310,N_9915,N_11419);
or U15311 (N_15311,N_11620,N_8083);
and U15312 (N_15312,N_10913,N_8165);
and U15313 (N_15313,N_10881,N_9810);
nor U15314 (N_15314,N_8077,N_9688);
and U15315 (N_15315,N_10339,N_10068);
nand U15316 (N_15316,N_9991,N_8492);
and U15317 (N_15317,N_8446,N_11769);
nand U15318 (N_15318,N_10036,N_11636);
nand U15319 (N_15319,N_11766,N_9151);
xnor U15320 (N_15320,N_9741,N_11668);
and U15321 (N_15321,N_8059,N_11980);
nor U15322 (N_15322,N_9522,N_8597);
or U15323 (N_15323,N_8298,N_8026);
nor U15324 (N_15324,N_8133,N_10882);
nor U15325 (N_15325,N_10330,N_8395);
or U15326 (N_15326,N_10436,N_11398);
nor U15327 (N_15327,N_11941,N_10064);
nor U15328 (N_15328,N_9301,N_8506);
or U15329 (N_15329,N_11841,N_8988);
nand U15330 (N_15330,N_9128,N_9232);
nand U15331 (N_15331,N_9401,N_9424);
or U15332 (N_15332,N_11163,N_10893);
nand U15333 (N_15333,N_9829,N_9154);
nand U15334 (N_15334,N_9019,N_10370);
nand U15335 (N_15335,N_9724,N_9191);
nand U15336 (N_15336,N_11368,N_8056);
nand U15337 (N_15337,N_8972,N_8398);
and U15338 (N_15338,N_11484,N_11882);
and U15339 (N_15339,N_10567,N_10171);
nor U15340 (N_15340,N_8310,N_8003);
and U15341 (N_15341,N_11052,N_11029);
nor U15342 (N_15342,N_10996,N_11276);
or U15343 (N_15343,N_10730,N_9006);
nand U15344 (N_15344,N_10650,N_8833);
and U15345 (N_15345,N_8459,N_9125);
nor U15346 (N_15346,N_9645,N_9373);
or U15347 (N_15347,N_8591,N_10287);
nand U15348 (N_15348,N_10059,N_8301);
or U15349 (N_15349,N_11626,N_11290);
nand U15350 (N_15350,N_9213,N_9683);
nand U15351 (N_15351,N_10454,N_11858);
nand U15352 (N_15352,N_10205,N_8687);
nor U15353 (N_15353,N_8027,N_9267);
and U15354 (N_15354,N_10475,N_11399);
and U15355 (N_15355,N_8211,N_8653);
nor U15356 (N_15356,N_10811,N_11993);
or U15357 (N_15357,N_8337,N_10985);
nand U15358 (N_15358,N_9513,N_10774);
or U15359 (N_15359,N_8877,N_10608);
and U15360 (N_15360,N_10981,N_8074);
nand U15361 (N_15361,N_11359,N_9808);
nor U15362 (N_15362,N_11733,N_9151);
and U15363 (N_15363,N_11126,N_9238);
nand U15364 (N_15364,N_9783,N_8500);
nand U15365 (N_15365,N_10977,N_10800);
or U15366 (N_15366,N_10818,N_8090);
xnor U15367 (N_15367,N_10310,N_9899);
and U15368 (N_15368,N_8061,N_10508);
nor U15369 (N_15369,N_9392,N_11564);
or U15370 (N_15370,N_11061,N_8083);
or U15371 (N_15371,N_10262,N_11233);
and U15372 (N_15372,N_8761,N_9708);
and U15373 (N_15373,N_11510,N_11421);
nand U15374 (N_15374,N_11986,N_9789);
nand U15375 (N_15375,N_11721,N_10389);
nand U15376 (N_15376,N_9290,N_11956);
nand U15377 (N_15377,N_10622,N_8423);
or U15378 (N_15378,N_8160,N_8302);
nand U15379 (N_15379,N_11653,N_8934);
nor U15380 (N_15380,N_10501,N_11639);
nand U15381 (N_15381,N_10005,N_11767);
and U15382 (N_15382,N_9182,N_10059);
and U15383 (N_15383,N_11452,N_11217);
and U15384 (N_15384,N_9421,N_11063);
and U15385 (N_15385,N_10632,N_10060);
nor U15386 (N_15386,N_11600,N_9418);
nand U15387 (N_15387,N_9374,N_10009);
and U15388 (N_15388,N_9402,N_9530);
nor U15389 (N_15389,N_10487,N_9410);
nand U15390 (N_15390,N_8434,N_10059);
and U15391 (N_15391,N_8690,N_11103);
or U15392 (N_15392,N_9329,N_10892);
and U15393 (N_15393,N_8572,N_9792);
and U15394 (N_15394,N_11522,N_8980);
nor U15395 (N_15395,N_9981,N_10301);
and U15396 (N_15396,N_9157,N_8332);
nor U15397 (N_15397,N_11729,N_9886);
nand U15398 (N_15398,N_10667,N_9730);
nand U15399 (N_15399,N_8016,N_9790);
or U15400 (N_15400,N_10129,N_8427);
nor U15401 (N_15401,N_8306,N_8816);
or U15402 (N_15402,N_10905,N_8936);
or U15403 (N_15403,N_9238,N_9071);
or U15404 (N_15404,N_10498,N_9303);
nor U15405 (N_15405,N_11450,N_10991);
nand U15406 (N_15406,N_8230,N_9222);
nand U15407 (N_15407,N_11788,N_9108);
and U15408 (N_15408,N_11794,N_11395);
nand U15409 (N_15409,N_8464,N_8884);
nand U15410 (N_15410,N_9172,N_8566);
nor U15411 (N_15411,N_11185,N_9020);
and U15412 (N_15412,N_10271,N_11569);
nand U15413 (N_15413,N_10542,N_11961);
nand U15414 (N_15414,N_8377,N_8829);
and U15415 (N_15415,N_11458,N_9052);
or U15416 (N_15416,N_9611,N_11086);
nor U15417 (N_15417,N_11344,N_9482);
nor U15418 (N_15418,N_10781,N_8510);
nand U15419 (N_15419,N_11079,N_9867);
nor U15420 (N_15420,N_10959,N_8280);
nor U15421 (N_15421,N_9861,N_11310);
and U15422 (N_15422,N_11748,N_10918);
nand U15423 (N_15423,N_10903,N_11492);
and U15424 (N_15424,N_11770,N_9824);
nor U15425 (N_15425,N_11747,N_9409);
nand U15426 (N_15426,N_11973,N_9730);
nand U15427 (N_15427,N_11841,N_9870);
and U15428 (N_15428,N_8788,N_11757);
nand U15429 (N_15429,N_11910,N_11603);
or U15430 (N_15430,N_11809,N_8143);
nor U15431 (N_15431,N_11835,N_8720);
nand U15432 (N_15432,N_10651,N_11137);
or U15433 (N_15433,N_10028,N_11838);
and U15434 (N_15434,N_9397,N_9807);
nand U15435 (N_15435,N_10493,N_11027);
nor U15436 (N_15436,N_10242,N_10033);
nor U15437 (N_15437,N_8071,N_9020);
nand U15438 (N_15438,N_8931,N_11209);
nor U15439 (N_15439,N_9196,N_10802);
nand U15440 (N_15440,N_11005,N_10544);
or U15441 (N_15441,N_11704,N_8448);
or U15442 (N_15442,N_11698,N_11108);
nand U15443 (N_15443,N_10806,N_11976);
nor U15444 (N_15444,N_11011,N_8075);
nand U15445 (N_15445,N_9761,N_9824);
nand U15446 (N_15446,N_9352,N_8139);
and U15447 (N_15447,N_10433,N_8551);
nand U15448 (N_15448,N_10438,N_10776);
and U15449 (N_15449,N_9052,N_9445);
xnor U15450 (N_15450,N_8041,N_10944);
and U15451 (N_15451,N_8422,N_11278);
or U15452 (N_15452,N_8073,N_9859);
nor U15453 (N_15453,N_10479,N_9306);
nor U15454 (N_15454,N_8578,N_10843);
nand U15455 (N_15455,N_8562,N_8061);
and U15456 (N_15456,N_9661,N_11861);
or U15457 (N_15457,N_11306,N_9013);
or U15458 (N_15458,N_10871,N_10055);
nand U15459 (N_15459,N_8369,N_11652);
nand U15460 (N_15460,N_9205,N_9387);
nand U15461 (N_15461,N_10845,N_10911);
and U15462 (N_15462,N_8415,N_9371);
nor U15463 (N_15463,N_8055,N_11400);
and U15464 (N_15464,N_11209,N_11782);
nand U15465 (N_15465,N_8602,N_11456);
and U15466 (N_15466,N_11929,N_10678);
or U15467 (N_15467,N_11663,N_9710);
nor U15468 (N_15468,N_10973,N_9309);
or U15469 (N_15469,N_8774,N_10463);
or U15470 (N_15470,N_10653,N_10009);
nor U15471 (N_15471,N_10239,N_8739);
and U15472 (N_15472,N_10342,N_10594);
and U15473 (N_15473,N_10198,N_8946);
nand U15474 (N_15474,N_10264,N_11925);
nor U15475 (N_15475,N_9792,N_8551);
or U15476 (N_15476,N_10740,N_11719);
nand U15477 (N_15477,N_8031,N_10922);
nor U15478 (N_15478,N_9081,N_10143);
and U15479 (N_15479,N_9438,N_8096);
or U15480 (N_15480,N_8786,N_10268);
nand U15481 (N_15481,N_9465,N_8439);
or U15482 (N_15482,N_8615,N_10198);
nor U15483 (N_15483,N_11995,N_11528);
or U15484 (N_15484,N_11108,N_9486);
and U15485 (N_15485,N_10986,N_10848);
or U15486 (N_15486,N_10244,N_8036);
nor U15487 (N_15487,N_11430,N_8593);
and U15488 (N_15488,N_9882,N_8872);
nand U15489 (N_15489,N_10872,N_11501);
and U15490 (N_15490,N_9198,N_8538);
nand U15491 (N_15491,N_10721,N_11626);
and U15492 (N_15492,N_9303,N_8811);
or U15493 (N_15493,N_10805,N_8539);
or U15494 (N_15494,N_11824,N_8823);
nor U15495 (N_15495,N_11663,N_9233);
nand U15496 (N_15496,N_9310,N_9179);
and U15497 (N_15497,N_10321,N_11090);
nor U15498 (N_15498,N_9555,N_10690);
nand U15499 (N_15499,N_10906,N_9603);
nand U15500 (N_15500,N_10772,N_9384);
nor U15501 (N_15501,N_11673,N_9585);
and U15502 (N_15502,N_8943,N_10079);
and U15503 (N_15503,N_8249,N_8115);
or U15504 (N_15504,N_8287,N_10048);
nor U15505 (N_15505,N_10932,N_8751);
nor U15506 (N_15506,N_10284,N_9318);
or U15507 (N_15507,N_10826,N_11744);
and U15508 (N_15508,N_11580,N_8814);
nand U15509 (N_15509,N_8064,N_9994);
nor U15510 (N_15510,N_8003,N_9745);
and U15511 (N_15511,N_10257,N_8658);
nor U15512 (N_15512,N_9171,N_10697);
and U15513 (N_15513,N_9466,N_9780);
nand U15514 (N_15514,N_8754,N_10260);
or U15515 (N_15515,N_11494,N_9663);
or U15516 (N_15516,N_11816,N_9898);
and U15517 (N_15517,N_10609,N_9911);
nor U15518 (N_15518,N_9062,N_11995);
nand U15519 (N_15519,N_9720,N_10226);
or U15520 (N_15520,N_8106,N_8244);
nor U15521 (N_15521,N_9793,N_9378);
nor U15522 (N_15522,N_9542,N_10802);
and U15523 (N_15523,N_11336,N_11736);
and U15524 (N_15524,N_9640,N_10080);
nand U15525 (N_15525,N_10904,N_10197);
nor U15526 (N_15526,N_9346,N_8550);
nand U15527 (N_15527,N_10225,N_11040);
and U15528 (N_15528,N_9130,N_11261);
and U15529 (N_15529,N_10206,N_8089);
or U15530 (N_15530,N_8313,N_8153);
and U15531 (N_15531,N_8488,N_8366);
and U15532 (N_15532,N_9649,N_9299);
and U15533 (N_15533,N_8311,N_8694);
and U15534 (N_15534,N_8485,N_10005);
and U15535 (N_15535,N_11825,N_10948);
or U15536 (N_15536,N_11038,N_8643);
nand U15537 (N_15537,N_9101,N_8328);
nand U15538 (N_15538,N_9916,N_10703);
and U15539 (N_15539,N_8696,N_10248);
nor U15540 (N_15540,N_11271,N_10520);
nand U15541 (N_15541,N_8373,N_10046);
nor U15542 (N_15542,N_10624,N_10491);
nand U15543 (N_15543,N_10021,N_9497);
or U15544 (N_15544,N_10543,N_10470);
or U15545 (N_15545,N_11460,N_8085);
nand U15546 (N_15546,N_8462,N_8325);
nand U15547 (N_15547,N_9877,N_9809);
nand U15548 (N_15548,N_11109,N_11072);
and U15549 (N_15549,N_9143,N_8618);
nand U15550 (N_15550,N_9564,N_10281);
nor U15551 (N_15551,N_11288,N_11920);
or U15552 (N_15552,N_10825,N_9191);
or U15553 (N_15553,N_8593,N_9841);
or U15554 (N_15554,N_11878,N_11732);
and U15555 (N_15555,N_9665,N_11264);
and U15556 (N_15556,N_9418,N_9927);
nor U15557 (N_15557,N_8251,N_8590);
or U15558 (N_15558,N_10982,N_8208);
and U15559 (N_15559,N_8112,N_11780);
and U15560 (N_15560,N_8531,N_10214);
nor U15561 (N_15561,N_10153,N_9489);
nor U15562 (N_15562,N_10211,N_8252);
and U15563 (N_15563,N_10925,N_9653);
nor U15564 (N_15564,N_9053,N_8273);
nand U15565 (N_15565,N_9383,N_10233);
nand U15566 (N_15566,N_9571,N_10402);
nand U15567 (N_15567,N_9962,N_8318);
or U15568 (N_15568,N_10929,N_9947);
and U15569 (N_15569,N_11970,N_8778);
nor U15570 (N_15570,N_8092,N_10184);
or U15571 (N_15571,N_11538,N_10096);
and U15572 (N_15572,N_10364,N_11756);
nand U15573 (N_15573,N_10457,N_9654);
and U15574 (N_15574,N_10775,N_10417);
or U15575 (N_15575,N_10657,N_11714);
nor U15576 (N_15576,N_11250,N_11206);
and U15577 (N_15577,N_10445,N_10780);
or U15578 (N_15578,N_11458,N_10391);
nor U15579 (N_15579,N_8516,N_11925);
or U15580 (N_15580,N_9105,N_10198);
and U15581 (N_15581,N_9462,N_10809);
xor U15582 (N_15582,N_11270,N_10936);
or U15583 (N_15583,N_8769,N_8103);
and U15584 (N_15584,N_10123,N_11402);
or U15585 (N_15585,N_10384,N_9941);
nor U15586 (N_15586,N_10338,N_9986);
and U15587 (N_15587,N_8373,N_11606);
and U15588 (N_15588,N_8910,N_9726);
and U15589 (N_15589,N_10652,N_10721);
and U15590 (N_15590,N_9509,N_9139);
nor U15591 (N_15591,N_9017,N_8226);
and U15592 (N_15592,N_11038,N_9125);
nand U15593 (N_15593,N_9500,N_9365);
or U15594 (N_15594,N_8596,N_11232);
nand U15595 (N_15595,N_9804,N_10973);
nand U15596 (N_15596,N_9066,N_10917);
nand U15597 (N_15597,N_10020,N_11327);
nor U15598 (N_15598,N_8488,N_10212);
nor U15599 (N_15599,N_11612,N_10889);
nor U15600 (N_15600,N_11859,N_11973);
nor U15601 (N_15601,N_8742,N_9880);
nand U15602 (N_15602,N_10027,N_9398);
nand U15603 (N_15603,N_11397,N_8603);
nor U15604 (N_15604,N_8389,N_8431);
nor U15605 (N_15605,N_8386,N_11015);
nand U15606 (N_15606,N_9967,N_11270);
nor U15607 (N_15607,N_11007,N_11888);
or U15608 (N_15608,N_9106,N_8547);
nand U15609 (N_15609,N_9941,N_9087);
nor U15610 (N_15610,N_10932,N_10789);
nand U15611 (N_15611,N_10152,N_9634);
and U15612 (N_15612,N_8834,N_11656);
nand U15613 (N_15613,N_9260,N_10141);
nand U15614 (N_15614,N_8197,N_11040);
or U15615 (N_15615,N_11655,N_8210);
or U15616 (N_15616,N_11328,N_8504);
nand U15617 (N_15617,N_11583,N_11664);
nor U15618 (N_15618,N_8227,N_8559);
or U15619 (N_15619,N_10788,N_9414);
and U15620 (N_15620,N_11477,N_11537);
and U15621 (N_15621,N_10870,N_11872);
nor U15622 (N_15622,N_10495,N_9873);
nand U15623 (N_15623,N_8091,N_9882);
or U15624 (N_15624,N_8014,N_9454);
or U15625 (N_15625,N_8828,N_9406);
and U15626 (N_15626,N_11247,N_11113);
nor U15627 (N_15627,N_11006,N_11104);
and U15628 (N_15628,N_10716,N_11653);
and U15629 (N_15629,N_8825,N_11186);
nand U15630 (N_15630,N_9805,N_9366);
or U15631 (N_15631,N_8415,N_8580);
nand U15632 (N_15632,N_11533,N_10267);
or U15633 (N_15633,N_8866,N_8405);
and U15634 (N_15634,N_9770,N_11306);
nor U15635 (N_15635,N_10338,N_10827);
nand U15636 (N_15636,N_11777,N_10075);
or U15637 (N_15637,N_8720,N_11475);
nor U15638 (N_15638,N_9234,N_11245);
nor U15639 (N_15639,N_11515,N_10549);
nand U15640 (N_15640,N_11098,N_11085);
nand U15641 (N_15641,N_9580,N_10991);
and U15642 (N_15642,N_9849,N_9784);
nand U15643 (N_15643,N_11544,N_10573);
nand U15644 (N_15644,N_11998,N_10603);
nand U15645 (N_15645,N_10162,N_9746);
or U15646 (N_15646,N_10777,N_9266);
or U15647 (N_15647,N_11944,N_10301);
and U15648 (N_15648,N_11522,N_8279);
and U15649 (N_15649,N_8425,N_8872);
nor U15650 (N_15650,N_9632,N_10352);
nor U15651 (N_15651,N_10543,N_8821);
and U15652 (N_15652,N_10148,N_8864);
nand U15653 (N_15653,N_11697,N_11653);
and U15654 (N_15654,N_8977,N_11233);
and U15655 (N_15655,N_10902,N_10562);
nand U15656 (N_15656,N_11188,N_11535);
and U15657 (N_15657,N_9923,N_11059);
nand U15658 (N_15658,N_11432,N_9313);
or U15659 (N_15659,N_10973,N_10193);
or U15660 (N_15660,N_10482,N_9315);
nor U15661 (N_15661,N_9056,N_11901);
nor U15662 (N_15662,N_9292,N_11306);
nor U15663 (N_15663,N_9005,N_9631);
nand U15664 (N_15664,N_9788,N_8284);
or U15665 (N_15665,N_9799,N_9343);
nand U15666 (N_15666,N_9374,N_10776);
nor U15667 (N_15667,N_11009,N_11668);
and U15668 (N_15668,N_11736,N_11092);
and U15669 (N_15669,N_11253,N_8446);
and U15670 (N_15670,N_10206,N_10850);
nand U15671 (N_15671,N_10819,N_9342);
and U15672 (N_15672,N_8787,N_11361);
or U15673 (N_15673,N_11583,N_9102);
nor U15674 (N_15674,N_10822,N_8904);
and U15675 (N_15675,N_9288,N_9355);
and U15676 (N_15676,N_10378,N_8623);
nand U15677 (N_15677,N_10440,N_11836);
nand U15678 (N_15678,N_10049,N_9325);
and U15679 (N_15679,N_8240,N_8486);
and U15680 (N_15680,N_8959,N_8681);
and U15681 (N_15681,N_10100,N_9519);
nand U15682 (N_15682,N_9408,N_11927);
nand U15683 (N_15683,N_11676,N_11273);
xnor U15684 (N_15684,N_9992,N_11006);
and U15685 (N_15685,N_11962,N_9537);
nand U15686 (N_15686,N_9904,N_11247);
nor U15687 (N_15687,N_10819,N_11070);
and U15688 (N_15688,N_9296,N_10758);
nand U15689 (N_15689,N_10338,N_8558);
nor U15690 (N_15690,N_10566,N_8619);
nand U15691 (N_15691,N_8656,N_11366);
nor U15692 (N_15692,N_8010,N_11283);
or U15693 (N_15693,N_8356,N_9592);
xor U15694 (N_15694,N_9063,N_8241);
nand U15695 (N_15695,N_10105,N_11455);
or U15696 (N_15696,N_10170,N_10388);
and U15697 (N_15697,N_11585,N_10930);
and U15698 (N_15698,N_10423,N_9070);
and U15699 (N_15699,N_10185,N_10153);
nand U15700 (N_15700,N_8680,N_9284);
nand U15701 (N_15701,N_8248,N_11503);
nor U15702 (N_15702,N_10009,N_9442);
and U15703 (N_15703,N_11535,N_11897);
and U15704 (N_15704,N_9301,N_8402);
nor U15705 (N_15705,N_10602,N_11861);
nor U15706 (N_15706,N_10419,N_11509);
nor U15707 (N_15707,N_11639,N_11673);
and U15708 (N_15708,N_8134,N_11672);
nor U15709 (N_15709,N_10182,N_10643);
nor U15710 (N_15710,N_11246,N_10278);
and U15711 (N_15711,N_8462,N_8715);
and U15712 (N_15712,N_11413,N_9951);
nor U15713 (N_15713,N_10626,N_8767);
and U15714 (N_15714,N_8014,N_9963);
nand U15715 (N_15715,N_8532,N_8708);
nor U15716 (N_15716,N_8030,N_8192);
or U15717 (N_15717,N_9903,N_10480);
or U15718 (N_15718,N_9154,N_11146);
nor U15719 (N_15719,N_11069,N_8006);
or U15720 (N_15720,N_10387,N_9725);
nand U15721 (N_15721,N_8514,N_10959);
nand U15722 (N_15722,N_10522,N_10499);
nand U15723 (N_15723,N_8728,N_8753);
or U15724 (N_15724,N_10754,N_9558);
nand U15725 (N_15725,N_10657,N_9045);
nor U15726 (N_15726,N_11760,N_10639);
and U15727 (N_15727,N_9400,N_11655);
or U15728 (N_15728,N_11339,N_8436);
nor U15729 (N_15729,N_10675,N_9345);
or U15730 (N_15730,N_8522,N_10530);
nand U15731 (N_15731,N_10378,N_11098);
and U15732 (N_15732,N_8125,N_10443);
and U15733 (N_15733,N_9112,N_9496);
and U15734 (N_15734,N_11683,N_10098);
nand U15735 (N_15735,N_9177,N_9060);
and U15736 (N_15736,N_8459,N_11107);
or U15737 (N_15737,N_9134,N_9669);
nor U15738 (N_15738,N_11763,N_8594);
or U15739 (N_15739,N_8245,N_10498);
or U15740 (N_15740,N_11085,N_10135);
nor U15741 (N_15741,N_10353,N_11197);
or U15742 (N_15742,N_11465,N_11708);
and U15743 (N_15743,N_10814,N_11933);
or U15744 (N_15744,N_10555,N_10739);
nor U15745 (N_15745,N_8744,N_10816);
xnor U15746 (N_15746,N_10459,N_11676);
and U15747 (N_15747,N_10217,N_9045);
or U15748 (N_15748,N_11270,N_8600);
nand U15749 (N_15749,N_8216,N_11494);
nand U15750 (N_15750,N_10776,N_8051);
nand U15751 (N_15751,N_8022,N_9014);
or U15752 (N_15752,N_9271,N_10279);
and U15753 (N_15753,N_11714,N_8717);
nand U15754 (N_15754,N_8490,N_8545);
or U15755 (N_15755,N_9548,N_10863);
and U15756 (N_15756,N_11010,N_11512);
nand U15757 (N_15757,N_9334,N_11081);
nand U15758 (N_15758,N_10769,N_8097);
nand U15759 (N_15759,N_11537,N_11628);
or U15760 (N_15760,N_9706,N_8830);
nor U15761 (N_15761,N_10926,N_11395);
or U15762 (N_15762,N_8702,N_9617);
nand U15763 (N_15763,N_10786,N_11227);
and U15764 (N_15764,N_8738,N_10710);
nor U15765 (N_15765,N_11160,N_9762);
xor U15766 (N_15766,N_9117,N_9500);
or U15767 (N_15767,N_11905,N_11285);
and U15768 (N_15768,N_9234,N_9089);
or U15769 (N_15769,N_8479,N_10245);
or U15770 (N_15770,N_8439,N_10210);
or U15771 (N_15771,N_11692,N_9475);
nand U15772 (N_15772,N_10178,N_11007);
and U15773 (N_15773,N_8974,N_10324);
and U15774 (N_15774,N_9613,N_10410);
or U15775 (N_15775,N_9741,N_8680);
nor U15776 (N_15776,N_10681,N_9380);
nor U15777 (N_15777,N_9096,N_8238);
nor U15778 (N_15778,N_9192,N_10145);
or U15779 (N_15779,N_9978,N_10578);
and U15780 (N_15780,N_8605,N_11291);
nand U15781 (N_15781,N_10990,N_10864);
and U15782 (N_15782,N_11218,N_11763);
or U15783 (N_15783,N_8751,N_10704);
xor U15784 (N_15784,N_8213,N_8099);
or U15785 (N_15785,N_10644,N_9216);
and U15786 (N_15786,N_10407,N_10537);
xnor U15787 (N_15787,N_11314,N_11459);
or U15788 (N_15788,N_9333,N_11122);
nor U15789 (N_15789,N_9449,N_11406);
nor U15790 (N_15790,N_9062,N_8113);
nor U15791 (N_15791,N_9245,N_11815);
and U15792 (N_15792,N_9577,N_8251);
nor U15793 (N_15793,N_11815,N_9446);
or U15794 (N_15794,N_8098,N_8584);
nand U15795 (N_15795,N_11563,N_11222);
nand U15796 (N_15796,N_10578,N_11287);
and U15797 (N_15797,N_8174,N_10303);
nand U15798 (N_15798,N_11737,N_8181);
nand U15799 (N_15799,N_11709,N_9997);
nor U15800 (N_15800,N_11604,N_11386);
nor U15801 (N_15801,N_8211,N_11817);
nand U15802 (N_15802,N_9413,N_8699);
nor U15803 (N_15803,N_10145,N_10648);
nand U15804 (N_15804,N_9115,N_10115);
nand U15805 (N_15805,N_9506,N_10717);
and U15806 (N_15806,N_11073,N_9896);
and U15807 (N_15807,N_10559,N_11489);
or U15808 (N_15808,N_9909,N_10871);
and U15809 (N_15809,N_9530,N_10500);
or U15810 (N_15810,N_9349,N_10800);
or U15811 (N_15811,N_8394,N_10051);
or U15812 (N_15812,N_11049,N_11885);
nand U15813 (N_15813,N_11713,N_9873);
xor U15814 (N_15814,N_9708,N_8368);
or U15815 (N_15815,N_8281,N_9026);
nor U15816 (N_15816,N_11974,N_9682);
nor U15817 (N_15817,N_9987,N_10100);
nor U15818 (N_15818,N_9390,N_10071);
nand U15819 (N_15819,N_9403,N_8292);
and U15820 (N_15820,N_9351,N_8395);
nor U15821 (N_15821,N_8025,N_10621);
nor U15822 (N_15822,N_9950,N_8562);
nand U15823 (N_15823,N_8204,N_10392);
xor U15824 (N_15824,N_11096,N_10198);
and U15825 (N_15825,N_9272,N_11274);
or U15826 (N_15826,N_11828,N_9848);
nand U15827 (N_15827,N_8324,N_11235);
and U15828 (N_15828,N_11393,N_9059);
nor U15829 (N_15829,N_8001,N_11438);
or U15830 (N_15830,N_9005,N_11244);
nor U15831 (N_15831,N_9297,N_10567);
or U15832 (N_15832,N_8790,N_10135);
nand U15833 (N_15833,N_10805,N_10638);
nor U15834 (N_15834,N_9345,N_8261);
nand U15835 (N_15835,N_11659,N_8653);
and U15836 (N_15836,N_8925,N_8020);
nor U15837 (N_15837,N_11060,N_10168);
nor U15838 (N_15838,N_11813,N_8523);
or U15839 (N_15839,N_9334,N_8092);
nor U15840 (N_15840,N_8287,N_10321);
and U15841 (N_15841,N_8243,N_11624);
and U15842 (N_15842,N_9678,N_10423);
or U15843 (N_15843,N_11856,N_10325);
or U15844 (N_15844,N_9866,N_9674);
nand U15845 (N_15845,N_9507,N_10550);
or U15846 (N_15846,N_8526,N_11000);
nand U15847 (N_15847,N_9553,N_8589);
and U15848 (N_15848,N_8007,N_8548);
or U15849 (N_15849,N_9127,N_10126);
nor U15850 (N_15850,N_9724,N_8825);
or U15851 (N_15851,N_9288,N_8199);
nand U15852 (N_15852,N_9203,N_11262);
nand U15853 (N_15853,N_8056,N_10470);
and U15854 (N_15854,N_10649,N_11692);
or U15855 (N_15855,N_8435,N_8720);
nand U15856 (N_15856,N_8324,N_10423);
nor U15857 (N_15857,N_10468,N_9548);
or U15858 (N_15858,N_11808,N_10641);
and U15859 (N_15859,N_11592,N_10676);
nand U15860 (N_15860,N_8981,N_11410);
nand U15861 (N_15861,N_10439,N_10620);
and U15862 (N_15862,N_10514,N_11513);
nand U15863 (N_15863,N_10115,N_9662);
and U15864 (N_15864,N_9163,N_10263);
and U15865 (N_15865,N_9158,N_9531);
nand U15866 (N_15866,N_8136,N_8628);
nand U15867 (N_15867,N_11544,N_8877);
and U15868 (N_15868,N_10878,N_11104);
nand U15869 (N_15869,N_9401,N_8637);
nand U15870 (N_15870,N_8956,N_11739);
nor U15871 (N_15871,N_10200,N_8040);
nand U15872 (N_15872,N_8288,N_11307);
or U15873 (N_15873,N_9643,N_10509);
and U15874 (N_15874,N_8417,N_8960);
or U15875 (N_15875,N_9113,N_10712);
nand U15876 (N_15876,N_10107,N_11416);
nor U15877 (N_15877,N_9454,N_8915);
nand U15878 (N_15878,N_8157,N_9413);
and U15879 (N_15879,N_10018,N_10642);
nor U15880 (N_15880,N_10064,N_10542);
or U15881 (N_15881,N_8387,N_11190);
nor U15882 (N_15882,N_8337,N_10522);
nor U15883 (N_15883,N_8986,N_11797);
or U15884 (N_15884,N_9998,N_10965);
or U15885 (N_15885,N_11958,N_9468);
and U15886 (N_15886,N_11316,N_10036);
or U15887 (N_15887,N_10432,N_8336);
and U15888 (N_15888,N_9106,N_8206);
nand U15889 (N_15889,N_8340,N_10789);
nor U15890 (N_15890,N_9285,N_10045);
nand U15891 (N_15891,N_10793,N_11742);
nand U15892 (N_15892,N_10194,N_8067);
nand U15893 (N_15893,N_8573,N_10541);
nand U15894 (N_15894,N_10201,N_8659);
nand U15895 (N_15895,N_10052,N_11307);
or U15896 (N_15896,N_10404,N_8548);
or U15897 (N_15897,N_8496,N_10672);
and U15898 (N_15898,N_8971,N_10702);
or U15899 (N_15899,N_11465,N_9273);
or U15900 (N_15900,N_9419,N_9276);
nor U15901 (N_15901,N_11880,N_8391);
nor U15902 (N_15902,N_9397,N_11532);
nand U15903 (N_15903,N_8594,N_10275);
nand U15904 (N_15904,N_9258,N_10759);
or U15905 (N_15905,N_9214,N_11688);
nor U15906 (N_15906,N_11416,N_10377);
nor U15907 (N_15907,N_10374,N_8930);
and U15908 (N_15908,N_9902,N_8830);
nor U15909 (N_15909,N_9291,N_11759);
or U15910 (N_15910,N_11734,N_10817);
xnor U15911 (N_15911,N_9715,N_8129);
and U15912 (N_15912,N_11115,N_8224);
or U15913 (N_15913,N_9067,N_10131);
or U15914 (N_15914,N_11324,N_9284);
or U15915 (N_15915,N_10822,N_8340);
nand U15916 (N_15916,N_10829,N_11222);
nor U15917 (N_15917,N_10810,N_9623);
nor U15918 (N_15918,N_11961,N_9243);
and U15919 (N_15919,N_8716,N_8481);
nand U15920 (N_15920,N_9922,N_10563);
nor U15921 (N_15921,N_11612,N_11313);
nor U15922 (N_15922,N_8251,N_10875);
nand U15923 (N_15923,N_11514,N_8173);
or U15924 (N_15924,N_10254,N_8327);
or U15925 (N_15925,N_9057,N_10816);
nor U15926 (N_15926,N_10416,N_8088);
and U15927 (N_15927,N_11639,N_11584);
and U15928 (N_15928,N_9919,N_10619);
nor U15929 (N_15929,N_10865,N_8147);
and U15930 (N_15930,N_11995,N_9040);
or U15931 (N_15931,N_8411,N_9821);
nor U15932 (N_15932,N_10750,N_8014);
or U15933 (N_15933,N_10002,N_11876);
nand U15934 (N_15934,N_10514,N_9895);
nor U15935 (N_15935,N_8561,N_8730);
or U15936 (N_15936,N_11349,N_9434);
nor U15937 (N_15937,N_8455,N_10468);
nand U15938 (N_15938,N_9659,N_8393);
or U15939 (N_15939,N_10681,N_8270);
xor U15940 (N_15940,N_8620,N_10342);
nand U15941 (N_15941,N_11301,N_8158);
nor U15942 (N_15942,N_9281,N_11602);
nand U15943 (N_15943,N_9801,N_10661);
nor U15944 (N_15944,N_9554,N_9081);
and U15945 (N_15945,N_9079,N_11435);
and U15946 (N_15946,N_11334,N_8024);
nor U15947 (N_15947,N_11257,N_11005);
nor U15948 (N_15948,N_9417,N_10087);
nand U15949 (N_15949,N_10082,N_9754);
nand U15950 (N_15950,N_8433,N_8462);
nor U15951 (N_15951,N_8880,N_9512);
nor U15952 (N_15952,N_10543,N_8635);
or U15953 (N_15953,N_11087,N_8116);
nand U15954 (N_15954,N_8147,N_9027);
and U15955 (N_15955,N_11599,N_11773);
nor U15956 (N_15956,N_8534,N_10027);
and U15957 (N_15957,N_10380,N_9655);
or U15958 (N_15958,N_8927,N_10208);
or U15959 (N_15959,N_10821,N_11812);
and U15960 (N_15960,N_11490,N_8318);
nand U15961 (N_15961,N_10675,N_11999);
nor U15962 (N_15962,N_10715,N_8074);
nand U15963 (N_15963,N_10732,N_9424);
nand U15964 (N_15964,N_10928,N_11500);
nor U15965 (N_15965,N_9035,N_9120);
or U15966 (N_15966,N_9196,N_10876);
and U15967 (N_15967,N_10331,N_10542);
and U15968 (N_15968,N_8577,N_10073);
nand U15969 (N_15969,N_11879,N_11306);
nor U15970 (N_15970,N_8033,N_8137);
and U15971 (N_15971,N_11490,N_11344);
nor U15972 (N_15972,N_11238,N_8063);
and U15973 (N_15973,N_9726,N_9513);
xnor U15974 (N_15974,N_9690,N_8107);
or U15975 (N_15975,N_10684,N_8666);
xnor U15976 (N_15976,N_8538,N_8774);
or U15977 (N_15977,N_10569,N_10126);
and U15978 (N_15978,N_11047,N_10798);
and U15979 (N_15979,N_8936,N_9372);
nand U15980 (N_15980,N_9368,N_11431);
nor U15981 (N_15981,N_11641,N_10185);
nand U15982 (N_15982,N_8479,N_11313);
nor U15983 (N_15983,N_8738,N_10190);
and U15984 (N_15984,N_10326,N_8201);
and U15985 (N_15985,N_9335,N_10970);
nand U15986 (N_15986,N_9087,N_9791);
nand U15987 (N_15987,N_10828,N_8224);
nand U15988 (N_15988,N_10494,N_9592);
and U15989 (N_15989,N_9079,N_8381);
nand U15990 (N_15990,N_9862,N_10855);
nand U15991 (N_15991,N_11295,N_11518);
nand U15992 (N_15992,N_11144,N_10274);
nand U15993 (N_15993,N_8987,N_8150);
nor U15994 (N_15994,N_10062,N_8527);
nand U15995 (N_15995,N_8086,N_11861);
and U15996 (N_15996,N_10548,N_9375);
nor U15997 (N_15997,N_8011,N_11060);
nand U15998 (N_15998,N_11177,N_11877);
nor U15999 (N_15999,N_10260,N_8749);
nor U16000 (N_16000,N_15176,N_13722);
nand U16001 (N_16001,N_15812,N_15454);
and U16002 (N_16002,N_15253,N_15047);
nand U16003 (N_16003,N_14299,N_15592);
nor U16004 (N_16004,N_12939,N_14185);
nand U16005 (N_16005,N_14300,N_15843);
nor U16006 (N_16006,N_15219,N_12750);
nor U16007 (N_16007,N_14787,N_13400);
and U16008 (N_16008,N_15094,N_13796);
or U16009 (N_16009,N_15603,N_12028);
and U16010 (N_16010,N_14292,N_15002);
or U16011 (N_16011,N_15408,N_13290);
nor U16012 (N_16012,N_15144,N_14397);
nor U16013 (N_16013,N_15652,N_12607);
nand U16014 (N_16014,N_12634,N_12370);
nand U16015 (N_16015,N_15245,N_14626);
or U16016 (N_16016,N_12139,N_13074);
and U16017 (N_16017,N_12424,N_12996);
and U16018 (N_16018,N_15829,N_12371);
and U16019 (N_16019,N_15528,N_12391);
nor U16020 (N_16020,N_13735,N_15788);
nand U16021 (N_16021,N_13712,N_12372);
or U16022 (N_16022,N_14865,N_12853);
nor U16023 (N_16023,N_15383,N_13416);
nand U16024 (N_16024,N_13525,N_13921);
and U16025 (N_16025,N_13833,N_13164);
nor U16026 (N_16026,N_15612,N_13345);
xor U16027 (N_16027,N_12809,N_13111);
nor U16028 (N_16028,N_15581,N_12074);
and U16029 (N_16029,N_15618,N_12163);
nand U16030 (N_16030,N_14301,N_15049);
and U16031 (N_16031,N_15388,N_14168);
nor U16032 (N_16032,N_13101,N_12116);
or U16033 (N_16033,N_12223,N_15835);
and U16034 (N_16034,N_12460,N_13113);
and U16035 (N_16035,N_15319,N_14765);
nor U16036 (N_16036,N_15071,N_12127);
nand U16037 (N_16037,N_15860,N_15923);
or U16038 (N_16038,N_13421,N_15789);
or U16039 (N_16039,N_14181,N_15819);
nand U16040 (N_16040,N_14536,N_12967);
nor U16041 (N_16041,N_12664,N_14226);
or U16042 (N_16042,N_13397,N_12350);
and U16043 (N_16043,N_12388,N_15839);
nand U16044 (N_16044,N_14955,N_14766);
nor U16045 (N_16045,N_14323,N_12494);
nor U16046 (N_16046,N_13570,N_13083);
or U16047 (N_16047,N_13269,N_14574);
nand U16048 (N_16048,N_12037,N_12616);
nor U16049 (N_16049,N_14072,N_14751);
nor U16050 (N_16050,N_15854,N_12364);
and U16051 (N_16051,N_15223,N_15595);
nand U16052 (N_16052,N_13087,N_14875);
nand U16053 (N_16053,N_14690,N_14704);
nor U16054 (N_16054,N_13254,N_12246);
or U16055 (N_16055,N_12457,N_13537);
nand U16056 (N_16056,N_14159,N_15302);
and U16057 (N_16057,N_15748,N_14519);
or U16058 (N_16058,N_15763,N_14268);
or U16059 (N_16059,N_14885,N_13190);
or U16060 (N_16060,N_13834,N_13612);
nor U16061 (N_16061,N_12896,N_13985);
or U16062 (N_16062,N_12727,N_14694);
or U16063 (N_16063,N_13774,N_13931);
nor U16064 (N_16064,N_13408,N_13470);
and U16065 (N_16065,N_14145,N_14763);
and U16066 (N_16066,N_12486,N_12373);
nor U16067 (N_16067,N_12908,N_15548);
nand U16068 (N_16068,N_13749,N_14971);
nor U16069 (N_16069,N_15869,N_12635);
nor U16070 (N_16070,N_12061,N_14812);
nand U16071 (N_16071,N_14054,N_12331);
or U16072 (N_16072,N_14647,N_12319);
or U16073 (N_16073,N_12324,N_15434);
or U16074 (N_16074,N_13285,N_13339);
and U16075 (N_16075,N_13468,N_12518);
nand U16076 (N_16076,N_14798,N_15879);
nand U16077 (N_16077,N_14102,N_12277);
and U16078 (N_16078,N_15042,N_14863);
or U16079 (N_16079,N_14628,N_12636);
or U16080 (N_16080,N_12320,N_12829);
and U16081 (N_16081,N_13532,N_14212);
nor U16082 (N_16082,N_14051,N_15754);
nor U16083 (N_16083,N_14516,N_15721);
or U16084 (N_16084,N_12733,N_12591);
and U16085 (N_16085,N_12304,N_14517);
or U16086 (N_16086,N_15944,N_15397);
nor U16087 (N_16087,N_15191,N_15582);
or U16088 (N_16088,N_14119,N_12793);
or U16089 (N_16089,N_13337,N_15145);
or U16090 (N_16090,N_13714,N_12870);
and U16091 (N_16091,N_13271,N_15705);
or U16092 (N_16092,N_12416,N_15289);
nor U16093 (N_16093,N_13179,N_15782);
or U16094 (N_16094,N_13205,N_13106);
and U16095 (N_16095,N_12489,N_14353);
and U16096 (N_16096,N_14316,N_12792);
nor U16097 (N_16097,N_14289,N_12479);
xor U16098 (N_16098,N_12260,N_14629);
nand U16099 (N_16099,N_15585,N_15804);
nand U16100 (N_16100,N_12671,N_12195);
and U16101 (N_16101,N_13255,N_14553);
or U16102 (N_16102,N_12004,N_13375);
nand U16103 (N_16103,N_15858,N_13218);
and U16104 (N_16104,N_15294,N_15960);
nand U16105 (N_16105,N_14393,N_13697);
nand U16106 (N_16106,N_14936,N_13309);
nand U16107 (N_16107,N_12578,N_12965);
or U16108 (N_16108,N_12643,N_14200);
or U16109 (N_16109,N_12267,N_14919);
and U16110 (N_16110,N_14350,N_12527);
nand U16111 (N_16111,N_14252,N_12913);
and U16112 (N_16112,N_15014,N_13303);
or U16113 (N_16113,N_13755,N_15363);
nor U16114 (N_16114,N_14201,N_14917);
or U16115 (N_16115,N_14696,N_14741);
nor U16116 (N_16116,N_14828,N_14439);
or U16117 (N_16117,N_13093,N_14387);
nand U16118 (N_16118,N_15416,N_13549);
or U16119 (N_16119,N_12042,N_14005);
nand U16120 (N_16120,N_14986,N_14213);
nand U16121 (N_16121,N_15221,N_13913);
nand U16122 (N_16122,N_14240,N_13778);
nor U16123 (N_16123,N_14153,N_15569);
and U16124 (N_16124,N_15951,N_14154);
xnor U16125 (N_16125,N_14758,N_15903);
nand U16126 (N_16126,N_15136,N_13431);
or U16127 (N_16127,N_14872,N_12014);
and U16128 (N_16128,N_13624,N_13464);
nor U16129 (N_16129,N_14110,N_13999);
and U16130 (N_16130,N_12013,N_12261);
nor U16131 (N_16131,N_15064,N_15532);
and U16132 (N_16132,N_12086,N_14882);
nand U16133 (N_16133,N_14113,N_14537);
nand U16134 (N_16134,N_14555,N_15072);
and U16135 (N_16135,N_14134,N_15674);
and U16136 (N_16136,N_14265,N_13601);
nand U16137 (N_16137,N_14898,N_13091);
and U16138 (N_16138,N_12642,N_15729);
nor U16139 (N_16139,N_14438,N_15965);
nor U16140 (N_16140,N_14379,N_15163);
nand U16141 (N_16141,N_13950,N_14480);
nand U16142 (N_16142,N_13306,N_12406);
nor U16143 (N_16143,N_14257,N_15719);
nand U16144 (N_16144,N_12748,N_15124);
or U16145 (N_16145,N_15432,N_13635);
nor U16146 (N_16146,N_12485,N_15076);
or U16147 (N_16147,N_15403,N_15392);
nand U16148 (N_16148,N_13591,N_12194);
or U16149 (N_16149,N_15095,N_14884);
nor U16150 (N_16150,N_15957,N_12933);
and U16151 (N_16151,N_15778,N_14707);
nor U16152 (N_16152,N_13890,N_14891);
and U16153 (N_16153,N_14640,N_13978);
nor U16154 (N_16154,N_14368,N_13895);
nor U16155 (N_16155,N_14067,N_14907);
and U16156 (N_16156,N_13391,N_13676);
nor U16157 (N_16157,N_14246,N_12492);
nor U16158 (N_16158,N_12383,N_13486);
nand U16159 (N_16159,N_15430,N_14311);
and U16160 (N_16160,N_13594,N_15650);
or U16161 (N_16161,N_15629,N_15779);
or U16162 (N_16162,N_13264,N_15620);
and U16163 (N_16163,N_13509,N_14006);
nor U16164 (N_16164,N_12926,N_12640);
or U16165 (N_16165,N_14395,N_12690);
nor U16166 (N_16166,N_13172,N_14278);
nand U16167 (N_16167,N_13905,N_15513);
nand U16168 (N_16168,N_15972,N_12230);
nand U16169 (N_16169,N_14254,N_14730);
or U16170 (N_16170,N_12624,N_14531);
or U16171 (N_16171,N_14981,N_12335);
nand U16172 (N_16172,N_12393,N_13744);
nor U16173 (N_16173,N_12120,N_12081);
nor U16174 (N_16174,N_15898,N_14927);
or U16175 (N_16175,N_14799,N_13129);
nor U16176 (N_16176,N_13283,N_15011);
or U16177 (N_16177,N_15060,N_15129);
and U16178 (N_16178,N_14992,N_14816);
nor U16179 (N_16179,N_15375,N_14792);
xnor U16180 (N_16180,N_12645,N_13387);
or U16181 (N_16181,N_15613,N_15417);
nor U16182 (N_16182,N_14048,N_15662);
or U16183 (N_16183,N_12265,N_15406);
or U16184 (N_16184,N_13515,N_15648);
nor U16185 (N_16185,N_15287,N_12274);
and U16186 (N_16186,N_12975,N_12715);
and U16187 (N_16187,N_14139,N_14859);
nand U16188 (N_16188,N_15596,N_12171);
nor U16189 (N_16189,N_15633,N_15006);
nor U16190 (N_16190,N_15797,N_13415);
or U16191 (N_16191,N_14222,N_12475);
nand U16192 (N_16192,N_15982,N_15916);
and U16193 (N_16193,N_15959,N_15946);
or U16194 (N_16194,N_12558,N_14564);
nand U16195 (N_16195,N_13148,N_15225);
or U16196 (N_16196,N_13210,N_14060);
and U16197 (N_16197,N_13141,N_15828);
nor U16198 (N_16198,N_15493,N_15050);
and U16199 (N_16199,N_13865,N_14235);
nand U16200 (N_16200,N_12576,N_12875);
nor U16201 (N_16201,N_12336,N_12509);
nor U16202 (N_16202,N_13260,N_14312);
or U16203 (N_16203,N_12654,N_14476);
or U16204 (N_16204,N_13144,N_15233);
and U16205 (N_16205,N_13351,N_15004);
and U16206 (N_16206,N_15267,N_15382);
nand U16207 (N_16207,N_12849,N_15504);
nor U16208 (N_16208,N_15669,N_14321);
nand U16209 (N_16209,N_15948,N_15731);
and U16210 (N_16210,N_15000,N_14520);
and U16211 (N_16211,N_13672,N_12556);
and U16212 (N_16212,N_13632,N_13114);
or U16213 (N_16213,N_15832,N_15987);
and U16214 (N_16214,N_14179,N_13763);
and U16215 (N_16215,N_15085,N_14893);
and U16216 (N_16216,N_14295,N_14877);
and U16217 (N_16217,N_15676,N_14601);
nand U16218 (N_16218,N_12621,N_12856);
and U16219 (N_16219,N_15553,N_13851);
or U16220 (N_16220,N_12029,N_13568);
nand U16221 (N_16221,N_12780,N_14967);
nand U16222 (N_16222,N_13495,N_14302);
and U16223 (N_16223,N_14774,N_12831);
nor U16224 (N_16224,N_14619,N_13687);
and U16225 (N_16225,N_12857,N_13282);
nand U16226 (N_16226,N_13108,N_13636);
nor U16227 (N_16227,N_13498,N_14495);
and U16228 (N_16228,N_12278,N_15706);
nand U16229 (N_16229,N_13385,N_13068);
and U16230 (N_16230,N_14053,N_13551);
nor U16231 (N_16231,N_12765,N_13473);
xor U16232 (N_16232,N_14627,N_13821);
or U16233 (N_16233,N_12135,N_15580);
and U16234 (N_16234,N_13906,N_14140);
and U16235 (N_16235,N_15475,N_14750);
nor U16236 (N_16236,N_15820,N_14988);
nand U16237 (N_16237,N_14572,N_12234);
nor U16238 (N_16238,N_13628,N_14016);
nand U16239 (N_16239,N_13945,N_12960);
nor U16240 (N_16240,N_13469,N_15758);
and U16241 (N_16241,N_14605,N_12840);
nand U16242 (N_16242,N_14160,N_15838);
nor U16243 (N_16243,N_14983,N_12145);
and U16244 (N_16244,N_14366,N_12667);
or U16245 (N_16245,N_12528,N_15378);
or U16246 (N_16246,N_13969,N_14015);
nand U16247 (N_16247,N_15907,N_13328);
nor U16248 (N_16248,N_12451,N_15542);
nand U16249 (N_16249,N_13747,N_14237);
nor U16250 (N_16250,N_12264,N_12893);
or U16251 (N_16251,N_13530,N_13586);
or U16252 (N_16252,N_14421,N_13758);
or U16253 (N_16253,N_14184,N_15703);
or U16254 (N_16254,N_13727,N_12892);
nand U16255 (N_16255,N_13364,N_12627);
and U16256 (N_16256,N_12103,N_15490);
nor U16257 (N_16257,N_12961,N_14683);
and U16258 (N_16258,N_14633,N_14271);
nand U16259 (N_16259,N_13948,N_15059);
and U16260 (N_16260,N_14337,N_14288);
and U16261 (N_16261,N_15340,N_13675);
nor U16262 (N_16262,N_12015,N_15936);
nand U16263 (N_16263,N_13152,N_14535);
xor U16264 (N_16264,N_15451,N_13317);
nor U16265 (N_16265,N_13053,N_12532);
nor U16266 (N_16266,N_12085,N_12186);
or U16267 (N_16267,N_13380,N_12844);
or U16268 (N_16268,N_12073,N_12589);
and U16269 (N_16269,N_12096,N_14611);
or U16270 (N_16270,N_13962,N_14442);
and U16271 (N_16271,N_12779,N_13867);
nor U16272 (N_16272,N_14786,N_14406);
nor U16273 (N_16273,N_14415,N_15376);
and U16274 (N_16274,N_12041,N_14563);
nor U16275 (N_16275,N_15154,N_12988);
nand U16276 (N_16276,N_14019,N_14597);
nor U16277 (N_16277,N_12531,N_14881);
or U16278 (N_16278,N_15529,N_13147);
nor U16279 (N_16279,N_13599,N_13668);
and U16280 (N_16280,N_12330,N_15237);
nor U16281 (N_16281,N_13573,N_13544);
and U16282 (N_16282,N_12858,N_15422);
nand U16283 (N_16283,N_13363,N_13926);
nand U16284 (N_16284,N_14229,N_14162);
and U16285 (N_16285,N_13811,N_12030);
nor U16286 (N_16286,N_13968,N_15764);
and U16287 (N_16287,N_13826,N_14959);
or U16288 (N_16288,N_14409,N_13557);
and U16289 (N_16289,N_14701,N_13349);
and U16290 (N_16290,N_14469,N_13428);
and U16291 (N_16291,N_15512,N_12266);
and U16292 (N_16292,N_15279,N_14042);
and U16293 (N_16293,N_15536,N_12498);
or U16294 (N_16294,N_12932,N_14194);
xnor U16295 (N_16295,N_14214,N_12409);
nand U16296 (N_16296,N_12429,N_12731);
and U16297 (N_16297,N_12414,N_12470);
or U16298 (N_16298,N_13889,N_12698);
xor U16299 (N_16299,N_12403,N_15332);
or U16300 (N_16300,N_13874,N_15455);
or U16301 (N_16301,N_12900,N_13578);
nor U16302 (N_16302,N_13281,N_14324);
nor U16303 (N_16303,N_14565,N_14455);
and U16304 (N_16304,N_13947,N_13606);
and U16305 (N_16305,N_15681,N_13278);
nor U16306 (N_16306,N_14192,N_14784);
or U16307 (N_16307,N_12365,N_12435);
or U16308 (N_16308,N_13572,N_15278);
and U16309 (N_16309,N_13063,N_12231);
nor U16310 (N_16310,N_14909,N_12174);
or U16311 (N_16311,N_15762,N_15414);
or U16312 (N_16312,N_13365,N_13604);
or U16313 (N_16313,N_15649,N_13453);
nand U16314 (N_16314,N_15808,N_13079);
nor U16315 (N_16315,N_12399,N_13237);
nor U16316 (N_16316,N_14720,N_12738);
nor U16317 (N_16317,N_13801,N_15105);
nand U16318 (N_16318,N_12024,N_13550);
nor U16319 (N_16319,N_15367,N_14030);
and U16320 (N_16320,N_12561,N_14270);
or U16321 (N_16321,N_13886,N_15335);
nand U16322 (N_16322,N_14583,N_13772);
or U16323 (N_16323,N_14167,N_13018);
nand U16324 (N_16324,N_12128,N_14620);
nand U16325 (N_16325,N_13773,N_12522);
nor U16326 (N_16326,N_15966,N_14835);
nor U16327 (N_16327,N_15990,N_14900);
or U16328 (N_16328,N_13992,N_15108);
nor U16329 (N_16329,N_15306,N_15074);
and U16330 (N_16330,N_14653,N_14526);
nor U16331 (N_16331,N_15549,N_15038);
nor U16332 (N_16332,N_15423,N_13994);
and U16333 (N_16333,N_12554,N_13643);
or U16334 (N_16334,N_13776,N_12196);
nand U16335 (N_16335,N_14025,N_13465);
nor U16336 (N_16336,N_13137,N_12818);
nand U16337 (N_16337,N_13173,N_15628);
and U16338 (N_16338,N_13983,N_14394);
or U16339 (N_16339,N_13312,N_14903);
nor U16340 (N_16340,N_12841,N_13374);
nor U16341 (N_16341,N_15089,N_12541);
nand U16342 (N_16342,N_12797,N_15458);
or U16343 (N_16343,N_15657,N_12091);
and U16344 (N_16344,N_13883,N_12390);
nand U16345 (N_16345,N_15167,N_13297);
nor U16346 (N_16346,N_13754,N_13619);
nor U16347 (N_16347,N_12010,N_13263);
nand U16348 (N_16348,N_13598,N_15498);
nor U16349 (N_16349,N_14498,N_12472);
nor U16350 (N_16350,N_12357,N_13903);
or U16351 (N_16351,N_12100,N_14255);
and U16352 (N_16352,N_14357,N_13630);
or U16353 (N_16353,N_13030,N_12550);
nor U16354 (N_16354,N_14326,N_14142);
or U16355 (N_16355,N_12751,N_14839);
xor U16356 (N_16356,N_12262,N_12072);
nand U16357 (N_16357,N_15939,N_15554);
or U16358 (N_16358,N_13574,N_14273);
or U16359 (N_16359,N_14883,N_14512);
nand U16360 (N_16360,N_12675,N_13181);
nand U16361 (N_16361,N_13177,N_15610);
nor U16362 (N_16362,N_12166,N_14441);
nor U16363 (N_16363,N_14592,N_12579);
nor U16364 (N_16364,N_12292,N_14026);
or U16365 (N_16365,N_13582,N_12680);
nand U16366 (N_16366,N_13812,N_13437);
or U16367 (N_16367,N_14735,N_13974);
nand U16368 (N_16368,N_13011,N_15453);
nor U16369 (N_16369,N_15815,N_14842);
nor U16370 (N_16370,N_15487,N_14714);
or U16371 (N_16371,N_13228,N_13910);
nand U16372 (N_16372,N_12843,N_13585);
nand U16373 (N_16373,N_13850,N_15785);
nor U16374 (N_16374,N_12069,N_12966);
nand U16375 (N_16375,N_14541,N_12876);
and U16376 (N_16376,N_12252,N_14376);
and U16377 (N_16377,N_12712,N_14958);
nand U16378 (N_16378,N_15550,N_12801);
and U16379 (N_16379,N_14550,N_13216);
and U16380 (N_16380,N_13357,N_12756);
or U16381 (N_16381,N_13249,N_15546);
and U16382 (N_16382,N_12814,N_12471);
xor U16383 (N_16383,N_13614,N_15096);
or U16384 (N_16384,N_14857,N_15895);
nor U16385 (N_16385,N_13679,N_12995);
nand U16386 (N_16386,N_13824,N_15911);
nor U16387 (N_16387,N_12218,N_14477);
nand U16388 (N_16388,N_13964,N_13793);
nand U16389 (N_16389,N_15343,N_12693);
nor U16390 (N_16390,N_14328,N_12920);
nor U16391 (N_16391,N_14845,N_12925);
and U16392 (N_16392,N_12948,N_14112);
nand U16393 (N_16393,N_15093,N_15645);
and U16394 (N_16394,N_13299,N_14259);
or U16395 (N_16395,N_14745,N_15924);
nand U16396 (N_16396,N_15373,N_15738);
and U16397 (N_16397,N_12413,N_13780);
nor U16398 (N_16398,N_13989,N_12321);
or U16399 (N_16399,N_12347,N_15057);
and U16400 (N_16400,N_14840,N_12235);
nand U16401 (N_16401,N_15502,N_14176);
or U16402 (N_16402,N_12059,N_15565);
nand U16403 (N_16403,N_13569,N_14780);
or U16404 (N_16404,N_12438,N_14059);
nor U16405 (N_16405,N_12417,N_14231);
and U16406 (N_16406,N_12696,N_12138);
nand U16407 (N_16407,N_13085,N_14396);
and U16408 (N_16408,N_14155,N_14841);
xnor U16409 (N_16409,N_14729,N_14020);
nor U16410 (N_16410,N_12396,N_15692);
and U16411 (N_16411,N_12592,N_13566);
or U16412 (N_16412,N_15992,N_15817);
and U16413 (N_16413,N_12563,N_14362);
nand U16414 (N_16414,N_13244,N_14807);
nor U16415 (N_16415,N_14449,N_14933);
nand U16416 (N_16416,N_15606,N_12172);
and U16417 (N_16417,N_12101,N_12758);
nand U16418 (N_16418,N_13155,N_13936);
nand U16419 (N_16419,N_12400,N_13224);
nand U16420 (N_16420,N_12703,N_15412);
and U16421 (N_16421,N_15372,N_13439);
nand U16422 (N_16422,N_12655,N_14669);
nand U16423 (N_16423,N_12520,N_12517);
or U16424 (N_16424,N_13422,N_14417);
nand U16425 (N_16425,N_13322,N_13836);
or U16426 (N_16426,N_12942,N_15130);
or U16427 (N_16427,N_12351,N_12297);
or U16428 (N_16428,N_15964,N_15391);
nor U16429 (N_16429,N_15583,N_14493);
and U16430 (N_16430,N_12067,N_13406);
nor U16431 (N_16431,N_12889,N_15651);
or U16432 (N_16432,N_15699,N_12628);
and U16433 (N_16433,N_13343,N_14528);
nor U16434 (N_16434,N_15418,N_13595);
nor U16435 (N_16435,N_14225,N_12318);
or U16436 (N_16436,N_15440,N_15709);
nand U16437 (N_16437,N_12983,N_15009);
nand U16438 (N_16438,N_14068,N_15141);
and U16439 (N_16439,N_13088,N_13478);
and U16440 (N_16440,N_12419,N_13314);
and U16441 (N_16441,N_14961,N_15698);
nor U16442 (N_16442,N_15464,N_15845);
or U16443 (N_16443,N_15848,N_12130);
and U16444 (N_16444,N_14105,N_14795);
and U16445 (N_16445,N_13878,N_12596);
and U16446 (N_16446,N_13132,N_14223);
nor U16447 (N_16447,N_13262,N_14461);
nor U16448 (N_16448,N_13590,N_13526);
and U16449 (N_16449,N_14910,N_14614);
or U16450 (N_16450,N_12169,N_12016);
nor U16451 (N_16451,N_12572,N_13392);
and U16452 (N_16452,N_15909,N_12011);
and U16453 (N_16453,N_13884,N_13045);
nand U16454 (N_16454,N_12156,N_15571);
nand U16455 (N_16455,N_14849,N_12917);
or U16456 (N_16456,N_13589,N_15197);
nor U16457 (N_16457,N_14475,N_12770);
and U16458 (N_16458,N_12648,N_14448);
or U16459 (N_16459,N_13295,N_13208);
nand U16460 (N_16460,N_14645,N_13165);
nand U16461 (N_16461,N_12200,N_15570);
or U16462 (N_16462,N_15524,N_13760);
nand U16463 (N_16463,N_13855,N_15426);
and U16464 (N_16464,N_12773,N_13008);
xor U16465 (N_16465,N_13332,N_13857);
and U16466 (N_16466,N_15022,N_15846);
and U16467 (N_16467,N_15280,N_15053);
or U16468 (N_16468,N_14269,N_15202);
nor U16469 (N_16469,N_12697,N_13841);
and U16470 (N_16470,N_13845,N_15780);
or U16471 (N_16471,N_13555,N_15996);
nand U16472 (N_16472,N_14125,N_15068);
or U16473 (N_16473,N_14979,N_12871);
and U16474 (N_16474,N_14291,N_12238);
or U16475 (N_16475,N_12997,N_13965);
and U16476 (N_16476,N_15617,N_13703);
or U16477 (N_16477,N_15930,N_15831);
and U16478 (N_16478,N_14658,N_12431);
and U16479 (N_16479,N_14494,N_13116);
and U16480 (N_16480,N_12237,N_12952);
and U16481 (N_16481,N_12583,N_14566);
or U16482 (N_16482,N_13513,N_13706);
or U16483 (N_16483,N_13440,N_15720);
nand U16484 (N_16484,N_12879,N_12381);
nand U16485 (N_16485,N_14062,N_13417);
nor U16486 (N_16486,N_15457,N_12389);
and U16487 (N_16487,N_13898,N_12302);
nor U16488 (N_16488,N_14771,N_14416);
or U16489 (N_16489,N_13117,N_12306);
and U16490 (N_16490,N_15230,N_15218);
nand U16491 (N_16491,N_12944,N_14670);
or U16492 (N_16492,N_14238,N_15467);
nor U16493 (N_16493,N_12865,N_13429);
nor U16494 (N_16494,N_14734,N_15404);
or U16495 (N_16495,N_15349,N_15465);
nor U16496 (N_16496,N_15041,N_15427);
and U16497 (N_16497,N_14636,N_12695);
nor U16498 (N_16498,N_15186,N_15252);
nor U16499 (N_16499,N_12106,N_12514);
nor U16500 (N_16500,N_15500,N_13702);
and U16501 (N_16501,N_14334,N_14610);
nor U16502 (N_16502,N_12193,N_12250);
or U16503 (N_16503,N_14728,N_15381);
and U16504 (N_16504,N_15021,N_13893);
nand U16505 (N_16505,N_12420,N_14769);
nand U16506 (N_16506,N_14659,N_14430);
nor U16507 (N_16507,N_14283,N_15675);
or U16508 (N_16508,N_13031,N_15045);
nand U16509 (N_16509,N_15161,N_14937);
and U16510 (N_16510,N_13831,N_12647);
and U16511 (N_16511,N_13970,N_13330);
or U16512 (N_16512,N_13504,N_13459);
nand U16513 (N_16513,N_12830,N_13122);
or U16514 (N_16514,N_15783,N_15935);
or U16515 (N_16515,N_14785,N_14128);
or U16516 (N_16516,N_13020,N_13274);
or U16517 (N_16517,N_15138,N_13105);
or U16518 (N_16518,N_14333,N_15097);
or U16519 (N_16519,N_12746,N_15485);
nor U16520 (N_16520,N_14363,N_15940);
nand U16521 (N_16521,N_12774,N_12003);
nor U16522 (N_16522,N_12826,N_15301);
nand U16523 (N_16523,N_13182,N_15505);
nor U16524 (N_16524,N_12084,N_15688);
or U16525 (N_16525,N_13853,N_13816);
or U16526 (N_16526,N_15887,N_15545);
or U16527 (N_16527,N_15339,N_15249);
and U16528 (N_16528,N_13562,N_12207);
nand U16529 (N_16529,N_13461,N_14485);
nor U16530 (N_16530,N_12141,N_15142);
or U16531 (N_16531,N_13159,N_13242);
nand U16532 (N_16532,N_12794,N_14513);
nor U16533 (N_16533,N_15162,N_14923);
nor U16534 (N_16534,N_15590,N_14146);
or U16535 (N_16535,N_15200,N_14715);
and U16536 (N_16536,N_14343,N_12651);
and U16537 (N_16537,N_15787,N_13308);
or U16538 (N_16538,N_14738,N_13937);
nor U16539 (N_16539,N_13871,N_12025);
nor U16540 (N_16540,N_15774,N_13502);
or U16541 (N_16541,N_12885,N_12775);
nor U16542 (N_16542,N_13823,N_13001);
nand U16543 (N_16543,N_14567,N_12157);
and U16544 (N_16544,N_12158,N_14319);
nand U16545 (N_16545,N_12982,N_12499);
or U16546 (N_16546,N_14191,N_15389);
nand U16547 (N_16547,N_12658,N_12287);
nor U16548 (N_16548,N_12614,N_12125);
nor U16549 (N_16549,N_13995,N_14850);
nand U16550 (N_16550,N_13756,N_14392);
nand U16551 (N_16551,N_12461,N_12567);
and U16552 (N_16552,N_12650,N_13815);
and U16553 (N_16553,N_12482,N_12462);
nor U16554 (N_16554,N_13003,N_14621);
and U16555 (N_16555,N_12604,N_13099);
or U16556 (N_16556,N_14742,N_12064);
nor U16557 (N_16557,N_12745,N_15429);
nand U16558 (N_16558,N_12544,N_13125);
xnor U16559 (N_16559,N_14317,N_13009);
nor U16560 (N_16560,N_14004,N_15063);
and U16561 (N_16561,N_15608,N_15007);
nand U16562 (N_16562,N_15480,N_15227);
or U16563 (N_16563,N_14248,N_14607);
nor U16564 (N_16564,N_14109,N_15150);
nand U16565 (N_16565,N_14652,N_15401);
nor U16566 (N_16566,N_14589,N_15874);
or U16567 (N_16567,N_14630,N_12363);
nand U16568 (N_16568,N_15474,N_14608);
or U16569 (N_16569,N_12862,N_14759);
and U16570 (N_16570,N_13956,N_15883);
and U16571 (N_16571,N_13734,N_13072);
and U16572 (N_16572,N_12863,N_15479);
and U16573 (N_16573,N_14892,N_12310);
and U16574 (N_16574,N_14141,N_13538);
nor U16575 (N_16575,N_15685,N_12440);
nand U16576 (N_16576,N_12049,N_15030);
nand U16577 (N_16577,N_12869,N_13684);
and U16578 (N_16578,N_13489,N_15438);
or U16579 (N_16579,N_15607,N_13136);
or U16580 (N_16580,N_14440,N_14717);
and U16581 (N_16581,N_13810,N_13069);
nand U16582 (N_16582,N_15170,N_15642);
nor U16583 (N_16583,N_13130,N_14086);
nand U16584 (N_16584,N_14939,N_14540);
nor U16585 (N_16585,N_12884,N_12822);
nand U16586 (N_16586,N_13933,N_15707);
nor U16587 (N_16587,N_12763,N_13298);
nor U16588 (N_16588,N_15523,N_12755);
or U16589 (N_16589,N_12071,N_12039);
or U16590 (N_16590,N_15103,N_15896);
or U16591 (N_16591,N_12160,N_12668);
and U16592 (N_16592,N_14280,N_14446);
and U16593 (N_16593,N_14508,N_13843);
or U16594 (N_16594,N_13745,N_13761);
or U16595 (N_16595,N_12283,N_13806);
and U16596 (N_16596,N_14827,N_15116);
nor U16597 (N_16597,N_13885,N_13174);
nand U16598 (N_16598,N_15722,N_12075);
or U16599 (N_16599,N_12911,N_15793);
nand U16600 (N_16600,N_12924,N_14800);
nand U16601 (N_16601,N_15061,N_14806);
or U16602 (N_16602,N_14447,N_15535);
nor U16603 (N_16603,N_12824,N_13656);
nor U16604 (N_16604,N_13446,N_13925);
or U16605 (N_16605,N_14340,N_13301);
and U16606 (N_16606,N_12378,N_14642);
nor U16607 (N_16607,N_13448,N_12386);
and U16608 (N_16608,N_12326,N_14093);
nor U16609 (N_16609,N_12959,N_12031);
or U16610 (N_16610,N_15634,N_13201);
nand U16611 (N_16611,N_15750,N_15320);
nand U16612 (N_16612,N_14993,N_12946);
and U16613 (N_16613,N_13809,N_13320);
or U16614 (N_16614,N_12446,N_15616);
nor U16615 (N_16615,N_13854,N_12897);
nand U16616 (N_16616,N_13396,N_15424);
or U16617 (N_16617,N_15212,N_14314);
nand U16618 (N_16618,N_12123,N_13187);
nor U16619 (N_16619,N_15684,N_14024);
and U16620 (N_16620,N_15099,N_12053);
nand U16621 (N_16621,N_12377,N_14984);
and U16622 (N_16622,N_15993,N_15286);
or U16623 (N_16623,N_15284,N_15156);
and U16624 (N_16624,N_15446,N_14533);
nand U16625 (N_16625,N_13957,N_13036);
nand U16626 (N_16626,N_14364,N_12087);
or U16627 (N_16627,N_12713,N_13296);
and U16628 (N_16628,N_12612,N_14358);
or U16629 (N_16629,N_15352,N_13613);
or U16630 (N_16630,N_15396,N_14169);
or U16631 (N_16631,N_12359,N_13753);
and U16632 (N_16632,N_15148,N_15949);
nor U16633 (N_16633,N_15661,N_14010);
and U16634 (N_16634,N_14901,N_13771);
and U16635 (N_16635,N_14612,N_14744);
nor U16636 (N_16636,N_15370,N_12361);
nand U16637 (N_16637,N_14370,N_13472);
nand U16638 (N_16638,N_13171,N_12183);
nand U16639 (N_16639,N_14178,N_12854);
and U16640 (N_16640,N_12192,N_15133);
and U16641 (N_16641,N_15271,N_12633);
nand U16642 (N_16642,N_13090,N_12002);
or U16643 (N_16643,N_15885,N_12006);
and U16644 (N_16644,N_13580,N_12813);
and U16645 (N_16645,N_12001,N_12850);
or U16646 (N_16646,N_12711,N_14497);
and U16647 (N_16647,N_12630,N_15979);
and U16648 (N_16648,N_12796,N_13888);
nor U16649 (N_16649,N_13622,N_13243);
or U16650 (N_16650,N_15912,N_14510);
and U16651 (N_16651,N_15888,N_14561);
and U16652 (N_16652,N_13371,N_14503);
and U16653 (N_16653,N_12761,N_14914);
nor U16654 (N_16654,N_15868,N_14228);
xnor U16655 (N_16655,N_13593,N_14138);
or U16656 (N_16656,N_14187,N_12922);
nand U16657 (N_16657,N_12971,N_12574);
or U16658 (N_16658,N_14968,N_15769);
nor U16659 (N_16659,N_15997,N_12466);
and U16660 (N_16660,N_13487,N_14468);
or U16661 (N_16661,N_12398,N_13663);
or U16662 (N_16662,N_14678,N_15254);
or U16663 (N_16663,N_14797,N_14926);
or U16664 (N_16664,N_15111,N_15755);
or U16665 (N_16665,N_15637,N_15265);
and U16666 (N_16666,N_14454,N_12962);
nand U16667 (N_16667,N_12760,N_12935);
or U16668 (N_16668,N_12559,N_15683);
nand U16669 (N_16669,N_13701,N_12434);
or U16670 (N_16670,N_12930,N_12392);
and U16671 (N_16671,N_12881,N_12730);
and U16672 (N_16672,N_14210,N_15666);
nand U16673 (N_16673,N_15256,N_13981);
nand U16674 (N_16674,N_15220,N_13261);
nor U16675 (N_16675,N_14781,N_13647);
and U16676 (N_16676,N_12190,N_15365);
nor U16677 (N_16677,N_14066,N_13247);
or U16678 (N_16678,N_15830,N_14133);
or U16679 (N_16679,N_14997,N_14718);
and U16680 (N_16680,N_14284,N_12410);
nand U16681 (N_16681,N_14211,N_12587);
or U16682 (N_16682,N_14320,N_15214);
nand U16683 (N_16683,N_14065,N_15555);
nor U16684 (N_16684,N_14496,N_13342);
nand U16685 (N_16685,N_12785,N_15488);
and U16686 (N_16686,N_12672,N_14753);
or U16687 (N_16687,N_12380,N_12595);
nor U16688 (N_16688,N_15521,N_15507);
nand U16689 (N_16689,N_12985,N_12411);
or U16690 (N_16690,N_14716,N_14413);
nand U16691 (N_16691,N_13897,N_12601);
and U16692 (N_16692,N_13418,N_13646);
and U16693 (N_16693,N_13779,N_13250);
xor U16694 (N_16694,N_14722,N_12241);
or U16695 (N_16695,N_12717,N_14293);
or U16696 (N_16696,N_15266,N_13017);
or U16697 (N_16697,N_14676,N_12443);
nand U16698 (N_16698,N_15342,N_14801);
nor U16699 (N_16699,N_15557,N_13196);
nand U16700 (N_16700,N_14925,N_14813);
nor U16701 (N_16701,N_15863,N_15496);
or U16702 (N_16702,N_14825,N_14205);
and U16703 (N_16703,N_13879,N_14890);
and U16704 (N_16704,N_15140,N_14584);
nor U16705 (N_16705,N_14656,N_13019);
and U16706 (N_16706,N_14556,N_12325);
nand U16707 (N_16707,N_12949,N_12827);
or U16708 (N_16708,N_12198,N_15541);
nand U16709 (N_16709,N_14402,N_14697);
nand U16710 (N_16710,N_12739,N_12248);
nor U16711 (N_16711,N_15663,N_12684);
nor U16712 (N_16712,N_15035,N_15180);
nor U16713 (N_16713,N_13880,N_15761);
or U16714 (N_16714,N_14499,N_13929);
nand U16715 (N_16715,N_14172,N_15889);
and U16716 (N_16716,N_12227,N_14341);
nor U16717 (N_16717,N_15781,N_15627);
nand U16718 (N_16718,N_14136,N_14639);
and U16719 (N_16719,N_12692,N_15058);
nor U16720 (N_16720,N_12291,N_12957);
nor U16721 (N_16721,N_14171,N_12253);
and U16722 (N_16722,N_14338,N_15501);
or U16723 (N_16723,N_15189,N_14838);
nand U16724 (N_16724,N_13151,N_12082);
nor U16725 (N_16725,N_13928,N_13863);
nor U16726 (N_16726,N_14055,N_15052);
or U16727 (N_16727,N_14585,N_14286);
and U16728 (N_16728,N_15723,N_14691);
and U16729 (N_16729,N_14646,N_12859);
nor U16730 (N_16730,N_13694,N_14805);
nand U16731 (N_16731,N_13168,N_12724);
and U16732 (N_16732,N_12815,N_12269);
and U16733 (N_16733,N_14970,N_15425);
or U16734 (N_16734,N_13649,N_13560);
or U16735 (N_16735,N_13225,N_14266);
nand U16736 (N_16736,N_13548,N_12249);
nor U16737 (N_16737,N_12851,N_12999);
nand U16738 (N_16738,N_13596,N_14602);
and U16739 (N_16739,N_12216,N_14873);
or U16740 (N_16740,N_13503,N_14664);
or U16741 (N_16741,N_13432,N_13102);
nand U16742 (N_16742,N_14164,N_12626);
nor U16743 (N_16743,N_13750,N_14788);
or U16744 (N_16744,N_13584,N_13134);
nor U16745 (N_16745,N_14783,N_15264);
nor U16746 (N_16746,N_15644,N_12901);
or U16747 (N_16747,N_12427,N_15822);
nor U16748 (N_16748,N_13163,N_12298);
and U16749 (N_16749,N_12009,N_12685);
nor U16750 (N_16750,N_13930,N_12538);
and U16751 (N_16751,N_14000,N_12093);
or U16752 (N_16752,N_14644,N_13752);
nand U16753 (N_16753,N_15520,N_14091);
nand U16754 (N_16754,N_14502,N_13661);
nor U16755 (N_16755,N_15020,N_13819);
nor U16756 (N_16756,N_12102,N_14796);
or U16757 (N_16757,N_12323,N_13565);
nor U16758 (N_16758,N_15098,N_15745);
nor U16759 (N_16759,N_15360,N_14023);
nand U16760 (N_16760,N_13534,N_14309);
and U16761 (N_16761,N_15701,N_13176);
nand U16762 (N_16762,N_14264,N_12990);
nor U16763 (N_16763,N_12228,N_14344);
and U16764 (N_16764,N_14808,N_14978);
and U16765 (N_16765,N_14770,N_15572);
nand U16766 (N_16766,N_12436,N_13154);
nand U16767 (N_16767,N_12119,N_15522);
or U16768 (N_16768,N_14727,N_15506);
and U16769 (N_16769,N_15747,N_14117);
or U16770 (N_16770,N_12021,N_15776);
nand U16771 (N_16771,N_15318,N_14380);
nor U16772 (N_16772,N_15348,N_12993);
or U16773 (N_16773,N_15811,N_15856);
nand U16774 (N_16774,N_12940,N_13873);
nor U16775 (N_16775,N_14427,N_12448);
nand U16776 (N_16776,N_12807,N_14327);
and U16777 (N_16777,N_14369,N_12259);
nand U16778 (N_16778,N_12054,N_15155);
and U16779 (N_16779,N_13167,N_15526);
and U16780 (N_16780,N_13430,N_13399);
and U16781 (N_16781,N_15902,N_15559);
and U16782 (N_16782,N_13790,N_12661);
nor U16783 (N_16783,N_14208,N_14552);
nand U16784 (N_16784,N_12463,N_13405);
and U16785 (N_16785,N_12020,N_15356);
nand U16786 (N_16786,N_14700,N_13623);
nand U16787 (N_16787,N_13556,N_14234);
or U16788 (N_16788,N_13015,N_13927);
and U16789 (N_16789,N_13543,N_14743);
and U16790 (N_16790,N_14132,N_13424);
nand U16791 (N_16791,N_13711,N_14218);
nand U16792 (N_16792,N_13839,N_13531);
or U16793 (N_16793,N_15667,N_14361);
or U16794 (N_16794,N_12706,N_12976);
nand U16795 (N_16795,N_12938,N_14124);
and U16796 (N_16796,N_12887,N_14507);
nand U16797 (N_16797,N_12439,N_15152);
nor U16798 (N_16798,N_15665,N_14782);
nand U16799 (N_16799,N_15244,N_15028);
and U16800 (N_16800,N_12906,N_14435);
nor U16801 (N_16801,N_13742,N_14410);
nand U16802 (N_16802,N_12508,N_13445);
nor U16803 (N_16803,N_13027,N_14764);
or U16804 (N_16804,N_13324,N_12133);
nand U16805 (N_16805,N_14131,N_13292);
nor U16806 (N_16806,N_14473,N_12421);
nand U16807 (N_16807,N_13539,N_13536);
nand U16808 (N_16808,N_13608,N_15806);
nor U16809 (N_16809,N_12530,N_15591);
and U16810 (N_16810,N_13082,N_14916);
or U16811 (N_16811,N_14836,N_14980);
nor U16812 (N_16812,N_13900,N_12033);
and U16813 (N_16813,N_14679,N_14374);
or U16814 (N_16814,N_12928,N_15864);
nand U16815 (N_16815,N_13961,N_15293);
nand U16816 (N_16816,N_13315,N_15913);
nand U16817 (N_16817,N_13782,N_14768);
nor U16818 (N_16818,N_13650,N_14071);
and U16819 (N_16819,N_14381,N_14115);
and U16820 (N_16820,N_12798,N_13497);
or U16821 (N_16821,N_14721,N_12987);
nand U16822 (N_16822,N_14027,N_14052);
and U16823 (N_16823,N_12566,N_13000);
or U16824 (N_16824,N_12062,N_14422);
and U16825 (N_16825,N_12702,N_14613);
nand U16826 (N_16826,N_12741,N_12045);
or U16827 (N_16827,N_12483,N_12110);
nand U16828 (N_16828,N_12257,N_14101);
and U16829 (N_16829,N_12783,N_13442);
nand U16830 (N_16830,N_13896,N_14562);
and U16831 (N_16831,N_14079,N_12118);
or U16832 (N_16832,N_13775,N_12121);
nor U16833 (N_16833,N_15671,N_13579);
nor U16834 (N_16834,N_15483,N_15728);
nor U16835 (N_16835,N_15881,N_12136);
and U16836 (N_16836,N_12212,N_13026);
nor U16837 (N_16837,N_14831,N_13481);
nor U16838 (N_16838,N_15697,N_14711);
and U16839 (N_16839,N_13037,N_15941);
and U16840 (N_16840,N_15345,N_14488);
nand U16841 (N_16841,N_15120,N_14772);
nor U16842 (N_16842,N_12251,N_14078);
and U16843 (N_16843,N_15088,N_12308);
and U16844 (N_16844,N_13577,N_13583);
or U16845 (N_16845,N_15643,N_15991);
and U16846 (N_16846,N_14046,N_15273);
nor U16847 (N_16847,N_13270,N_14313);
nor U16848 (N_16848,N_15563,N_14277);
or U16849 (N_16849,N_14405,N_12213);
nand U16850 (N_16850,N_12442,N_12065);
nand U16851 (N_16851,N_15379,N_12529);
or U16852 (N_16852,N_15873,N_13491);
nor U16853 (N_16853,N_14013,N_13131);
nand U16854 (N_16854,N_14386,N_12833);
and U16855 (N_16855,N_12670,N_12099);
and U16856 (N_16856,N_12980,N_14236);
nor U16857 (N_16857,N_12705,N_12521);
nand U16858 (N_16858,N_14665,N_12787);
nor U16859 (N_16859,N_15882,N_14858);
or U16860 (N_16860,N_12534,N_14870);
nor U16861 (N_16861,N_12239,N_14463);
and U16862 (N_16862,N_15201,N_15304);
and U16863 (N_16863,N_14069,N_12159);
xnor U16864 (N_16864,N_13273,N_15246);
or U16865 (N_16865,N_13805,N_15849);
nor U16866 (N_16866,N_14896,N_15187);
nand U16867 (N_16867,N_14830,N_13362);
nand U16868 (N_16868,N_14242,N_14408);
and U16869 (N_16869,N_14149,N_15067);
and U16870 (N_16870,N_14948,N_12104);
or U16871 (N_16871,N_12955,N_14643);
nand U16872 (N_16872,N_13847,N_13802);
nand U16873 (N_16873,N_12784,N_12094);
or U16874 (N_16874,N_14045,N_15371);
nand U16875 (N_16875,N_12043,N_14118);
and U16876 (N_16876,N_14360,N_14199);
nand U16877 (N_16877,N_12943,N_13160);
nor U16878 (N_16878,N_15986,N_14084);
nor U16879 (N_16879,N_14123,N_13056);
nand U16880 (N_16880,N_15786,N_15824);
or U16881 (N_16881,N_12282,N_12496);
nand U16882 (N_16882,N_15325,N_14594);
and U16883 (N_16883,N_13138,N_13333);
and U16884 (N_16884,N_12970,N_13955);
nand U16885 (N_16885,N_13103,N_12464);
or U16886 (N_16886,N_13143,N_12426);
nor U16887 (N_16887,N_12203,N_15359);
or U16888 (N_16888,N_14569,N_14746);
nand U16889 (N_16889,N_12184,N_13038);
nor U16890 (N_16890,N_15118,N_12484);
or U16891 (N_16891,N_13146,N_13207);
or U16892 (N_16892,N_15090,N_15017);
nand U16893 (N_16893,N_15866,N_12232);
and U16894 (N_16894,N_13409,N_14654);
nor U16895 (N_16895,N_15037,N_14147);
nand U16896 (N_16896,N_12474,N_12340);
nor U16897 (N_16897,N_13600,N_12222);
nand U16898 (N_16898,N_13629,N_13717);
nor U16899 (N_16899,N_14920,N_15482);
and U16900 (N_16900,N_13441,N_12842);
or U16901 (N_16901,N_15449,N_14481);
and U16902 (N_16902,N_13726,N_12077);
nand U16903 (N_16903,N_14180,N_12929);
and U16904 (N_16904,N_15622,N_13546);
and U16905 (N_16905,N_14625,N_12221);
nand U16906 (N_16906,N_14021,N_13784);
and U16907 (N_16907,N_13033,N_13696);
nand U16908 (N_16908,N_14790,N_14482);
nor U16909 (N_16909,N_12752,N_12931);
nor U16910 (N_16910,N_13658,N_14479);
or U16911 (N_16911,N_15751,N_15241);
nand U16912 (N_16912,N_14817,N_12972);
and U16913 (N_16913,N_13724,N_14260);
or U16914 (N_16914,N_13140,N_13954);
nor U16915 (N_16915,N_13368,N_15922);
or U16916 (N_16916,N_13450,N_14018);
xnor U16917 (N_16917,N_12852,N_13700);
or U16918 (N_16918,N_12477,N_13617);
or U16919 (N_16919,N_14008,N_14708);
nand U16920 (N_16920,N_12301,N_13276);
nand U16921 (N_16921,N_13275,N_12836);
nand U16922 (N_16922,N_14219,N_13916);
or U16923 (N_16923,N_14692,N_13355);
and U16924 (N_16924,N_14732,N_13528);
nand U16925 (N_16925,N_15013,N_15102);
and U16926 (N_16926,N_12937,N_12047);
nand U16927 (N_16927,N_15217,N_12070);
nor U16928 (N_16928,N_15576,N_15840);
nor U16929 (N_16929,N_15177,N_13321);
nand U16930 (N_16930,N_13231,N_12872);
nand U16931 (N_16931,N_13220,N_13563);
and U16932 (N_16932,N_12300,N_13677);
and U16933 (N_16933,N_13523,N_12111);
nor U16934 (N_16934,N_12404,N_13178);
and U16935 (N_16935,N_15599,N_13976);
nand U16936 (N_16936,N_12332,N_15510);
or U16937 (N_16937,N_15851,N_15324);
nand U16938 (N_16938,N_13859,N_15183);
and U16939 (N_16939,N_12089,N_15646);
and U16940 (N_16940,N_15471,N_14748);
nor U16941 (N_16941,N_15310,N_12891);
nand U16942 (N_16942,N_15696,N_13239);
nand U16943 (N_16943,N_12454,N_14511);
or U16944 (N_16944,N_15203,N_13545);
nand U16945 (N_16945,N_14220,N_12215);
nand U16946 (N_16946,N_14650,N_15691);
nand U16947 (N_16947,N_14963,N_15802);
and U16948 (N_16948,N_12430,N_12618);
nand U16949 (N_16949,N_13413,N_14459);
or U16950 (N_16950,N_12515,N_13547);
and U16951 (N_16951,N_13862,N_14591);
nand U16952 (N_16952,N_12777,N_15519);
and U16953 (N_16953,N_12720,N_12354);
and U16954 (N_16954,N_15525,N_14315);
nand U16955 (N_16955,N_14256,N_15491);
or U16956 (N_16956,N_15561,N_13733);
or U16957 (N_16957,N_12142,N_14239);
nand U16958 (N_16958,N_12977,N_13286);
nand U16959 (N_16959,N_12032,N_13792);
nand U16960 (N_16960,N_15900,N_14976);
or U16961 (N_16961,N_15579,N_12134);
nand U16962 (N_16962,N_15190,N_13704);
and U16963 (N_16963,N_12395,N_12682);
nor U16964 (N_16964,N_15243,N_14855);
nor U16965 (N_16965,N_14505,N_13028);
or U16966 (N_16966,N_13185,N_12547);
nand U16967 (N_16967,N_14641,N_12771);
nand U16968 (N_16968,N_13625,N_15655);
nand U16969 (N_16969,N_15794,N_14582);
or U16970 (N_16970,N_15543,N_12909);
nor U16971 (N_16971,N_14945,N_13611);
nor U16972 (N_16972,N_13748,N_15055);
or U16973 (N_16973,N_13336,N_15847);
or U16974 (N_16974,N_12281,N_14174);
nor U16975 (N_16975,N_12144,N_13104);
and U16976 (N_16976,N_12468,N_14977);
and U16977 (N_16977,N_12907,N_15687);
and U16978 (N_16978,N_14869,N_12740);
and U16979 (N_16979,N_15961,N_15078);
or U16980 (N_16980,N_13621,N_14012);
nor U16981 (N_16981,N_12747,N_15604);
nor U16982 (N_16982,N_12847,N_15814);
nor U16983 (N_16983,N_14310,N_12714);
or U16984 (N_16984,N_15193,N_15734);
or U16985 (N_16985,N_15478,N_12811);
and U16986 (N_16986,N_12405,N_15082);
nand U16987 (N_16987,N_15906,N_13737);
and U16988 (N_16988,N_12744,N_15631);
or U16989 (N_16989,N_13667,N_12603);
nand U16990 (N_16990,N_14940,N_13466);
nor U16991 (N_16991,N_12641,N_14151);
nand U16992 (N_16992,N_15952,N_13678);
and U16993 (N_16993,N_13710,N_14515);
and U16994 (N_16994,N_15330,N_15462);
xor U16995 (N_16995,N_15973,N_15967);
nor U16996 (N_16996,N_14349,N_13963);
and U16997 (N_16997,N_15208,N_12516);
or U16998 (N_16998,N_12776,N_12376);
or U16999 (N_16999,N_12057,N_13300);
nor U17000 (N_17000,N_13248,N_14244);
or U17001 (N_17001,N_15693,N_14851);
or U17002 (N_17002,N_12124,N_13200);
or U17003 (N_17003,N_14539,N_15573);
xnor U17004 (N_17004,N_13454,N_14177);
or U17005 (N_17005,N_15611,N_14398);
and U17006 (N_17006,N_13081,N_14022);
and U17007 (N_17007,N_15770,N_14011);
and U17008 (N_17008,N_12678,N_13652);
nor U17009 (N_17009,N_14888,N_15736);
or U17010 (N_17010,N_14521,N_13691);
nor U17011 (N_17011,N_12519,N_15364);
or U17012 (N_17012,N_15614,N_13506);
and U17013 (N_17013,N_15768,N_12998);
nor U17014 (N_17014,N_13360,N_13032);
and U17015 (N_17015,N_15641,N_13025);
and U17016 (N_17016,N_14985,N_14532);
nand U17017 (N_17017,N_14325,N_12565);
nand U17018 (N_17018,N_14822,N_15547);
nor U17019 (N_17019,N_13971,N_13347);
nand U17020 (N_17020,N_14157,N_12346);
nor U17021 (N_17021,N_14452,N_15210);
or U17022 (N_17022,N_13084,N_12586);
nand U17023 (N_17023,N_14061,N_15402);
and U17024 (N_17024,N_15127,N_13757);
nor U17025 (N_17025,N_14725,N_12432);
nand U17026 (N_17026,N_12548,N_13517);
nor U17027 (N_17027,N_15357,N_13223);
and U17028 (N_17028,N_15322,N_14272);
and U17029 (N_17029,N_14703,N_12536);
nor U17030 (N_17030,N_15974,N_15198);
nor U17031 (N_17031,N_13323,N_12375);
nor U17032 (N_17032,N_13049,N_12832);
nor U17033 (N_17033,N_15715,N_13660);
nor U17034 (N_17034,N_13067,N_15800);
or U17035 (N_17035,N_13804,N_13291);
nand U17036 (N_17036,N_13952,N_12622);
xnor U17037 (N_17037,N_12800,N_14378);
nand U17038 (N_17038,N_14570,N_14603);
and U17039 (N_17039,N_15635,N_13765);
nor U17040 (N_17040,N_14837,N_13919);
nand U17041 (N_17041,N_13770,N_13078);
nor U17042 (N_17042,N_12191,N_12506);
nand U17043 (N_17043,N_14609,N_13370);
nor U17044 (N_17044,N_15660,N_13356);
nor U17045 (N_17045,N_15248,N_12979);
and U17046 (N_17046,N_12126,N_14853);
or U17047 (N_17047,N_15016,N_15005);
nor U17048 (N_17048,N_12611,N_12994);
nor U17049 (N_17049,N_12208,N_14075);
nor U17050 (N_17050,N_14693,N_14216);
and U17051 (N_17051,N_13554,N_12764);
or U17052 (N_17052,N_13827,N_13935);
nand U17053 (N_17053,N_12535,N_14709);
nor U17054 (N_17054,N_13039,N_15704);
nand U17055 (N_17055,N_13662,N_12867);
and U17056 (N_17056,N_14994,N_13055);
nor U17057 (N_17057,N_14241,N_13183);
xnor U17058 (N_17058,N_14346,N_13488);
and U17059 (N_17059,N_13681,N_15407);
or U17060 (N_17060,N_13567,N_14947);
and U17061 (N_17061,N_13311,N_12728);
and U17062 (N_17062,N_13115,N_12704);
nand U17063 (N_17063,N_15329,N_12914);
nor U17064 (N_17064,N_13064,N_14547);
and U17065 (N_17065,N_13318,N_14009);
and U17066 (N_17066,N_12902,N_15481);
and U17067 (N_17067,N_15509,N_12716);
nor U17068 (N_17068,N_13875,N_15695);
nor U17069 (N_17069,N_15178,N_15001);
nor U17070 (N_17070,N_13384,N_14778);
nor U17071 (N_17071,N_15387,N_13980);
and U17072 (N_17072,N_15270,N_13066);
nor U17073 (N_17073,N_12035,N_15169);
and U17074 (N_17074,N_13840,N_14329);
nand U17075 (N_17075,N_12619,N_15717);
nor U17076 (N_17076,N_13041,N_13800);
or U17077 (N_17077,N_15173,N_13917);
or U17078 (N_17078,N_12638,N_13123);
or U17079 (N_17079,N_15772,N_13738);
nor U17080 (N_17080,N_15552,N_13746);
and U17081 (N_17081,N_14557,N_14789);
nor U17082 (N_17082,N_15384,N_12545);
nor U17083 (N_17083,N_15578,N_12401);
nor U17084 (N_17084,N_14258,N_12353);
or U17085 (N_17085,N_15514,N_15333);
and U17086 (N_17086,N_15447,N_13759);
or U17087 (N_17087,N_13674,N_12769);
or U17088 (N_17088,N_12105,N_15368);
nor U17089 (N_17089,N_12293,N_13510);
nor U17090 (N_17090,N_14035,N_15366);
nor U17091 (N_17091,N_12540,N_15238);
nand U17092 (N_17092,N_14262,N_14663);
and U17093 (N_17093,N_14935,N_14548);
or U17094 (N_17094,N_15131,N_12941);
nor U17095 (N_17095,N_15714,N_14549);
and U17096 (N_17096,N_13245,N_15915);
nand U17097 (N_17097,N_13482,N_13803);
or U17098 (N_17098,N_12557,N_14634);
nor U17099 (N_17099,N_13685,N_13427);
and U17100 (N_17100,N_15153,N_14460);
nor U17101 (N_17101,N_12441,N_15884);
and U17102 (N_17102,N_15347,N_13075);
nand U17103 (N_17103,N_15399,N_13313);
nand U17104 (N_17104,N_15393,N_14586);
nor U17105 (N_17105,N_15901,N_12500);
nand U17106 (N_17106,N_12285,N_14946);
nor U17107 (N_17107,N_15308,N_12095);
nor U17108 (N_17108,N_14606,N_12873);
nand U17109 (N_17109,N_15128,N_15516);
and U17110 (N_17110,N_12963,N_13393);
nor U17111 (N_17111,N_14969,N_12735);
nor U17112 (N_17112,N_14197,N_12076);
and U17113 (N_17113,N_12185,N_15792);
nor U17114 (N_17114,N_14854,N_12445);
and U17115 (N_17115,N_15107,N_13213);
and U17116 (N_17116,N_13419,N_15291);
nor U17117 (N_17117,N_13197,N_15234);
and U17118 (N_17118,N_15313,N_14886);
and U17119 (N_17119,N_13204,N_15624);
or U17120 (N_17120,N_13868,N_12539);
nand U17121 (N_17121,N_13139,N_13690);
and U17122 (N_17122,N_12311,N_14617);
nor U17123 (N_17123,N_12609,N_15725);
or U17124 (N_17124,N_14204,N_14196);
or U17125 (N_17125,N_14832,N_13561);
and U17126 (N_17126,N_15998,N_15823);
nand U17127 (N_17127,N_15362,N_13736);
and U17128 (N_17128,N_14538,N_13943);
and U17129 (N_17129,N_14815,N_12349);
nor U17130 (N_17130,N_15269,N_14829);
nand U17131 (N_17131,N_13219,N_12247);
nor U17132 (N_17132,N_15718,N_15328);
and U17133 (N_17133,N_14504,N_12606);
nor U17134 (N_17134,N_13112,N_13378);
and U17135 (N_17135,N_15168,N_15497);
or U17136 (N_17136,N_14874,N_14616);
nand U17137 (N_17137,N_13655,N_12245);
and U17138 (N_17138,N_15261,N_14087);
and U17139 (N_17139,N_14710,N_13209);
or U17140 (N_17140,N_14173,N_12895);
nand U17141 (N_17141,N_15999,N_12568);
or U17142 (N_17142,N_12224,N_14017);
nand U17143 (N_17143,N_12510,N_13436);
and U17144 (N_17144,N_15679,N_14966);
nor U17145 (N_17145,N_15943,N_14593);
and U17146 (N_17146,N_14974,N_12052);
and U17147 (N_17147,N_12743,N_13212);
nand U17148 (N_17148,N_14043,N_14267);
nand U17149 (N_17149,N_14190,N_15861);
nand U17150 (N_17150,N_13002,N_15821);
nand U17151 (N_17151,N_15989,N_12487);
xnor U17152 (N_17152,N_13899,N_12012);
nand U17153 (N_17153,N_13798,N_14982);
nand U17154 (N_17154,N_14675,N_14298);
or U17155 (N_17155,N_13829,N_13721);
nor U17156 (N_17156,N_14749,N_12339);
nor U17157 (N_17157,N_15702,N_15272);
nor U17158 (N_17158,N_14972,N_13639);
nor U17159 (N_17159,N_12788,N_13086);
xnor U17160 (N_17160,N_13825,N_15795);
and U17161 (N_17161,N_14819,N_12367);
nor U17162 (N_17162,N_14034,N_14215);
or U17163 (N_17163,N_12689,N_13887);
nor U17164 (N_17164,N_14462,N_13006);
and U17165 (N_17165,N_13817,N_12280);
and U17166 (N_17166,N_14662,N_14209);
nor U17167 (N_17167,N_12973,N_12786);
and U17168 (N_17168,N_14107,N_12877);
or U17169 (N_17169,N_14483,N_15746);
and U17170 (N_17170,N_15609,N_12894);
or U17171 (N_17171,N_15615,N_15299);
nor U17172 (N_17172,N_15436,N_15184);
or U17173 (N_17173,N_13346,N_15215);
nand U17174 (N_17174,N_13835,N_14092);
nor U17175 (N_17175,N_14514,N_12290);
nor U17176 (N_17176,N_13353,N_14037);
or U17177 (N_17177,N_14754,N_15346);
nand U17178 (N_17178,N_12284,N_15113);
nor U17179 (N_17179,N_14247,N_14761);
and U17180 (N_17180,N_13476,N_15194);
nand U17181 (N_17181,N_14166,N_12560);
nand U17182 (N_17182,N_15236,N_12113);
nand U17183 (N_17183,N_12617,N_13664);
nor U17184 (N_17184,N_15338,N_14944);
or U17185 (N_17185,N_14365,N_13246);
nor U17186 (N_17186,N_14122,N_14673);
and U17187 (N_17187,N_15377,N_14028);
nor U17188 (N_17188,N_14894,N_13975);
or U17189 (N_17189,N_15400,N_14635);
and U17190 (N_17190,N_13052,N_14261);
or U17191 (N_17191,N_13864,N_14686);
nor U17192 (N_17192,N_15586,N_14044);
and U17193 (N_17193,N_15222,N_14451);
xnor U17194 (N_17194,N_12162,N_14198);
and U17195 (N_17195,N_12677,N_14719);
nand U17196 (N_17196,N_13034,N_12459);
and U17197 (N_17197,N_13327,N_13860);
nand U17198 (N_17198,N_12958,N_14100);
nor U17199 (N_17199,N_12151,N_14450);
and U17200 (N_17200,N_13688,N_12473);
and U17201 (N_17201,N_14090,N_15540);
nand U17202 (N_17202,N_12552,N_14472);
nand U17203 (N_17203,N_15307,N_13142);
and U17204 (N_17204,N_15826,N_14165);
and U17205 (N_17205,N_12088,N_13426);
nor U17206 (N_17206,N_13358,N_15654);
or U17207 (N_17207,N_14305,N_15341);
nand U17208 (N_17208,N_15260,N_15195);
nand U17209 (N_17209,N_15231,N_15876);
nand U17210 (N_17210,N_15026,N_14524);
nand U17211 (N_17211,N_13789,N_13743);
or U17212 (N_17212,N_13251,N_12806);
or U17213 (N_17213,N_13169,N_12631);
and U17214 (N_17214,N_14810,N_15213);
nand U17215 (N_17215,N_12757,N_13195);
or U17216 (N_17216,N_14120,N_14484);
or U17217 (N_17217,N_13128,N_15934);
and U17218 (N_17218,N_13715,N_12969);
and U17219 (N_17219,N_13076,N_12038);
nand U17220 (N_17220,N_14918,N_14954);
nand U17221 (N_17221,N_15938,N_15630);
nor U17222 (N_17222,N_14401,N_12407);
and U17223 (N_17223,N_15262,N_13618);
nand U17224 (N_17224,N_14057,N_15737);
nor U17225 (N_17225,N_12533,N_12187);
nor U17226 (N_17226,N_14478,N_13951);
nand U17227 (N_17227,N_12729,N_14871);
and U17228 (N_17228,N_14638,N_13194);
and U17229 (N_17229,N_14375,N_15353);
and U17230 (N_17230,N_13587,N_13682);
or U17231 (N_17231,N_14862,N_14070);
and U17232 (N_17232,N_13610,N_13180);
nand U17233 (N_17233,N_12817,N_15065);
and U17234 (N_17234,N_13848,N_14390);
and U17235 (N_17235,N_12188,N_15159);
nor U17236 (N_17236,N_15626,N_12263);
and U17237 (N_17237,N_15850,N_13170);
nor U17238 (N_17238,N_13379,N_14002);
nand U17239 (N_17239,N_12594,N_15689);
nand U17240 (N_17240,N_14576,N_12722);
nand U17241 (N_17241,N_15531,N_12083);
nand U17242 (N_17242,N_15314,N_12180);
nand U17243 (N_17243,N_12299,N_13411);
xor U17244 (N_17244,N_13638,N_15968);
or U17245 (N_17245,N_14354,N_15955);
nand U17246 (N_17246,N_15211,N_13404);
nand U17247 (N_17247,N_15494,N_15331);
or U17248 (N_17248,N_14649,N_15477);
and U17249 (N_17249,N_15147,N_15872);
and U17250 (N_17250,N_15019,N_15066);
or U17251 (N_17251,N_15257,N_14400);
nand U17252 (N_17252,N_15994,N_15710);
or U17253 (N_17253,N_15079,N_12258);
nor U17254 (N_17254,N_13923,N_14137);
and U17255 (N_17255,N_12243,N_13741);
nor U17256 (N_17256,N_15929,N_14731);
or U17257 (N_17257,N_12097,N_12637);
nor U17258 (N_17258,N_13226,N_15771);
or U17259 (N_17259,N_12945,N_14632);
nand U17260 (N_17260,N_15515,N_12137);
nand U17261 (N_17261,N_14667,N_13512);
or U17262 (N_17262,N_13359,N_15100);
and U17263 (N_17263,N_15827,N_13777);
or U17264 (N_17264,N_14588,N_13837);
nand U17265 (N_17265,N_13153,N_13463);
nor U17266 (N_17266,N_14348,N_12819);
or U17267 (N_17267,N_13708,N_15101);
nor U17268 (N_17268,N_12412,N_14527);
nand U17269 (N_17269,N_15926,N_13941);
or U17270 (N_17270,N_14031,N_12575);
and U17271 (N_17271,N_13022,N_13120);
and U17272 (N_17272,N_12465,N_13942);
or U17273 (N_17273,N_13227,N_14367);
and U17274 (N_17274,N_12915,N_15534);
nor U17275 (N_17275,N_12217,N_14672);
and U17276 (N_17276,N_14443,N_13830);
or U17277 (N_17277,N_14296,N_14975);
nand U17278 (N_17278,N_12978,N_14906);
or U17279 (N_17279,N_12570,N_13634);
nor U17280 (N_17280,N_13516,N_15894);
and U17281 (N_17281,N_12242,N_15921);
and U17282 (N_17282,N_12537,N_15206);
or U17283 (N_17283,N_13048,N_14762);
nor U17284 (N_17284,N_12478,N_13984);
and U17285 (N_17285,N_12233,N_12147);
nor U17286 (N_17286,N_14403,N_13766);
xnor U17287 (N_17287,N_15757,N_12328);
nand U17288 (N_17288,N_15012,N_14207);
nand U17289 (N_17289,N_12802,N_14868);
nor U17290 (N_17290,N_13521,N_12210);
nor U17291 (N_17291,N_12918,N_14878);
and U17292 (N_17292,N_14928,N_13211);
nand U17293 (N_17293,N_14509,N_12687);
nand U17294 (N_17294,N_12352,N_15239);
and U17295 (N_17295,N_13458,N_13740);
and U17296 (N_17296,N_14085,N_12546);
nand U17297 (N_17297,N_15029,N_12882);
and U17298 (N_17298,N_14545,N_12513);
nand U17299 (N_17299,N_15945,N_12008);
nand U17300 (N_17300,N_12450,N_14860);
and U17301 (N_17301,N_14183,N_12662);
nand U17302 (N_17302,N_12936,N_12768);
nand U17303 (N_17303,N_13241,N_15925);
nor U17304 (N_17304,N_13149,N_12327);
nor U17305 (N_17305,N_14600,N_15355);
or U17306 (N_17306,N_15708,N_15836);
or U17307 (N_17307,N_15841,N_14206);
nand U17308 (N_17308,N_14377,N_15733);
nor U17309 (N_17309,N_14224,N_13986);
nand U17310 (N_17310,N_15752,N_14615);
nor U17311 (N_17311,N_15024,N_12580);
nand U17312 (N_17312,N_14036,N_13192);
nor U17313 (N_17313,N_12112,N_15137);
and U17314 (N_17314,N_12066,N_14879);
or U17315 (N_17315,N_13507,N_12288);
or U17316 (N_17316,N_12000,N_12178);
nand U17317 (N_17317,N_12480,N_15875);
nand U17318 (N_17318,N_13615,N_12456);
or U17319 (N_17319,N_15395,N_13869);
nand U17320 (N_17320,N_12964,N_12289);
nand U17321 (N_17321,N_14294,N_14922);
nor U17322 (N_17322,N_14657,N_13258);
nand U17323 (N_17323,N_15410,N_14773);
nand U17324 (N_17324,N_13914,N_15749);
or U17325 (N_17325,N_15411,N_13098);
and U17326 (N_17326,N_13198,N_14429);
and U17327 (N_17327,N_15880,N_15905);
or U17328 (N_17328,N_13719,N_13524);
or U17329 (N_17329,N_14623,N_12912);
or U17330 (N_17330,N_13150,N_12721);
or U17331 (N_17331,N_12337,N_12444);
and U17332 (N_17332,N_13781,N_15682);
nor U17333 (N_17333,N_13447,N_13716);
nand U17334 (N_17334,N_13121,N_13222);
and U17335 (N_17335,N_14492,N_13966);
nor U17336 (N_17336,N_12543,N_15756);
or U17337 (N_17337,N_14099,N_12899);
nand U17338 (N_17338,N_14779,N_13206);
and U17339 (N_17339,N_13235,N_15209);
nor U17340 (N_17340,N_15533,N_13233);
or U17341 (N_17341,N_14501,N_15537);
nor U17342 (N_17342,N_12481,N_12526);
nand U17343 (N_17343,N_13325,N_12107);
or U17344 (N_17344,N_14930,N_12709);
and U17345 (N_17345,N_13386,N_13861);
and U17346 (N_17346,N_12742,N_12504);
or U17347 (N_17347,N_12653,N_14551);
nand U17348 (N_17348,N_14960,N_13581);
nand U17349 (N_17349,N_15623,N_13294);
nor U17350 (N_17350,N_14826,N_15092);
and U17351 (N_17351,N_13511,N_13044);
xnor U17352 (N_17352,N_13670,N_15859);
nand U17353 (N_17353,N_12625,N_15226);
or U17354 (N_17354,N_15334,N_15087);
and U17355 (N_17355,N_15647,N_15598);
nor U17356 (N_17356,N_12795,N_12256);
or U17357 (N_17357,N_14351,N_14637);
and U17358 (N_17358,N_15164,N_15656);
nor U17359 (N_17359,N_12051,N_12060);
or U17360 (N_17360,N_14962,N_14322);
nand U17361 (N_17361,N_12584,N_15539);
and U17362 (N_17362,N_12950,N_12726);
or U17363 (N_17363,N_14143,N_15740);
and U17364 (N_17364,N_13016,N_12694);
or U17365 (N_17365,N_15825,N_12649);
nand U17366 (N_17366,N_15867,N_15268);
or U17367 (N_17367,N_15914,N_13377);
and U17368 (N_17368,N_15673,N_15463);
nor U17369 (N_17369,N_15468,N_15503);
and U17370 (N_17370,N_12040,N_12523);
nand U17371 (N_17371,N_12345,N_13731);
nand U17372 (N_17372,N_13828,N_12150);
and U17373 (N_17373,N_15369,N_15048);
and U17374 (N_17374,N_15904,N_12490);
nand U17375 (N_17375,N_12910,N_13529);
or U17376 (N_17376,N_13423,N_13135);
and U17377 (N_17377,N_15281,N_15295);
and U17378 (N_17378,N_14950,N_15386);
or U17379 (N_17379,N_15784,N_15556);
nand U17380 (N_17380,N_12175,N_15350);
or U17381 (N_17381,N_13319,N_15171);
xnor U17382 (N_17382,N_12329,N_15303);
nand U17383 (N_17383,N_14331,N_14821);
nand U17384 (N_17384,N_14175,N_13354);
or U17385 (N_17385,N_15080,N_13005);
or U17386 (N_17386,N_12140,N_15046);
nor U17387 (N_17387,N_12652,N_15439);
and U17388 (N_17388,N_15694,N_12577);
and U17389 (N_17389,N_14424,N_15584);
nor U17390 (N_17390,N_12803,N_15250);
or U17391 (N_17391,N_15954,N_14251);
and U17392 (N_17392,N_15354,N_15842);
or U17393 (N_17393,N_15664,N_13344);
and U17394 (N_17394,N_15594,N_14431);
nor U17395 (N_17395,N_12270,N_15766);
nor U17396 (N_17396,N_13508,N_15321);
and U17397 (N_17397,N_12597,N_12505);
or U17398 (N_17398,N_15639,N_14097);
and U17399 (N_17399,N_14671,N_14575);
nand U17400 (N_17400,N_13161,N_13553);
or U17401 (N_17401,N_13004,N_12954);
and U17402 (N_17402,N_13645,N_12394);
xnor U17403 (N_17403,N_14689,N_15484);
nor U17404 (N_17404,N_12581,N_12916);
and U17405 (N_17405,N_14736,N_14089);
and U17406 (N_17406,N_13382,N_15632);
nand U17407 (N_17407,N_14897,N_14245);
nor U17408 (N_17408,N_15473,N_15224);
or U17409 (N_17409,N_12956,N_12501);
and U17410 (N_17410,N_15980,N_12179);
nand U17411 (N_17411,N_13007,N_14458);
xnor U17412 (N_17412,N_13073,N_14308);
nor U17413 (N_17413,N_15932,N_13059);
nand U17414 (N_17414,N_12718,N_15123);
or U17415 (N_17415,N_13340,N_13124);
and U17416 (N_17416,N_15855,N_12129);
nand U17417 (N_17417,N_14757,N_14073);
nor U17418 (N_17418,N_13918,N_12864);
nand U17419 (N_17419,N_14924,N_15470);
or U17420 (N_17420,N_13189,N_15121);
nand U17421 (N_17421,N_13485,N_12148);
and U17422 (N_17422,N_12762,N_14776);
and U17423 (N_17423,N_13051,N_13533);
and U17424 (N_17424,N_13452,N_15686);
and U17425 (N_17425,N_13266,N_14705);
nor U17426 (N_17426,N_14058,N_13852);
or U17427 (N_17427,N_15073,N_14389);
or U17428 (N_17428,N_14404,N_15890);
and U17429 (N_17429,N_13403,N_13214);
nor U17430 (N_17430,N_14818,N_14414);
nor U17431 (N_17431,N_12108,N_14253);
or U17432 (N_17432,N_14342,N_15274);
nor U17433 (N_17433,N_15920,N_15810);
nor U17434 (N_17434,N_12068,N_13096);
nand U17435 (N_17435,N_14491,N_15765);
or U17436 (N_17436,N_15928,N_15374);
nand U17437 (N_17437,N_14263,N_15139);
or U17438 (N_17438,N_14487,N_13279);
and U17439 (N_17439,N_15431,N_14056);
and U17440 (N_17440,N_15179,N_13797);
nor U17441 (N_17441,N_12385,N_14391);
or U17442 (N_17442,N_14106,N_14793);
nor U17443 (N_17443,N_12674,N_13683);
nand U17444 (N_17444,N_14559,N_15833);
or U17445 (N_17445,N_13338,N_15818);
or U17446 (N_17446,N_14755,N_13288);
and U17447 (N_17447,N_13657,N_14573);
and U17448 (N_17448,N_12379,N_13990);
nand U17449 (N_17449,N_14760,N_13987);
or U17450 (N_17450,N_14794,N_13785);
nand U17451 (N_17451,N_14739,N_14418);
or U17452 (N_17452,N_12555,N_15893);
nor U17453 (N_17453,N_13236,N_14063);
and U17454 (N_17454,N_14964,N_14651);
nor U17455 (N_17455,N_12927,N_14470);
nand U17456 (N_17456,N_15976,N_13475);
nor U17457 (N_17457,N_15259,N_12046);
or U17458 (N_17458,N_15008,N_13071);
nand U17459 (N_17459,N_14677,N_13631);
or U17460 (N_17460,N_12334,N_13014);
or U17461 (N_17461,N_12423,N_15727);
or U17462 (N_17462,N_12360,N_14457);
nand U17463 (N_17463,N_13725,N_13361);
nand U17464 (N_17464,N_12027,N_14631);
or U17465 (N_17465,N_15420,N_13414);
or U17466 (N_17466,N_13818,N_15601);
nand U17467 (N_17467,N_12620,N_13047);
nor U17468 (N_17468,N_14595,N_13366);
nand U17469 (N_17469,N_14465,N_15796);
nand U17470 (N_17470,N_13023,N_15110);
and U17471 (N_17471,N_15942,N_12374);
or U17472 (N_17472,N_13234,N_14303);
and U17473 (N_17473,N_12673,N_12165);
nand U17474 (N_17474,N_15958,N_13972);
nor U17475 (N_17475,N_12984,N_13390);
and U17476 (N_17476,N_15732,N_12683);
and U17477 (N_17477,N_13934,N_13648);
nand U17478 (N_17478,N_12173,N_14544);
nor U17479 (N_17479,N_12992,N_14121);
and U17480 (N_17480,N_13592,N_15175);
and U17481 (N_17481,N_12317,N_13061);
or U17482 (N_17482,N_12878,N_12605);
nand U17483 (N_17483,N_14581,N_12181);
or U17484 (N_17484,N_13229,N_13402);
nand U17485 (N_17485,N_15205,N_13267);
nand U17486 (N_17486,N_13527,N_12564);
and U17487 (N_17487,N_14921,N_14580);
nand U17488 (N_17488,N_15476,N_15309);
or U17489 (N_17489,N_15978,N_13988);
or U17490 (N_17490,N_13070,N_12453);
nand U17491 (N_17491,N_13265,N_12883);
and U17492 (N_17492,N_12177,N_15448);
nor U17493 (N_17493,N_15361,N_13277);
nor U17494 (N_17494,N_13832,N_14530);
and U17495 (N_17495,N_12199,N_12968);
or U17496 (N_17496,N_15871,N_15277);
nor U17497 (N_17497,N_15135,N_13156);
and U17498 (N_17498,N_14578,N_12657);
or U17499 (N_17499,N_12312,N_13973);
or U17500 (N_17500,N_13238,N_14803);
and U17501 (N_17501,N_15344,N_15311);
nand U17502 (N_17502,N_13302,N_14811);
nand U17503 (N_17503,N_14973,N_14931);
or U17504 (N_17504,N_15947,N_14542);
or U17505 (N_17505,N_15305,N_15204);
or U17506 (N_17506,N_15040,N_12656);
nand U17507 (N_17507,N_14929,N_12358);
or U17508 (N_17508,N_12356,N_14525);
xnor U17509 (N_17509,N_15700,N_15621);
and U17510 (N_17510,N_15126,N_14895);
nand U17511 (N_17511,N_13881,N_14152);
and U17512 (N_17512,N_12991,N_12812);
xor U17513 (N_17513,N_12422,N_15791);
and U17514 (N_17514,N_13518,N_14230);
nand U17515 (N_17515,N_14336,N_13145);
nor U17516 (N_17516,N_13369,N_14843);
nor U17517 (N_17517,N_12725,N_15023);
or U17518 (N_17518,N_12825,N_15712);
nand U17519 (N_17519,N_14307,N_12268);
nand U17520 (N_17520,N_13982,N_15805);
nor U17521 (N_17521,N_15216,N_14436);
nand U17522 (N_17522,N_14956,N_15834);
or U17523 (N_17523,N_13953,N_13813);
nand U17524 (N_17524,N_14047,N_13705);
nand U17525 (N_17525,N_12117,N_15877);
nor U17526 (N_17526,N_13065,N_12767);
or U17527 (N_17527,N_14952,N_12305);
nor U17528 (N_17528,N_12719,N_15288);
or U17529 (N_17529,N_14304,N_12220);
nor U17530 (N_17530,N_14648,N_14546);
nand U17531 (N_17531,N_15538,N_12511);
nor U17532 (N_17532,N_14695,N_15199);
nand U17533 (N_17533,N_12114,N_14411);
nor U17534 (N_17534,N_13603,N_14941);
nand U17535 (N_17535,N_12781,N_14359);
or U17536 (N_17536,N_13535,N_13221);
and U17537 (N_17537,N_14726,N_12737);
nand U17538 (N_17538,N_14227,N_15816);
or U17539 (N_17539,N_12593,N_14347);
and U17540 (N_17540,N_15119,N_12452);
nor U17541 (N_17541,N_12382,N_15963);
and U17542 (N_17542,N_15917,N_14330);
or U17543 (N_17543,N_13451,N_12341);
nor U17544 (N_17544,N_15056,N_12834);
nand U17545 (N_17545,N_12458,N_15143);
and U17546 (N_17546,N_12153,N_14332);
nor U17547 (N_17547,N_13967,N_13559);
nor U17548 (N_17548,N_13126,N_14949);
nand U17549 (N_17549,N_14355,N_12152);
and U17550 (N_17550,N_13230,N_13435);
nand U17551 (N_17551,N_14661,N_13912);
nor U17552 (N_17552,N_14522,N_15472);
or U17553 (N_17553,N_12805,N_12502);
nand U17554 (N_17554,N_15166,N_14723);
or U17555 (N_17555,N_12146,N_14217);
nand U17556 (N_17556,N_12205,N_12272);
nor U17557 (N_17557,N_12701,N_12974);
nor U17558 (N_17558,N_13268,N_12835);
nand U17559 (N_17559,N_12090,N_15777);
nor U17560 (N_17560,N_14666,N_12855);
nor U17561 (N_17561,N_12455,N_13376);
and U17562 (N_17562,N_13133,N_12449);
or U17563 (N_17563,N_12366,N_14156);
nor U17564 (N_17564,N_13483,N_12681);
nand U17565 (N_17565,N_14996,N_13844);
and U17566 (N_17566,N_13698,N_15865);
and U17567 (N_17567,N_15530,N_12369);
or U17568 (N_17568,N_12058,N_13998);
or U17569 (N_17569,N_12275,N_15870);
nand U17570 (N_17570,N_13199,N_15456);
nand U17571 (N_17571,N_15953,N_15015);
nor U17572 (N_17572,N_13882,N_12397);
or U17573 (N_17573,N_13519,N_14687);
or U17574 (N_17574,N_12669,N_14598);
and U17575 (N_17575,N_15192,N_14911);
and U17576 (N_17576,N_12018,N_12582);
nor U17577 (N_17577,N_14823,N_14064);
nand U17578 (N_17578,N_13494,N_13693);
and U17579 (N_17579,N_14814,N_14489);
and U17580 (N_17580,N_12428,N_15051);
nand U17581 (N_17581,N_13689,N_12467);
nand U17582 (N_17582,N_12700,N_13109);
and U17583 (N_17583,N_14908,N_15185);
nand U17584 (N_17584,N_14942,N_14426);
and U17585 (N_17585,N_14558,N_13977);
nor U17586 (N_17586,N_13013,N_15574);
nand U17587 (N_17587,N_14074,N_15247);
and U17588 (N_17588,N_15327,N_15316);
nor U17589 (N_17589,N_14880,N_15034);
nand U17590 (N_17590,N_12947,N_13467);
and U17591 (N_17591,N_14384,N_15117);
or U17592 (N_17592,N_13849,N_14474);
nand U17593 (N_17593,N_15390,N_15809);
nor U17594 (N_17594,N_13060,N_13256);
nand U17595 (N_17595,N_15837,N_15445);
or U17596 (N_17596,N_12092,N_14938);
nand U17597 (N_17597,N_15413,N_12686);
nor U17598 (N_17598,N_14804,N_12903);
nand U17599 (N_17599,N_13707,N_12273);
nand U17600 (N_17600,N_15469,N_12823);
nand U17601 (N_17601,N_14193,N_12017);
and U17602 (N_17602,N_12307,N_15931);
or U17603 (N_17603,N_14486,N_12688);
nor U17604 (N_17604,N_15977,N_15878);
and U17605 (N_17605,N_12204,N_14096);
and U17606 (N_17606,N_14590,N_13728);
or U17607 (N_17607,N_15160,N_13637);
and U17608 (N_17608,N_13024,N_13046);
or U17609 (N_17609,N_13991,N_14618);
nand U17610 (N_17610,N_13443,N_13651);
and U17611 (N_17611,N_13398,N_14383);
nand U17612 (N_17612,N_13686,N_14007);
or U17613 (N_17613,N_14464,N_12615);
or U17614 (N_17614,N_14466,N_14733);
nor U17615 (N_17615,N_15151,N_13520);
nand U17616 (N_17616,N_13012,N_14604);
or U17617 (N_17617,N_13762,N_13997);
xor U17618 (N_17618,N_14335,N_14523);
xnor U17619 (N_17619,N_12839,N_14233);
and U17620 (N_17620,N_14103,N_15018);
or U17621 (N_17621,N_14756,N_13924);
and U17622 (N_17622,N_13444,N_12821);
or U17623 (N_17623,N_14560,N_13304);
nor U17624 (N_17624,N_14861,N_14388);
or U17625 (N_17625,N_14094,N_15104);
nand U17626 (N_17626,N_12846,N_15228);
nor U17627 (N_17627,N_13080,N_12837);
nor U17628 (N_17628,N_14077,N_14202);
and U17629 (N_17629,N_15207,N_15112);
xor U17630 (N_17630,N_14029,N_13822);
or U17631 (N_17631,N_13310,N_12313);
or U17632 (N_17632,N_13373,N_15711);
nand U17633 (N_17633,N_13642,N_15419);
nor U17634 (N_17634,N_13326,N_13838);
xnor U17635 (N_17635,N_15568,N_15442);
nor U17636 (N_17636,N_15492,N_15950);
or U17637 (N_17637,N_13764,N_12880);
nor U17638 (N_17638,N_14249,N_14724);
or U17639 (N_17639,N_15125,N_15844);
nand U17640 (N_17640,N_14889,N_12507);
nand U17641 (N_17641,N_14150,N_12338);
and U17642 (N_17642,N_14680,N_13605);
xnor U17643 (N_17643,N_12921,N_13434);
nor U17644 (N_17644,N_14221,N_13202);
and U17645 (N_17645,N_13858,N_12782);
nor U17646 (N_17646,N_12600,N_15918);
nand U17647 (N_17647,N_15033,N_15300);
nor U17648 (N_17648,N_14902,N_12888);
or U17649 (N_17649,N_12525,N_15593);
and U17650 (N_17650,N_12229,N_14543);
or U17651 (N_17651,N_15337,N_12495);
nand U17652 (N_17652,N_13877,N_14467);
nand U17653 (N_17653,N_14668,N_12005);
and U17654 (N_17654,N_15134,N_15229);
or U17655 (N_17655,N_12322,N_12333);
nand U17656 (N_17656,N_13455,N_14285);
and U17657 (N_17657,N_13609,N_13499);
nor U17658 (N_17658,N_15083,N_13949);
or U17659 (N_17659,N_12934,N_15739);
and U17660 (N_17660,N_14682,N_12026);
or U17661 (N_17661,N_13062,N_15862);
or U17662 (N_17662,N_15444,N_12048);
or U17663 (N_17663,N_15044,N_14752);
nand U17664 (N_17664,N_15315,N_13381);
or U17665 (N_17665,N_14385,N_15433);
nand U17666 (N_17666,N_12663,N_13480);
nor U17667 (N_17667,N_13666,N_12314);
nor U17668 (N_17668,N_12791,N_15678);
xnor U17669 (N_17669,N_13876,N_13054);
nand U17670 (N_17670,N_15235,N_12080);
and U17671 (N_17671,N_15172,N_14740);
nor U17672 (N_17672,N_13627,N_13820);
or U17673 (N_17673,N_15927,N_13257);
and U17674 (N_17674,N_15511,N_13870);
or U17675 (N_17675,N_13383,N_14082);
nor U17676 (N_17676,N_13901,N_13767);
nand U17677 (N_17677,N_12986,N_12007);
nand U17678 (N_17678,N_15567,N_13751);
nand U17679 (N_17679,N_13944,N_15638);
nand U17680 (N_17680,N_14737,N_13329);
nand U17681 (N_17681,N_15460,N_12469);
nand U17682 (N_17682,N_12613,N_12749);
nand U17683 (N_17683,N_12055,N_15670);
or U17684 (N_17684,N_14428,N_15677);
nand U17685 (N_17685,N_12838,N_15910);
or U17686 (N_17686,N_15081,N_15276);
or U17687 (N_17687,N_15886,N_12772);
and U17688 (N_17688,N_13438,N_13433);
and U17689 (N_17689,N_13287,N_13490);
nor U17690 (N_17690,N_15985,N_14195);
or U17691 (N_17691,N_15577,N_12122);
nand U17692 (N_17692,N_12808,N_14660);
and U17693 (N_17693,N_15625,N_13786);
nor U17694 (N_17694,N_13284,N_12820);
nand U17695 (N_17695,N_15380,N_15394);
or U17696 (N_17696,N_14444,N_15459);
nand U17697 (N_17697,N_14001,N_15285);
and U17698 (N_17698,N_12362,N_12164);
and U17699 (N_17699,N_13866,N_14596);
or U17700 (N_17700,N_15149,N_15713);
or U17701 (N_17701,N_13791,N_12447);
and U17702 (N_17702,N_13732,N_15619);
nand U17703 (N_17703,N_13058,N_12154);
or U17704 (N_17704,N_15054,N_13892);
and U17705 (N_17705,N_15970,N_14279);
xnor U17706 (N_17706,N_14777,N_13808);
nor U17707 (N_17707,N_15499,N_13939);
and U17708 (N_17708,N_12904,N_12659);
or U17709 (N_17709,N_15027,N_15653);
or U17710 (N_17710,N_13040,N_13456);
nor U17711 (N_17711,N_12211,N_13232);
and U17712 (N_17712,N_12036,N_12491);
nor U17713 (N_17713,N_12953,N_12707);
and U17714 (N_17714,N_14281,N_13669);
nand U17715 (N_17715,N_13729,N_12623);
nand U17716 (N_17716,N_15544,N_12551);
nor U17717 (N_17717,N_13695,N_13305);
and U17718 (N_17718,N_13640,N_12295);
or U17719 (N_17719,N_14571,N_13907);
nand U17720 (N_17720,N_12132,N_13394);
or U17721 (N_17721,N_14624,N_12286);
nor U17722 (N_17722,N_15495,N_13673);
or U17723 (N_17723,N_13118,N_15659);
nand U17724 (N_17724,N_13938,N_13787);
xnor U17725 (N_17725,N_12402,N_13993);
nand U17726 (N_17726,N_14490,N_13042);
nand U17727 (N_17727,N_12355,N_15799);
or U17728 (N_17728,N_14820,N_14747);
and U17729 (N_17729,N_14306,N_14040);
nand U17730 (N_17730,N_12610,N_13633);
or U17731 (N_17731,N_14083,N_15452);
nor U17732 (N_17732,N_14014,N_12433);
nor U17733 (N_17733,N_13021,N_15283);
nor U17734 (N_17734,N_13412,N_13558);
or U17735 (N_17735,N_13166,N_14135);
nor U17736 (N_17736,N_15069,N_13540);
nor U17737 (N_17737,N_15807,N_13960);
nand U17738 (N_17738,N_14371,N_12710);
nand U17739 (N_17739,N_14352,N_14399);
or U17740 (N_17740,N_15326,N_12886);
and U17741 (N_17741,N_14848,N_13940);
nor U17742 (N_17742,N_13449,N_14844);
or U17743 (N_17743,N_15003,N_13904);
nor U17744 (N_17744,N_13500,N_13462);
and U17745 (N_17745,N_14290,N_14186);
nand U17746 (N_17746,N_14864,N_15415);
nor U17747 (N_17747,N_13807,N_15658);
nor U17748 (N_17748,N_12271,N_15759);
nor U17749 (N_17749,N_15036,N_15240);
nor U17750 (N_17750,N_13367,N_13094);
nor U17751 (N_17751,N_12209,N_15084);
nor U17752 (N_17752,N_13564,N_15767);
nor U17753 (N_17753,N_15962,N_12598);
nor U17754 (N_17754,N_13571,N_12816);
and U17755 (N_17755,N_13110,N_14423);
or U17756 (N_17756,N_14108,N_13644);
nand U17757 (N_17757,N_15937,N_14033);
or U17758 (N_17758,N_15743,N_15466);
and U17759 (N_17759,N_15775,N_15690);
and U17760 (N_17760,N_12989,N_13186);
and U17761 (N_17761,N_13193,N_15672);
nor U17762 (N_17762,N_12309,N_15351);
and U17763 (N_17763,N_12766,N_13911);
nand U17764 (N_17764,N_15428,N_14282);
nor U17765 (N_17765,N_15518,N_13188);
nand U17766 (N_17766,N_14287,N_14111);
nor U17767 (N_17767,N_15988,N_14999);
xnor U17768 (N_17768,N_13894,N_12149);
and U17769 (N_17769,N_15588,N_13100);
and U17770 (N_17770,N_12022,N_12734);
and U17771 (N_17771,N_12240,N_14163);
nand U17772 (N_17772,N_14681,N_14622);
and U17773 (N_17773,N_14425,N_12476);
nand U17774 (N_17774,N_14767,N_14577);
or U17775 (N_17775,N_14148,N_13492);
and U17776 (N_17776,N_12343,N_15031);
or U17777 (N_17777,N_12898,N_15421);
and U17778 (N_17778,N_14987,N_14129);
and U17779 (N_17779,N_13713,N_12736);
nand U17780 (N_17780,N_13471,N_15132);
nand U17781 (N_17781,N_14373,N_12981);
or U17782 (N_17782,N_15726,N_13709);
or U17783 (N_17783,N_15760,N_12078);
xnor U17784 (N_17784,N_12549,N_15181);
and U17785 (N_17785,N_13252,N_15813);
or U17786 (N_17786,N_14852,N_15317);
and U17787 (N_17787,N_14995,N_14943);
or U17788 (N_17788,N_14445,N_14934);
nor U17789 (N_17789,N_12206,N_15441);
nand U17790 (N_17790,N_14356,N_12488);
nand U17791 (N_17791,N_15437,N_12599);
and U17792 (N_17792,N_14453,N_13788);
nand U17793 (N_17793,N_15551,N_14081);
and U17794 (N_17794,N_14998,N_13092);
nor U17795 (N_17795,N_12754,N_14420);
nor U17796 (N_17796,N_15508,N_13341);
and U17797 (N_17797,N_14554,N_12056);
nor U17798 (N_17798,N_12790,N_15852);
nor U17799 (N_17799,N_12666,N_14712);
or U17800 (N_17800,N_15744,N_14412);
or U17801 (N_17801,N_15077,N_12019);
or U17802 (N_17802,N_13407,N_15983);
or U17803 (N_17803,N_14915,N_14144);
or U17804 (N_17804,N_15984,N_13293);
nor U17805 (N_17805,N_15010,N_13307);
or U17806 (N_17806,N_15242,N_14706);
nor U17807 (N_17807,N_12845,N_12644);
nand U17808 (N_17808,N_15182,N_13191);
or U17809 (N_17809,N_12197,N_14599);
and U17810 (N_17810,N_14041,N_13720);
nand U17811 (N_17811,N_13514,N_14104);
and U17812 (N_17812,N_15106,N_12418);
or U17813 (N_17813,N_12176,N_13654);
nor U17814 (N_17814,N_13289,N_15801);
or U17815 (N_17815,N_13626,N_14127);
or U17816 (N_17816,N_15640,N_13420);
and U17817 (N_17817,N_14876,N_13607);
or U17818 (N_17818,N_14702,N_15919);
or U17819 (N_17819,N_13331,N_14965);
or U17820 (N_17820,N_12890,N_15636);
or U17821 (N_17821,N_12848,N_15258);
and U17822 (N_17822,N_15897,N_14116);
nand U17823 (N_17823,N_13814,N_13505);
nor U17824 (N_17824,N_13410,N_15165);
nand U17825 (N_17825,N_12951,N_15146);
nor U17826 (N_17826,N_15450,N_15114);
or U17827 (N_17827,N_15443,N_13389);
nand U17828 (N_17828,N_13922,N_15312);
nor U17829 (N_17829,N_14791,N_13522);
or U17830 (N_17830,N_12753,N_13493);
nand U17831 (N_17831,N_14775,N_13909);
and U17832 (N_17832,N_14579,N_13979);
or U17833 (N_17833,N_13946,N_13316);
nand U17834 (N_17834,N_12415,N_13127);
nor U17835 (N_17835,N_15275,N_14990);
and U17836 (N_17836,N_12063,N_14685);
and U17837 (N_17837,N_12044,N_12219);
nand U17838 (N_17838,N_13035,N_14991);
and U17839 (N_17839,N_13029,N_14049);
nand U17840 (N_17840,N_12866,N_12384);
nor U17841 (N_17841,N_13077,N_12408);
and U17842 (N_17842,N_12828,N_14076);
nand U17843 (N_17843,N_13184,N_14905);
or U17844 (N_17844,N_15803,N_15251);
nand U17845 (N_17845,N_14953,N_14203);
nand U17846 (N_17846,N_13496,N_12131);
or U17847 (N_17847,N_14437,N_15435);
nand U17848 (N_17848,N_13915,N_15263);
nor U17849 (N_17849,N_12493,N_12759);
or U17850 (N_17850,N_12789,N_13501);
nand U17851 (N_17851,N_12608,N_14080);
nor U17852 (N_17852,N_14098,N_15115);
nand U17853 (N_17853,N_12919,N_14518);
nand U17854 (N_17854,N_13783,N_14904);
or U17855 (N_17855,N_15724,N_13575);
nor U17856 (N_17856,N_13799,N_13350);
nand U17857 (N_17857,N_12316,N_14957);
or U17858 (N_17858,N_12553,N_14088);
nor U17859 (N_17859,N_12569,N_13335);
nor U17860 (N_17860,N_14802,N_14932);
and U17861 (N_17861,N_15070,N_12588);
and U17862 (N_17862,N_15025,N_15336);
and U17863 (N_17863,N_15290,N_13616);
or U17864 (N_17864,N_14846,N_14456);
nand U17865 (N_17865,N_14032,N_15971);
nor U17866 (N_17866,N_14899,N_12524);
nor U17867 (N_17867,N_15742,N_12170);
and U17868 (N_17868,N_14339,N_12868);
or U17869 (N_17869,N_12874,N_15600);
and U17870 (N_17870,N_15798,N_12699);
or U17871 (N_17871,N_13542,N_15282);
nand U17872 (N_17872,N_13641,N_15730);
nand U17873 (N_17873,N_13602,N_12632);
nand U17874 (N_17874,N_15486,N_14471);
nor U17875 (N_17875,N_14833,N_15892);
and U17876 (N_17876,N_12639,N_15122);
nand U17877 (N_17877,N_14188,N_14913);
and U17878 (N_17878,N_14250,N_12804);
nand U17879 (N_17879,N_13588,N_15587);
and U17880 (N_17880,N_14232,N_12905);
and U17881 (N_17881,N_15908,N_13217);
nor U17882 (N_17882,N_13680,N_14297);
or U17883 (N_17883,N_13474,N_14866);
or U17884 (N_17884,N_12254,N_13158);
nand U17885 (N_17885,N_13050,N_13043);
and U17886 (N_17886,N_12708,N_12155);
or U17887 (N_17887,N_12182,N_15680);
xnor U17888 (N_17888,N_13902,N_13334);
nor U17889 (N_17889,N_13932,N_14182);
or U17890 (N_17890,N_15188,N_14050);
nand U17891 (N_17891,N_15489,N_15668);
nor U17892 (N_17892,N_13846,N_15981);
or U17893 (N_17893,N_15575,N_13372);
nand U17894 (N_17894,N_14243,N_15956);
nand U17895 (N_17895,N_13597,N_15589);
nor U17896 (N_17896,N_13920,N_15517);
or U17897 (N_17897,N_12387,N_12296);
or U17898 (N_17898,N_12344,N_15564);
and U17899 (N_17899,N_14847,N_15358);
nor U17900 (N_17900,N_15255,N_14003);
and U17901 (N_17901,N_14407,N_15086);
nor U17902 (N_17902,N_14318,N_13280);
nor U17903 (N_17903,N_12189,N_13425);
nand U17904 (N_17904,N_12315,N_15385);
nor U17905 (N_17905,N_13401,N_12143);
nor U17906 (N_17906,N_14655,N_12225);
nor U17907 (N_17907,N_13272,N_15298);
nand U17908 (N_17908,N_15296,N_14382);
xnor U17909 (N_17909,N_13959,N_15995);
or U17910 (N_17910,N_13162,N_13541);
nor U17911 (N_17911,N_14506,N_14568);
nor U17912 (N_17912,N_15043,N_12023);
nand U17913 (N_17913,N_15562,N_13095);
nand U17914 (N_17914,N_15969,N_14534);
or U17915 (N_17915,N_12778,N_15527);
nand U17916 (N_17916,N_14433,N_13723);
nand U17917 (N_17917,N_15790,N_14095);
and U17918 (N_17918,N_12348,N_12861);
or U17919 (N_17919,N_13794,N_14856);
nand U17920 (N_17920,N_12542,N_12342);
or U17921 (N_17921,N_15566,N_12799);
or U17922 (N_17922,N_12602,N_12723);
or U17923 (N_17923,N_13908,N_15297);
nor U17924 (N_17924,N_13157,N_13958);
or U17925 (N_17925,N_14688,N_12276);
or U17926 (N_17926,N_13460,N_13253);
nor U17927 (N_17927,N_15602,N_15853);
nor U17928 (N_17928,N_12255,N_13856);
nand U17929 (N_17929,N_12590,N_15933);
and U17930 (N_17930,N_14867,N_12294);
or U17931 (N_17931,N_15753,N_12244);
nor U17932 (N_17932,N_15232,N_14912);
nand U17933 (N_17933,N_14130,N_13671);
nand U17934 (N_17934,N_12202,N_14824);
nor U17935 (N_17935,N_15891,N_13653);
or U17936 (N_17936,N_12167,N_14038);
or U17937 (N_17937,N_13659,N_12079);
or U17938 (N_17938,N_15560,N_13692);
nand U17939 (N_17939,N_12109,N_15735);
nand U17940 (N_17940,N_12573,N_13107);
xor U17941 (N_17941,N_14274,N_14276);
and U17942 (N_17942,N_13352,N_13215);
or U17943 (N_17943,N_15597,N_15558);
or U17944 (N_17944,N_14834,N_12679);
and U17945 (N_17945,N_15975,N_14500);
and U17946 (N_17946,N_12437,N_12810);
nor U17947 (N_17947,N_12098,N_15409);
or U17948 (N_17948,N_15292,N_15899);
and U17949 (N_17949,N_12665,N_12497);
or U17950 (N_17950,N_13768,N_12732);
or U17951 (N_17951,N_13259,N_13842);
and U17952 (N_17952,N_13119,N_13010);
nand U17953 (N_17953,N_14698,N_15109);
nor U17954 (N_17954,N_13240,N_14114);
or U17955 (N_17955,N_12236,N_12425);
or U17956 (N_17956,N_12860,N_13795);
nand U17957 (N_17957,N_15773,N_12226);
or U17958 (N_17958,N_14887,N_12201);
nor U17959 (N_17959,N_15741,N_14158);
and U17960 (N_17960,N_14713,N_14809);
or U17961 (N_17961,N_14189,N_13395);
nand U17962 (N_17962,N_14989,N_14372);
nor U17963 (N_17963,N_12660,N_14432);
nand U17964 (N_17964,N_15091,N_14126);
nand U17965 (N_17965,N_12034,N_12691);
nor U17966 (N_17966,N_13479,N_13739);
and U17967 (N_17967,N_12512,N_13457);
nand U17968 (N_17968,N_15158,N_12115);
nor U17969 (N_17969,N_12646,N_12368);
and U17970 (N_17970,N_14951,N_13620);
and U17971 (N_17971,N_15605,N_12303);
nand U17972 (N_17972,N_14275,N_15323);
nand U17973 (N_17973,N_12629,N_12676);
nand U17974 (N_17974,N_12562,N_12585);
nor U17975 (N_17975,N_12279,N_15857);
and U17976 (N_17976,N_13891,N_14587);
and U17977 (N_17977,N_13665,N_12214);
or U17978 (N_17978,N_15196,N_14699);
or U17979 (N_17979,N_15039,N_14419);
and U17980 (N_17980,N_13089,N_12571);
nand U17981 (N_17981,N_14170,N_14684);
nor U17982 (N_17982,N_15157,N_13097);
or U17983 (N_17983,N_14345,N_15405);
nand U17984 (N_17984,N_13769,N_13477);
nor U17985 (N_17985,N_12923,N_13552);
nand U17986 (N_17986,N_13730,N_13175);
or U17987 (N_17987,N_13699,N_13348);
and U17988 (N_17988,N_13996,N_13576);
nor U17989 (N_17989,N_15461,N_14674);
or U17990 (N_17990,N_13203,N_12503);
nor U17991 (N_17991,N_13718,N_12161);
nand U17992 (N_17992,N_13872,N_15174);
and U17993 (N_17993,N_13057,N_14529);
xor U17994 (N_17994,N_15716,N_15398);
or U17995 (N_17995,N_15032,N_15062);
or U17996 (N_17996,N_14434,N_15075);
and U17997 (N_17997,N_13484,N_14039);
nor U17998 (N_17998,N_12050,N_14161);
and U17999 (N_17999,N_13388,N_12168);
or U18000 (N_18000,N_12350,N_15769);
and U18001 (N_18001,N_14261,N_12398);
or U18002 (N_18002,N_12523,N_15618);
nor U18003 (N_18003,N_15534,N_14614);
and U18004 (N_18004,N_12471,N_14921);
or U18005 (N_18005,N_14843,N_12284);
nand U18006 (N_18006,N_14701,N_12063);
nand U18007 (N_18007,N_14482,N_14856);
or U18008 (N_18008,N_14631,N_14331);
nand U18009 (N_18009,N_13772,N_14875);
or U18010 (N_18010,N_13507,N_13789);
or U18011 (N_18011,N_14167,N_15623);
or U18012 (N_18012,N_12555,N_12639);
nand U18013 (N_18013,N_12475,N_14646);
or U18014 (N_18014,N_14286,N_15606);
or U18015 (N_18015,N_12618,N_14473);
nand U18016 (N_18016,N_14695,N_15631);
or U18017 (N_18017,N_13894,N_15488);
or U18018 (N_18018,N_15973,N_12885);
or U18019 (N_18019,N_13602,N_12375);
or U18020 (N_18020,N_15566,N_14083);
nand U18021 (N_18021,N_12866,N_13424);
or U18022 (N_18022,N_12561,N_14994);
or U18023 (N_18023,N_14078,N_14625);
or U18024 (N_18024,N_14262,N_13328);
or U18025 (N_18025,N_13516,N_13947);
and U18026 (N_18026,N_15355,N_12181);
nor U18027 (N_18027,N_13670,N_15664);
nor U18028 (N_18028,N_13839,N_15320);
nor U18029 (N_18029,N_13106,N_12233);
nand U18030 (N_18030,N_13541,N_12814);
or U18031 (N_18031,N_15845,N_14544);
and U18032 (N_18032,N_13043,N_13925);
and U18033 (N_18033,N_12634,N_14702);
nand U18034 (N_18034,N_14561,N_13686);
and U18035 (N_18035,N_15439,N_15741);
nor U18036 (N_18036,N_14228,N_15367);
nor U18037 (N_18037,N_14044,N_12317);
and U18038 (N_18038,N_14743,N_12036);
nor U18039 (N_18039,N_14255,N_12363);
nor U18040 (N_18040,N_14870,N_13144);
nor U18041 (N_18041,N_15164,N_15659);
or U18042 (N_18042,N_13217,N_15432);
or U18043 (N_18043,N_15238,N_12100);
and U18044 (N_18044,N_14839,N_14466);
nand U18045 (N_18045,N_15809,N_15012);
nor U18046 (N_18046,N_12394,N_15858);
and U18047 (N_18047,N_15149,N_14536);
or U18048 (N_18048,N_15928,N_14333);
nor U18049 (N_18049,N_14608,N_14739);
or U18050 (N_18050,N_15377,N_14283);
nor U18051 (N_18051,N_13998,N_13810);
nand U18052 (N_18052,N_12413,N_13482);
nor U18053 (N_18053,N_13836,N_14586);
or U18054 (N_18054,N_15092,N_15301);
nand U18055 (N_18055,N_13622,N_13465);
nand U18056 (N_18056,N_13177,N_15136);
or U18057 (N_18057,N_15498,N_14829);
nor U18058 (N_18058,N_14263,N_14813);
nand U18059 (N_18059,N_12623,N_14027);
nand U18060 (N_18060,N_14779,N_12734);
and U18061 (N_18061,N_14351,N_15640);
nand U18062 (N_18062,N_13599,N_12492);
nor U18063 (N_18063,N_15667,N_15779);
and U18064 (N_18064,N_15275,N_13437);
or U18065 (N_18065,N_14221,N_14459);
or U18066 (N_18066,N_15544,N_14119);
and U18067 (N_18067,N_13800,N_13168);
and U18068 (N_18068,N_14476,N_12489);
nand U18069 (N_18069,N_14015,N_15319);
and U18070 (N_18070,N_12778,N_12694);
nor U18071 (N_18071,N_14032,N_13311);
nand U18072 (N_18072,N_15431,N_15215);
or U18073 (N_18073,N_12090,N_12887);
nor U18074 (N_18074,N_14306,N_13840);
or U18075 (N_18075,N_13959,N_15661);
or U18076 (N_18076,N_15736,N_15544);
nor U18077 (N_18077,N_15960,N_14734);
nor U18078 (N_18078,N_15327,N_15638);
or U18079 (N_18079,N_14873,N_15881);
nand U18080 (N_18080,N_15300,N_12406);
or U18081 (N_18081,N_14698,N_13119);
or U18082 (N_18082,N_12460,N_13943);
or U18083 (N_18083,N_15481,N_12211);
nor U18084 (N_18084,N_13806,N_12299);
and U18085 (N_18085,N_14452,N_13965);
or U18086 (N_18086,N_15134,N_13117);
nand U18087 (N_18087,N_13946,N_15829);
and U18088 (N_18088,N_12755,N_13367);
nand U18089 (N_18089,N_14622,N_15186);
or U18090 (N_18090,N_14995,N_13611);
nor U18091 (N_18091,N_13094,N_15249);
nand U18092 (N_18092,N_13266,N_13590);
nor U18093 (N_18093,N_14833,N_14673);
nand U18094 (N_18094,N_14338,N_13764);
and U18095 (N_18095,N_15246,N_12065);
and U18096 (N_18096,N_14325,N_14756);
and U18097 (N_18097,N_13420,N_15834);
nand U18098 (N_18098,N_13135,N_13262);
or U18099 (N_18099,N_12029,N_14190);
or U18100 (N_18100,N_14605,N_12148);
nand U18101 (N_18101,N_15418,N_13862);
or U18102 (N_18102,N_15246,N_15153);
and U18103 (N_18103,N_12049,N_15694);
nor U18104 (N_18104,N_15534,N_15179);
nand U18105 (N_18105,N_15430,N_14112);
nand U18106 (N_18106,N_14327,N_12776);
and U18107 (N_18107,N_13278,N_13883);
nor U18108 (N_18108,N_15620,N_14063);
nor U18109 (N_18109,N_12455,N_14001);
nand U18110 (N_18110,N_13534,N_12809);
nor U18111 (N_18111,N_13949,N_13060);
or U18112 (N_18112,N_14944,N_14649);
and U18113 (N_18113,N_13249,N_12840);
and U18114 (N_18114,N_14610,N_13480);
nand U18115 (N_18115,N_13720,N_12278);
nand U18116 (N_18116,N_15648,N_13800);
nand U18117 (N_18117,N_13494,N_14977);
nand U18118 (N_18118,N_14650,N_14617);
and U18119 (N_18119,N_15804,N_14628);
and U18120 (N_18120,N_13658,N_12354);
nor U18121 (N_18121,N_15979,N_14140);
nand U18122 (N_18122,N_13657,N_15742);
and U18123 (N_18123,N_13050,N_14239);
or U18124 (N_18124,N_15473,N_12021);
nor U18125 (N_18125,N_13090,N_14902);
and U18126 (N_18126,N_13592,N_12515);
and U18127 (N_18127,N_14027,N_13872);
nor U18128 (N_18128,N_13892,N_13416);
nor U18129 (N_18129,N_12340,N_15019);
nand U18130 (N_18130,N_12066,N_14116);
nand U18131 (N_18131,N_13471,N_14698);
or U18132 (N_18132,N_12184,N_13041);
or U18133 (N_18133,N_13716,N_12859);
or U18134 (N_18134,N_15243,N_14435);
or U18135 (N_18135,N_14951,N_15279);
nand U18136 (N_18136,N_12948,N_15201);
and U18137 (N_18137,N_13235,N_15597);
nand U18138 (N_18138,N_15802,N_12217);
nand U18139 (N_18139,N_13018,N_12806);
nand U18140 (N_18140,N_14203,N_13699);
or U18141 (N_18141,N_12074,N_13040);
nand U18142 (N_18142,N_12100,N_12932);
nand U18143 (N_18143,N_15551,N_15008);
nand U18144 (N_18144,N_13822,N_13733);
nor U18145 (N_18145,N_15638,N_13762);
nand U18146 (N_18146,N_14514,N_15566);
and U18147 (N_18147,N_14977,N_13241);
nand U18148 (N_18148,N_15348,N_13346);
or U18149 (N_18149,N_12727,N_14341);
or U18150 (N_18150,N_15216,N_13743);
or U18151 (N_18151,N_12542,N_12158);
or U18152 (N_18152,N_14919,N_12487);
and U18153 (N_18153,N_12215,N_14599);
or U18154 (N_18154,N_12060,N_14958);
and U18155 (N_18155,N_14474,N_12781);
or U18156 (N_18156,N_13632,N_12459);
or U18157 (N_18157,N_12733,N_12678);
and U18158 (N_18158,N_12573,N_14795);
and U18159 (N_18159,N_12042,N_15044);
and U18160 (N_18160,N_15367,N_13805);
nand U18161 (N_18161,N_12728,N_13497);
nor U18162 (N_18162,N_13504,N_15322);
nor U18163 (N_18163,N_14849,N_13401);
nand U18164 (N_18164,N_14966,N_12031);
and U18165 (N_18165,N_15552,N_13156);
nor U18166 (N_18166,N_14685,N_15041);
nor U18167 (N_18167,N_12755,N_12442);
and U18168 (N_18168,N_14896,N_12098);
nor U18169 (N_18169,N_14772,N_14261);
and U18170 (N_18170,N_14091,N_15676);
and U18171 (N_18171,N_15912,N_15081);
nand U18172 (N_18172,N_15939,N_14375);
nor U18173 (N_18173,N_12515,N_14484);
or U18174 (N_18174,N_13389,N_15996);
and U18175 (N_18175,N_13336,N_13375);
and U18176 (N_18176,N_15881,N_15164);
nor U18177 (N_18177,N_14061,N_14431);
and U18178 (N_18178,N_13794,N_13241);
or U18179 (N_18179,N_13641,N_13687);
and U18180 (N_18180,N_13922,N_15330);
and U18181 (N_18181,N_12513,N_12589);
nand U18182 (N_18182,N_12735,N_12236);
or U18183 (N_18183,N_12984,N_14036);
and U18184 (N_18184,N_14113,N_14446);
or U18185 (N_18185,N_15047,N_14110);
and U18186 (N_18186,N_12912,N_15665);
nand U18187 (N_18187,N_12069,N_15647);
nand U18188 (N_18188,N_12137,N_12096);
and U18189 (N_18189,N_14310,N_12809);
and U18190 (N_18190,N_13593,N_12293);
or U18191 (N_18191,N_14504,N_13332);
nand U18192 (N_18192,N_13391,N_15472);
or U18193 (N_18193,N_13285,N_15426);
nor U18194 (N_18194,N_14231,N_15055);
nand U18195 (N_18195,N_14589,N_13325);
or U18196 (N_18196,N_13283,N_13807);
and U18197 (N_18197,N_14543,N_12385);
or U18198 (N_18198,N_13197,N_14114);
nor U18199 (N_18199,N_14999,N_12890);
or U18200 (N_18200,N_15039,N_15394);
or U18201 (N_18201,N_15802,N_15654);
and U18202 (N_18202,N_15703,N_13257);
and U18203 (N_18203,N_13209,N_13372);
and U18204 (N_18204,N_15309,N_15478);
nor U18205 (N_18205,N_14321,N_14175);
nand U18206 (N_18206,N_12867,N_14618);
and U18207 (N_18207,N_13927,N_13819);
nor U18208 (N_18208,N_12055,N_15715);
or U18209 (N_18209,N_14623,N_15326);
or U18210 (N_18210,N_13845,N_13366);
nor U18211 (N_18211,N_15914,N_12678);
and U18212 (N_18212,N_13362,N_14477);
or U18213 (N_18213,N_15144,N_15236);
and U18214 (N_18214,N_15096,N_15976);
or U18215 (N_18215,N_12445,N_13672);
nor U18216 (N_18216,N_14293,N_14424);
and U18217 (N_18217,N_12720,N_15752);
nor U18218 (N_18218,N_12531,N_15991);
and U18219 (N_18219,N_15846,N_13705);
xor U18220 (N_18220,N_12522,N_13182);
and U18221 (N_18221,N_12740,N_12553);
nand U18222 (N_18222,N_14695,N_15799);
or U18223 (N_18223,N_15735,N_14820);
nand U18224 (N_18224,N_12311,N_12424);
nand U18225 (N_18225,N_14563,N_15528);
and U18226 (N_18226,N_15839,N_14614);
nor U18227 (N_18227,N_15074,N_15790);
or U18228 (N_18228,N_13654,N_12426);
nor U18229 (N_18229,N_15196,N_12107);
and U18230 (N_18230,N_12027,N_15217);
and U18231 (N_18231,N_13547,N_15262);
nand U18232 (N_18232,N_15655,N_15161);
and U18233 (N_18233,N_12617,N_13554);
and U18234 (N_18234,N_13391,N_15711);
nand U18235 (N_18235,N_12827,N_13977);
or U18236 (N_18236,N_15354,N_13128);
and U18237 (N_18237,N_15864,N_15716);
and U18238 (N_18238,N_12969,N_15883);
nor U18239 (N_18239,N_12781,N_12615);
or U18240 (N_18240,N_13114,N_13796);
or U18241 (N_18241,N_13680,N_12210);
or U18242 (N_18242,N_13069,N_15376);
nor U18243 (N_18243,N_15502,N_15476);
and U18244 (N_18244,N_12176,N_15642);
and U18245 (N_18245,N_13504,N_12230);
or U18246 (N_18246,N_14233,N_13762);
nor U18247 (N_18247,N_15037,N_15912);
or U18248 (N_18248,N_12775,N_14300);
nand U18249 (N_18249,N_12778,N_15549);
and U18250 (N_18250,N_15707,N_13795);
nand U18251 (N_18251,N_12355,N_12735);
nand U18252 (N_18252,N_14834,N_15172);
nor U18253 (N_18253,N_13656,N_13874);
and U18254 (N_18254,N_13996,N_15725);
and U18255 (N_18255,N_12068,N_12926);
nor U18256 (N_18256,N_14018,N_13977);
and U18257 (N_18257,N_14903,N_15695);
and U18258 (N_18258,N_13009,N_15092);
and U18259 (N_18259,N_15604,N_14756);
or U18260 (N_18260,N_15573,N_15482);
nor U18261 (N_18261,N_13094,N_13032);
nand U18262 (N_18262,N_12038,N_15225);
or U18263 (N_18263,N_14989,N_12716);
nor U18264 (N_18264,N_12058,N_14019);
or U18265 (N_18265,N_13780,N_15404);
or U18266 (N_18266,N_15199,N_15194);
nor U18267 (N_18267,N_13750,N_12203);
or U18268 (N_18268,N_13238,N_13460);
nor U18269 (N_18269,N_12293,N_13461);
xor U18270 (N_18270,N_13190,N_15390);
nor U18271 (N_18271,N_15321,N_15961);
or U18272 (N_18272,N_15111,N_13512);
or U18273 (N_18273,N_13467,N_12687);
and U18274 (N_18274,N_13176,N_13201);
nor U18275 (N_18275,N_12061,N_13796);
and U18276 (N_18276,N_15109,N_13549);
nand U18277 (N_18277,N_15127,N_14318);
or U18278 (N_18278,N_13737,N_14302);
nor U18279 (N_18279,N_12272,N_14779);
nor U18280 (N_18280,N_13388,N_14752);
and U18281 (N_18281,N_15537,N_15671);
nand U18282 (N_18282,N_13654,N_15870);
and U18283 (N_18283,N_14723,N_15746);
or U18284 (N_18284,N_13592,N_13523);
and U18285 (N_18285,N_15970,N_15915);
nand U18286 (N_18286,N_13768,N_13681);
nand U18287 (N_18287,N_13153,N_15426);
nor U18288 (N_18288,N_13456,N_13307);
nor U18289 (N_18289,N_13981,N_13199);
or U18290 (N_18290,N_15702,N_15319);
or U18291 (N_18291,N_14190,N_12990);
nand U18292 (N_18292,N_15293,N_12691);
or U18293 (N_18293,N_15504,N_12498);
and U18294 (N_18294,N_15789,N_15282);
and U18295 (N_18295,N_13480,N_12585);
or U18296 (N_18296,N_14733,N_12968);
nor U18297 (N_18297,N_12159,N_14211);
or U18298 (N_18298,N_13741,N_15970);
nand U18299 (N_18299,N_15232,N_14117);
nand U18300 (N_18300,N_12189,N_15623);
and U18301 (N_18301,N_15852,N_15942);
nand U18302 (N_18302,N_15593,N_13987);
or U18303 (N_18303,N_14931,N_14863);
and U18304 (N_18304,N_14459,N_15033);
nor U18305 (N_18305,N_13719,N_13982);
nor U18306 (N_18306,N_13281,N_15888);
or U18307 (N_18307,N_14373,N_13877);
nand U18308 (N_18308,N_15161,N_13330);
and U18309 (N_18309,N_12082,N_14820);
and U18310 (N_18310,N_12899,N_12885);
nor U18311 (N_18311,N_12071,N_15850);
nor U18312 (N_18312,N_15254,N_12349);
and U18313 (N_18313,N_14602,N_13747);
nand U18314 (N_18314,N_15277,N_13121);
nand U18315 (N_18315,N_15376,N_12474);
nor U18316 (N_18316,N_15824,N_13061);
and U18317 (N_18317,N_14700,N_12459);
and U18318 (N_18318,N_13631,N_15552);
nor U18319 (N_18319,N_12198,N_15860);
nor U18320 (N_18320,N_12965,N_12707);
nor U18321 (N_18321,N_15225,N_14024);
and U18322 (N_18322,N_13721,N_13027);
or U18323 (N_18323,N_14147,N_13977);
or U18324 (N_18324,N_15185,N_12286);
and U18325 (N_18325,N_12256,N_13044);
or U18326 (N_18326,N_15902,N_14338);
and U18327 (N_18327,N_13629,N_12187);
nand U18328 (N_18328,N_12166,N_15770);
or U18329 (N_18329,N_12555,N_12916);
nor U18330 (N_18330,N_15052,N_13946);
or U18331 (N_18331,N_13078,N_13156);
and U18332 (N_18332,N_14246,N_12607);
nand U18333 (N_18333,N_15614,N_13975);
nor U18334 (N_18334,N_14330,N_13479);
and U18335 (N_18335,N_15215,N_15074);
nor U18336 (N_18336,N_14264,N_14772);
or U18337 (N_18337,N_12113,N_15168);
and U18338 (N_18338,N_12785,N_15552);
and U18339 (N_18339,N_12321,N_14055);
and U18340 (N_18340,N_15664,N_14175);
or U18341 (N_18341,N_12841,N_15787);
or U18342 (N_18342,N_14141,N_12666);
nand U18343 (N_18343,N_13997,N_12458);
or U18344 (N_18344,N_12041,N_15717);
nor U18345 (N_18345,N_13468,N_15962);
and U18346 (N_18346,N_15817,N_14290);
or U18347 (N_18347,N_14195,N_14850);
nand U18348 (N_18348,N_12530,N_13937);
and U18349 (N_18349,N_12812,N_15841);
nor U18350 (N_18350,N_12119,N_14237);
or U18351 (N_18351,N_14988,N_15646);
or U18352 (N_18352,N_12302,N_15115);
or U18353 (N_18353,N_15160,N_12188);
and U18354 (N_18354,N_14472,N_15614);
nor U18355 (N_18355,N_13700,N_12058);
nor U18356 (N_18356,N_13875,N_13656);
nor U18357 (N_18357,N_14400,N_12475);
and U18358 (N_18358,N_12211,N_15717);
or U18359 (N_18359,N_13576,N_12966);
and U18360 (N_18360,N_13837,N_14544);
nand U18361 (N_18361,N_15641,N_14677);
or U18362 (N_18362,N_13807,N_14653);
nor U18363 (N_18363,N_14181,N_15620);
and U18364 (N_18364,N_13481,N_13682);
nand U18365 (N_18365,N_14162,N_14699);
and U18366 (N_18366,N_13127,N_13176);
nor U18367 (N_18367,N_13379,N_13266);
nand U18368 (N_18368,N_15983,N_15871);
nor U18369 (N_18369,N_14273,N_14665);
nor U18370 (N_18370,N_15819,N_15612);
nand U18371 (N_18371,N_13376,N_12364);
and U18372 (N_18372,N_13568,N_13501);
nor U18373 (N_18373,N_12946,N_15192);
and U18374 (N_18374,N_14398,N_15352);
or U18375 (N_18375,N_12302,N_15521);
xnor U18376 (N_18376,N_12900,N_15983);
nor U18377 (N_18377,N_13834,N_14743);
nand U18378 (N_18378,N_13776,N_13541);
nand U18379 (N_18379,N_15370,N_14991);
nand U18380 (N_18380,N_12535,N_14572);
nand U18381 (N_18381,N_12273,N_12190);
and U18382 (N_18382,N_12891,N_14047);
or U18383 (N_18383,N_14447,N_14707);
or U18384 (N_18384,N_12101,N_12525);
nand U18385 (N_18385,N_13413,N_13019);
nor U18386 (N_18386,N_12894,N_12568);
nor U18387 (N_18387,N_12162,N_14365);
nand U18388 (N_18388,N_12588,N_14126);
and U18389 (N_18389,N_12049,N_14868);
or U18390 (N_18390,N_15781,N_12464);
and U18391 (N_18391,N_14287,N_15684);
nor U18392 (N_18392,N_14875,N_13316);
and U18393 (N_18393,N_12488,N_15445);
or U18394 (N_18394,N_14067,N_14728);
and U18395 (N_18395,N_13222,N_13841);
or U18396 (N_18396,N_15210,N_13554);
nand U18397 (N_18397,N_15344,N_12757);
nand U18398 (N_18398,N_14538,N_15035);
nor U18399 (N_18399,N_15849,N_15709);
nand U18400 (N_18400,N_13976,N_14420);
xor U18401 (N_18401,N_13811,N_13048);
nor U18402 (N_18402,N_14391,N_14953);
nand U18403 (N_18403,N_15558,N_14456);
and U18404 (N_18404,N_14053,N_13838);
nand U18405 (N_18405,N_15659,N_13435);
or U18406 (N_18406,N_13284,N_14564);
or U18407 (N_18407,N_14292,N_13290);
nand U18408 (N_18408,N_13218,N_13571);
and U18409 (N_18409,N_13367,N_13942);
nand U18410 (N_18410,N_12254,N_15371);
or U18411 (N_18411,N_13936,N_15927);
or U18412 (N_18412,N_15606,N_12189);
nor U18413 (N_18413,N_12653,N_13780);
nor U18414 (N_18414,N_12609,N_13346);
or U18415 (N_18415,N_12782,N_13879);
or U18416 (N_18416,N_12626,N_14661);
and U18417 (N_18417,N_12310,N_12918);
or U18418 (N_18418,N_12666,N_13862);
nand U18419 (N_18419,N_12197,N_14972);
nand U18420 (N_18420,N_14238,N_13318);
or U18421 (N_18421,N_12402,N_12907);
nor U18422 (N_18422,N_14581,N_12001);
nor U18423 (N_18423,N_12818,N_14880);
and U18424 (N_18424,N_15194,N_12252);
and U18425 (N_18425,N_14987,N_15612);
nand U18426 (N_18426,N_15107,N_14395);
nand U18427 (N_18427,N_13808,N_13106);
and U18428 (N_18428,N_14192,N_14793);
and U18429 (N_18429,N_12964,N_14186);
nand U18430 (N_18430,N_13085,N_13301);
nor U18431 (N_18431,N_15230,N_12380);
nand U18432 (N_18432,N_15159,N_12572);
or U18433 (N_18433,N_14587,N_15021);
nor U18434 (N_18434,N_12495,N_15921);
or U18435 (N_18435,N_15740,N_13669);
nand U18436 (N_18436,N_14334,N_13548);
nor U18437 (N_18437,N_13201,N_14306);
and U18438 (N_18438,N_14523,N_14518);
nand U18439 (N_18439,N_12923,N_12927);
nor U18440 (N_18440,N_14905,N_15548);
or U18441 (N_18441,N_14822,N_15120);
or U18442 (N_18442,N_15568,N_14010);
nor U18443 (N_18443,N_13179,N_14696);
and U18444 (N_18444,N_15297,N_13496);
and U18445 (N_18445,N_13275,N_15850);
nand U18446 (N_18446,N_12750,N_14281);
nand U18447 (N_18447,N_12250,N_14431);
and U18448 (N_18448,N_12459,N_13366);
nand U18449 (N_18449,N_15333,N_13015);
nor U18450 (N_18450,N_15478,N_15222);
nand U18451 (N_18451,N_13913,N_14314);
or U18452 (N_18452,N_14805,N_12563);
or U18453 (N_18453,N_13145,N_15122);
nand U18454 (N_18454,N_12028,N_12497);
or U18455 (N_18455,N_14844,N_13856);
and U18456 (N_18456,N_13821,N_12758);
or U18457 (N_18457,N_15986,N_15082);
nor U18458 (N_18458,N_12006,N_14482);
or U18459 (N_18459,N_12065,N_14258);
nand U18460 (N_18460,N_13709,N_12119);
nand U18461 (N_18461,N_15415,N_14914);
nand U18462 (N_18462,N_12706,N_12074);
and U18463 (N_18463,N_12195,N_13935);
nand U18464 (N_18464,N_12633,N_12204);
nand U18465 (N_18465,N_15957,N_12619);
or U18466 (N_18466,N_14569,N_15581);
nor U18467 (N_18467,N_12385,N_12745);
and U18468 (N_18468,N_12648,N_13477);
nand U18469 (N_18469,N_13793,N_12188);
or U18470 (N_18470,N_14470,N_15627);
nand U18471 (N_18471,N_13191,N_12463);
or U18472 (N_18472,N_15978,N_15228);
and U18473 (N_18473,N_15392,N_13630);
nor U18474 (N_18474,N_12603,N_12189);
and U18475 (N_18475,N_14547,N_15354);
and U18476 (N_18476,N_15425,N_13592);
and U18477 (N_18477,N_14693,N_14515);
or U18478 (N_18478,N_15259,N_14614);
and U18479 (N_18479,N_14580,N_14210);
nand U18480 (N_18480,N_15612,N_13504);
nor U18481 (N_18481,N_12780,N_15634);
nand U18482 (N_18482,N_12713,N_15784);
nor U18483 (N_18483,N_15632,N_12408);
nand U18484 (N_18484,N_13667,N_12445);
and U18485 (N_18485,N_14333,N_13036);
or U18486 (N_18486,N_12667,N_14849);
or U18487 (N_18487,N_14677,N_13152);
or U18488 (N_18488,N_15374,N_14862);
nor U18489 (N_18489,N_14148,N_14702);
nand U18490 (N_18490,N_12222,N_15027);
nand U18491 (N_18491,N_13732,N_14108);
nand U18492 (N_18492,N_15600,N_12357);
or U18493 (N_18493,N_14436,N_14627);
or U18494 (N_18494,N_14968,N_14964);
and U18495 (N_18495,N_15724,N_13906);
and U18496 (N_18496,N_12931,N_14899);
nand U18497 (N_18497,N_14110,N_13065);
and U18498 (N_18498,N_15785,N_14642);
and U18499 (N_18499,N_13895,N_14566);
nor U18500 (N_18500,N_13557,N_14672);
and U18501 (N_18501,N_15763,N_12932);
and U18502 (N_18502,N_14568,N_14166);
or U18503 (N_18503,N_13569,N_15278);
nand U18504 (N_18504,N_13472,N_15663);
and U18505 (N_18505,N_15373,N_15692);
nand U18506 (N_18506,N_12310,N_13314);
nand U18507 (N_18507,N_15747,N_14457);
nor U18508 (N_18508,N_13303,N_12182);
and U18509 (N_18509,N_13369,N_13810);
nand U18510 (N_18510,N_14355,N_12016);
and U18511 (N_18511,N_13345,N_12409);
nand U18512 (N_18512,N_15452,N_15507);
nor U18513 (N_18513,N_12844,N_13311);
and U18514 (N_18514,N_15779,N_12387);
nor U18515 (N_18515,N_15604,N_12063);
and U18516 (N_18516,N_12682,N_12337);
or U18517 (N_18517,N_15577,N_13478);
nand U18518 (N_18518,N_14868,N_12624);
nand U18519 (N_18519,N_14290,N_14040);
nor U18520 (N_18520,N_14683,N_13691);
nor U18521 (N_18521,N_13650,N_13070);
or U18522 (N_18522,N_14536,N_13387);
and U18523 (N_18523,N_13069,N_12332);
or U18524 (N_18524,N_12371,N_15591);
or U18525 (N_18525,N_14653,N_12054);
nor U18526 (N_18526,N_15079,N_14158);
or U18527 (N_18527,N_13502,N_14340);
or U18528 (N_18528,N_12176,N_12471);
and U18529 (N_18529,N_14959,N_15174);
and U18530 (N_18530,N_15264,N_14841);
nand U18531 (N_18531,N_12014,N_15176);
nand U18532 (N_18532,N_14908,N_15109);
or U18533 (N_18533,N_12831,N_12072);
nor U18534 (N_18534,N_15062,N_15419);
nor U18535 (N_18535,N_13169,N_13209);
and U18536 (N_18536,N_12240,N_14344);
or U18537 (N_18537,N_13742,N_13284);
xor U18538 (N_18538,N_13145,N_15999);
or U18539 (N_18539,N_13748,N_15651);
nor U18540 (N_18540,N_15583,N_15410);
or U18541 (N_18541,N_15445,N_13274);
and U18542 (N_18542,N_15596,N_13365);
nand U18543 (N_18543,N_14731,N_13876);
nand U18544 (N_18544,N_14240,N_12278);
and U18545 (N_18545,N_12680,N_14372);
nand U18546 (N_18546,N_12274,N_15901);
nor U18547 (N_18547,N_12362,N_15963);
nand U18548 (N_18548,N_13017,N_13042);
nand U18549 (N_18549,N_15016,N_12620);
and U18550 (N_18550,N_12767,N_12096);
nand U18551 (N_18551,N_13437,N_12006);
nand U18552 (N_18552,N_14852,N_14017);
nand U18553 (N_18553,N_12119,N_15088);
or U18554 (N_18554,N_15901,N_12706);
nor U18555 (N_18555,N_14178,N_14762);
nand U18556 (N_18556,N_13390,N_12617);
nor U18557 (N_18557,N_14519,N_14148);
nor U18558 (N_18558,N_13156,N_12880);
and U18559 (N_18559,N_13470,N_15007);
and U18560 (N_18560,N_12604,N_13187);
or U18561 (N_18561,N_15367,N_12537);
nor U18562 (N_18562,N_13750,N_15093);
and U18563 (N_18563,N_13923,N_15059);
nand U18564 (N_18564,N_15997,N_14571);
nor U18565 (N_18565,N_15455,N_15953);
nor U18566 (N_18566,N_13067,N_13700);
and U18567 (N_18567,N_12008,N_15246);
nand U18568 (N_18568,N_13154,N_12281);
nor U18569 (N_18569,N_12712,N_14527);
nand U18570 (N_18570,N_15028,N_13592);
nand U18571 (N_18571,N_13194,N_14331);
nand U18572 (N_18572,N_14873,N_12961);
nor U18573 (N_18573,N_13282,N_12996);
and U18574 (N_18574,N_14155,N_13141);
and U18575 (N_18575,N_13366,N_15539);
nor U18576 (N_18576,N_15897,N_12509);
and U18577 (N_18577,N_15506,N_13930);
nor U18578 (N_18578,N_14922,N_12344);
or U18579 (N_18579,N_14439,N_14139);
nor U18580 (N_18580,N_14788,N_13563);
nor U18581 (N_18581,N_12708,N_15426);
or U18582 (N_18582,N_14635,N_14238);
nor U18583 (N_18583,N_13828,N_14129);
or U18584 (N_18584,N_12510,N_14231);
nor U18585 (N_18585,N_13039,N_13625);
or U18586 (N_18586,N_14472,N_12151);
nand U18587 (N_18587,N_15583,N_12811);
and U18588 (N_18588,N_12388,N_12967);
and U18589 (N_18589,N_15237,N_13732);
nand U18590 (N_18590,N_12096,N_14157);
nor U18591 (N_18591,N_13679,N_12753);
and U18592 (N_18592,N_12515,N_15278);
nor U18593 (N_18593,N_12788,N_14812);
nand U18594 (N_18594,N_14164,N_13109);
or U18595 (N_18595,N_14217,N_13185);
nand U18596 (N_18596,N_15733,N_12994);
nor U18597 (N_18597,N_13527,N_15173);
nand U18598 (N_18598,N_14287,N_15028);
and U18599 (N_18599,N_14009,N_13474);
nor U18600 (N_18600,N_12829,N_15649);
nand U18601 (N_18601,N_13536,N_15358);
nand U18602 (N_18602,N_13703,N_13278);
and U18603 (N_18603,N_12926,N_15793);
nor U18604 (N_18604,N_14886,N_14687);
nor U18605 (N_18605,N_14385,N_14978);
or U18606 (N_18606,N_15305,N_14271);
nor U18607 (N_18607,N_12241,N_14827);
or U18608 (N_18608,N_14881,N_14335);
nor U18609 (N_18609,N_12618,N_12465);
or U18610 (N_18610,N_15773,N_13309);
or U18611 (N_18611,N_13009,N_14239);
and U18612 (N_18612,N_15808,N_12052);
nand U18613 (N_18613,N_13307,N_12571);
and U18614 (N_18614,N_13761,N_13645);
or U18615 (N_18615,N_13277,N_13045);
or U18616 (N_18616,N_14155,N_12393);
nor U18617 (N_18617,N_13561,N_12214);
nor U18618 (N_18618,N_12559,N_12801);
and U18619 (N_18619,N_12271,N_12111);
nand U18620 (N_18620,N_12998,N_12218);
nor U18621 (N_18621,N_13256,N_14203);
nor U18622 (N_18622,N_12495,N_15967);
and U18623 (N_18623,N_13030,N_14996);
nor U18624 (N_18624,N_13673,N_12956);
nand U18625 (N_18625,N_14397,N_12447);
nand U18626 (N_18626,N_15051,N_15857);
nor U18627 (N_18627,N_14628,N_12861);
or U18628 (N_18628,N_13295,N_15425);
or U18629 (N_18629,N_14519,N_12415);
nor U18630 (N_18630,N_12575,N_15905);
or U18631 (N_18631,N_13192,N_12384);
nand U18632 (N_18632,N_15877,N_15532);
nand U18633 (N_18633,N_14591,N_13643);
or U18634 (N_18634,N_13626,N_12690);
and U18635 (N_18635,N_12941,N_14527);
and U18636 (N_18636,N_13984,N_14742);
nand U18637 (N_18637,N_15894,N_13801);
or U18638 (N_18638,N_14056,N_14664);
nor U18639 (N_18639,N_15145,N_13617);
nand U18640 (N_18640,N_15216,N_12131);
nand U18641 (N_18641,N_13531,N_15139);
nand U18642 (N_18642,N_12877,N_14468);
nand U18643 (N_18643,N_13131,N_12939);
nand U18644 (N_18644,N_14652,N_12248);
or U18645 (N_18645,N_13676,N_15095);
and U18646 (N_18646,N_13122,N_13055);
nand U18647 (N_18647,N_14897,N_14434);
nor U18648 (N_18648,N_13790,N_15489);
or U18649 (N_18649,N_13292,N_15940);
and U18650 (N_18650,N_12032,N_14479);
nand U18651 (N_18651,N_15262,N_13536);
or U18652 (N_18652,N_13976,N_14625);
nor U18653 (N_18653,N_15703,N_15692);
and U18654 (N_18654,N_12941,N_14059);
nand U18655 (N_18655,N_13383,N_15700);
and U18656 (N_18656,N_13098,N_15755);
nor U18657 (N_18657,N_15418,N_15681);
or U18658 (N_18658,N_13717,N_15740);
nand U18659 (N_18659,N_12476,N_12201);
nor U18660 (N_18660,N_13258,N_14206);
nand U18661 (N_18661,N_13488,N_14132);
or U18662 (N_18662,N_14690,N_12047);
or U18663 (N_18663,N_15816,N_12146);
nor U18664 (N_18664,N_12080,N_15067);
and U18665 (N_18665,N_14111,N_13870);
nor U18666 (N_18666,N_13688,N_12566);
nand U18667 (N_18667,N_15946,N_14817);
nor U18668 (N_18668,N_13019,N_12523);
nand U18669 (N_18669,N_15577,N_13812);
nand U18670 (N_18670,N_15145,N_13998);
nor U18671 (N_18671,N_14017,N_15197);
nor U18672 (N_18672,N_14484,N_14137);
or U18673 (N_18673,N_14850,N_13286);
or U18674 (N_18674,N_13189,N_13818);
or U18675 (N_18675,N_13678,N_12661);
nor U18676 (N_18676,N_14789,N_14396);
and U18677 (N_18677,N_15234,N_15913);
and U18678 (N_18678,N_13141,N_15691);
nor U18679 (N_18679,N_14864,N_13789);
or U18680 (N_18680,N_15883,N_12368);
nor U18681 (N_18681,N_15876,N_12400);
nor U18682 (N_18682,N_12816,N_13182);
or U18683 (N_18683,N_15499,N_15684);
nor U18684 (N_18684,N_14251,N_13894);
nor U18685 (N_18685,N_15769,N_14548);
nand U18686 (N_18686,N_12986,N_14333);
and U18687 (N_18687,N_14663,N_13114);
and U18688 (N_18688,N_12572,N_15757);
nand U18689 (N_18689,N_15112,N_13965);
nand U18690 (N_18690,N_12193,N_14957);
and U18691 (N_18691,N_15321,N_15221);
or U18692 (N_18692,N_13016,N_13304);
and U18693 (N_18693,N_12248,N_15775);
nor U18694 (N_18694,N_12111,N_12719);
nor U18695 (N_18695,N_15353,N_12959);
or U18696 (N_18696,N_12565,N_14062);
or U18697 (N_18697,N_12861,N_14633);
nand U18698 (N_18698,N_13818,N_13002);
or U18699 (N_18699,N_12935,N_14125);
nand U18700 (N_18700,N_13444,N_13534);
nand U18701 (N_18701,N_13050,N_12593);
or U18702 (N_18702,N_15537,N_12477);
and U18703 (N_18703,N_15984,N_13767);
and U18704 (N_18704,N_12414,N_13373);
nor U18705 (N_18705,N_13735,N_14511);
and U18706 (N_18706,N_14169,N_12447);
nand U18707 (N_18707,N_13688,N_14476);
or U18708 (N_18708,N_15069,N_15180);
or U18709 (N_18709,N_13595,N_13953);
nor U18710 (N_18710,N_15908,N_12595);
nor U18711 (N_18711,N_15709,N_12158);
nand U18712 (N_18712,N_12732,N_15626);
or U18713 (N_18713,N_12112,N_13833);
or U18714 (N_18714,N_12082,N_13499);
nor U18715 (N_18715,N_14934,N_15689);
or U18716 (N_18716,N_13232,N_13545);
and U18717 (N_18717,N_13626,N_13632);
and U18718 (N_18718,N_13467,N_13268);
nor U18719 (N_18719,N_14740,N_12932);
or U18720 (N_18720,N_15964,N_15853);
nand U18721 (N_18721,N_14023,N_15217);
nor U18722 (N_18722,N_13961,N_15026);
nor U18723 (N_18723,N_12950,N_14056);
and U18724 (N_18724,N_14087,N_12723);
or U18725 (N_18725,N_15596,N_12352);
nand U18726 (N_18726,N_13902,N_12139);
xor U18727 (N_18727,N_14984,N_13562);
nand U18728 (N_18728,N_12286,N_15542);
nand U18729 (N_18729,N_13751,N_12890);
or U18730 (N_18730,N_13149,N_13257);
and U18731 (N_18731,N_14211,N_14127);
and U18732 (N_18732,N_14600,N_15360);
nand U18733 (N_18733,N_15183,N_14556);
or U18734 (N_18734,N_13948,N_12668);
nand U18735 (N_18735,N_13229,N_15022);
nor U18736 (N_18736,N_12335,N_14581);
nand U18737 (N_18737,N_12766,N_15947);
nand U18738 (N_18738,N_13980,N_15772);
and U18739 (N_18739,N_15196,N_13688);
or U18740 (N_18740,N_15307,N_12803);
nand U18741 (N_18741,N_13791,N_14258);
nor U18742 (N_18742,N_13256,N_14869);
or U18743 (N_18743,N_15791,N_12688);
and U18744 (N_18744,N_13034,N_12625);
nand U18745 (N_18745,N_12172,N_14692);
nand U18746 (N_18746,N_13925,N_13763);
nand U18747 (N_18747,N_12354,N_12932);
and U18748 (N_18748,N_12395,N_13604);
or U18749 (N_18749,N_15067,N_13913);
or U18750 (N_18750,N_14867,N_15150);
and U18751 (N_18751,N_14163,N_13356);
or U18752 (N_18752,N_12267,N_13382);
xnor U18753 (N_18753,N_12009,N_12523);
or U18754 (N_18754,N_13414,N_15164);
nor U18755 (N_18755,N_13649,N_15261);
or U18756 (N_18756,N_14134,N_14839);
nor U18757 (N_18757,N_12080,N_14627);
or U18758 (N_18758,N_13122,N_14585);
or U18759 (N_18759,N_13522,N_14638);
or U18760 (N_18760,N_13193,N_14631);
nor U18761 (N_18761,N_13313,N_12453);
or U18762 (N_18762,N_14086,N_14856);
nor U18763 (N_18763,N_13987,N_12350);
xor U18764 (N_18764,N_13165,N_12131);
or U18765 (N_18765,N_13774,N_13326);
and U18766 (N_18766,N_12932,N_14902);
nand U18767 (N_18767,N_14030,N_15772);
and U18768 (N_18768,N_13076,N_12367);
and U18769 (N_18769,N_12878,N_12768);
nor U18770 (N_18770,N_14350,N_15775);
nor U18771 (N_18771,N_13561,N_12330);
or U18772 (N_18772,N_15303,N_13506);
and U18773 (N_18773,N_12033,N_13627);
nor U18774 (N_18774,N_14767,N_13581);
nand U18775 (N_18775,N_12122,N_13297);
and U18776 (N_18776,N_12630,N_13990);
and U18777 (N_18777,N_12189,N_15739);
or U18778 (N_18778,N_13713,N_12439);
nand U18779 (N_18779,N_15469,N_14032);
or U18780 (N_18780,N_14065,N_15156);
nor U18781 (N_18781,N_13472,N_12102);
nor U18782 (N_18782,N_14132,N_15203);
or U18783 (N_18783,N_13636,N_13030);
nor U18784 (N_18784,N_14375,N_14106);
and U18785 (N_18785,N_14677,N_14570);
and U18786 (N_18786,N_12724,N_15065);
nand U18787 (N_18787,N_14238,N_15637);
and U18788 (N_18788,N_15667,N_14749);
nor U18789 (N_18789,N_13644,N_12555);
nand U18790 (N_18790,N_12486,N_13641);
or U18791 (N_18791,N_14884,N_15852);
nand U18792 (N_18792,N_14925,N_12814);
nand U18793 (N_18793,N_13028,N_12651);
and U18794 (N_18794,N_12227,N_14286);
and U18795 (N_18795,N_15686,N_14127);
and U18796 (N_18796,N_15980,N_15055);
nand U18797 (N_18797,N_13976,N_15231);
and U18798 (N_18798,N_15241,N_14878);
or U18799 (N_18799,N_12665,N_14881);
and U18800 (N_18800,N_14663,N_15783);
nand U18801 (N_18801,N_13451,N_12860);
nor U18802 (N_18802,N_15879,N_12411);
or U18803 (N_18803,N_14028,N_13203);
nor U18804 (N_18804,N_12818,N_13117);
nor U18805 (N_18805,N_12084,N_15473);
and U18806 (N_18806,N_14821,N_14897);
nand U18807 (N_18807,N_14729,N_15265);
and U18808 (N_18808,N_13620,N_13504);
or U18809 (N_18809,N_15769,N_13021);
nand U18810 (N_18810,N_12072,N_12377);
and U18811 (N_18811,N_14768,N_12369);
nand U18812 (N_18812,N_12990,N_12897);
nand U18813 (N_18813,N_13411,N_15227);
nor U18814 (N_18814,N_13072,N_12430);
nor U18815 (N_18815,N_15954,N_15010);
or U18816 (N_18816,N_12437,N_15397);
nand U18817 (N_18817,N_13297,N_15290);
nor U18818 (N_18818,N_15295,N_15422);
nand U18819 (N_18819,N_13024,N_12491);
or U18820 (N_18820,N_14947,N_12236);
nor U18821 (N_18821,N_13388,N_15811);
nor U18822 (N_18822,N_13504,N_15843);
nand U18823 (N_18823,N_12296,N_13307);
nor U18824 (N_18824,N_13152,N_12925);
nand U18825 (N_18825,N_13107,N_15571);
or U18826 (N_18826,N_13890,N_13053);
nand U18827 (N_18827,N_15255,N_14341);
and U18828 (N_18828,N_14978,N_13786);
nand U18829 (N_18829,N_12321,N_12649);
or U18830 (N_18830,N_14336,N_13768);
and U18831 (N_18831,N_14420,N_15475);
and U18832 (N_18832,N_14576,N_12545);
nand U18833 (N_18833,N_12287,N_13402);
nand U18834 (N_18834,N_13836,N_15784);
and U18835 (N_18835,N_12967,N_14891);
nor U18836 (N_18836,N_13757,N_13113);
or U18837 (N_18837,N_13130,N_14749);
nand U18838 (N_18838,N_15657,N_14156);
nand U18839 (N_18839,N_13549,N_15127);
and U18840 (N_18840,N_14401,N_13893);
nand U18841 (N_18841,N_12951,N_12740);
nor U18842 (N_18842,N_14134,N_13540);
nand U18843 (N_18843,N_13841,N_13268);
or U18844 (N_18844,N_15265,N_14645);
nand U18845 (N_18845,N_12594,N_12886);
or U18846 (N_18846,N_14906,N_14289);
nand U18847 (N_18847,N_13794,N_13335);
nor U18848 (N_18848,N_14948,N_13528);
or U18849 (N_18849,N_14742,N_12666);
and U18850 (N_18850,N_15611,N_13135);
nor U18851 (N_18851,N_13990,N_12925);
nand U18852 (N_18852,N_13995,N_13882);
and U18853 (N_18853,N_14212,N_13571);
or U18854 (N_18854,N_14387,N_13762);
nand U18855 (N_18855,N_14240,N_12337);
and U18856 (N_18856,N_12188,N_13554);
or U18857 (N_18857,N_14049,N_14762);
or U18858 (N_18858,N_14253,N_13783);
and U18859 (N_18859,N_15659,N_14988);
and U18860 (N_18860,N_13038,N_13428);
and U18861 (N_18861,N_15848,N_13875);
nor U18862 (N_18862,N_13172,N_12786);
and U18863 (N_18863,N_14154,N_14163);
xnor U18864 (N_18864,N_13958,N_13565);
or U18865 (N_18865,N_13780,N_13938);
and U18866 (N_18866,N_12157,N_13918);
or U18867 (N_18867,N_15712,N_13349);
nor U18868 (N_18868,N_12363,N_14731);
or U18869 (N_18869,N_14737,N_15274);
and U18870 (N_18870,N_15114,N_14912);
nor U18871 (N_18871,N_15526,N_12276);
and U18872 (N_18872,N_12891,N_14634);
nor U18873 (N_18873,N_14966,N_14417);
nor U18874 (N_18874,N_14771,N_13707);
nor U18875 (N_18875,N_12501,N_14579);
xnor U18876 (N_18876,N_12357,N_13310);
nand U18877 (N_18877,N_14477,N_13000);
nor U18878 (N_18878,N_15730,N_13034);
or U18879 (N_18879,N_15981,N_12656);
or U18880 (N_18880,N_13847,N_13178);
and U18881 (N_18881,N_13345,N_12398);
or U18882 (N_18882,N_15996,N_14200);
and U18883 (N_18883,N_14015,N_14242);
or U18884 (N_18884,N_14668,N_15776);
and U18885 (N_18885,N_13634,N_14609);
or U18886 (N_18886,N_15271,N_15678);
nand U18887 (N_18887,N_14078,N_15304);
nor U18888 (N_18888,N_13441,N_12846);
or U18889 (N_18889,N_12170,N_12620);
nor U18890 (N_18890,N_12935,N_12051);
and U18891 (N_18891,N_13077,N_12690);
nor U18892 (N_18892,N_15925,N_12373);
or U18893 (N_18893,N_13860,N_14827);
nor U18894 (N_18894,N_14505,N_13522);
and U18895 (N_18895,N_15654,N_15101);
nand U18896 (N_18896,N_12754,N_13229);
xor U18897 (N_18897,N_14903,N_15477);
and U18898 (N_18898,N_14732,N_14883);
and U18899 (N_18899,N_13684,N_15331);
nor U18900 (N_18900,N_12382,N_15322);
nand U18901 (N_18901,N_14840,N_14604);
nand U18902 (N_18902,N_14719,N_12358);
nand U18903 (N_18903,N_12462,N_13518);
xnor U18904 (N_18904,N_15953,N_14717);
nand U18905 (N_18905,N_14080,N_12895);
or U18906 (N_18906,N_15702,N_15517);
nor U18907 (N_18907,N_13282,N_13920);
nand U18908 (N_18908,N_14646,N_13108);
or U18909 (N_18909,N_13661,N_15773);
and U18910 (N_18910,N_15450,N_15730);
or U18911 (N_18911,N_13838,N_14668);
or U18912 (N_18912,N_13622,N_12025);
nor U18913 (N_18913,N_13561,N_15620);
or U18914 (N_18914,N_14370,N_14799);
or U18915 (N_18915,N_13074,N_12964);
nor U18916 (N_18916,N_15319,N_14467);
and U18917 (N_18917,N_13774,N_12487);
or U18918 (N_18918,N_12542,N_14012);
and U18919 (N_18919,N_12659,N_13084);
nand U18920 (N_18920,N_12004,N_13556);
or U18921 (N_18921,N_12855,N_14131);
nand U18922 (N_18922,N_14993,N_13413);
or U18923 (N_18923,N_13357,N_13338);
nand U18924 (N_18924,N_15832,N_14386);
nor U18925 (N_18925,N_14856,N_14305);
and U18926 (N_18926,N_12410,N_14305);
or U18927 (N_18927,N_14564,N_14598);
nand U18928 (N_18928,N_15731,N_14614);
nand U18929 (N_18929,N_14459,N_12603);
nand U18930 (N_18930,N_13322,N_12011);
nand U18931 (N_18931,N_13574,N_13564);
nor U18932 (N_18932,N_14972,N_14997);
nor U18933 (N_18933,N_13878,N_15571);
nand U18934 (N_18934,N_13365,N_13342);
nand U18935 (N_18935,N_13354,N_14986);
or U18936 (N_18936,N_12017,N_14960);
nor U18937 (N_18937,N_12761,N_14109);
or U18938 (N_18938,N_13259,N_15398);
nand U18939 (N_18939,N_15213,N_14659);
nand U18940 (N_18940,N_15570,N_13209);
or U18941 (N_18941,N_15033,N_13122);
nand U18942 (N_18942,N_15589,N_15571);
or U18943 (N_18943,N_14362,N_14455);
and U18944 (N_18944,N_15294,N_13828);
or U18945 (N_18945,N_14585,N_13544);
nand U18946 (N_18946,N_15782,N_12978);
nor U18947 (N_18947,N_15652,N_14727);
nor U18948 (N_18948,N_12210,N_13352);
nor U18949 (N_18949,N_12102,N_13947);
nor U18950 (N_18950,N_13301,N_12358);
nor U18951 (N_18951,N_13119,N_12185);
and U18952 (N_18952,N_15793,N_14377);
and U18953 (N_18953,N_15433,N_12992);
nor U18954 (N_18954,N_13252,N_14086);
or U18955 (N_18955,N_15375,N_13467);
or U18956 (N_18956,N_14329,N_13897);
nand U18957 (N_18957,N_15134,N_15446);
and U18958 (N_18958,N_15552,N_14738);
and U18959 (N_18959,N_14029,N_14284);
nor U18960 (N_18960,N_15193,N_12603);
nand U18961 (N_18961,N_13278,N_13216);
nor U18962 (N_18962,N_13886,N_15880);
nor U18963 (N_18963,N_12220,N_14567);
or U18964 (N_18964,N_14045,N_12510);
nor U18965 (N_18965,N_13968,N_13638);
or U18966 (N_18966,N_15050,N_13189);
or U18967 (N_18967,N_13843,N_13879);
nand U18968 (N_18968,N_15239,N_13203);
and U18969 (N_18969,N_15050,N_14197);
nand U18970 (N_18970,N_15216,N_13195);
and U18971 (N_18971,N_15109,N_12718);
or U18972 (N_18972,N_14281,N_12818);
nor U18973 (N_18973,N_12847,N_15381);
nor U18974 (N_18974,N_14070,N_13549);
nor U18975 (N_18975,N_13309,N_13844);
nand U18976 (N_18976,N_15785,N_15684);
nand U18977 (N_18977,N_13622,N_14469);
and U18978 (N_18978,N_15200,N_14574);
or U18979 (N_18979,N_15638,N_15068);
nand U18980 (N_18980,N_13605,N_14454);
and U18981 (N_18981,N_15991,N_12430);
and U18982 (N_18982,N_12530,N_12586);
nor U18983 (N_18983,N_12836,N_12968);
nor U18984 (N_18984,N_15076,N_15147);
or U18985 (N_18985,N_13387,N_12428);
or U18986 (N_18986,N_15337,N_14445);
and U18987 (N_18987,N_14903,N_15111);
and U18988 (N_18988,N_14657,N_14924);
nand U18989 (N_18989,N_14450,N_15344);
nand U18990 (N_18990,N_15640,N_12719);
and U18991 (N_18991,N_15997,N_14251);
or U18992 (N_18992,N_12786,N_14675);
nor U18993 (N_18993,N_15397,N_12924);
or U18994 (N_18994,N_14916,N_13333);
nor U18995 (N_18995,N_12473,N_14767);
or U18996 (N_18996,N_14311,N_13924);
or U18997 (N_18997,N_12631,N_13141);
nand U18998 (N_18998,N_15259,N_12977);
nand U18999 (N_18999,N_15077,N_12697);
and U19000 (N_19000,N_14499,N_15738);
and U19001 (N_19001,N_12939,N_13438);
nor U19002 (N_19002,N_12370,N_14203);
nand U19003 (N_19003,N_12356,N_12581);
nor U19004 (N_19004,N_12450,N_15330);
and U19005 (N_19005,N_12511,N_14672);
xor U19006 (N_19006,N_12934,N_14228);
nand U19007 (N_19007,N_12676,N_15123);
nor U19008 (N_19008,N_12628,N_14502);
and U19009 (N_19009,N_15522,N_12555);
and U19010 (N_19010,N_15664,N_15709);
nor U19011 (N_19011,N_15756,N_14384);
and U19012 (N_19012,N_14671,N_15463);
and U19013 (N_19013,N_12482,N_13626);
and U19014 (N_19014,N_14872,N_15109);
or U19015 (N_19015,N_13697,N_12123);
xnor U19016 (N_19016,N_14272,N_13522);
and U19017 (N_19017,N_13889,N_13563);
nand U19018 (N_19018,N_13702,N_12010);
or U19019 (N_19019,N_14748,N_13765);
or U19020 (N_19020,N_12672,N_14014);
and U19021 (N_19021,N_14506,N_14770);
nand U19022 (N_19022,N_15482,N_15552);
nand U19023 (N_19023,N_15013,N_13797);
nor U19024 (N_19024,N_12359,N_12271);
nor U19025 (N_19025,N_15996,N_15692);
and U19026 (N_19026,N_12035,N_15634);
or U19027 (N_19027,N_14452,N_14057);
and U19028 (N_19028,N_13479,N_13781);
and U19029 (N_19029,N_15222,N_12967);
nor U19030 (N_19030,N_14226,N_12692);
nor U19031 (N_19031,N_14727,N_12678);
nand U19032 (N_19032,N_14111,N_13449);
or U19033 (N_19033,N_14814,N_12077);
and U19034 (N_19034,N_14342,N_15768);
nor U19035 (N_19035,N_13009,N_13053);
or U19036 (N_19036,N_12404,N_12396);
or U19037 (N_19037,N_14984,N_14974);
and U19038 (N_19038,N_13042,N_12148);
nand U19039 (N_19039,N_13600,N_13834);
nor U19040 (N_19040,N_13167,N_14215);
nor U19041 (N_19041,N_13084,N_14933);
nor U19042 (N_19042,N_12438,N_12891);
or U19043 (N_19043,N_15628,N_15992);
nand U19044 (N_19044,N_15838,N_12304);
and U19045 (N_19045,N_14485,N_13049);
nor U19046 (N_19046,N_13079,N_12388);
or U19047 (N_19047,N_13799,N_12647);
nor U19048 (N_19048,N_15800,N_14717);
and U19049 (N_19049,N_13848,N_13366);
and U19050 (N_19050,N_14158,N_13277);
nor U19051 (N_19051,N_13550,N_14692);
nor U19052 (N_19052,N_15132,N_15993);
nand U19053 (N_19053,N_14959,N_14193);
nor U19054 (N_19054,N_13691,N_12155);
nor U19055 (N_19055,N_12410,N_12527);
nand U19056 (N_19056,N_15763,N_15454);
nand U19057 (N_19057,N_14342,N_14889);
or U19058 (N_19058,N_13861,N_14412);
and U19059 (N_19059,N_14909,N_15658);
and U19060 (N_19060,N_15444,N_13533);
nor U19061 (N_19061,N_12878,N_13787);
and U19062 (N_19062,N_15805,N_13346);
or U19063 (N_19063,N_13554,N_12829);
nor U19064 (N_19064,N_12088,N_14891);
and U19065 (N_19065,N_13195,N_12411);
nand U19066 (N_19066,N_12235,N_15823);
or U19067 (N_19067,N_13698,N_13756);
and U19068 (N_19068,N_14343,N_14079);
or U19069 (N_19069,N_15871,N_12863);
nand U19070 (N_19070,N_12768,N_13167);
or U19071 (N_19071,N_13135,N_13958);
nor U19072 (N_19072,N_12738,N_13994);
nor U19073 (N_19073,N_12142,N_15405);
or U19074 (N_19074,N_14357,N_13736);
and U19075 (N_19075,N_13830,N_12034);
nor U19076 (N_19076,N_14091,N_15596);
or U19077 (N_19077,N_14528,N_15727);
nor U19078 (N_19078,N_12234,N_14095);
nand U19079 (N_19079,N_15378,N_14391);
nor U19080 (N_19080,N_14733,N_12876);
and U19081 (N_19081,N_14126,N_14518);
and U19082 (N_19082,N_15562,N_14495);
and U19083 (N_19083,N_15879,N_15156);
nor U19084 (N_19084,N_15571,N_12813);
and U19085 (N_19085,N_12684,N_12031);
and U19086 (N_19086,N_12370,N_13619);
and U19087 (N_19087,N_15437,N_15027);
nand U19088 (N_19088,N_14920,N_14822);
and U19089 (N_19089,N_15545,N_14336);
nor U19090 (N_19090,N_12295,N_14311);
and U19091 (N_19091,N_14513,N_14179);
or U19092 (N_19092,N_12776,N_13869);
nand U19093 (N_19093,N_13347,N_13337);
nand U19094 (N_19094,N_14104,N_12352);
nor U19095 (N_19095,N_13583,N_15015);
or U19096 (N_19096,N_14519,N_13207);
and U19097 (N_19097,N_13174,N_14928);
nand U19098 (N_19098,N_13107,N_13595);
and U19099 (N_19099,N_15148,N_15113);
nor U19100 (N_19100,N_14520,N_13921);
nor U19101 (N_19101,N_15022,N_13362);
nor U19102 (N_19102,N_12489,N_14933);
nand U19103 (N_19103,N_15262,N_12660);
or U19104 (N_19104,N_15359,N_12295);
nor U19105 (N_19105,N_13077,N_12647);
and U19106 (N_19106,N_12258,N_14539);
or U19107 (N_19107,N_12618,N_15667);
or U19108 (N_19108,N_12238,N_14105);
and U19109 (N_19109,N_12550,N_14349);
nor U19110 (N_19110,N_12117,N_14095);
or U19111 (N_19111,N_14524,N_13453);
or U19112 (N_19112,N_15673,N_15364);
nor U19113 (N_19113,N_14773,N_12822);
or U19114 (N_19114,N_15278,N_14119);
and U19115 (N_19115,N_14251,N_13327);
nor U19116 (N_19116,N_15062,N_12714);
or U19117 (N_19117,N_13224,N_13965);
nand U19118 (N_19118,N_14022,N_12376);
nand U19119 (N_19119,N_12007,N_13568);
xnor U19120 (N_19120,N_15845,N_14391);
or U19121 (N_19121,N_15611,N_14947);
nand U19122 (N_19122,N_13187,N_15690);
and U19123 (N_19123,N_14149,N_15294);
or U19124 (N_19124,N_14932,N_12134);
or U19125 (N_19125,N_12967,N_13085);
nand U19126 (N_19126,N_12864,N_15857);
or U19127 (N_19127,N_15033,N_13571);
and U19128 (N_19128,N_15733,N_14423);
nand U19129 (N_19129,N_15859,N_13692);
and U19130 (N_19130,N_12211,N_12954);
nor U19131 (N_19131,N_15557,N_13889);
and U19132 (N_19132,N_15397,N_14430);
and U19133 (N_19133,N_13134,N_15874);
nor U19134 (N_19134,N_13125,N_14867);
nor U19135 (N_19135,N_14603,N_13886);
or U19136 (N_19136,N_14444,N_14854);
or U19137 (N_19137,N_13482,N_14261);
nor U19138 (N_19138,N_12662,N_14152);
nand U19139 (N_19139,N_15942,N_15763);
nand U19140 (N_19140,N_15821,N_15754);
nor U19141 (N_19141,N_13573,N_14211);
and U19142 (N_19142,N_13911,N_13389);
or U19143 (N_19143,N_13919,N_13982);
nor U19144 (N_19144,N_14301,N_14486);
and U19145 (N_19145,N_15220,N_15939);
nand U19146 (N_19146,N_12088,N_14304);
or U19147 (N_19147,N_13883,N_14735);
nand U19148 (N_19148,N_14650,N_14691);
nor U19149 (N_19149,N_15594,N_13005);
nor U19150 (N_19150,N_13783,N_14691);
and U19151 (N_19151,N_14930,N_12695);
nor U19152 (N_19152,N_14527,N_13427);
nor U19153 (N_19153,N_14408,N_12369);
nor U19154 (N_19154,N_14000,N_13507);
nor U19155 (N_19155,N_14338,N_12949);
or U19156 (N_19156,N_15009,N_15205);
or U19157 (N_19157,N_13107,N_15926);
or U19158 (N_19158,N_14835,N_13705);
nor U19159 (N_19159,N_15576,N_13859);
nand U19160 (N_19160,N_15232,N_12325);
nand U19161 (N_19161,N_15919,N_13062);
and U19162 (N_19162,N_15297,N_14049);
nand U19163 (N_19163,N_14904,N_15996);
or U19164 (N_19164,N_15320,N_12606);
or U19165 (N_19165,N_14487,N_12022);
nor U19166 (N_19166,N_12210,N_15356);
nor U19167 (N_19167,N_14980,N_13621);
or U19168 (N_19168,N_13050,N_14819);
or U19169 (N_19169,N_13165,N_14960);
nor U19170 (N_19170,N_13589,N_14746);
nor U19171 (N_19171,N_14577,N_15296);
or U19172 (N_19172,N_13755,N_13242);
or U19173 (N_19173,N_13252,N_12224);
or U19174 (N_19174,N_13028,N_14419);
and U19175 (N_19175,N_13708,N_14571);
nor U19176 (N_19176,N_14366,N_13917);
and U19177 (N_19177,N_14389,N_15854);
nor U19178 (N_19178,N_14219,N_12698);
and U19179 (N_19179,N_12883,N_14377);
nand U19180 (N_19180,N_13249,N_14871);
nand U19181 (N_19181,N_15141,N_13085);
nor U19182 (N_19182,N_14278,N_14975);
or U19183 (N_19183,N_14960,N_15542);
nand U19184 (N_19184,N_12318,N_15958);
nand U19185 (N_19185,N_15919,N_15880);
and U19186 (N_19186,N_15619,N_14874);
nand U19187 (N_19187,N_13432,N_14063);
and U19188 (N_19188,N_13835,N_14878);
or U19189 (N_19189,N_15165,N_13445);
nor U19190 (N_19190,N_12719,N_14630);
or U19191 (N_19191,N_12633,N_14338);
or U19192 (N_19192,N_13882,N_14931);
or U19193 (N_19193,N_12660,N_15025);
or U19194 (N_19194,N_12411,N_13041);
or U19195 (N_19195,N_12371,N_12826);
or U19196 (N_19196,N_13237,N_13401);
and U19197 (N_19197,N_14888,N_12529);
nand U19198 (N_19198,N_13564,N_13535);
nor U19199 (N_19199,N_13132,N_12086);
or U19200 (N_19200,N_14122,N_12939);
nor U19201 (N_19201,N_13535,N_15724);
and U19202 (N_19202,N_14636,N_13277);
or U19203 (N_19203,N_15779,N_14280);
nand U19204 (N_19204,N_14077,N_13793);
and U19205 (N_19205,N_13778,N_15448);
nand U19206 (N_19206,N_12862,N_13252);
nand U19207 (N_19207,N_12600,N_12645);
and U19208 (N_19208,N_14002,N_14413);
nand U19209 (N_19209,N_12861,N_12692);
or U19210 (N_19210,N_12822,N_14918);
or U19211 (N_19211,N_13582,N_14454);
nand U19212 (N_19212,N_14140,N_14930);
nand U19213 (N_19213,N_14180,N_13156);
nor U19214 (N_19214,N_13289,N_15752);
nor U19215 (N_19215,N_12715,N_12795);
nand U19216 (N_19216,N_13509,N_15226);
nand U19217 (N_19217,N_13797,N_14240);
nor U19218 (N_19218,N_13614,N_12585);
or U19219 (N_19219,N_13113,N_12220);
or U19220 (N_19220,N_13869,N_13360);
and U19221 (N_19221,N_12195,N_12205);
or U19222 (N_19222,N_14895,N_14533);
and U19223 (N_19223,N_15595,N_14255);
nor U19224 (N_19224,N_12621,N_12235);
and U19225 (N_19225,N_12777,N_14332);
nor U19226 (N_19226,N_13506,N_12618);
and U19227 (N_19227,N_13949,N_12615);
nor U19228 (N_19228,N_13508,N_14121);
nor U19229 (N_19229,N_12546,N_13502);
or U19230 (N_19230,N_12773,N_15282);
and U19231 (N_19231,N_12130,N_12963);
and U19232 (N_19232,N_12906,N_15558);
or U19233 (N_19233,N_14785,N_15315);
nand U19234 (N_19234,N_14548,N_12954);
nand U19235 (N_19235,N_12961,N_14003);
nor U19236 (N_19236,N_12421,N_12185);
or U19237 (N_19237,N_14284,N_13182);
and U19238 (N_19238,N_12840,N_15249);
nor U19239 (N_19239,N_12972,N_14169);
and U19240 (N_19240,N_15809,N_15687);
and U19241 (N_19241,N_14852,N_14047);
nor U19242 (N_19242,N_14976,N_12349);
nand U19243 (N_19243,N_15126,N_15693);
nand U19244 (N_19244,N_12449,N_14442);
nand U19245 (N_19245,N_12268,N_15595);
and U19246 (N_19246,N_13569,N_15222);
nor U19247 (N_19247,N_12488,N_14374);
or U19248 (N_19248,N_14131,N_14582);
and U19249 (N_19249,N_14745,N_13126);
nand U19250 (N_19250,N_12702,N_12320);
and U19251 (N_19251,N_15189,N_12774);
or U19252 (N_19252,N_13125,N_14661);
nor U19253 (N_19253,N_12284,N_13180);
nand U19254 (N_19254,N_14875,N_12139);
nand U19255 (N_19255,N_13796,N_14551);
or U19256 (N_19256,N_12475,N_14919);
or U19257 (N_19257,N_13696,N_13728);
nand U19258 (N_19258,N_12192,N_13256);
and U19259 (N_19259,N_14081,N_14978);
and U19260 (N_19260,N_13629,N_14740);
and U19261 (N_19261,N_13384,N_13884);
nor U19262 (N_19262,N_12534,N_12779);
nor U19263 (N_19263,N_12526,N_13978);
nand U19264 (N_19264,N_15897,N_13805);
and U19265 (N_19265,N_12865,N_15573);
xor U19266 (N_19266,N_12890,N_13058);
nor U19267 (N_19267,N_12630,N_13028);
nor U19268 (N_19268,N_12022,N_14628);
nor U19269 (N_19269,N_15482,N_12490);
nand U19270 (N_19270,N_14972,N_13171);
nand U19271 (N_19271,N_13694,N_14579);
nor U19272 (N_19272,N_13789,N_12994);
or U19273 (N_19273,N_12331,N_15413);
or U19274 (N_19274,N_12626,N_13139);
xor U19275 (N_19275,N_13095,N_15282);
and U19276 (N_19276,N_15386,N_15347);
nor U19277 (N_19277,N_13518,N_13153);
and U19278 (N_19278,N_12430,N_15687);
nor U19279 (N_19279,N_14476,N_14157);
nor U19280 (N_19280,N_14217,N_14733);
xor U19281 (N_19281,N_13147,N_13001);
and U19282 (N_19282,N_13762,N_14605);
nand U19283 (N_19283,N_13669,N_14622);
or U19284 (N_19284,N_12732,N_15751);
nand U19285 (N_19285,N_13506,N_15587);
and U19286 (N_19286,N_14813,N_13866);
and U19287 (N_19287,N_14776,N_13401);
nor U19288 (N_19288,N_12625,N_13391);
nand U19289 (N_19289,N_12200,N_14850);
or U19290 (N_19290,N_15509,N_14520);
or U19291 (N_19291,N_13511,N_13202);
and U19292 (N_19292,N_15325,N_13311);
and U19293 (N_19293,N_15103,N_13980);
nand U19294 (N_19294,N_15852,N_14700);
or U19295 (N_19295,N_14056,N_14430);
and U19296 (N_19296,N_15777,N_14468);
nand U19297 (N_19297,N_13320,N_15763);
nand U19298 (N_19298,N_13039,N_12086);
and U19299 (N_19299,N_13700,N_12976);
or U19300 (N_19300,N_12861,N_15699);
nand U19301 (N_19301,N_14548,N_14960);
nor U19302 (N_19302,N_15548,N_12981);
or U19303 (N_19303,N_13195,N_15428);
nand U19304 (N_19304,N_14896,N_15991);
or U19305 (N_19305,N_13856,N_13883);
or U19306 (N_19306,N_15392,N_12675);
and U19307 (N_19307,N_15848,N_13322);
nor U19308 (N_19308,N_13035,N_12601);
or U19309 (N_19309,N_13595,N_14221);
nand U19310 (N_19310,N_12226,N_13409);
or U19311 (N_19311,N_15791,N_13077);
nor U19312 (N_19312,N_13482,N_14158);
nor U19313 (N_19313,N_15311,N_13658);
nor U19314 (N_19314,N_15482,N_14797);
nand U19315 (N_19315,N_15451,N_15356);
nand U19316 (N_19316,N_12014,N_12927);
nor U19317 (N_19317,N_12032,N_15468);
and U19318 (N_19318,N_13768,N_15785);
nor U19319 (N_19319,N_15203,N_15395);
or U19320 (N_19320,N_12193,N_14547);
nor U19321 (N_19321,N_12547,N_15622);
and U19322 (N_19322,N_13718,N_13733);
and U19323 (N_19323,N_14019,N_14686);
and U19324 (N_19324,N_14306,N_15223);
nand U19325 (N_19325,N_14242,N_13177);
nor U19326 (N_19326,N_15232,N_12167);
nand U19327 (N_19327,N_15438,N_13309);
nand U19328 (N_19328,N_14404,N_15345);
nand U19329 (N_19329,N_14425,N_13594);
and U19330 (N_19330,N_14786,N_15211);
and U19331 (N_19331,N_15312,N_12594);
and U19332 (N_19332,N_12496,N_12933);
nor U19333 (N_19333,N_14464,N_15167);
xnor U19334 (N_19334,N_15950,N_13803);
or U19335 (N_19335,N_14479,N_15435);
nor U19336 (N_19336,N_13235,N_13007);
nor U19337 (N_19337,N_13218,N_15033);
and U19338 (N_19338,N_15327,N_13390);
nand U19339 (N_19339,N_14731,N_15720);
nor U19340 (N_19340,N_14779,N_14998);
nand U19341 (N_19341,N_13542,N_15305);
and U19342 (N_19342,N_15926,N_12613);
nand U19343 (N_19343,N_13627,N_15364);
nor U19344 (N_19344,N_13935,N_12365);
nor U19345 (N_19345,N_14953,N_13573);
and U19346 (N_19346,N_15952,N_13773);
and U19347 (N_19347,N_15139,N_12406);
nor U19348 (N_19348,N_13346,N_13434);
nand U19349 (N_19349,N_12316,N_13657);
or U19350 (N_19350,N_14926,N_13330);
nand U19351 (N_19351,N_14119,N_12679);
nor U19352 (N_19352,N_14090,N_15015);
or U19353 (N_19353,N_15664,N_14907);
nor U19354 (N_19354,N_12490,N_13199);
and U19355 (N_19355,N_15984,N_14457);
nor U19356 (N_19356,N_15082,N_13004);
nor U19357 (N_19357,N_13198,N_14802);
nor U19358 (N_19358,N_15238,N_12710);
or U19359 (N_19359,N_12187,N_13560);
or U19360 (N_19360,N_14007,N_15748);
nand U19361 (N_19361,N_13081,N_12587);
nand U19362 (N_19362,N_13799,N_12236);
nor U19363 (N_19363,N_12793,N_12330);
nor U19364 (N_19364,N_13504,N_14158);
or U19365 (N_19365,N_14609,N_15812);
and U19366 (N_19366,N_14535,N_15262);
nor U19367 (N_19367,N_14099,N_12541);
or U19368 (N_19368,N_15463,N_15118);
and U19369 (N_19369,N_13207,N_13310);
nand U19370 (N_19370,N_14517,N_14518);
nor U19371 (N_19371,N_12499,N_14659);
nor U19372 (N_19372,N_12544,N_12716);
and U19373 (N_19373,N_14335,N_15911);
or U19374 (N_19374,N_14050,N_12179);
nor U19375 (N_19375,N_14604,N_12356);
or U19376 (N_19376,N_12811,N_12422);
or U19377 (N_19377,N_15480,N_12178);
or U19378 (N_19378,N_14972,N_15139);
nand U19379 (N_19379,N_12269,N_15832);
or U19380 (N_19380,N_14180,N_12826);
nand U19381 (N_19381,N_12869,N_15048);
nor U19382 (N_19382,N_12745,N_12668);
nand U19383 (N_19383,N_12505,N_14634);
nor U19384 (N_19384,N_13418,N_12988);
or U19385 (N_19385,N_15794,N_15956);
nor U19386 (N_19386,N_12691,N_15374);
or U19387 (N_19387,N_14037,N_13663);
and U19388 (N_19388,N_15891,N_13410);
nand U19389 (N_19389,N_13252,N_13258);
or U19390 (N_19390,N_15837,N_14063);
or U19391 (N_19391,N_12594,N_14791);
and U19392 (N_19392,N_15617,N_13603);
or U19393 (N_19393,N_12666,N_12828);
xor U19394 (N_19394,N_15338,N_14478);
and U19395 (N_19395,N_12255,N_12298);
or U19396 (N_19396,N_12528,N_15001);
nand U19397 (N_19397,N_12680,N_12878);
or U19398 (N_19398,N_13903,N_15987);
or U19399 (N_19399,N_14205,N_13221);
or U19400 (N_19400,N_15368,N_15271);
xor U19401 (N_19401,N_14600,N_12233);
and U19402 (N_19402,N_15858,N_14220);
and U19403 (N_19403,N_12407,N_13305);
nand U19404 (N_19404,N_14420,N_12073);
or U19405 (N_19405,N_15407,N_12890);
or U19406 (N_19406,N_12587,N_12647);
or U19407 (N_19407,N_12117,N_12645);
or U19408 (N_19408,N_14907,N_13706);
or U19409 (N_19409,N_15219,N_12463);
nor U19410 (N_19410,N_13715,N_14003);
or U19411 (N_19411,N_13120,N_15390);
nor U19412 (N_19412,N_14513,N_12948);
or U19413 (N_19413,N_14313,N_14084);
or U19414 (N_19414,N_13589,N_13732);
and U19415 (N_19415,N_12278,N_15894);
and U19416 (N_19416,N_15901,N_15433);
and U19417 (N_19417,N_13327,N_13475);
nor U19418 (N_19418,N_15537,N_13537);
or U19419 (N_19419,N_13949,N_13367);
nor U19420 (N_19420,N_12650,N_13495);
nand U19421 (N_19421,N_15890,N_12114);
nand U19422 (N_19422,N_14769,N_12121);
nand U19423 (N_19423,N_13122,N_15295);
or U19424 (N_19424,N_13130,N_12707);
nand U19425 (N_19425,N_15538,N_15264);
xnor U19426 (N_19426,N_12881,N_13562);
and U19427 (N_19427,N_12269,N_12944);
or U19428 (N_19428,N_12459,N_12971);
and U19429 (N_19429,N_15283,N_15696);
nor U19430 (N_19430,N_13076,N_14541);
or U19431 (N_19431,N_12503,N_13936);
nor U19432 (N_19432,N_14396,N_13543);
or U19433 (N_19433,N_14368,N_13079);
and U19434 (N_19434,N_12384,N_12999);
or U19435 (N_19435,N_15292,N_12907);
or U19436 (N_19436,N_13357,N_14174);
nand U19437 (N_19437,N_14763,N_13082);
or U19438 (N_19438,N_13951,N_14449);
nor U19439 (N_19439,N_13709,N_15639);
and U19440 (N_19440,N_14655,N_13218);
nand U19441 (N_19441,N_12156,N_12517);
nand U19442 (N_19442,N_14938,N_15459);
or U19443 (N_19443,N_13089,N_14032);
nand U19444 (N_19444,N_13414,N_15575);
or U19445 (N_19445,N_14703,N_13362);
nor U19446 (N_19446,N_15024,N_13142);
nor U19447 (N_19447,N_15349,N_13569);
nor U19448 (N_19448,N_13206,N_13409);
or U19449 (N_19449,N_14712,N_13333);
nand U19450 (N_19450,N_13799,N_12107);
or U19451 (N_19451,N_15895,N_14091);
and U19452 (N_19452,N_14388,N_14375);
or U19453 (N_19453,N_12576,N_14721);
nand U19454 (N_19454,N_15950,N_12838);
nand U19455 (N_19455,N_13192,N_14444);
nor U19456 (N_19456,N_15022,N_13292);
nor U19457 (N_19457,N_14579,N_15127);
and U19458 (N_19458,N_15255,N_13396);
and U19459 (N_19459,N_12013,N_15877);
or U19460 (N_19460,N_14933,N_12419);
and U19461 (N_19461,N_14982,N_13420);
and U19462 (N_19462,N_14600,N_13496);
xor U19463 (N_19463,N_15777,N_15202);
or U19464 (N_19464,N_14956,N_13972);
nand U19465 (N_19465,N_15659,N_15149);
nor U19466 (N_19466,N_14135,N_12207);
nand U19467 (N_19467,N_15087,N_14874);
and U19468 (N_19468,N_12255,N_15091);
nor U19469 (N_19469,N_14239,N_14887);
nor U19470 (N_19470,N_12286,N_12063);
or U19471 (N_19471,N_13204,N_13833);
nor U19472 (N_19472,N_12389,N_14908);
nand U19473 (N_19473,N_12558,N_12542);
nand U19474 (N_19474,N_13835,N_12828);
nor U19475 (N_19475,N_13888,N_14365);
xor U19476 (N_19476,N_13174,N_13548);
nand U19477 (N_19477,N_12734,N_12283);
nand U19478 (N_19478,N_13512,N_13662);
and U19479 (N_19479,N_14290,N_15078);
and U19480 (N_19480,N_15012,N_12406);
nor U19481 (N_19481,N_13589,N_15752);
and U19482 (N_19482,N_15799,N_12909);
nor U19483 (N_19483,N_13528,N_15748);
nor U19484 (N_19484,N_13633,N_13775);
and U19485 (N_19485,N_13358,N_13796);
nand U19486 (N_19486,N_12080,N_15834);
or U19487 (N_19487,N_12414,N_14709);
nor U19488 (N_19488,N_14415,N_15202);
or U19489 (N_19489,N_13905,N_12300);
or U19490 (N_19490,N_12675,N_13741);
and U19491 (N_19491,N_15343,N_14231);
nor U19492 (N_19492,N_15698,N_14972);
or U19493 (N_19493,N_12754,N_15720);
nor U19494 (N_19494,N_14514,N_12055);
nand U19495 (N_19495,N_15717,N_14681);
nor U19496 (N_19496,N_13694,N_13956);
and U19497 (N_19497,N_14633,N_12404);
nand U19498 (N_19498,N_12419,N_12898);
xor U19499 (N_19499,N_12321,N_15929);
and U19500 (N_19500,N_15198,N_12978);
or U19501 (N_19501,N_12503,N_13327);
nor U19502 (N_19502,N_12649,N_13221);
nor U19503 (N_19503,N_14421,N_14398);
and U19504 (N_19504,N_14206,N_12887);
and U19505 (N_19505,N_13348,N_15812);
or U19506 (N_19506,N_13701,N_14410);
or U19507 (N_19507,N_12831,N_12958);
nor U19508 (N_19508,N_14434,N_12502);
xnor U19509 (N_19509,N_15763,N_13353);
nor U19510 (N_19510,N_14632,N_13951);
or U19511 (N_19511,N_12775,N_13177);
nand U19512 (N_19512,N_15206,N_15932);
or U19513 (N_19513,N_13832,N_12609);
nand U19514 (N_19514,N_14389,N_12739);
and U19515 (N_19515,N_15585,N_13209);
or U19516 (N_19516,N_13458,N_14488);
nand U19517 (N_19517,N_14123,N_13710);
and U19518 (N_19518,N_15032,N_12199);
and U19519 (N_19519,N_13087,N_12066);
nor U19520 (N_19520,N_15285,N_14409);
nor U19521 (N_19521,N_12262,N_12123);
nand U19522 (N_19522,N_14984,N_12200);
nand U19523 (N_19523,N_15333,N_13780);
or U19524 (N_19524,N_15222,N_15397);
and U19525 (N_19525,N_13807,N_12691);
nand U19526 (N_19526,N_12616,N_15946);
nor U19527 (N_19527,N_12771,N_15201);
nand U19528 (N_19528,N_15312,N_15902);
nor U19529 (N_19529,N_15721,N_13809);
and U19530 (N_19530,N_14964,N_15040);
nor U19531 (N_19531,N_13273,N_14002);
or U19532 (N_19532,N_14836,N_15033);
or U19533 (N_19533,N_12448,N_14571);
nor U19534 (N_19534,N_14625,N_14396);
nand U19535 (N_19535,N_12385,N_12163);
nor U19536 (N_19536,N_14270,N_14287);
or U19537 (N_19537,N_15068,N_13994);
nor U19538 (N_19538,N_13436,N_13190);
and U19539 (N_19539,N_14094,N_15298);
and U19540 (N_19540,N_14796,N_13380);
and U19541 (N_19541,N_13299,N_13157);
nor U19542 (N_19542,N_15949,N_15616);
or U19543 (N_19543,N_15676,N_15668);
or U19544 (N_19544,N_13389,N_12258);
or U19545 (N_19545,N_15723,N_13238);
nor U19546 (N_19546,N_15772,N_14175);
nor U19547 (N_19547,N_14798,N_15319);
nor U19548 (N_19548,N_15150,N_13775);
nand U19549 (N_19549,N_13653,N_15441);
nor U19550 (N_19550,N_14298,N_13630);
nand U19551 (N_19551,N_13066,N_12450);
nand U19552 (N_19552,N_13586,N_13673);
or U19553 (N_19553,N_13299,N_14861);
and U19554 (N_19554,N_14330,N_12446);
nor U19555 (N_19555,N_15062,N_12718);
nand U19556 (N_19556,N_13477,N_15771);
or U19557 (N_19557,N_12196,N_15570);
nand U19558 (N_19558,N_15942,N_14709);
nor U19559 (N_19559,N_12581,N_15967);
nand U19560 (N_19560,N_13114,N_14015);
nor U19561 (N_19561,N_14614,N_15058);
nor U19562 (N_19562,N_13913,N_15241);
nand U19563 (N_19563,N_13686,N_15506);
nor U19564 (N_19564,N_14277,N_13672);
nor U19565 (N_19565,N_12380,N_15813);
nor U19566 (N_19566,N_12552,N_13313);
nand U19567 (N_19567,N_12493,N_15406);
nor U19568 (N_19568,N_12096,N_12049);
nand U19569 (N_19569,N_12230,N_12258);
xnor U19570 (N_19570,N_14944,N_15597);
nor U19571 (N_19571,N_12424,N_15972);
and U19572 (N_19572,N_13699,N_13080);
and U19573 (N_19573,N_14653,N_14921);
nor U19574 (N_19574,N_13402,N_12923);
nand U19575 (N_19575,N_14017,N_14626);
nand U19576 (N_19576,N_13010,N_12587);
and U19577 (N_19577,N_14772,N_15678);
or U19578 (N_19578,N_15297,N_13751);
and U19579 (N_19579,N_12491,N_14775);
or U19580 (N_19580,N_14365,N_13926);
or U19581 (N_19581,N_13318,N_12489);
nand U19582 (N_19582,N_13812,N_13599);
and U19583 (N_19583,N_15177,N_14811);
nand U19584 (N_19584,N_12365,N_15696);
nor U19585 (N_19585,N_13746,N_15358);
and U19586 (N_19586,N_14438,N_12469);
and U19587 (N_19587,N_13587,N_15684);
nand U19588 (N_19588,N_12327,N_15934);
nor U19589 (N_19589,N_12055,N_14846);
nor U19590 (N_19590,N_15814,N_13568);
nor U19591 (N_19591,N_14243,N_15507);
nand U19592 (N_19592,N_13249,N_12930);
and U19593 (N_19593,N_13423,N_15980);
nand U19594 (N_19594,N_12721,N_15537);
and U19595 (N_19595,N_13790,N_13236);
and U19596 (N_19596,N_12253,N_12206);
and U19597 (N_19597,N_14502,N_14148);
nand U19598 (N_19598,N_15967,N_12742);
nand U19599 (N_19599,N_14300,N_15546);
nand U19600 (N_19600,N_12975,N_15329);
nor U19601 (N_19601,N_13447,N_12607);
and U19602 (N_19602,N_12050,N_14026);
or U19603 (N_19603,N_14223,N_15921);
nor U19604 (N_19604,N_12698,N_12779);
and U19605 (N_19605,N_14156,N_15420);
or U19606 (N_19606,N_13669,N_13484);
nor U19607 (N_19607,N_14141,N_14030);
and U19608 (N_19608,N_15984,N_13328);
or U19609 (N_19609,N_13781,N_12908);
and U19610 (N_19610,N_13114,N_13270);
or U19611 (N_19611,N_12916,N_13013);
or U19612 (N_19612,N_12687,N_14662);
nor U19613 (N_19613,N_13839,N_12900);
and U19614 (N_19614,N_13331,N_13144);
xor U19615 (N_19615,N_14474,N_15252);
and U19616 (N_19616,N_14655,N_15847);
nand U19617 (N_19617,N_13637,N_14346);
nor U19618 (N_19618,N_14731,N_13685);
or U19619 (N_19619,N_14360,N_12595);
and U19620 (N_19620,N_13235,N_13219);
nor U19621 (N_19621,N_12834,N_13044);
or U19622 (N_19622,N_13594,N_12166);
or U19623 (N_19623,N_13720,N_12867);
and U19624 (N_19624,N_15994,N_13840);
or U19625 (N_19625,N_14302,N_14260);
nor U19626 (N_19626,N_14077,N_14750);
nand U19627 (N_19627,N_14165,N_15956);
nand U19628 (N_19628,N_15700,N_15851);
and U19629 (N_19629,N_15898,N_15001);
nor U19630 (N_19630,N_12209,N_13258);
and U19631 (N_19631,N_15899,N_15032);
nand U19632 (N_19632,N_13539,N_13860);
or U19633 (N_19633,N_15360,N_15046);
and U19634 (N_19634,N_14967,N_12437);
or U19635 (N_19635,N_12659,N_15213);
and U19636 (N_19636,N_14027,N_13796);
or U19637 (N_19637,N_12570,N_13151);
or U19638 (N_19638,N_14685,N_15477);
and U19639 (N_19639,N_13053,N_12884);
or U19640 (N_19640,N_14911,N_15807);
nand U19641 (N_19641,N_15245,N_12342);
nand U19642 (N_19642,N_14121,N_13335);
nand U19643 (N_19643,N_15731,N_15985);
and U19644 (N_19644,N_13960,N_15833);
nor U19645 (N_19645,N_12208,N_14453);
nor U19646 (N_19646,N_14168,N_14803);
nor U19647 (N_19647,N_13221,N_15701);
and U19648 (N_19648,N_14644,N_14662);
and U19649 (N_19649,N_13286,N_12778);
or U19650 (N_19650,N_12365,N_12839);
nor U19651 (N_19651,N_13607,N_13453);
or U19652 (N_19652,N_15168,N_14890);
or U19653 (N_19653,N_13068,N_15592);
nand U19654 (N_19654,N_12420,N_12902);
or U19655 (N_19655,N_15617,N_14617);
or U19656 (N_19656,N_12697,N_13761);
and U19657 (N_19657,N_13605,N_14663);
nand U19658 (N_19658,N_15894,N_15825);
nor U19659 (N_19659,N_13953,N_12648);
nor U19660 (N_19660,N_13406,N_14272);
and U19661 (N_19661,N_12497,N_13089);
nor U19662 (N_19662,N_15223,N_15144);
nor U19663 (N_19663,N_14555,N_15631);
nand U19664 (N_19664,N_15838,N_14270);
or U19665 (N_19665,N_12726,N_15543);
or U19666 (N_19666,N_12767,N_14902);
and U19667 (N_19667,N_12048,N_12884);
or U19668 (N_19668,N_15366,N_13596);
and U19669 (N_19669,N_13155,N_14107);
nand U19670 (N_19670,N_15204,N_13281);
nand U19671 (N_19671,N_15794,N_13029);
nor U19672 (N_19672,N_15286,N_15779);
or U19673 (N_19673,N_14269,N_14061);
or U19674 (N_19674,N_13107,N_13460);
or U19675 (N_19675,N_15689,N_12115);
or U19676 (N_19676,N_13672,N_13036);
nor U19677 (N_19677,N_14369,N_14857);
or U19678 (N_19678,N_12483,N_15814);
nor U19679 (N_19679,N_14953,N_14736);
and U19680 (N_19680,N_14052,N_13407);
nand U19681 (N_19681,N_14162,N_15855);
and U19682 (N_19682,N_14337,N_12267);
nand U19683 (N_19683,N_12988,N_15651);
nor U19684 (N_19684,N_12020,N_12155);
or U19685 (N_19685,N_14772,N_13430);
or U19686 (N_19686,N_13778,N_12610);
or U19687 (N_19687,N_15946,N_13791);
or U19688 (N_19688,N_13023,N_14012);
or U19689 (N_19689,N_12588,N_15753);
and U19690 (N_19690,N_12788,N_12577);
or U19691 (N_19691,N_14493,N_13053);
nand U19692 (N_19692,N_14537,N_14779);
nand U19693 (N_19693,N_15703,N_13073);
nor U19694 (N_19694,N_14446,N_14413);
nand U19695 (N_19695,N_12505,N_15488);
or U19696 (N_19696,N_14976,N_12140);
or U19697 (N_19697,N_13104,N_14197);
nor U19698 (N_19698,N_12927,N_14071);
or U19699 (N_19699,N_13483,N_12588);
and U19700 (N_19700,N_13945,N_15420);
nor U19701 (N_19701,N_15388,N_15077);
or U19702 (N_19702,N_15664,N_14178);
and U19703 (N_19703,N_13073,N_12969);
or U19704 (N_19704,N_15927,N_15713);
nand U19705 (N_19705,N_12612,N_14144);
and U19706 (N_19706,N_13567,N_12409);
nor U19707 (N_19707,N_14337,N_12127);
nor U19708 (N_19708,N_12285,N_12415);
or U19709 (N_19709,N_13869,N_13933);
and U19710 (N_19710,N_13658,N_12612);
nor U19711 (N_19711,N_12141,N_12005);
and U19712 (N_19712,N_15384,N_12578);
or U19713 (N_19713,N_14515,N_15816);
or U19714 (N_19714,N_15981,N_13680);
or U19715 (N_19715,N_13496,N_13039);
or U19716 (N_19716,N_13342,N_15362);
or U19717 (N_19717,N_14335,N_14095);
nand U19718 (N_19718,N_13311,N_15184);
or U19719 (N_19719,N_12993,N_14876);
and U19720 (N_19720,N_15686,N_13857);
nor U19721 (N_19721,N_12768,N_12839);
nor U19722 (N_19722,N_14231,N_13761);
and U19723 (N_19723,N_14157,N_14191);
and U19724 (N_19724,N_14606,N_12081);
nor U19725 (N_19725,N_12938,N_15739);
and U19726 (N_19726,N_13245,N_14374);
and U19727 (N_19727,N_12256,N_14810);
nand U19728 (N_19728,N_14279,N_14551);
or U19729 (N_19729,N_12934,N_15388);
nor U19730 (N_19730,N_12830,N_13974);
and U19731 (N_19731,N_15028,N_14162);
nor U19732 (N_19732,N_13642,N_13014);
nand U19733 (N_19733,N_14577,N_14257);
or U19734 (N_19734,N_12716,N_14966);
and U19735 (N_19735,N_13961,N_15653);
or U19736 (N_19736,N_12543,N_15201);
and U19737 (N_19737,N_12716,N_14752);
nand U19738 (N_19738,N_13638,N_13407);
nand U19739 (N_19739,N_12650,N_15947);
and U19740 (N_19740,N_15238,N_13489);
nand U19741 (N_19741,N_14015,N_14647);
and U19742 (N_19742,N_12387,N_15438);
and U19743 (N_19743,N_12006,N_12658);
nand U19744 (N_19744,N_15517,N_15117);
or U19745 (N_19745,N_14645,N_14791);
nor U19746 (N_19746,N_13758,N_15274);
nor U19747 (N_19747,N_14858,N_13232);
xor U19748 (N_19748,N_13407,N_15649);
and U19749 (N_19749,N_15542,N_12785);
nand U19750 (N_19750,N_14572,N_15312);
nor U19751 (N_19751,N_12618,N_13859);
nor U19752 (N_19752,N_14060,N_14435);
and U19753 (N_19753,N_13484,N_15986);
and U19754 (N_19754,N_15829,N_12222);
nand U19755 (N_19755,N_14855,N_12094);
nand U19756 (N_19756,N_13082,N_12261);
nand U19757 (N_19757,N_12185,N_13571);
or U19758 (N_19758,N_12753,N_15234);
nand U19759 (N_19759,N_12828,N_15635);
or U19760 (N_19760,N_13230,N_14285);
or U19761 (N_19761,N_12042,N_14235);
nor U19762 (N_19762,N_13538,N_12550);
nand U19763 (N_19763,N_13502,N_13677);
and U19764 (N_19764,N_15627,N_12007);
and U19765 (N_19765,N_13634,N_14114);
and U19766 (N_19766,N_15074,N_15576);
nand U19767 (N_19767,N_14229,N_15381);
or U19768 (N_19768,N_12514,N_12097);
or U19769 (N_19769,N_12799,N_13528);
or U19770 (N_19770,N_12844,N_13537);
or U19771 (N_19771,N_15609,N_12904);
or U19772 (N_19772,N_15810,N_15671);
and U19773 (N_19773,N_15597,N_12257);
nand U19774 (N_19774,N_15274,N_13936);
and U19775 (N_19775,N_14168,N_15694);
nor U19776 (N_19776,N_12242,N_12421);
nor U19777 (N_19777,N_12798,N_13762);
and U19778 (N_19778,N_14967,N_15627);
and U19779 (N_19779,N_15881,N_13820);
and U19780 (N_19780,N_13170,N_15325);
nand U19781 (N_19781,N_12697,N_13916);
nand U19782 (N_19782,N_12366,N_13886);
nor U19783 (N_19783,N_13966,N_14346);
and U19784 (N_19784,N_12288,N_13885);
or U19785 (N_19785,N_14868,N_15927);
and U19786 (N_19786,N_15444,N_12020);
or U19787 (N_19787,N_14583,N_12068);
and U19788 (N_19788,N_14901,N_14297);
nor U19789 (N_19789,N_15872,N_15288);
nand U19790 (N_19790,N_15675,N_15392);
nor U19791 (N_19791,N_14472,N_14688);
or U19792 (N_19792,N_12031,N_13227);
nand U19793 (N_19793,N_12640,N_14397);
nand U19794 (N_19794,N_14244,N_14860);
and U19795 (N_19795,N_13546,N_13890);
nand U19796 (N_19796,N_14061,N_14610);
nand U19797 (N_19797,N_13384,N_12225);
xnor U19798 (N_19798,N_14866,N_13810);
or U19799 (N_19799,N_12991,N_12720);
or U19800 (N_19800,N_12261,N_13625);
nand U19801 (N_19801,N_14355,N_15544);
nor U19802 (N_19802,N_13925,N_12590);
and U19803 (N_19803,N_15027,N_12364);
and U19804 (N_19804,N_12513,N_14784);
and U19805 (N_19805,N_12479,N_13967);
and U19806 (N_19806,N_15261,N_12252);
nor U19807 (N_19807,N_15569,N_13315);
or U19808 (N_19808,N_15691,N_14621);
or U19809 (N_19809,N_12085,N_15105);
or U19810 (N_19810,N_12058,N_14871);
and U19811 (N_19811,N_12064,N_12867);
or U19812 (N_19812,N_15200,N_12975);
nand U19813 (N_19813,N_13071,N_14220);
nor U19814 (N_19814,N_14187,N_14505);
and U19815 (N_19815,N_12768,N_12288);
or U19816 (N_19816,N_12679,N_15982);
or U19817 (N_19817,N_12132,N_15052);
nor U19818 (N_19818,N_12555,N_14069);
or U19819 (N_19819,N_14486,N_13248);
and U19820 (N_19820,N_15611,N_15016);
nor U19821 (N_19821,N_12632,N_15440);
or U19822 (N_19822,N_14105,N_13569);
or U19823 (N_19823,N_14656,N_13963);
nor U19824 (N_19824,N_12637,N_13393);
nor U19825 (N_19825,N_13848,N_13089);
nand U19826 (N_19826,N_12735,N_15654);
nand U19827 (N_19827,N_14527,N_14622);
and U19828 (N_19828,N_13294,N_14955);
nand U19829 (N_19829,N_13451,N_15427);
and U19830 (N_19830,N_14593,N_12996);
nand U19831 (N_19831,N_14263,N_13887);
or U19832 (N_19832,N_13248,N_13318);
or U19833 (N_19833,N_12007,N_13350);
nand U19834 (N_19834,N_15420,N_12697);
or U19835 (N_19835,N_12361,N_15613);
or U19836 (N_19836,N_14934,N_12957);
nor U19837 (N_19837,N_13031,N_13331);
or U19838 (N_19838,N_15037,N_14324);
nor U19839 (N_19839,N_12864,N_12250);
nand U19840 (N_19840,N_13976,N_14404);
or U19841 (N_19841,N_14974,N_15018);
nor U19842 (N_19842,N_12904,N_14506);
nor U19843 (N_19843,N_14221,N_15430);
nand U19844 (N_19844,N_13765,N_12028);
or U19845 (N_19845,N_12265,N_14014);
nand U19846 (N_19846,N_13488,N_13231);
nor U19847 (N_19847,N_13091,N_14487);
and U19848 (N_19848,N_12524,N_14538);
nor U19849 (N_19849,N_15124,N_14545);
and U19850 (N_19850,N_15802,N_12173);
nand U19851 (N_19851,N_13429,N_14995);
nand U19852 (N_19852,N_15808,N_15321);
or U19853 (N_19853,N_15571,N_13806);
nand U19854 (N_19854,N_13358,N_12718);
nand U19855 (N_19855,N_14248,N_14527);
nor U19856 (N_19856,N_15363,N_15600);
or U19857 (N_19857,N_15579,N_14632);
nor U19858 (N_19858,N_12497,N_15921);
nor U19859 (N_19859,N_12899,N_15306);
nor U19860 (N_19860,N_14816,N_12792);
xor U19861 (N_19861,N_15874,N_14784);
nor U19862 (N_19862,N_15631,N_14901);
and U19863 (N_19863,N_14907,N_15460);
or U19864 (N_19864,N_14853,N_13969);
or U19865 (N_19865,N_12477,N_13311);
and U19866 (N_19866,N_14929,N_15754);
or U19867 (N_19867,N_14834,N_12529);
and U19868 (N_19868,N_14773,N_12613);
and U19869 (N_19869,N_14874,N_14404);
nor U19870 (N_19870,N_12714,N_14969);
nand U19871 (N_19871,N_15480,N_15343);
nor U19872 (N_19872,N_15475,N_15666);
nand U19873 (N_19873,N_15482,N_15483);
nand U19874 (N_19874,N_15031,N_15427);
nand U19875 (N_19875,N_12116,N_15292);
nor U19876 (N_19876,N_15051,N_14318);
nand U19877 (N_19877,N_15978,N_14801);
nand U19878 (N_19878,N_14579,N_13103);
nor U19879 (N_19879,N_15386,N_15596);
nor U19880 (N_19880,N_12030,N_13556);
xnor U19881 (N_19881,N_14808,N_14216);
and U19882 (N_19882,N_13464,N_14533);
and U19883 (N_19883,N_13599,N_14853);
nand U19884 (N_19884,N_12430,N_15899);
and U19885 (N_19885,N_15783,N_14771);
and U19886 (N_19886,N_14311,N_14127);
and U19887 (N_19887,N_15354,N_14195);
nor U19888 (N_19888,N_12136,N_12878);
nand U19889 (N_19889,N_14930,N_15139);
nand U19890 (N_19890,N_15281,N_12890);
nand U19891 (N_19891,N_13481,N_13870);
or U19892 (N_19892,N_14907,N_14666);
nor U19893 (N_19893,N_13580,N_12318);
and U19894 (N_19894,N_14260,N_13796);
and U19895 (N_19895,N_13665,N_12159);
and U19896 (N_19896,N_12767,N_14520);
or U19897 (N_19897,N_14057,N_13837);
or U19898 (N_19898,N_15972,N_13365);
or U19899 (N_19899,N_13049,N_12359);
nand U19900 (N_19900,N_14771,N_12017);
nand U19901 (N_19901,N_12900,N_15301);
nor U19902 (N_19902,N_14759,N_14867);
or U19903 (N_19903,N_15643,N_14594);
nor U19904 (N_19904,N_15919,N_13613);
nand U19905 (N_19905,N_14231,N_14144);
and U19906 (N_19906,N_13912,N_14351);
nand U19907 (N_19907,N_13843,N_15356);
nor U19908 (N_19908,N_14322,N_12632);
and U19909 (N_19909,N_12330,N_15764);
nor U19910 (N_19910,N_13712,N_15333);
nor U19911 (N_19911,N_15691,N_15657);
nor U19912 (N_19912,N_14542,N_15328);
nand U19913 (N_19913,N_12847,N_12368);
and U19914 (N_19914,N_12050,N_12336);
nor U19915 (N_19915,N_14349,N_15386);
nand U19916 (N_19916,N_13232,N_14821);
nand U19917 (N_19917,N_15070,N_12019);
or U19918 (N_19918,N_14670,N_12141);
nand U19919 (N_19919,N_13116,N_12936);
nand U19920 (N_19920,N_13306,N_15879);
or U19921 (N_19921,N_14720,N_12257);
and U19922 (N_19922,N_13363,N_13016);
and U19923 (N_19923,N_14154,N_15887);
or U19924 (N_19924,N_15798,N_12782);
or U19925 (N_19925,N_13052,N_12602);
and U19926 (N_19926,N_12599,N_15718);
or U19927 (N_19927,N_13626,N_15076);
or U19928 (N_19928,N_15827,N_13275);
and U19929 (N_19929,N_15770,N_14118);
nand U19930 (N_19930,N_15667,N_15781);
or U19931 (N_19931,N_12089,N_12823);
nand U19932 (N_19932,N_13061,N_13901);
or U19933 (N_19933,N_15625,N_15417);
nand U19934 (N_19934,N_15485,N_15972);
and U19935 (N_19935,N_13278,N_12106);
or U19936 (N_19936,N_12367,N_12300);
or U19937 (N_19937,N_14993,N_13215);
nor U19938 (N_19938,N_15037,N_15072);
and U19939 (N_19939,N_13036,N_12628);
and U19940 (N_19940,N_14399,N_13973);
nand U19941 (N_19941,N_13682,N_14511);
nand U19942 (N_19942,N_13564,N_13337);
and U19943 (N_19943,N_15612,N_12464);
and U19944 (N_19944,N_14053,N_12219);
and U19945 (N_19945,N_12222,N_13275);
nor U19946 (N_19946,N_12533,N_15555);
and U19947 (N_19947,N_13597,N_14503);
or U19948 (N_19948,N_12267,N_12019);
or U19949 (N_19949,N_12260,N_13261);
or U19950 (N_19950,N_13083,N_15045);
nand U19951 (N_19951,N_12184,N_12740);
nor U19952 (N_19952,N_14571,N_15017);
and U19953 (N_19953,N_12327,N_13741);
or U19954 (N_19954,N_13806,N_14944);
or U19955 (N_19955,N_12489,N_12581);
nand U19956 (N_19956,N_12290,N_12703);
nand U19957 (N_19957,N_15219,N_15095);
nand U19958 (N_19958,N_12949,N_14281);
or U19959 (N_19959,N_15074,N_15771);
or U19960 (N_19960,N_15458,N_13528);
nand U19961 (N_19961,N_12674,N_14311);
nand U19962 (N_19962,N_13436,N_15398);
nor U19963 (N_19963,N_14155,N_15408);
or U19964 (N_19964,N_12653,N_14673);
nor U19965 (N_19965,N_15633,N_12296);
nor U19966 (N_19966,N_13597,N_12754);
or U19967 (N_19967,N_14753,N_12502);
and U19968 (N_19968,N_12979,N_13504);
nor U19969 (N_19969,N_14172,N_14542);
and U19970 (N_19970,N_14359,N_13348);
or U19971 (N_19971,N_14457,N_13894);
nor U19972 (N_19972,N_15031,N_15017);
or U19973 (N_19973,N_14101,N_12151);
and U19974 (N_19974,N_14971,N_12295);
or U19975 (N_19975,N_13176,N_13119);
and U19976 (N_19976,N_13015,N_13330);
and U19977 (N_19977,N_13726,N_14376);
nor U19978 (N_19978,N_13535,N_14002);
and U19979 (N_19979,N_12889,N_12876);
or U19980 (N_19980,N_15031,N_13995);
or U19981 (N_19981,N_15503,N_13866);
and U19982 (N_19982,N_14873,N_14767);
nand U19983 (N_19983,N_12077,N_13499);
xnor U19984 (N_19984,N_15979,N_12977);
nand U19985 (N_19985,N_12732,N_13888);
nor U19986 (N_19986,N_15100,N_14161);
and U19987 (N_19987,N_14422,N_13366);
nand U19988 (N_19988,N_15495,N_13314);
and U19989 (N_19989,N_13361,N_12686);
nand U19990 (N_19990,N_13758,N_12300);
nand U19991 (N_19991,N_14368,N_12335);
and U19992 (N_19992,N_12657,N_12460);
and U19993 (N_19993,N_12015,N_15568);
or U19994 (N_19994,N_13464,N_12649);
nand U19995 (N_19995,N_12022,N_14394);
nor U19996 (N_19996,N_15521,N_15138);
or U19997 (N_19997,N_15684,N_14077);
nand U19998 (N_19998,N_12131,N_13596);
xnor U19999 (N_19999,N_12332,N_13215);
or UO_0 (O_0,N_19109,N_16825);
and UO_1 (O_1,N_17641,N_16093);
and UO_2 (O_2,N_16740,N_16896);
xnor UO_3 (O_3,N_17833,N_17254);
nor UO_4 (O_4,N_19269,N_17984);
nand UO_5 (O_5,N_18647,N_19210);
nor UO_6 (O_6,N_16866,N_17938);
nor UO_7 (O_7,N_19317,N_16432);
or UO_8 (O_8,N_19534,N_17924);
nand UO_9 (O_9,N_18544,N_17502);
and UO_10 (O_10,N_19642,N_18917);
or UO_11 (O_11,N_17644,N_19896);
or UO_12 (O_12,N_19571,N_18916);
and UO_13 (O_13,N_16722,N_18008);
or UO_14 (O_14,N_16876,N_17554);
nor UO_15 (O_15,N_18998,N_19915);
nor UO_16 (O_16,N_19004,N_17677);
nand UO_17 (O_17,N_16552,N_18040);
and UO_18 (O_18,N_16182,N_17671);
nor UO_19 (O_19,N_17031,N_19715);
nand UO_20 (O_20,N_19398,N_17816);
or UO_21 (O_21,N_16021,N_17224);
and UO_22 (O_22,N_16696,N_19339);
nand UO_23 (O_23,N_18278,N_17615);
nand UO_24 (O_24,N_16675,N_19048);
nand UO_25 (O_25,N_18273,N_17587);
nand UO_26 (O_26,N_19789,N_17464);
nand UO_27 (O_27,N_16512,N_18759);
nor UO_28 (O_28,N_16116,N_19712);
nor UO_29 (O_29,N_17434,N_19679);
nor UO_30 (O_30,N_17424,N_19652);
or UO_31 (O_31,N_17474,N_19047);
and UO_32 (O_32,N_17949,N_16090);
nand UO_33 (O_33,N_16530,N_17020);
or UO_34 (O_34,N_19201,N_16578);
nand UO_35 (O_35,N_16789,N_16726);
nand UO_36 (O_36,N_16461,N_17828);
and UO_37 (O_37,N_16854,N_18626);
or UO_38 (O_38,N_19344,N_16306);
and UO_39 (O_39,N_17163,N_19010);
nor UO_40 (O_40,N_17574,N_17704);
nand UO_41 (O_41,N_18932,N_19887);
and UO_42 (O_42,N_19076,N_16573);
xnor UO_43 (O_43,N_19550,N_19877);
nand UO_44 (O_44,N_16074,N_16155);
nand UO_45 (O_45,N_18120,N_16180);
or UO_46 (O_46,N_19916,N_16503);
or UO_47 (O_47,N_16786,N_19893);
or UO_48 (O_48,N_17810,N_18638);
or UO_49 (O_49,N_18750,N_18337);
and UO_50 (O_50,N_17981,N_19529);
nor UO_51 (O_51,N_16707,N_19346);
or UO_52 (O_52,N_19666,N_18828);
nand UO_53 (O_53,N_19836,N_19357);
nand UO_54 (O_54,N_19116,N_18241);
nand UO_55 (O_55,N_17771,N_16792);
or UO_56 (O_56,N_18509,N_17097);
or UO_57 (O_57,N_16905,N_19886);
or UO_58 (O_58,N_16625,N_19823);
and UO_59 (O_59,N_19145,N_18595);
and UO_60 (O_60,N_16001,N_16233);
and UO_61 (O_61,N_19178,N_19502);
nor UO_62 (O_62,N_17272,N_19921);
nand UO_63 (O_63,N_18719,N_17011);
nand UO_64 (O_64,N_16504,N_18801);
xnor UO_65 (O_65,N_19544,N_16641);
nand UO_66 (O_66,N_19624,N_16010);
nor UO_67 (O_67,N_16126,N_19997);
nand UO_68 (O_68,N_17923,N_19956);
nand UO_69 (O_69,N_16351,N_18649);
nand UO_70 (O_70,N_17822,N_16883);
nand UO_71 (O_71,N_18812,N_16867);
nand UO_72 (O_72,N_19373,N_19432);
nand UO_73 (O_73,N_18028,N_18648);
nor UO_74 (O_74,N_17630,N_18347);
or UO_75 (O_75,N_16066,N_18063);
or UO_76 (O_76,N_19288,N_17631);
nor UO_77 (O_77,N_17387,N_18836);
nor UO_78 (O_78,N_16215,N_17479);
and UO_79 (O_79,N_19598,N_16365);
or UO_80 (O_80,N_16421,N_16743);
nor UO_81 (O_81,N_19707,N_17779);
xnor UO_82 (O_82,N_16541,N_16255);
nor UO_83 (O_83,N_17935,N_18152);
nand UO_84 (O_84,N_19929,N_17957);
and UO_85 (O_85,N_19845,N_19858);
nor UO_86 (O_86,N_16647,N_18733);
or UO_87 (O_87,N_16293,N_17660);
nand UO_88 (O_88,N_16906,N_16645);
nand UO_89 (O_89,N_19170,N_17967);
nand UO_90 (O_90,N_17307,N_17512);
and UO_91 (O_91,N_18309,N_19358);
or UO_92 (O_92,N_17766,N_17746);
nor UO_93 (O_93,N_17226,N_18013);
nand UO_94 (O_94,N_16030,N_18054);
and UO_95 (O_95,N_17802,N_17475);
nor UO_96 (O_96,N_18275,N_18789);
nand UO_97 (O_97,N_16847,N_17157);
or UO_98 (O_98,N_19903,N_18955);
and UO_99 (O_99,N_17528,N_18671);
nand UO_100 (O_100,N_16763,N_16484);
and UO_101 (O_101,N_18543,N_19521);
nand UO_102 (O_102,N_19644,N_17296);
and UO_103 (O_103,N_19000,N_16810);
nand UO_104 (O_104,N_18491,N_18195);
nor UO_105 (O_105,N_16655,N_16472);
nor UO_106 (O_106,N_18823,N_17262);
and UO_107 (O_107,N_16976,N_18147);
nand UO_108 (O_108,N_19214,N_17971);
nor UO_109 (O_109,N_17009,N_16188);
or UO_110 (O_110,N_18257,N_18798);
or UO_111 (O_111,N_16542,N_19276);
or UO_112 (O_112,N_18310,N_18230);
or UO_113 (O_113,N_16547,N_18997);
nand UO_114 (O_114,N_18334,N_18482);
nor UO_115 (O_115,N_19452,N_16413);
and UO_116 (O_116,N_19393,N_19950);
nor UO_117 (O_117,N_18353,N_16238);
nor UO_118 (O_118,N_16540,N_16449);
nand UO_119 (O_119,N_19466,N_18048);
nor UO_120 (O_120,N_18285,N_18531);
nor UO_121 (O_121,N_18617,N_18426);
or UO_122 (O_122,N_17683,N_19904);
or UO_123 (O_123,N_17666,N_17743);
nor UO_124 (O_124,N_19427,N_19198);
nor UO_125 (O_125,N_16756,N_17113);
nand UO_126 (O_126,N_18322,N_17370);
or UO_127 (O_127,N_16209,N_17565);
nor UO_128 (O_128,N_18066,N_17039);
nor UO_129 (O_129,N_16428,N_19295);
and UO_130 (O_130,N_19699,N_19142);
nor UO_131 (O_131,N_16782,N_17385);
and UO_132 (O_132,N_18592,N_18663);
nand UO_133 (O_133,N_16612,N_18236);
nand UO_134 (O_134,N_17170,N_19273);
or UO_135 (O_135,N_17592,N_17614);
or UO_136 (O_136,N_17008,N_16137);
nand UO_137 (O_137,N_16550,N_19923);
nand UO_138 (O_138,N_16244,N_16834);
and UO_139 (O_139,N_16523,N_16049);
and UO_140 (O_140,N_19447,N_19077);
nand UO_141 (O_141,N_17278,N_17872);
and UO_142 (O_142,N_16460,N_19404);
nor UO_143 (O_143,N_17289,N_17140);
or UO_144 (O_144,N_16135,N_17827);
nand UO_145 (O_145,N_19918,N_19575);
and UO_146 (O_146,N_17636,N_16916);
nand UO_147 (O_147,N_18866,N_17438);
or UO_148 (O_148,N_19875,N_19949);
nand UO_149 (O_149,N_17798,N_19730);
nor UO_150 (O_150,N_18042,N_18556);
or UO_151 (O_151,N_17996,N_18291);
and UO_152 (O_152,N_16636,N_18511);
xor UO_153 (O_153,N_19675,N_18151);
or UO_154 (O_154,N_17159,N_19134);
or UO_155 (O_155,N_17580,N_17247);
nand UO_156 (O_156,N_19342,N_17514);
nor UO_157 (O_157,N_17190,N_18657);
or UO_158 (O_158,N_18739,N_18465);
or UO_159 (O_159,N_17764,N_16242);
or UO_160 (O_160,N_18969,N_17790);
and UO_161 (O_161,N_16628,N_16200);
or UO_162 (O_162,N_16249,N_16517);
nand UO_163 (O_163,N_19113,N_18442);
or UO_164 (O_164,N_16173,N_17467);
nand UO_165 (O_165,N_16761,N_19121);
or UO_166 (O_166,N_17330,N_16379);
or UO_167 (O_167,N_16603,N_16687);
nor UO_168 (O_168,N_19922,N_18365);
and UO_169 (O_169,N_16462,N_19580);
and UO_170 (O_170,N_16206,N_19017);
and UO_171 (O_171,N_17072,N_16246);
or UO_172 (O_172,N_19764,N_18603);
xnor UO_173 (O_173,N_19488,N_17657);
and UO_174 (O_174,N_19321,N_19453);
or UO_175 (O_175,N_18171,N_17102);
nor UO_176 (O_176,N_16390,N_19628);
nor UO_177 (O_177,N_16548,N_16493);
nor UO_178 (O_178,N_18794,N_16836);
or UO_179 (O_179,N_19979,N_18914);
nor UO_180 (O_180,N_18587,N_16909);
and UO_181 (O_181,N_17193,N_19869);
nand UO_182 (O_182,N_18102,N_18316);
or UO_183 (O_183,N_17044,N_19767);
nand UO_184 (O_184,N_16471,N_17391);
or UO_185 (O_185,N_19531,N_18039);
nor UO_186 (O_186,N_17059,N_19481);
nand UO_187 (O_187,N_17210,N_18877);
and UO_188 (O_188,N_18747,N_18565);
nand UO_189 (O_189,N_19567,N_19822);
or UO_190 (O_190,N_16737,N_18148);
xnor UO_191 (O_191,N_16746,N_19479);
nor UO_192 (O_192,N_19640,N_17122);
nor UO_193 (O_193,N_17322,N_19503);
nor UO_194 (O_194,N_18317,N_19927);
nand UO_195 (O_195,N_16608,N_16869);
nand UO_196 (O_196,N_17856,N_17087);
or UO_197 (O_197,N_18047,N_16168);
nand UO_198 (O_198,N_17914,N_16760);
nand UO_199 (O_199,N_17845,N_19176);
and UO_200 (O_200,N_18486,N_19302);
or UO_201 (O_201,N_16564,N_19805);
nor UO_202 (O_202,N_18443,N_19648);
nor UO_203 (O_203,N_19191,N_17042);
or UO_204 (O_204,N_17842,N_18608);
and UO_205 (O_205,N_18986,N_19464);
nand UO_206 (O_206,N_18600,N_16739);
nor UO_207 (O_207,N_16557,N_19797);
nand UO_208 (O_208,N_19055,N_18264);
and UO_209 (O_209,N_17147,N_16447);
and UO_210 (O_210,N_17369,N_18912);
nand UO_211 (O_211,N_17741,N_16827);
nand UO_212 (O_212,N_18384,N_18566);
nand UO_213 (O_213,N_18176,N_19171);
nand UO_214 (O_214,N_16348,N_17136);
nor UO_215 (O_215,N_18425,N_18643);
nor UO_216 (O_216,N_17498,N_16497);
and UO_217 (O_217,N_17941,N_16654);
nand UO_218 (O_218,N_18835,N_19414);
nor UO_219 (O_219,N_16820,N_18646);
and UO_220 (O_220,N_18072,N_18406);
nand UO_221 (O_221,N_19959,N_18618);
nor UO_222 (O_222,N_19800,N_16940);
nor UO_223 (O_223,N_16361,N_16014);
and UO_224 (O_224,N_19755,N_16527);
nor UO_225 (O_225,N_18819,N_17055);
nand UO_226 (O_226,N_16585,N_18286);
and UO_227 (O_227,N_17586,N_19381);
nand UO_228 (O_228,N_18075,N_16691);
nor UO_229 (O_229,N_19029,N_18050);
nor UO_230 (O_230,N_18175,N_17890);
and UO_231 (O_231,N_19538,N_19131);
nand UO_232 (O_232,N_18161,N_18242);
or UO_233 (O_233,N_17619,N_19265);
and UO_234 (O_234,N_16828,N_16167);
or UO_235 (O_235,N_16230,N_17187);
nor UO_236 (O_236,N_18748,N_17543);
or UO_237 (O_237,N_17846,N_17211);
and UO_238 (O_238,N_17668,N_18266);
nand UO_239 (O_239,N_17000,N_17742);
nand UO_240 (O_240,N_16294,N_19693);
or UO_241 (O_241,N_16424,N_16323);
nand UO_242 (O_242,N_16910,N_19833);
and UO_243 (O_243,N_19743,N_19555);
nor UO_244 (O_244,N_17319,N_18745);
nand UO_245 (O_245,N_18321,N_16485);
nand UO_246 (O_246,N_17001,N_19924);
or UO_247 (O_247,N_18762,N_17598);
and UO_248 (O_248,N_16218,N_19603);
nor UO_249 (O_249,N_16721,N_16035);
nor UO_250 (O_250,N_19011,N_16026);
or UO_251 (O_251,N_18628,N_19401);
nand UO_252 (O_252,N_16849,N_17905);
nor UO_253 (O_253,N_16858,N_16742);
or UO_254 (O_254,N_17973,N_17682);
or UO_255 (O_255,N_19331,N_17976);
and UO_256 (O_256,N_16235,N_16873);
nand UO_257 (O_257,N_18298,N_19704);
nor UO_258 (O_258,N_18934,N_16618);
or UO_259 (O_259,N_18696,N_19849);
or UO_260 (O_260,N_19083,N_19971);
nand UO_261 (O_261,N_16054,N_17333);
or UO_262 (O_262,N_16963,N_19165);
or UO_263 (O_263,N_16699,N_19527);
nand UO_264 (O_264,N_17379,N_17392);
and UO_265 (O_265,N_18729,N_19277);
or UO_266 (O_266,N_17160,N_16772);
nor UO_267 (O_267,N_19721,N_19155);
nor UO_268 (O_268,N_16490,N_18112);
and UO_269 (O_269,N_19554,N_17911);
and UO_270 (O_270,N_17745,N_16016);
and UO_271 (O_271,N_16892,N_19200);
and UO_272 (O_272,N_18031,N_19219);
nand UO_273 (O_273,N_19016,N_17071);
or UO_274 (O_274,N_19036,N_18407);
and UO_275 (O_275,N_17215,N_16749);
and UO_276 (O_276,N_17687,N_17904);
nand UO_277 (O_277,N_19287,N_19574);
and UO_278 (O_278,N_18280,N_18928);
or UO_279 (O_279,N_19596,N_18036);
or UO_280 (O_280,N_17478,N_18207);
nor UO_281 (O_281,N_18668,N_16708);
or UO_282 (O_282,N_16544,N_19749);
or UO_283 (O_283,N_19211,N_17110);
and UO_284 (O_284,N_16444,N_16520);
and UO_285 (O_285,N_18666,N_19551);
nand UO_286 (O_286,N_17046,N_16702);
or UO_287 (O_287,N_19347,N_19156);
nand UO_288 (O_288,N_19478,N_16214);
nor UO_289 (O_289,N_17246,N_17584);
nor UO_290 (O_290,N_16566,N_18272);
or UO_291 (O_291,N_19750,N_16446);
and UO_292 (O_292,N_17133,N_16770);
nor UO_293 (O_293,N_18771,N_17466);
nand UO_294 (O_294,N_17866,N_17026);
nor UO_295 (O_295,N_19543,N_17583);
and UO_296 (O_296,N_17383,N_17639);
or UO_297 (O_297,N_18067,N_19760);
nand UO_298 (O_298,N_19561,N_18698);
or UO_299 (O_299,N_17678,N_17540);
nor UO_300 (O_300,N_18205,N_16689);
or UO_301 (O_301,N_17092,N_18709);
and UO_302 (O_302,N_18640,N_18078);
or UO_303 (O_303,N_16104,N_19966);
nor UO_304 (O_304,N_17198,N_16279);
or UO_305 (O_305,N_18179,N_18623);
and UO_306 (O_306,N_16673,N_17117);
and UO_307 (O_307,N_16656,N_18213);
or UO_308 (O_308,N_17993,N_19152);
nand UO_309 (O_309,N_18740,N_17441);
nand UO_310 (O_310,N_16060,N_16859);
nand UO_311 (O_311,N_16989,N_19172);
or UO_312 (O_312,N_18715,N_19999);
xor UO_313 (O_313,N_19238,N_16939);
nand UO_314 (O_314,N_19089,N_19233);
or UO_315 (O_315,N_16166,N_19565);
nand UO_316 (O_316,N_18597,N_17793);
and UO_317 (O_317,N_17916,N_19197);
or UO_318 (O_318,N_18447,N_19313);
or UO_319 (O_319,N_17068,N_19448);
nor UO_320 (O_320,N_16328,N_17653);
nor UO_321 (O_321,N_16960,N_18956);
and UO_322 (O_322,N_18989,N_17130);
xnor UO_323 (O_323,N_17899,N_18034);
or UO_324 (O_324,N_16437,N_16677);
or UO_325 (O_325,N_16481,N_17393);
nor UO_326 (O_326,N_19043,N_19147);
and UO_327 (O_327,N_16213,N_16394);
nor UO_328 (O_328,N_18826,N_17267);
nand UO_329 (O_329,N_18383,N_16013);
or UO_330 (O_330,N_16052,N_19286);
or UO_331 (O_331,N_19280,N_19117);
and UO_332 (O_332,N_19292,N_17564);
nand UO_333 (O_333,N_17294,N_18742);
and UO_334 (O_334,N_18265,N_18253);
nand UO_335 (O_335,N_17123,N_18009);
and UO_336 (O_336,N_18950,N_16931);
nand UO_337 (O_337,N_16952,N_16871);
and UO_338 (O_338,N_17964,N_17052);
nor UO_339 (O_339,N_17538,N_17406);
or UO_340 (O_340,N_16095,N_17354);
nand UO_341 (O_341,N_17504,N_19973);
and UO_342 (O_342,N_19240,N_19144);
nor UO_343 (O_343,N_17222,N_16046);
and UO_344 (O_344,N_16451,N_16565);
and UO_345 (O_345,N_17633,N_18159);
nor UO_346 (O_346,N_19952,N_18844);
nor UO_347 (O_347,N_19363,N_17548);
and UO_348 (O_348,N_17617,N_19057);
and UO_349 (O_349,N_19780,N_19412);
nand UO_350 (O_350,N_18217,N_16070);
or UO_351 (O_351,N_16253,N_18356);
nor UO_352 (O_352,N_16833,N_18899);
nand UO_353 (O_353,N_16368,N_16041);
and UO_354 (O_354,N_16968,N_18735);
nor UO_355 (O_355,N_18457,N_18341);
nand UO_356 (O_356,N_19119,N_18111);
or UO_357 (O_357,N_16217,N_16672);
nor UO_358 (O_358,N_16690,N_19088);
and UO_359 (O_359,N_18061,N_16105);
or UO_360 (O_360,N_16221,N_19647);
nor UO_361 (O_361,N_18460,N_19824);
and UO_362 (O_362,N_18585,N_17536);
nand UO_363 (O_363,N_19355,N_18182);
nor UO_364 (O_364,N_18708,N_19455);
and UO_365 (O_365,N_16899,N_17344);
and UO_366 (O_366,N_19963,N_18228);
and UO_367 (O_367,N_16767,N_18032);
nor UO_368 (O_368,N_18279,N_16818);
nand UO_369 (O_369,N_18687,N_18086);
or UO_370 (O_370,N_17847,N_18343);
nor UO_371 (O_371,N_19852,N_18029);
or UO_372 (O_372,N_18114,N_19935);
nand UO_373 (O_373,N_19705,N_17304);
nor UO_374 (O_374,N_17231,N_19670);
nor UO_375 (O_375,N_17882,N_18418);
nand UO_376 (O_376,N_17212,N_18252);
nor UO_377 (O_377,N_18725,N_17851);
nor UO_378 (O_378,N_16913,N_18791);
and UO_379 (O_379,N_19524,N_16031);
and UO_380 (O_380,N_16947,N_18021);
and UO_381 (O_381,N_17273,N_16057);
xor UO_382 (O_382,N_18327,N_19851);
and UO_383 (O_383,N_19941,N_16048);
nor UO_384 (O_384,N_18832,N_17883);
and UO_385 (O_385,N_19032,N_16056);
and UO_386 (O_386,N_17950,N_18606);
nand UO_387 (O_387,N_18017,N_17423);
nand UO_388 (O_388,N_16546,N_19847);
and UO_389 (O_389,N_19898,N_19892);
nand UO_390 (O_390,N_17107,N_17820);
nor UO_391 (O_391,N_17365,N_18372);
nand UO_392 (O_392,N_18436,N_16456);
nand UO_393 (O_393,N_19508,N_17956);
nor UO_394 (O_394,N_17195,N_17298);
nor UO_395 (O_395,N_17713,N_18233);
nand UO_396 (O_396,N_18658,N_17709);
or UO_397 (O_397,N_18221,N_19362);
nand UO_398 (O_398,N_16357,N_19774);
or UO_399 (O_399,N_18463,N_16649);
or UO_400 (O_400,N_19862,N_19964);
nor UO_401 (O_401,N_16814,N_19872);
nand UO_402 (O_402,N_19635,N_19977);
nand UO_403 (O_403,N_16304,N_17388);
and UO_404 (O_404,N_16441,N_16103);
nand UO_405 (O_405,N_19799,N_19878);
and UO_406 (O_406,N_19843,N_19808);
or UO_407 (O_407,N_16353,N_17537);
nor UO_408 (O_408,N_18644,N_19190);
or UO_409 (O_409,N_17091,N_19001);
nor UO_410 (O_410,N_19783,N_17208);
and UO_411 (O_411,N_18222,N_16698);
nand UO_412 (O_412,N_16982,N_19469);
nor UO_413 (O_413,N_19166,N_17098);
and UO_414 (O_414,N_17864,N_17038);
nand UO_415 (O_415,N_16538,N_17295);
or UO_416 (O_416,N_17643,N_17237);
or UO_417 (O_417,N_18350,N_16848);
or UO_418 (O_418,N_17989,N_18726);
nand UO_419 (O_419,N_16219,N_16296);
nor UO_420 (O_420,N_18097,N_17754);
nor UO_421 (O_421,N_18216,N_19994);
and UO_422 (O_422,N_19316,N_17016);
or UO_423 (O_423,N_19422,N_18464);
nand UO_424 (O_424,N_18810,N_17185);
and UO_425 (O_425,N_16384,N_18429);
nor UO_426 (O_426,N_18115,N_19650);
nand UO_427 (O_427,N_16904,N_18943);
nand UO_428 (O_428,N_16685,N_16668);
or UO_429 (O_429,N_18790,N_18631);
or UO_430 (O_430,N_19560,N_19739);
nand UO_431 (O_431,N_16400,N_19337);
nand UO_432 (O_432,N_18192,N_16985);
or UO_433 (O_433,N_19687,N_16494);
or UO_434 (O_434,N_19035,N_19992);
nand UO_435 (O_435,N_17378,N_18376);
nor UO_436 (O_436,N_16266,N_16592);
nor UO_437 (O_437,N_16156,N_16452);
or UO_438 (O_438,N_16222,N_16747);
nor UO_439 (O_439,N_17599,N_19821);
and UO_440 (O_440,N_19585,N_16897);
or UO_441 (O_441,N_19046,N_18804);
and UO_442 (O_442,N_17658,N_17638);
nor UO_443 (O_443,N_16912,N_18201);
or UO_444 (O_444,N_18449,N_19418);
nor UO_445 (O_445,N_16777,N_16034);
and UO_446 (O_446,N_16997,N_18226);
nand UO_447 (O_447,N_18753,N_16513);
nor UO_448 (O_448,N_18563,N_18168);
nor UO_449 (O_449,N_17966,N_16040);
nand UO_450 (O_450,N_19435,N_19577);
or UO_451 (O_451,N_19136,N_18968);
nand UO_452 (O_452,N_18038,N_17985);
and UO_453 (O_453,N_19075,N_17721);
and UO_454 (O_454,N_19279,N_16055);
or UO_455 (O_455,N_18288,N_17214);
and UO_456 (O_456,N_19492,N_17917);
or UO_457 (O_457,N_17659,N_16455);
or UO_458 (O_458,N_18417,N_18692);
and UO_459 (O_459,N_17610,N_19626);
nand UO_460 (O_460,N_16559,N_17189);
nor UO_461 (O_461,N_17446,N_18374);
nand UO_462 (O_462,N_17255,N_18076);
nor UO_463 (O_463,N_18554,N_18044);
or UO_464 (O_464,N_16987,N_16796);
nor UO_465 (O_465,N_18604,N_19135);
and UO_466 (O_466,N_17581,N_16694);
nand UO_467 (O_467,N_18331,N_19070);
or UO_468 (O_468,N_17862,N_19221);
or UO_469 (O_469,N_16744,N_17414);
nand UO_470 (O_470,N_16729,N_19763);
and UO_471 (O_471,N_17358,N_16995);
xor UO_472 (O_472,N_19868,N_17080);
nor UO_473 (O_473,N_19052,N_18143);
and UO_474 (O_474,N_18307,N_17250);
nand UO_475 (O_475,N_17332,N_16106);
nor UO_476 (O_476,N_19672,N_19270);
nor UO_477 (O_477,N_19753,N_16583);
or UO_478 (O_478,N_18037,N_16004);
and UO_479 (O_479,N_18688,N_16278);
nand UO_480 (O_480,N_19998,N_16301);
nand UO_481 (O_481,N_16369,N_19223);
nand UO_482 (O_482,N_16377,N_18905);
nor UO_483 (O_483,N_16596,N_16732);
or UO_484 (O_484,N_19110,N_16545);
nand UO_485 (O_485,N_18945,N_18555);
nand UO_486 (O_486,N_18548,N_18420);
nand UO_487 (O_487,N_19968,N_18277);
nor UO_488 (O_488,N_19741,N_17256);
nand UO_489 (O_489,N_16092,N_16844);
nand UO_490 (O_490,N_17735,N_16949);
and UO_491 (O_491,N_19600,N_19366);
or UO_492 (O_492,N_19445,N_18567);
or UO_493 (O_493,N_16574,N_16652);
or UO_494 (O_494,N_18510,N_19622);
nor UO_495 (O_495,N_17532,N_19193);
or UO_496 (O_496,N_18676,N_17323);
and UO_497 (O_497,N_16131,N_19752);
nor UO_498 (O_498,N_16581,N_18396);
nand UO_499 (O_499,N_18453,N_18974);
or UO_500 (O_500,N_16483,N_17232);
or UO_501 (O_501,N_16996,N_17179);
or UO_502 (O_502,N_17539,N_19336);
nand UO_503 (O_503,N_19243,N_16329);
nand UO_504 (O_504,N_18732,N_16374);
or UO_505 (O_505,N_19978,N_18189);
and UO_506 (O_506,N_17421,N_17868);
and UO_507 (O_507,N_18255,N_17591);
and UO_508 (O_508,N_18320,N_17929);
or UO_509 (O_509,N_17127,N_16616);
or UO_510 (O_510,N_19536,N_17576);
and UO_511 (O_511,N_17487,N_18833);
or UO_512 (O_512,N_16686,N_17048);
nand UO_513 (O_513,N_17762,N_19726);
and UO_514 (O_514,N_19607,N_16781);
nand UO_515 (O_515,N_18990,N_17955);
or UO_516 (O_516,N_16161,N_19573);
or UO_517 (O_517,N_16599,N_18413);
and UO_518 (O_518,N_17081,N_16479);
nor UO_519 (O_519,N_16298,N_19060);
or UO_520 (O_520,N_18596,N_18975);
or UO_521 (O_521,N_16395,N_18512);
nand UO_522 (O_522,N_18873,N_16674);
nor UO_523 (O_523,N_16247,N_18952);
nand UO_524 (O_524,N_18158,N_16524);
nand UO_525 (O_525,N_17252,N_16887);
nand UO_526 (O_526,N_16227,N_16389);
and UO_527 (O_527,N_19308,N_18223);
nor UO_528 (O_528,N_19128,N_19397);
or UO_529 (O_529,N_18760,N_18366);
and UO_530 (O_530,N_17166,N_19505);
or UO_531 (O_531,N_18730,N_19244);
or UO_532 (O_532,N_18691,N_16000);
nor UO_533 (O_533,N_17395,N_17535);
nor UO_534 (O_534,N_17715,N_16431);
nand UO_535 (O_535,N_19804,N_16332);
and UO_536 (O_536,N_19151,N_18910);
nand UO_537 (O_537,N_18870,N_16932);
or UO_538 (O_538,N_16558,N_19926);
nor UO_539 (O_539,N_18859,N_18918);
and UO_540 (O_540,N_18935,N_16148);
nand UO_541 (O_541,N_19439,N_16231);
nor UO_542 (O_542,N_18224,N_18843);
nand UO_543 (O_543,N_18766,N_17014);
nand UO_544 (O_544,N_16129,N_18987);
and UO_545 (O_545,N_16570,N_17470);
or UO_546 (O_546,N_19361,N_17748);
or UO_547 (O_547,N_16102,N_17120);
nor UO_548 (O_548,N_18939,N_18141);
or UO_549 (O_549,N_18551,N_18962);
nand UO_550 (O_550,N_18808,N_16267);
or UO_551 (O_551,N_17400,N_19578);
xor UO_552 (O_552,N_19264,N_19974);
and UO_553 (O_553,N_18445,N_18673);
or UO_554 (O_554,N_18202,N_18099);
or UO_555 (O_555,N_18164,N_17213);
nand UO_556 (O_556,N_16713,N_16458);
nor UO_557 (O_557,N_17274,N_18492);
nor UO_558 (O_558,N_18330,N_16514);
nand UO_559 (O_559,N_18414,N_16959);
or UO_560 (O_560,N_19746,N_19127);
or UO_561 (O_561,N_19078,N_18260);
and UO_562 (O_562,N_18476,N_16216);
nand UO_563 (O_563,N_16147,N_18336);
nand UO_564 (O_564,N_18199,N_16277);
and UO_565 (O_565,N_18909,N_19021);
nor UO_566 (O_566,N_17309,N_16276);
or UO_567 (O_567,N_16037,N_16604);
or UO_568 (O_568,N_17151,N_16633);
nor UO_569 (O_569,N_17381,N_19444);
or UO_570 (O_570,N_19993,N_17230);
and UO_571 (O_571,N_18624,N_19251);
or UO_572 (O_572,N_16634,N_18090);
or UO_573 (O_573,N_16920,N_18879);
nor UO_574 (O_574,N_16252,N_17263);
and UO_575 (O_575,N_17338,N_19085);
nor UO_576 (O_576,N_18387,N_17062);
xnor UO_577 (O_577,N_19962,N_18549);
or UO_578 (O_578,N_16181,N_16831);
nor UO_579 (O_579,N_18428,N_18838);
nand UO_580 (O_580,N_19643,N_18981);
nor UO_581 (O_581,N_16184,N_18295);
nand UO_582 (O_582,N_16498,N_19785);
nand UO_583 (O_583,N_16325,N_16631);
nor UO_584 (O_584,N_18024,N_19325);
nand UO_585 (O_585,N_17288,N_17088);
and UO_586 (O_586,N_19689,N_16927);
nand UO_587 (O_587,N_16426,N_17337);
or UO_588 (O_588,N_17472,N_18672);
nand UO_589 (O_589,N_19349,N_19825);
and UO_590 (O_590,N_16011,N_19917);
nor UO_591 (O_591,N_19456,N_16084);
or UO_592 (O_592,N_16127,N_16101);
and UO_593 (O_593,N_17264,N_16577);
and UO_594 (O_594,N_17998,N_18979);
nand UO_595 (O_595,N_19936,N_16640);
nor UO_596 (O_596,N_18964,N_18985);
nor UO_597 (O_597,N_19249,N_17753);
nand UO_598 (O_598,N_17769,N_18390);
or UO_599 (O_599,N_19734,N_16990);
nor UO_600 (O_600,N_16467,N_16984);
and UO_601 (O_601,N_19458,N_16754);
and UO_602 (O_602,N_17836,N_19934);
nor UO_603 (O_603,N_18340,N_18682);
nand UO_604 (O_604,N_16191,N_18232);
nor UO_605 (O_605,N_18058,N_18797);
nor UO_606 (O_606,N_19593,N_18062);
nor UO_607 (O_607,N_16648,N_19987);
nand UO_608 (O_608,N_19946,N_18129);
nand UO_609 (O_609,N_18922,N_16955);
and UO_610 (O_610,N_16282,N_16327);
or UO_611 (O_611,N_17010,N_17169);
nand UO_612 (O_612,N_17066,N_17429);
and UO_613 (O_613,N_17765,N_18104);
xnor UO_614 (O_614,N_18809,N_19681);
nor UO_615 (O_615,N_19039,N_17558);
nor UO_616 (O_616,N_16307,N_19415);
nor UO_617 (O_617,N_17436,N_19235);
nand UO_618 (O_618,N_17622,N_19291);
or UO_619 (O_619,N_19008,N_17997);
and UO_620 (O_620,N_17328,N_16863);
nor UO_621 (O_621,N_19133,N_17757);
nand UO_622 (O_622,N_18538,N_19129);
nand UO_623 (O_623,N_16032,N_17720);
nand UO_624 (O_624,N_19819,N_18088);
and UO_625 (O_625,N_18852,N_18025);
and UO_626 (O_626,N_16409,N_17410);
nand UO_627 (O_627,N_19208,N_17182);
or UO_628 (O_628,N_17690,N_16944);
nor UO_629 (O_629,N_19063,N_19438);
or UO_630 (O_630,N_18364,N_19382);
nor UO_631 (O_631,N_16478,N_17427);
or UO_632 (O_632,N_19476,N_17083);
nor UO_633 (O_633,N_18456,N_19449);
nor UO_634 (O_634,N_16715,N_18720);
or UO_635 (O_635,N_16024,N_18610);
and UO_636 (O_636,N_19972,N_16089);
nand UO_637 (O_637,N_18053,N_19482);
and UO_638 (O_638,N_16270,N_16720);
or UO_639 (O_639,N_17707,N_18145);
nand UO_640 (O_640,N_18612,N_19218);
or UO_641 (O_641,N_19913,N_16607);
and UO_642 (O_642,N_19123,N_18524);
or UO_643 (O_643,N_17838,N_17520);
nor UO_644 (O_644,N_16983,N_17927);
nand UO_645 (O_645,N_18611,N_16948);
and UO_646 (O_646,N_18527,N_17153);
nand UO_647 (O_647,N_18399,N_19697);
nand UO_648 (O_648,N_19920,N_17832);
or UO_649 (O_649,N_19192,N_16532);
nand UO_650 (O_650,N_18860,N_18769);
or UO_651 (O_651,N_19104,N_19161);
xnor UO_652 (O_652,N_19441,N_18686);
nor UO_653 (O_653,N_16802,N_17605);
nor UO_654 (O_654,N_18006,N_17428);
nand UO_655 (O_655,N_18166,N_19111);
nor UO_656 (O_656,N_19766,N_17484);
nor UO_657 (O_657,N_18949,N_17649);
nand UO_658 (O_658,N_17105,N_17749);
and UO_659 (O_659,N_19983,N_18581);
or UO_660 (O_660,N_16176,N_16643);
or UO_661 (O_661,N_19322,N_19654);
or UO_662 (O_662,N_17898,N_18427);
and UO_663 (O_663,N_19541,N_19623);
nand UO_664 (O_664,N_18765,N_16385);
nand UO_665 (O_665,N_17386,N_18533);
nand UO_666 (O_666,N_19056,N_17728);
nor UO_667 (O_667,N_18580,N_18016);
or UO_668 (O_668,N_18522,N_18746);
nand UO_669 (O_669,N_16396,N_16835);
nand UO_670 (O_670,N_17350,N_16438);
nand UO_671 (O_671,N_19827,N_18026);
nand UO_672 (O_672,N_18539,N_17855);
nand UO_673 (O_673,N_17148,N_19034);
nand UO_674 (O_674,N_16232,N_19787);
nor UO_675 (O_675,N_17499,N_19873);
nand UO_676 (O_676,N_18401,N_16164);
and UO_677 (O_677,N_16058,N_18625);
nand UO_678 (O_678,N_17221,N_16254);
nor UO_679 (O_679,N_16100,N_19118);
and UO_680 (O_680,N_16153,N_16516);
xor UO_681 (O_681,N_16028,N_18173);
or UO_682 (O_682,N_17718,N_18571);
or UO_683 (O_683,N_17522,N_18259);
and UO_684 (O_684,N_18530,N_18706);
nor UO_685 (O_685,N_18227,N_17341);
nand UO_686 (O_686,N_16515,N_17518);
nand UO_687 (O_687,N_19633,N_16480);
nor UO_688 (O_688,N_19025,N_16250);
and UO_689 (O_689,N_16891,N_18889);
nor UO_690 (O_690,N_16870,N_19369);
nor UO_691 (O_691,N_16158,N_19586);
nand UO_692 (O_692,N_17612,N_18520);
nand UO_693 (O_693,N_16042,N_17403);
nor UO_694 (O_694,N_16096,N_17821);
or UO_695 (O_695,N_19990,N_17547);
nand UO_696 (O_696,N_17513,N_16440);
and UO_697 (O_697,N_18896,N_19595);
nor UO_698 (O_698,N_18046,N_16531);
or UO_699 (O_699,N_19940,N_17389);
and UO_700 (O_700,N_19283,N_16998);
and UO_701 (O_701,N_19779,N_17106);
and UO_702 (O_702,N_17139,N_17186);
nor UO_703 (O_703,N_17944,N_19153);
and UO_704 (O_704,N_19720,N_19006);
nand UO_705 (O_705,N_17995,N_19744);
or UO_706 (O_706,N_16068,N_19710);
and UO_707 (O_707,N_17575,N_17355);
nand UO_708 (O_708,N_16839,N_18684);
and UO_709 (O_709,N_19801,N_17303);
or UO_710 (O_710,N_17181,N_18466);
xnor UO_711 (O_711,N_18575,N_17837);
nor UO_712 (O_712,N_18982,N_19061);
nor UO_713 (O_713,N_19533,N_17034);
nand UO_714 (O_714,N_19777,N_18160);
nor UO_715 (O_715,N_18290,N_19717);
nand UO_716 (O_716,N_19087,N_17632);
nor UO_717 (O_717,N_16284,N_18422);
and UO_718 (O_718,N_16717,N_18489);
nand UO_719 (O_719,N_16669,N_16539);
and UO_720 (O_720,N_16363,N_16391);
nor UO_721 (O_721,N_17667,N_16179);
nor UO_722 (O_722,N_19703,N_16376);
or UO_723 (O_723,N_16853,N_17590);
nand UO_724 (O_724,N_17542,N_17033);
nor UO_725 (O_725,N_16597,N_18149);
and UO_726 (O_726,N_16956,N_17351);
or UO_727 (O_727,N_16311,N_19005);
and UO_728 (O_728,N_16108,N_17596);
and UO_729 (O_729,N_16350,N_17077);
or UO_730 (O_730,N_17808,N_16468);
nand UO_731 (O_731,N_18313,N_16174);
nor UO_732 (O_732,N_17979,N_17780);
and UO_733 (O_733,N_19157,N_16555);
nand UO_734 (O_734,N_17336,N_16525);
nor UO_735 (O_735,N_18497,N_19301);
nor UO_736 (O_736,N_18319,N_18655);
nor UO_737 (O_737,N_19772,N_16274);
nand UO_738 (O_738,N_19669,N_18867);
nor UO_739 (O_739,N_19677,N_19082);
nor UO_740 (O_740,N_19173,N_19568);
nor UO_741 (O_741,N_18599,N_18978);
nand UO_742 (O_742,N_19379,N_19486);
nor UO_743 (O_743,N_17124,N_17594);
nand UO_744 (O_744,N_17708,N_19108);
or UO_745 (O_745,N_19564,N_17367);
or UO_746 (O_746,N_19947,N_16664);
or UO_747 (O_747,N_17076,N_18281);
or UO_748 (O_748,N_16975,N_17364);
nor UO_749 (O_749,N_19673,N_17946);
or UO_750 (O_750,N_19662,N_16808);
or UO_751 (O_751,N_16787,N_19320);
and UO_752 (O_752,N_19220,N_16022);
and UO_753 (O_753,N_18848,N_18206);
or UO_754 (O_754,N_17047,N_18444);
and UO_755 (O_755,N_18751,N_16336);
or UO_756 (O_756,N_18641,N_18540);
nand UO_757 (O_757,N_18537,N_17178);
or UO_758 (O_758,N_16355,N_19101);
and UO_759 (O_759,N_18096,N_19319);
or UO_760 (O_760,N_18204,N_18887);
nand UO_761 (O_761,N_17141,N_16387);
nand UO_762 (O_762,N_17265,N_19646);
nand UO_763 (O_763,N_16718,N_19409);
and UO_764 (O_764,N_16228,N_16132);
nor UO_765 (O_765,N_16805,N_19013);
nand UO_766 (O_766,N_17290,N_19436);
or UO_767 (O_767,N_17396,N_19740);
and UO_768 (O_768,N_19552,N_17219);
or UO_769 (O_769,N_16050,N_17647);
nand UO_770 (O_770,N_18764,N_17791);
or UO_771 (O_771,N_16338,N_18680);
nand UO_772 (O_772,N_18930,N_16752);
nor UO_773 (O_773,N_16860,N_18513);
and UO_774 (O_774,N_17453,N_18162);
or UO_775 (O_775,N_19899,N_19542);
nor UO_776 (O_776,N_17559,N_18965);
and UO_777 (O_777,N_19098,N_19985);
and UO_778 (O_778,N_19095,N_16418);
nor UO_779 (O_779,N_17480,N_17853);
and UO_780 (O_780,N_19305,N_19548);
or UO_781 (O_781,N_16688,N_19919);
nor UO_782 (O_782,N_16259,N_16627);
nor UO_783 (O_783,N_19257,N_17197);
or UO_784 (O_784,N_17501,N_17380);
and UO_785 (O_785,N_17161,N_19810);
nand UO_786 (O_786,N_18020,N_16018);
nand UO_787 (O_787,N_18659,N_19146);
and UO_788 (O_788,N_16043,N_17960);
and UO_789 (O_789,N_16366,N_18561);
or UO_790 (O_790,N_18452,N_16507);
or UO_791 (O_791,N_19154,N_19189);
or UO_792 (O_792,N_19518,N_18891);
nand UO_793 (O_793,N_17017,N_16302);
nand UO_794 (O_794,N_16878,N_17132);
or UO_795 (O_795,N_17819,N_16008);
or UO_796 (O_796,N_17593,N_18528);
nor UO_797 (O_797,N_17943,N_19645);
nor UO_798 (O_798,N_16519,N_16657);
nor UO_799 (O_799,N_17404,N_18854);
and UO_800 (O_800,N_19250,N_16114);
or UO_801 (O_801,N_19248,N_16261);
and UO_802 (O_802,N_19584,N_18139);
nor UO_803 (O_803,N_17149,N_18328);
and UO_804 (O_804,N_19975,N_18471);
or UO_805 (O_805,N_18736,N_17300);
or UO_806 (O_806,N_19148,N_18582);
and UO_807 (O_807,N_16930,N_17797);
and UO_808 (O_808,N_18231,N_19582);
or UO_809 (O_809,N_18087,N_18363);
nor UO_810 (O_810,N_19205,N_18358);
and UO_811 (O_811,N_17881,N_19483);
or UO_812 (O_812,N_18455,N_17570);
nor UO_813 (O_813,N_19421,N_16629);
nand UO_814 (O_814,N_16710,N_16741);
nor UO_815 (O_815,N_16915,N_18578);
and UO_816 (O_816,N_17411,N_18197);
nand UO_817 (O_817,N_16196,N_16572);
nor UO_818 (O_818,N_16773,N_17248);
or UO_819 (O_819,N_19107,N_16791);
or UO_820 (O_820,N_16033,N_18027);
nor UO_821 (O_821,N_17607,N_17782);
nand UO_822 (O_822,N_16433,N_17618);
nand UO_823 (O_823,N_19776,N_18354);
and UO_824 (O_824,N_19513,N_16371);
and UO_825 (O_825,N_18616,N_18000);
nor UO_826 (O_826,N_17843,N_17937);
and UO_827 (O_827,N_19514,N_16407);
xor UO_828 (O_828,N_19184,N_16412);
and UO_829 (O_829,N_16946,N_16234);
nand UO_830 (O_830,N_16124,N_17419);
nand UO_831 (O_831,N_17019,N_19649);
nand UO_832 (O_832,N_19185,N_19079);
nor UO_833 (O_833,N_17893,N_19365);
nand UO_834 (O_834,N_18738,N_18602);
and UO_835 (O_835,N_18133,N_19932);
xor UO_836 (O_836,N_19890,N_18815);
and UO_837 (O_837,N_18920,N_16047);
nor UO_838 (O_838,N_18109,N_18861);
and UO_839 (O_839,N_19343,N_17902);
nor UO_840 (O_840,N_17486,N_18440);
nor UO_841 (O_841,N_16569,N_18634);
or UO_842 (O_842,N_19086,N_16473);
nand UO_843 (O_843,N_16638,N_17415);
nand UO_844 (O_844,N_16921,N_17529);
and UO_845 (O_845,N_16333,N_16061);
nor UO_846 (O_846,N_17804,N_17865);
nand UO_847 (O_847,N_16408,N_17597);
nor UO_848 (O_848,N_17533,N_18991);
nor UO_849 (O_849,N_19402,N_18718);
or UO_850 (O_850,N_19031,N_17366);
nand UO_851 (O_851,N_16029,N_19125);
or UO_852 (O_852,N_18795,N_18057);
and UO_853 (O_853,N_19446,N_18886);
nor UO_854 (O_854,N_19442,N_16415);
and UO_855 (O_855,N_18924,N_17552);
or UO_856 (O_856,N_16798,N_16258);
nor UO_857 (O_857,N_17236,N_18621);
nor UO_858 (O_858,N_16728,N_17814);
nor UO_859 (O_859,N_19698,N_16679);
nor UO_860 (O_860,N_16149,N_18408);
nand UO_861 (O_861,N_17348,N_16881);
nand UO_862 (O_862,N_16993,N_18296);
nand UO_863 (O_863,N_16120,N_16775);
nand UO_864 (O_864,N_18342,N_17308);
nand UO_865 (O_865,N_18927,N_17489);
and UO_866 (O_866,N_17245,N_18881);
or UO_867 (O_867,N_16895,N_19050);
nand UO_868 (O_868,N_16651,N_16466);
and UO_869 (O_869,N_18636,N_18258);
and UO_870 (O_870,N_16806,N_17340);
and UO_871 (O_871,N_17420,N_16845);
nor UO_872 (O_872,N_17439,N_16207);
and UO_873 (O_873,N_19888,N_16457);
nor UO_874 (O_874,N_17209,N_19451);
and UO_875 (O_875,N_17963,N_19499);
nand UO_876 (O_876,N_18373,N_18690);
and UO_877 (O_877,N_18630,N_19206);
or UO_878 (O_878,N_17803,N_19627);
and UO_879 (O_879,N_17712,N_18778);
nor UO_880 (O_880,N_18071,N_17523);
or UO_881 (O_881,N_19706,N_18136);
or UO_882 (O_882,N_19213,N_18523);
and UO_883 (O_883,N_17870,N_17444);
and UO_884 (O_884,N_18305,N_16454);
nor UO_885 (O_885,N_17430,N_16936);
or UO_886 (O_886,N_18925,N_19341);
nor UO_887 (O_887,N_19690,N_19396);
nor UO_888 (O_888,N_19617,N_17954);
nor UO_889 (O_889,N_18919,N_19641);
or UO_890 (O_890,N_17114,N_17476);
and UO_891 (O_891,N_16724,N_18394);
nand UO_892 (O_892,N_17817,N_16397);
or UO_893 (O_893,N_19954,N_19581);
nand UO_894 (O_894,N_18411,N_19254);
nand UO_895 (O_895,N_18142,N_18271);
or UO_896 (O_896,N_18593,N_16553);
and UO_897 (O_897,N_17624,N_17717);
or UO_898 (O_898,N_19535,N_16109);
and UO_899 (O_899,N_18712,N_16551);
or UO_900 (O_900,N_17752,N_19630);
and UO_901 (O_901,N_19525,N_17061);
nand UO_902 (O_902,N_19266,N_19738);
nand UO_903 (O_903,N_16069,N_18763);
or UO_904 (O_904,N_17488,N_16506);
nand UO_905 (O_905,N_18303,N_16719);
nand UO_906 (O_906,N_16882,N_19986);
and UO_907 (O_907,N_17049,N_19509);
or UO_908 (O_908,N_19084,N_19405);
nand UO_909 (O_909,N_19995,N_18506);
and UO_910 (O_910,N_19081,N_17390);
nand UO_911 (O_911,N_16434,N_18113);
nand UO_912 (O_912,N_16243,N_19140);
nor UO_913 (O_913,N_18404,N_16800);
nor UO_914 (O_914,N_17697,N_16482);
or UO_915 (O_915,N_17377,N_19590);
and UO_916 (O_916,N_16183,N_16194);
and UO_917 (O_917,N_18379,N_16352);
or UO_918 (O_918,N_17795,N_19390);
nor UO_919 (O_919,N_19130,N_16321);
nand UO_920 (O_920,N_17731,N_18839);
nor UO_921 (O_921,N_17751,N_17701);
nor UO_922 (O_922,N_19811,N_17352);
or UO_923 (O_923,N_19387,N_17078);
nand UO_924 (O_924,N_16225,N_17922);
and UO_925 (O_925,N_18505,N_19895);
or UO_926 (O_926,N_18716,N_17880);
nor UO_927 (O_927,N_17942,N_17588);
nand UO_928 (O_928,N_19980,N_17194);
nand UO_929 (O_929,N_18254,N_19834);
or UO_930 (O_930,N_18240,N_17990);
and UO_931 (O_931,N_17435,N_18970);
nand UO_932 (O_932,N_18487,N_16356);
or UO_933 (O_933,N_16119,N_19324);
nor UO_934 (O_934,N_18300,N_18091);
nand UO_935 (O_935,N_16223,N_18882);
and UO_936 (O_936,N_19867,N_19981);
nand UO_937 (O_937,N_18140,N_17977);
nand UO_938 (O_938,N_19258,N_17458);
nor UO_939 (O_939,N_18190,N_18892);
or UO_940 (O_940,N_19522,N_18014);
nor UO_941 (O_941,N_17021,N_18484);
or UO_942 (O_942,N_16241,N_18678);
or UO_943 (O_943,N_16197,N_16141);
or UO_944 (O_944,N_17229,N_19471);
nand UO_945 (O_945,N_17270,N_16723);
or UO_946 (O_946,N_18783,N_16065);
and UO_947 (O_947,N_17202,N_17869);
and UO_948 (O_948,N_16240,N_19761);
or UO_949 (O_949,N_17726,N_18494);
or UO_950 (O_950,N_18126,N_17347);
nor UO_951 (O_951,N_18239,N_16730);
or UO_952 (O_952,N_17402,N_17702);
nand UO_953 (O_953,N_16518,N_18094);
nor UO_954 (O_954,N_18212,N_18817);
nor UO_955 (O_955,N_19806,N_18508);
and UO_956 (O_956,N_17602,N_17553);
and UO_957 (O_957,N_19758,N_16846);
and UO_958 (O_958,N_16053,N_17172);
or UO_959 (O_959,N_17906,N_17648);
or UO_960 (O_960,N_17947,N_18065);
nor UO_961 (O_961,N_18059,N_18845);
and UO_962 (O_962,N_19335,N_16335);
nand UO_963 (O_963,N_18876,N_16704);
and UO_964 (O_964,N_18574,N_19659);
and UO_965 (O_965,N_17646,N_17889);
or UO_966 (O_966,N_16822,N_16879);
and UO_967 (O_967,N_17164,N_16671);
nor UO_968 (O_968,N_16665,N_17756);
or UO_969 (O_969,N_16561,N_16610);
nand UO_970 (O_970,N_16682,N_17655);
xnor UO_971 (O_971,N_17284,N_16594);
nand UO_972 (O_972,N_19866,N_18335);
nor UO_973 (O_973,N_16938,N_16568);
or UO_974 (O_974,N_19771,N_19556);
nand UO_975 (O_975,N_17090,N_16125);
nand UO_976 (O_976,N_17679,N_18570);
or UO_977 (O_977,N_16038,N_19770);
nor UO_978 (O_978,N_16163,N_17999);
or UO_979 (O_979,N_19275,N_16186);
and UO_980 (O_980,N_18885,N_16423);
nand UO_981 (O_981,N_16986,N_19207);
and UO_982 (O_982,N_18633,N_16198);
or UO_983 (O_983,N_19431,N_17065);
nand UO_984 (O_984,N_16023,N_18073);
nand UO_985 (O_985,N_19665,N_17831);
and UO_986 (O_986,N_17654,N_16496);
and UO_987 (O_987,N_19723,N_18814);
and UO_988 (O_988,N_19501,N_17103);
and UO_989 (O_989,N_16399,N_19040);
and UO_990 (O_990,N_18699,N_17778);
nand UO_991 (O_991,N_17987,N_17952);
or UO_992 (O_992,N_16701,N_18082);
and UO_993 (O_993,N_18392,N_16508);
xor UO_994 (O_994,N_18983,N_16642);
and UO_995 (O_995,N_16880,N_19660);
or UO_996 (O_996,N_18514,N_18229);
or UO_997 (O_997,N_17073,N_18834);
and UO_998 (O_998,N_18813,N_17220);
and UO_999 (O_999,N_19880,N_19263);
nor UO_1000 (O_1000,N_18069,N_17623);
or UO_1001 (O_1001,N_16272,N_17541);
or UO_1002 (O_1002,N_18884,N_16961);
nor UO_1003 (O_1003,N_18700,N_18338);
nor UO_1004 (O_1004,N_16417,N_17544);
or UO_1005 (O_1005,N_18403,N_18894);
nand UO_1006 (O_1006,N_18857,N_18329);
or UO_1007 (O_1007,N_16121,N_19850);
nand UO_1008 (O_1008,N_16487,N_18619);
nor UO_1009 (O_1009,N_18770,N_19682);
and UO_1010 (O_1010,N_19367,N_19820);
or UO_1011 (O_1011,N_19709,N_19493);
nor UO_1012 (O_1012,N_19612,N_16410);
and UO_1013 (O_1013,N_17852,N_19559);
nand UO_1014 (O_1014,N_17500,N_19874);
nor UO_1015 (O_1015,N_19472,N_17627);
nand UO_1016 (O_1016,N_16571,N_16098);
nor UO_1017 (O_1017,N_19745,N_17375);
nor UO_1018 (O_1018,N_18409,N_16265);
or UO_1019 (O_1019,N_19228,N_17867);
and UO_1020 (O_1020,N_16420,N_16826);
nor UO_1021 (O_1021,N_18547,N_17432);
or UO_1022 (O_1022,N_18874,N_16591);
nor UO_1023 (O_1023,N_17907,N_17670);
or UO_1024 (O_1024,N_17111,N_18734);
nor UO_1025 (O_1025,N_18806,N_17811);
nand UO_1026 (O_1026,N_16044,N_17261);
nand UO_1027 (O_1027,N_16605,N_19164);
nor UO_1028 (O_1028,N_17885,N_16175);
nand UO_1029 (O_1029,N_18045,N_19430);
nand UO_1030 (O_1030,N_19368,N_19989);
and UO_1031 (O_1031,N_18326,N_19297);
and UO_1032 (O_1032,N_18004,N_19460);
nand UO_1033 (O_1033,N_19828,N_18052);
and UO_1034 (O_1034,N_16007,N_16974);
xor UO_1035 (O_1035,N_18402,N_19686);
nor UO_1036 (O_1036,N_17054,N_16602);
nor UO_1037 (O_1037,N_19395,N_16799);
and UO_1038 (O_1038,N_17125,N_17119);
or UO_1039 (O_1039,N_19030,N_18591);
nand UO_1040 (O_1040,N_19855,N_19814);
nor UO_1041 (O_1041,N_17903,N_19229);
nand UO_1042 (O_1042,N_16981,N_16459);
or UO_1043 (O_1043,N_18639,N_16264);
nand UO_1044 (O_1044,N_18137,N_18723);
or UO_1045 (O_1045,N_19137,N_18665);
nand UO_1046 (O_1046,N_19323,N_19692);
nor UO_1047 (O_1047,N_18685,N_17578);
nand UO_1048 (O_1048,N_17825,N_18490);
nand UO_1049 (O_1049,N_17302,N_18960);
or UO_1050 (O_1050,N_17918,N_18043);
or UO_1051 (O_1051,N_19786,N_18781);
or UO_1052 (O_1052,N_17884,N_16549);
nor UO_1053 (O_1053,N_16122,N_17184);
or UO_1054 (O_1054,N_16381,N_17689);
and UO_1055 (O_1055,N_19328,N_17259);
and UO_1056 (O_1056,N_16663,N_17975);
or UO_1057 (O_1057,N_17988,N_19859);
xnor UO_1058 (O_1058,N_18448,N_19897);
xnor UO_1059 (O_1059,N_16117,N_19732);
nand UO_1060 (O_1060,N_17768,N_17312);
or UO_1061 (O_1061,N_16877,N_18458);
nand UO_1062 (O_1062,N_17258,N_17912);
or UO_1063 (O_1063,N_16589,N_16855);
nand UO_1064 (O_1064,N_17849,N_18163);
nor UO_1065 (O_1065,N_17784,N_17096);
nand UO_1066 (O_1066,N_16872,N_19498);
nor UO_1067 (O_1067,N_16662,N_19604);
nor UO_1068 (O_1068,N_19380,N_19067);
nand UO_1069 (O_1069,N_18651,N_17408);
or UO_1070 (O_1070,N_17785,N_18724);
or UO_1071 (O_1071,N_16697,N_19948);
nor UO_1072 (O_1072,N_16170,N_17279);
nor UO_1073 (O_1073,N_16692,N_19711);
nand UO_1074 (O_1074,N_16988,N_18807);
and UO_1075 (O_1075,N_17551,N_18756);
or UO_1076 (O_1076,N_18799,N_17691);
nand UO_1077 (O_1077,N_16318,N_18780);
nor UO_1078 (O_1078,N_19838,N_17834);
and UO_1079 (O_1079,N_18774,N_17826);
nor UO_1080 (O_1080,N_16926,N_17775);
nand UO_1081 (O_1081,N_19694,N_18667);
nand UO_1082 (O_1082,N_17376,N_17152);
nand UO_1083 (O_1083,N_18134,N_18963);
nand UO_1084 (O_1084,N_18424,N_16632);
and UO_1085 (O_1085,N_18525,N_17306);
or UO_1086 (O_1086,N_17368,N_16445);
nor UO_1087 (O_1087,N_18410,N_19312);
or UO_1088 (O_1088,N_17527,N_16918);
and UO_1089 (O_1089,N_16821,N_18681);
and UO_1090 (O_1090,N_17940,N_18893);
or UO_1091 (O_1091,N_18802,N_19889);
nor UO_1092 (O_1092,N_19212,N_16139);
and UO_1093 (O_1093,N_19685,N_18620);
or UO_1094 (O_1094,N_19066,N_18292);
and UO_1095 (O_1095,N_18454,N_16346);
nand UO_1096 (O_1096,N_18314,N_17732);
and UO_1097 (O_1097,N_19619,N_18131);
and UO_1098 (O_1098,N_16943,N_18060);
nand UO_1099 (O_1099,N_19618,N_19203);
xnor UO_1100 (O_1100,N_18664,N_18901);
or UO_1101 (O_1101,N_19232,N_18958);
nand UO_1102 (O_1102,N_16152,N_19695);
or UO_1103 (O_1103,N_17968,N_17167);
or UO_1104 (O_1104,N_18683,N_18474);
nor UO_1105 (O_1105,N_17425,N_17437);
nor UO_1106 (O_1106,N_17281,N_17962);
nand UO_1107 (O_1107,N_17363,N_16793);
nand UO_1108 (O_1108,N_17074,N_17477);
or UO_1109 (O_1109,N_19976,N_16509);
nand UO_1110 (O_1110,N_16815,N_18416);
or UO_1111 (O_1111,N_18395,N_17445);
and UO_1112 (O_1112,N_19386,N_18711);
or UO_1113 (O_1113,N_17734,N_18423);
nor UO_1114 (O_1114,N_17801,N_19663);
or UO_1115 (O_1115,N_18361,N_19429);
nand UO_1116 (O_1116,N_17027,N_16080);
and UO_1117 (O_1117,N_17095,N_19674);
nor UO_1118 (O_1118,N_16195,N_16644);
and UO_1119 (O_1119,N_18412,N_16187);
nand UO_1120 (O_1120,N_19394,N_19007);
nor UO_1121 (O_1121,N_17253,N_17888);
or UO_1122 (O_1122,N_17449,N_19610);
or UO_1123 (O_1123,N_19237,N_17507);
nand UO_1124 (O_1124,N_17482,N_18613);
nor UO_1125 (O_1125,N_18318,N_17490);
nor UO_1126 (O_1126,N_19902,N_17469);
or UO_1127 (O_1127,N_18389,N_18468);
nand UO_1128 (O_1128,N_18030,N_17050);
and UO_1129 (O_1129,N_18947,N_16020);
xnor UO_1130 (O_1130,N_19356,N_16885);
nor UO_1131 (O_1131,N_19360,N_18614);
or UO_1132 (O_1132,N_19661,N_18493);
and UO_1133 (O_1133,N_16263,N_18352);
and UO_1134 (O_1134,N_19668,N_19225);
or UO_1135 (O_1135,N_19247,N_17492);
or UO_1136 (O_1136,N_17339,N_17025);
nand UO_1137 (O_1137,N_18895,N_18386);
nor UO_1138 (O_1138,N_17524,N_19629);
nand UO_1139 (O_1139,N_18940,N_18519);
nand UO_1140 (O_1140,N_18553,N_16924);
or UO_1141 (O_1141,N_17349,N_17664);
nand UO_1142 (O_1142,N_16192,N_19655);
nand UO_1143 (O_1143,N_19256,N_18101);
and UO_1144 (O_1144,N_18521,N_17154);
nand UO_1145 (O_1145,N_18850,N_19290);
or UO_1146 (O_1146,N_17268,N_18541);
and UO_1147 (O_1147,N_17608,N_19634);
nand UO_1148 (O_1148,N_19158,N_17037);
nor UO_1149 (O_1149,N_18157,N_16958);
nand UO_1150 (O_1150,N_16809,N_18472);
or UO_1151 (O_1151,N_18515,N_17863);
and UO_1152 (O_1152,N_18117,N_17299);
nor UO_1153 (O_1153,N_17958,N_18573);
or UO_1154 (O_1154,N_17799,N_19376);
or UO_1155 (O_1155,N_19434,N_19433);
and UO_1156 (O_1156,N_18459,N_16343);
nand UO_1157 (O_1157,N_17461,N_19303);
nand UO_1158 (O_1158,N_17249,N_17177);
or UO_1159 (O_1159,N_18381,N_16416);
and UO_1160 (O_1160,N_17606,N_19454);
nor UO_1161 (O_1161,N_17431,N_18988);
and UO_1162 (O_1162,N_16758,N_19865);
nor UO_1163 (O_1163,N_16630,N_17063);
and UO_1164 (O_1164,N_17573,N_17013);
or UO_1165 (O_1165,N_17282,N_19684);
nand UO_1166 (O_1166,N_17443,N_18357);
and UO_1167 (O_1167,N_19497,N_16502);
and UO_1168 (O_1168,N_18186,N_18446);
nand UO_1169 (O_1169,N_18064,N_16165);
and UO_1170 (O_1170,N_19735,N_17218);
nor UO_1171 (O_1171,N_16474,N_17491);
nand UO_1172 (O_1172,N_19883,N_18351);
nor UO_1173 (O_1173,N_17813,N_17634);
and UO_1174 (O_1174,N_18480,N_16683);
nand UO_1175 (O_1175,N_17233,N_16962);
nor UO_1176 (O_1176,N_16464,N_16083);
nand UO_1177 (O_1177,N_17982,N_18011);
nor UO_1178 (O_1178,N_18785,N_18098);
and UO_1179 (O_1179,N_16430,N_17244);
nor UO_1180 (O_1180,N_18921,N_16373);
nor UO_1181 (O_1181,N_17318,N_16972);
and UO_1182 (O_1182,N_17601,N_18607);
nand UO_1183 (O_1183,N_19637,N_17830);
nand UO_1184 (O_1184,N_16712,N_16626);
xor UO_1185 (O_1185,N_19407,N_16812);
nand UO_1186 (O_1186,N_17675,N_18103);
xor UO_1187 (O_1187,N_16765,N_19278);
and UO_1188 (O_1188,N_17568,N_19485);
or UO_1189 (O_1189,N_16829,N_16868);
nand UO_1190 (O_1190,N_18405,N_17695);
and UO_1191 (O_1191,N_19982,N_19019);
nor UO_1192 (O_1192,N_16966,N_18105);
and UO_1193 (O_1193,N_17910,N_18432);
or UO_1194 (O_1194,N_17736,N_19911);
and UO_1195 (O_1195,N_18155,N_17604);
and UO_1196 (O_1196,N_17471,N_17525);
and UO_1197 (O_1197,N_16140,N_16143);
and UO_1198 (O_1198,N_17099,N_16189);
and UO_1199 (O_1199,N_19714,N_18961);
nand UO_1200 (O_1200,N_16991,N_16079);
and UO_1201 (O_1201,N_19428,N_17345);
and UO_1202 (O_1202,N_17024,N_18911);
or UO_1203 (O_1203,N_19480,N_18999);
nor UO_1204 (O_1204,N_18559,N_16245);
or UO_1205 (O_1205,N_19318,N_19289);
or UO_1206 (O_1206,N_18360,N_17313);
or UO_1207 (O_1207,N_17729,N_18500);
nand UO_1208 (O_1208,N_19988,N_19271);
nand UO_1209 (O_1209,N_17959,N_19658);
or UO_1210 (O_1210,N_16159,N_19864);
nor UO_1211 (O_1211,N_18994,N_18225);
nor UO_1212 (O_1212,N_19589,N_17418);
or UO_1213 (O_1213,N_17663,N_16439);
nand UO_1214 (O_1214,N_18652,N_16375);
nand UO_1215 (O_1215,N_18863,N_17468);
and UO_1216 (O_1216,N_16714,N_16401);
nand UO_1217 (O_1217,N_18518,N_19372);
and UO_1218 (O_1218,N_16778,N_19099);
nand UO_1219 (O_1219,N_18601,N_18074);
nor UO_1220 (O_1220,N_18243,N_16780);
nor UO_1221 (O_1221,N_17786,N_17145);
nand UO_1222 (O_1222,N_19881,N_19495);
and UO_1223 (O_1223,N_19625,N_18695);
nor UO_1224 (O_1224,N_19352,N_17176);
nor UO_1225 (O_1225,N_18324,N_17104);
nand UO_1226 (O_1226,N_19609,N_17892);
nand UO_1227 (O_1227,N_18598,N_19621);
nand UO_1228 (O_1228,N_17311,N_18437);
nand UO_1229 (O_1229,N_17932,N_17251);
and UO_1230 (O_1230,N_17382,N_19870);
nor UO_1231 (O_1231,N_17495,N_18776);
and UO_1232 (O_1232,N_18200,N_19676);
xnor UO_1233 (O_1233,N_17227,N_18586);
nor UO_1234 (O_1234,N_18752,N_16289);
nand UO_1235 (O_1235,N_18694,N_17562);
nand UO_1236 (O_1236,N_17510,N_19657);
nand UO_1237 (O_1237,N_17018,N_17064);
nor UO_1238 (O_1238,N_18888,N_19796);
and UO_1239 (O_1239,N_18871,N_16950);
and UO_1240 (O_1240,N_18842,N_19440);
nand UO_1241 (O_1241,N_16291,N_17521);
or UO_1242 (O_1242,N_16453,N_19293);
and UO_1243 (O_1243,N_18282,N_18858);
nand UO_1244 (O_1244,N_19072,N_16314);
nor UO_1245 (O_1245,N_19613,N_16536);
and UO_1246 (O_1246,N_16220,N_17991);
or UO_1247 (O_1247,N_19174,N_18713);
or UO_1248 (O_1248,N_17792,N_16378);
nand UO_1249 (O_1249,N_16804,N_16015);
nand UO_1250 (O_1250,N_18677,N_16727);
and UO_1251 (O_1251,N_16486,N_16681);
nand UO_1252 (O_1252,N_19045,N_19159);
nor UO_1253 (O_1253,N_17915,N_16039);
or UO_1254 (O_1254,N_18793,N_16954);
nand UO_1255 (O_1255,N_16992,N_16528);
nand UO_1256 (O_1256,N_16208,N_18068);
and UO_1257 (O_1257,N_19177,N_17275);
nand UO_1258 (O_1258,N_17913,N_19423);
nand UO_1259 (O_1259,N_16239,N_18503);
or UO_1260 (O_1260,N_16347,N_19579);
nand UO_1261 (O_1261,N_18344,N_19572);
or UO_1262 (O_1262,N_18890,N_17763);
nand UO_1263 (O_1263,N_17465,N_17134);
nor UO_1264 (O_1264,N_17454,N_17895);
nor UO_1265 (O_1265,N_17109,N_19884);
nand UO_1266 (O_1266,N_19231,N_19064);
or UO_1267 (O_1267,N_17800,N_17002);
or UO_1268 (O_1268,N_19411,N_17669);
nand UO_1269 (O_1269,N_17891,N_19861);
nor UO_1270 (O_1270,N_17737,N_18297);
nor UO_1271 (O_1271,N_18315,N_16753);
nand UO_1272 (O_1272,N_18023,N_17875);
nand UO_1273 (O_1273,N_17101,N_16299);
nor UO_1274 (O_1274,N_18012,N_16788);
nor UO_1275 (O_1275,N_19300,N_19817);
or UO_1276 (O_1276,N_19239,N_18907);
nand UO_1277 (O_1277,N_18831,N_19384);
or UO_1278 (O_1278,N_16017,N_19093);
and UO_1279 (O_1279,N_19802,N_17401);
nor UO_1280 (O_1280,N_17374,N_16488);
and UO_1281 (O_1281,N_19425,N_19139);
and UO_1282 (O_1282,N_18749,N_19096);
nor UO_1283 (O_1283,N_18092,N_18211);
and UO_1284 (O_1284,N_16320,N_18577);
or UO_1285 (O_1285,N_18782,N_16999);
and UO_1286 (O_1286,N_16852,N_17310);
or UO_1287 (O_1287,N_18367,N_18209);
nor UO_1288 (O_1288,N_17405,N_18238);
nor UO_1289 (O_1289,N_19731,N_17201);
xnor UO_1290 (O_1290,N_17483,N_17953);
or UO_1291 (O_1291,N_19955,N_19733);
and UO_1292 (O_1292,N_17242,N_19553);
xor UO_1293 (O_1293,N_18055,N_18106);
nor UO_1294 (O_1294,N_16469,N_17156);
nand UO_1295 (O_1295,N_17519,N_19751);
nand UO_1296 (O_1296,N_16529,N_16292);
and UO_1297 (O_1297,N_18256,N_17459);
nand UO_1298 (O_1298,N_17146,N_18419);
and UO_1299 (O_1299,N_16862,N_17854);
nor UO_1300 (O_1300,N_17896,N_19832);
nor UO_1301 (O_1301,N_16287,N_17200);
or UO_1302 (O_1302,N_17595,N_18800);
and UO_1303 (O_1303,N_16251,N_19727);
or UO_1304 (O_1304,N_16340,N_18654);
and UO_1305 (O_1305,N_16118,N_19517);
and UO_1306 (O_1306,N_19701,N_16766);
xnor UO_1307 (O_1307,N_18875,N_19842);
and UO_1308 (O_1308,N_18461,N_19591);
nand UO_1309 (O_1309,N_19215,N_17060);
and UO_1310 (O_1310,N_17509,N_18532);
or UO_1311 (O_1311,N_19639,N_17877);
and UO_1312 (O_1312,N_18767,N_17807);
xnor UO_1313 (O_1313,N_18865,N_17696);
nand UO_1314 (O_1314,N_19274,N_18481);
and UO_1315 (O_1315,N_16435,N_17859);
nor UO_1316 (O_1316,N_19653,N_17725);
and UO_1317 (O_1317,N_19281,N_19261);
or UO_1318 (O_1318,N_18188,N_16150);
or UO_1319 (O_1319,N_17930,N_17609);
nand UO_1320 (O_1320,N_18721,N_17360);
and UO_1321 (O_1321,N_16404,N_16620);
or UO_1322 (O_1322,N_18755,N_18467);
nand UO_1323 (O_1323,N_19100,N_17285);
and UO_1324 (O_1324,N_18816,N_16275);
xor UO_1325 (O_1325,N_19122,N_19226);
nand UO_1326 (O_1326,N_17100,N_16646);
nor UO_1327 (O_1327,N_19038,N_19222);
and UO_1328 (O_1328,N_17223,N_17045);
nor UO_1329 (O_1329,N_17260,N_18557);
nor UO_1330 (O_1330,N_16521,N_17496);
or UO_1331 (O_1331,N_16850,N_16088);
nor UO_1332 (O_1332,N_17665,N_19632);
or UO_1333 (O_1333,N_18670,N_17493);
nor UO_1334 (O_1334,N_16650,N_17266);
nand UO_1335 (O_1335,N_19826,N_18936);
or UO_1336 (O_1336,N_19718,N_16002);
or UO_1337 (O_1337,N_17359,N_19528);
and UO_1338 (O_1338,N_17384,N_18193);
nor UO_1339 (O_1339,N_18903,N_18995);
xor UO_1340 (O_1340,N_18469,N_19333);
or UO_1341 (O_1341,N_19332,N_17041);
and UO_1342 (O_1342,N_19359,N_19124);
nor UO_1343 (O_1343,N_18435,N_18773);
and UO_1344 (O_1344,N_18304,N_19126);
nand UO_1345 (O_1345,N_18433,N_16738);
and UO_1346 (O_1346,N_17371,N_18079);
and UO_1347 (O_1347,N_17447,N_17286);
or UO_1348 (O_1348,N_16319,N_19377);
nand UO_1349 (O_1349,N_18946,N_16598);
nor UO_1350 (O_1350,N_18187,N_18653);
nor UO_1351 (O_1351,N_16190,N_16151);
nor UO_1352 (O_1352,N_18430,N_18872);
nand UO_1353 (O_1353,N_18311,N_16823);
nand UO_1354 (O_1354,N_19424,N_17789);
nor UO_1355 (O_1355,N_16450,N_19461);
nand UO_1356 (O_1356,N_17191,N_18089);
and UO_1357 (O_1357,N_18900,N_17116);
nand UO_1358 (O_1358,N_17776,N_16925);
nand UO_1359 (O_1359,N_17781,N_16204);
or UO_1360 (O_1360,N_19296,N_16771);
nor UO_1361 (O_1361,N_18897,N_17271);
nand UO_1362 (O_1362,N_17567,N_18355);
nand UO_1363 (O_1363,N_18015,N_17291);
and UO_1364 (O_1364,N_19419,N_17972);
or UO_1365 (O_1365,N_16505,N_19912);
or UO_1366 (O_1366,N_16146,N_18397);
or UO_1367 (O_1367,N_19051,N_19018);
nand UO_1368 (O_1368,N_19500,N_18529);
nand UO_1369 (O_1369,N_17563,N_19558);
nor UO_1370 (O_1370,N_17920,N_17861);
nand UO_1371 (O_1371,N_17758,N_18825);
nor UO_1372 (O_1372,N_19326,N_19879);
or UO_1373 (O_1373,N_19374,N_18714);
nor UO_1374 (O_1374,N_16199,N_19583);
and UO_1375 (O_1375,N_16706,N_18169);
nand UO_1376 (O_1376,N_17777,N_18041);
and UO_1377 (O_1377,N_18261,N_19848);
and UO_1378 (O_1378,N_16622,N_17788);
nand UO_1379 (O_1379,N_19620,N_19370);
and UO_1380 (O_1380,N_18840,N_18824);
nor UO_1381 (O_1381,N_17485,N_18584);
nor UO_1382 (O_1382,N_19262,N_16326);
and UO_1383 (O_1383,N_17680,N_18208);
nor UO_1384 (O_1384,N_16075,N_18637);
or UO_1385 (O_1385,N_16463,N_17334);
nor UO_1386 (O_1386,N_17970,N_18703);
xor UO_1387 (O_1387,N_19914,N_18977);
or UO_1388 (O_1388,N_17625,N_16819);
and UO_1389 (O_1389,N_18674,N_18132);
nor UO_1390 (O_1390,N_16840,N_16977);
or UO_1391 (O_1391,N_19299,N_18786);
or UO_1392 (O_1392,N_17129,N_16637);
nor UO_1393 (O_1393,N_16372,N_17407);
xnor UO_1394 (O_1394,N_16308,N_18542);
or UO_1395 (O_1395,N_17481,N_19102);
xnor UO_1396 (O_1396,N_17934,N_17645);
nand UO_1397 (O_1397,N_19562,N_19511);
nor UO_1398 (O_1398,N_18796,N_19537);
nand UO_1399 (O_1399,N_17948,N_19906);
and UO_1400 (O_1400,N_16951,N_16824);
and UO_1401 (O_1401,N_17874,N_17457);
or UO_1402 (O_1402,N_17901,N_19762);
nand UO_1403 (O_1403,N_18156,N_19150);
or UO_1404 (O_1404,N_18550,N_18908);
nand UO_1405 (O_1405,N_19942,N_16874);
xor UO_1406 (O_1406,N_16367,N_18267);
nor UO_1407 (O_1407,N_16382,N_16889);
or UO_1408 (O_1408,N_17992,N_16660);
and UO_1409 (O_1409,N_19765,N_19953);
or UO_1410 (O_1410,N_18110,N_18849);
nor UO_1411 (O_1411,N_17069,N_17331);
and UO_1412 (O_1412,N_18479,N_19058);
nor UO_1413 (O_1413,N_19651,N_18121);
nor UO_1414 (O_1414,N_17860,N_17566);
nand UO_1415 (O_1415,N_16162,N_17030);
nand UO_1416 (O_1416,N_19143,N_18821);
or UO_1417 (O_1417,N_16059,N_19163);
and UO_1418 (O_1418,N_17283,N_18772);
and UO_1419 (O_1419,N_19457,N_16969);
nor UO_1420 (O_1420,N_18244,N_18880);
and UO_1421 (O_1421,N_18526,N_18722);
and UO_1422 (O_1422,N_18153,N_17269);
or UO_1423 (O_1423,N_19410,N_19930);
nand UO_1424 (O_1424,N_18274,N_16757);
or UO_1425 (O_1425,N_17494,N_17057);
nor UO_1426 (O_1426,N_17876,N_17006);
and UO_1427 (O_1427,N_16448,N_16025);
or UO_1428 (O_1428,N_16971,N_17585);
nand UO_1429 (O_1429,N_16160,N_17508);
or UO_1430 (O_1430,N_16731,N_16893);
or UO_1431 (O_1431,N_17362,N_19683);
nand UO_1432 (O_1432,N_18146,N_18906);
and UO_1433 (O_1433,N_16888,N_16593);
and UO_1434 (O_1434,N_16784,N_19080);
or UO_1435 (O_1435,N_18944,N_16624);
nand UO_1436 (O_1436,N_17239,N_19636);
nor UO_1437 (O_1437,N_18827,N_17806);
nand UO_1438 (O_1438,N_18393,N_16864);
and UO_1439 (O_1439,N_16785,N_16288);
or UO_1440 (O_1440,N_19747,N_17204);
nand UO_1441 (O_1441,N_18325,N_19241);
and UO_1442 (O_1442,N_18629,N_18473);
or UO_1443 (O_1443,N_19074,N_18251);
and UO_1444 (O_1444,N_18118,N_17878);
nor UO_1445 (O_1445,N_19945,N_16967);
nand UO_1446 (O_1446,N_17463,N_19068);
and UO_1447 (O_1447,N_16269,N_16262);
and UO_1448 (O_1448,N_17324,N_16476);
or UO_1449 (O_1449,N_17613,N_19961);
nand UO_1450 (O_1450,N_17277,N_16584);
and UO_1451 (O_1451,N_18784,N_16705);
and UO_1452 (O_1452,N_18496,N_16734);
nand UO_1453 (O_1453,N_19187,N_19631);
nand UO_1454 (O_1454,N_17085,N_17939);
nor UO_1455 (O_1455,N_16816,N_16894);
nand UO_1456 (O_1456,N_17662,N_17144);
and UO_1457 (O_1457,N_18662,N_17550);
nor UO_1458 (O_1458,N_16062,N_19002);
nor UO_1459 (O_1459,N_18116,N_17216);
nor UO_1460 (O_1460,N_18246,N_18996);
nor UO_1461 (O_1461,N_18184,N_19815);
or UO_1462 (O_1462,N_17651,N_19268);
or UO_1463 (O_1463,N_18841,N_16902);
and UO_1464 (O_1464,N_19778,N_19015);
nor UO_1465 (O_1465,N_16567,N_18108);
nand UO_1466 (O_1466,N_16345,N_16510);
nand UO_1467 (O_1467,N_16491,N_19901);
nand UO_1468 (O_1468,N_19951,N_17969);
nor UO_1469 (O_1469,N_17199,N_17131);
or UO_1470 (O_1470,N_18485,N_18385);
nand UO_1471 (O_1471,N_19491,N_17398);
or UO_1472 (O_1472,N_17412,N_17399);
nor UO_1473 (O_1473,N_16283,N_19391);
or UO_1474 (O_1474,N_16429,N_16861);
nor UO_1475 (O_1475,N_16994,N_18339);
nand UO_1476 (O_1476,N_18830,N_17205);
nor UO_1477 (O_1477,N_17727,N_17422);
and UO_1478 (O_1478,N_19742,N_16383);
and UO_1479 (O_1479,N_19856,N_19775);
nand UO_1480 (O_1480,N_19540,N_17023);
or UO_1481 (O_1481,N_19437,N_19202);
nor UO_1482 (O_1482,N_19385,N_17450);
or UO_1483 (O_1483,N_16006,N_18822);
nand UO_1484 (O_1484,N_16680,N_16945);
and UO_1485 (O_1485,N_16586,N_16937);
and UO_1486 (O_1486,N_19294,N_19700);
or UO_1487 (O_1487,N_18967,N_18308);
nand UO_1488 (O_1488,N_19071,N_19716);
nand UO_1489 (O_1489,N_19614,N_17028);
or UO_1490 (O_1490,N_19022,N_19162);
nor UO_1491 (O_1491,N_16475,N_18154);
nor UO_1492 (O_1492,N_19310,N_17635);
nand UO_1493 (O_1493,N_18362,N_17965);
and UO_1494 (O_1494,N_16370,N_19928);
nor UO_1495 (O_1495,N_16380,N_17572);
and UO_1496 (O_1496,N_19757,N_19931);
and UO_1497 (O_1497,N_16133,N_19656);
nand UO_1498 (O_1498,N_18100,N_17346);
and UO_1499 (O_1499,N_19069,N_16842);
or UO_1500 (O_1500,N_16843,N_19576);
or UO_1501 (O_1501,N_18203,N_19885);
and UO_1502 (O_1502,N_16562,N_16260);
nor UO_1503 (O_1503,N_16639,N_17945);
nor UO_1504 (O_1504,N_19120,N_19304);
nand UO_1505 (O_1505,N_19378,N_18470);
and UO_1506 (O_1506,N_19795,N_17043);
nor UO_1507 (O_1507,N_17900,N_17629);
nor UO_1508 (O_1508,N_17093,N_16979);
or UO_1509 (O_1509,N_17203,N_16145);
nor UO_1510 (O_1510,N_16112,N_17086);
or UO_1511 (O_1511,N_16492,N_17320);
or UO_1512 (O_1512,N_16224,N_17356);
and UO_1513 (O_1513,N_19028,N_16768);
or UO_1514 (O_1514,N_19330,N_18421);
nor UO_1515 (O_1515,N_18980,N_18181);
nor UO_1516 (O_1516,N_19245,N_16113);
and UO_1517 (O_1517,N_19894,N_16837);
and UO_1518 (O_1518,N_16832,N_17672);
and UO_1519 (O_1519,N_17206,N_19702);
nor UO_1520 (O_1520,N_19781,N_16534);
or UO_1521 (O_1521,N_17526,N_19196);
nand UO_1522 (O_1522,N_19991,N_17394);
or UO_1523 (O_1523,N_19389,N_18263);
nand UO_1524 (O_1524,N_16297,N_16443);
nor UO_1525 (O_1525,N_18284,N_16436);
or UO_1526 (O_1526,N_18003,N_17115);
nor UO_1527 (O_1527,N_17926,N_19059);
or UO_1528 (O_1528,N_16178,N_19199);
nand UO_1529 (O_1529,N_19754,N_19520);
nor UO_1530 (O_1530,N_17505,N_17022);
and UO_1531 (O_1531,N_16776,N_17772);
or UO_1532 (O_1532,N_18546,N_17739);
and UO_1533 (O_1533,N_18937,N_16406);
or UO_1534 (O_1534,N_19638,N_19925);
or UO_1535 (O_1535,N_17809,N_16142);
nand UO_1536 (O_1536,N_19309,N_16271);
and UO_1537 (O_1537,N_18183,N_18669);
and UO_1538 (O_1538,N_18938,N_19194);
and UO_1539 (O_1539,N_17238,N_16533);
or UO_1540 (O_1540,N_17600,N_16211);
nor UO_1541 (O_1541,N_19091,N_18093);
or UO_1542 (O_1542,N_18971,N_18177);
nand UO_1543 (O_1543,N_16317,N_17142);
and UO_1544 (O_1544,N_16402,N_16623);
nand UO_1545 (O_1545,N_16354,N_16779);
nor UO_1546 (O_1546,N_17036,N_17555);
nand UO_1547 (O_1547,N_18002,N_17243);
and UO_1548 (O_1548,N_17174,N_17089);
nand UO_1549 (O_1549,N_17056,N_19062);
or UO_1550 (O_1550,N_16774,N_18400);
nor UO_1551 (O_1551,N_18033,N_18215);
or UO_1552 (O_1552,N_19601,N_18898);
nand UO_1553 (O_1553,N_17112,N_19490);
nor UO_1554 (O_1554,N_18642,N_17835);
or UO_1555 (O_1555,N_17257,N_18931);
or UO_1556 (O_1556,N_17426,N_18594);
nor UO_1557 (O_1557,N_17440,N_19132);
nor UO_1558 (O_1558,N_19216,N_19969);
and UO_1559 (O_1559,N_17225,N_16898);
and UO_1560 (O_1560,N_18847,N_16973);
or UO_1561 (O_1561,N_17722,N_19519);
nor UO_1562 (O_1562,N_19587,N_16134);
or UO_1563 (O_1563,N_17673,N_17188);
or UO_1564 (O_1564,N_16073,N_17029);
nor UO_1565 (O_1565,N_18235,N_19484);
or UO_1566 (O_1566,N_19532,N_18679);
or UO_1567 (O_1567,N_16003,N_18380);
and UO_1568 (O_1568,N_17700,N_18779);
and UO_1569 (O_1569,N_19354,N_17325);
or UO_1570 (O_1570,N_16411,N_19967);
and UO_1571 (O_1571,N_17719,N_18590);
nand UO_1572 (O_1572,N_16759,N_16477);
and UO_1573 (O_1573,N_17035,N_18144);
nand UO_1574 (O_1574,N_19713,N_19526);
or UO_1575 (O_1575,N_19807,N_18083);
and UO_1576 (O_1576,N_16522,N_18862);
nand UO_1577 (O_1577,N_19688,N_19462);
nand UO_1578 (O_1578,N_16576,N_19759);
or UO_1579 (O_1579,N_19041,N_17343);
or UO_1580 (O_1580,N_18247,N_16903);
nor UO_1581 (O_1581,N_18787,N_17812);
or UO_1582 (O_1582,N_18301,N_17983);
and UO_1583 (O_1583,N_18788,N_18761);
nor UO_1584 (O_1584,N_19049,N_19255);
or UO_1585 (O_1585,N_19791,N_19965);
and UO_1586 (O_1586,N_17314,N_16580);
nand UO_1587 (O_1587,N_16619,N_16185);
nor UO_1588 (O_1588,N_18777,N_16501);
and UO_1589 (O_1589,N_19236,N_19680);
and UO_1590 (O_1590,N_16362,N_19782);
or UO_1591 (O_1591,N_16601,N_18661);
nor UO_1592 (O_1592,N_18507,N_18846);
nand UO_1593 (O_1593,N_17361,N_19012);
and UO_1594 (O_1594,N_16813,N_17569);
nand UO_1595 (O_1595,N_19516,N_17829);
and UO_1596 (O_1596,N_17684,N_16144);
and UO_1597 (O_1597,N_16923,N_17511);
nand UO_1598 (O_1598,N_19037,N_16005);
or UO_1599 (O_1599,N_17497,N_16177);
and UO_1600 (O_1600,N_17207,N_18450);
or UO_1601 (O_1601,N_18727,N_17857);
nand UO_1602 (O_1602,N_19413,N_17783);
nand UO_1603 (O_1603,N_19033,N_18993);
nand UO_1604 (O_1604,N_18864,N_16670);
xnor UO_1605 (O_1605,N_16803,N_19510);
nor UO_1606 (O_1606,N_18589,N_18951);
and UO_1607 (O_1607,N_19876,N_19443);
xor UO_1608 (O_1608,N_18710,N_16919);
nor UO_1609 (O_1609,N_19282,N_16341);
nand UO_1610 (O_1610,N_18306,N_18517);
and UO_1611 (O_1611,N_17315,N_16229);
nor UO_1612 (O_1612,N_19539,N_18007);
and UO_1613 (O_1613,N_16543,N_19835);
and UO_1614 (O_1614,N_18346,N_19348);
nor UO_1615 (O_1615,N_16201,N_16322);
or UO_1616 (O_1616,N_17162,N_17240);
nor UO_1617 (O_1617,N_17652,N_16427);
or UO_1618 (O_1618,N_16358,N_18948);
or UO_1619 (O_1619,N_16838,N_17409);
nand UO_1620 (O_1620,N_16716,N_17925);
or UO_1621 (O_1621,N_19943,N_17887);
or UO_1622 (O_1622,N_16856,N_17372);
nor UO_1623 (O_1623,N_17079,N_18431);
and UO_1624 (O_1624,N_18754,N_18180);
or UO_1625 (O_1625,N_17534,N_18851);
nand UO_1626 (O_1626,N_17007,N_16935);
nor UO_1627 (O_1627,N_16884,N_18501);
or UO_1628 (O_1628,N_18382,N_17158);
nand UO_1629 (O_1629,N_19338,N_18135);
nor UO_1630 (O_1630,N_18534,N_17373);
or UO_1631 (O_1631,N_16790,N_17589);
nand UO_1632 (O_1632,N_16465,N_16324);
nand UO_1633 (O_1633,N_18818,N_19473);
and UO_1634 (O_1634,N_16313,N_16582);
nand UO_1635 (O_1635,N_18249,N_16285);
or UO_1636 (O_1636,N_16554,N_16764);
or UO_1637 (O_1637,N_18913,N_18707);
nor UO_1638 (O_1638,N_16045,N_19284);
nor UO_1639 (O_1639,N_17711,N_19506);
nand UO_1640 (O_1640,N_17824,N_19691);
nand UO_1641 (O_1641,N_19958,N_17755);
or UO_1642 (O_1642,N_16865,N_17473);
nor UO_1643 (O_1643,N_17760,N_16107);
or UO_1644 (O_1644,N_19515,N_17560);
or UO_1645 (O_1645,N_18299,N_19399);
nand UO_1646 (O_1646,N_18245,N_18312);
nor UO_1647 (O_1647,N_17723,N_18294);
and UO_1648 (O_1648,N_19097,N_18174);
and UO_1649 (O_1649,N_17961,N_16203);
and UO_1650 (O_1650,N_18792,N_19667);
nand UO_1651 (O_1651,N_18635,N_16635);
nand UO_1652 (O_1652,N_19599,N_18056);
nor UO_1653 (O_1653,N_16653,N_16316);
nor UO_1654 (O_1654,N_17706,N_18923);
or UO_1655 (O_1655,N_19788,N_18504);
nand UO_1656 (O_1656,N_16941,N_16736);
nand UO_1657 (O_1657,N_18237,N_17603);
and UO_1658 (O_1658,N_19114,N_17699);
and UO_1659 (O_1659,N_16312,N_19044);
nor UO_1660 (O_1660,N_18095,N_19530);
nand UO_1661 (O_1661,N_17744,N_18130);
nand UO_1662 (O_1662,N_16613,N_19267);
or UO_1663 (O_1663,N_19314,N_18289);
nor UO_1664 (O_1664,N_19597,N_18609);
nand UO_1665 (O_1665,N_17327,N_18853);
and UO_1666 (O_1666,N_16067,N_19209);
or UO_1667 (O_1667,N_17357,N_19615);
nor UO_1668 (O_1668,N_19307,N_16750);
nor UO_1669 (O_1669,N_16556,N_16248);
nand UO_1670 (O_1670,N_16914,N_18302);
and UO_1671 (O_1671,N_18693,N_18564);
nor UO_1672 (O_1672,N_18478,N_16666);
nor UO_1673 (O_1673,N_16755,N_17650);
nand UO_1674 (O_1674,N_19938,N_18829);
or UO_1675 (O_1675,N_17640,N_18705);
and UO_1676 (O_1676,N_16575,N_18250);
nor UO_1677 (O_1677,N_17909,N_19487);
nor UO_1678 (O_1678,N_17321,N_16099);
or UO_1679 (O_1679,N_17858,N_19329);
and UO_1680 (O_1680,N_19939,N_16537);
and UO_1681 (O_1681,N_19306,N_18536);
or UO_1682 (O_1682,N_17531,N_17703);
or UO_1683 (O_1683,N_19094,N_16091);
and UO_1684 (O_1684,N_18349,N_16360);
nor UO_1685 (O_1685,N_18622,N_19813);
and UO_1686 (O_1686,N_18803,N_19315);
nand UO_1687 (O_1687,N_19846,N_18869);
or UO_1688 (O_1688,N_17611,N_19724);
nand UO_1689 (O_1689,N_16659,N_17951);
nor UO_1690 (O_1690,N_16138,N_17698);
nor UO_1691 (O_1691,N_16128,N_17456);
and UO_1692 (O_1692,N_19204,N_17873);
and UO_1693 (O_1693,N_18915,N_19195);
and UO_1694 (O_1694,N_18010,N_17171);
or UO_1695 (O_1695,N_17844,N_18495);
and UO_1696 (O_1696,N_18579,N_18731);
and UO_1697 (O_1697,N_19854,N_19984);
and UO_1698 (O_1698,N_18287,N_19259);
or UO_1699 (O_1699,N_17986,N_16364);
and UO_1700 (O_1700,N_16600,N_18502);
nand UO_1701 (O_1701,N_18124,N_17128);
nor UO_1702 (O_1702,N_18572,N_19470);
or UO_1703 (O_1703,N_17416,N_19569);
and UO_1704 (O_1704,N_17012,N_19970);
nand UO_1705 (O_1705,N_16700,N_17773);
nand UO_1706 (O_1706,N_17067,N_19857);
or UO_1707 (O_1707,N_17058,N_16130);
or UO_1708 (O_1708,N_18576,N_16076);
nand UO_1709 (O_1709,N_16392,N_17329);
nand UO_1710 (O_1710,N_18323,N_16615);
nand UO_1711 (O_1711,N_16442,N_18370);
and UO_1712 (O_1712,N_19729,N_19406);
nand UO_1713 (O_1713,N_16315,N_18167);
nand UO_1714 (O_1714,N_17234,N_16281);
or UO_1715 (O_1715,N_17674,N_16172);
and UO_1716 (O_1716,N_19863,N_18441);
or UO_1717 (O_1717,N_18019,N_19468);
nor UO_1718 (O_1718,N_19840,N_17840);
and UO_1719 (O_1719,N_19252,N_16349);
nand UO_1720 (O_1720,N_17301,N_17241);
nand UO_1721 (O_1721,N_16414,N_16964);
nand UO_1722 (O_1722,N_18984,N_18902);
nand UO_1723 (O_1723,N_16425,N_18728);
or UO_1724 (O_1724,N_17342,N_16875);
nor UO_1725 (O_1725,N_17335,N_16419);
and UO_1726 (O_1726,N_16595,N_17805);
nor UO_1727 (O_1727,N_16535,N_19512);
or UO_1728 (O_1728,N_19115,N_18775);
nand UO_1729 (O_1729,N_17685,N_16733);
nand UO_1730 (O_1730,N_18954,N_16280);
nand UO_1731 (O_1731,N_19416,N_18837);
nand UO_1732 (O_1732,N_17517,N_17442);
and UO_1733 (O_1733,N_19809,N_17150);
and UO_1734 (O_1734,N_19141,N_17787);
and UO_1735 (O_1735,N_18001,N_17175);
or UO_1736 (O_1736,N_19792,N_18856);
and UO_1737 (O_1737,N_16667,N_19909);
or UO_1738 (O_1738,N_16386,N_16036);
nand UO_1739 (O_1739,N_17919,N_17546);
nor UO_1740 (O_1740,N_17841,N_18345);
nand UO_1741 (O_1741,N_16290,N_19594);
or UO_1742 (O_1742,N_17316,N_16676);
nor UO_1743 (O_1743,N_17897,N_19260);
xnor UO_1744 (O_1744,N_17693,N_16205);
and UO_1745 (O_1745,N_17287,N_19053);
xor UO_1746 (O_1746,N_17637,N_18929);
or UO_1747 (O_1747,N_17681,N_16851);
nand UO_1748 (O_1748,N_19803,N_19900);
nand UO_1749 (O_1749,N_18941,N_18388);
and UO_1750 (O_1750,N_18293,N_19090);
and UO_1751 (O_1751,N_17850,N_18198);
nor UO_1752 (O_1752,N_19736,N_17908);
nor UO_1753 (O_1753,N_16210,N_18689);
nor UO_1754 (O_1754,N_18332,N_16495);
nor UO_1755 (O_1755,N_17738,N_19224);
nor UO_1756 (O_1756,N_18049,N_19298);
or UO_1757 (O_1757,N_19907,N_18660);
nor UO_1758 (O_1758,N_17506,N_16857);
or UO_1759 (O_1759,N_18348,N_16922);
and UO_1760 (O_1760,N_17173,N_18656);
and UO_1761 (O_1761,N_19841,N_17276);
nor UO_1762 (O_1762,N_18196,N_17761);
nor UO_1763 (O_1763,N_16405,N_19181);
nand UO_1764 (O_1764,N_16115,N_19944);
or UO_1765 (O_1765,N_16890,N_16303);
and UO_1766 (O_1766,N_16588,N_18701);
and UO_1767 (O_1767,N_19784,N_16917);
nand UO_1768 (O_1768,N_18248,N_17108);
nand UO_1769 (O_1769,N_18992,N_19375);
nor UO_1770 (O_1770,N_19494,N_19549);
or UO_1771 (O_1771,N_16500,N_17126);
and UO_1772 (O_1772,N_19106,N_17978);
nand UO_1773 (O_1773,N_19719,N_16678);
or UO_1774 (O_1774,N_18276,N_19334);
and UO_1775 (O_1775,N_16193,N_18234);
or UO_1776 (O_1776,N_19790,N_16236);
nand UO_1777 (O_1777,N_17747,N_19180);
nand UO_1778 (O_1778,N_19230,N_16422);
nand UO_1779 (O_1779,N_19463,N_18080);
or UO_1780 (O_1780,N_16295,N_19773);
nor UO_1781 (O_1781,N_17305,N_16110);
and UO_1782 (O_1782,N_16063,N_17839);
or UO_1783 (O_1783,N_17516,N_16339);
nor UO_1784 (O_1784,N_19465,N_16009);
and UO_1785 (O_1785,N_17075,N_18172);
nand UO_1786 (O_1786,N_16330,N_19725);
nor UO_1787 (O_1787,N_17121,N_16019);
nor UO_1788 (O_1788,N_17082,N_19475);
and UO_1789 (O_1789,N_18368,N_17818);
nand UO_1790 (O_1790,N_19496,N_17317);
nor UO_1791 (O_1791,N_18498,N_16658);
nor UO_1792 (O_1792,N_19065,N_19523);
or UO_1793 (O_1793,N_19246,N_19253);
and UO_1794 (O_1794,N_17936,N_18283);
or UO_1795 (O_1795,N_18070,N_17894);
or UO_1796 (O_1796,N_16609,N_17556);
or UO_1797 (O_1797,N_19186,N_17676);
nor UO_1798 (O_1798,N_17455,N_18499);
or UO_1799 (O_1799,N_18926,N_16087);
nor UO_1800 (O_1800,N_17353,N_16393);
and UO_1801 (O_1801,N_17015,N_16082);
and UO_1802 (O_1802,N_19477,N_19003);
or UO_1803 (O_1803,N_19227,N_17180);
nand UO_1804 (O_1804,N_17053,N_19507);
nor UO_1805 (O_1805,N_17871,N_18632);
nor UO_1806 (O_1806,N_16300,N_18219);
nor UO_1807 (O_1807,N_18022,N_19546);
nand UO_1808 (O_1808,N_18220,N_18150);
and UO_1809 (O_1809,N_19179,N_19054);
nor UO_1810 (O_1810,N_19149,N_16703);
or UO_1811 (O_1811,N_19588,N_17192);
nor UO_1812 (O_1812,N_18878,N_16077);
and UO_1813 (O_1813,N_17767,N_19608);
and UO_1814 (O_1814,N_17974,N_19183);
nand UO_1815 (O_1815,N_17451,N_16511);
nor UO_1816 (O_1816,N_18051,N_17503);
or UO_1817 (O_1817,N_18462,N_17561);
nor UO_1818 (O_1818,N_18717,N_17094);
nand UO_1819 (O_1819,N_17621,N_19616);
nand UO_1820 (O_1820,N_18369,N_17397);
or UO_1821 (O_1821,N_18645,N_19371);
nor UO_1822 (O_1822,N_18084,N_19167);
nor UO_1823 (O_1823,N_18959,N_19234);
and UO_1824 (O_1824,N_18165,N_17661);
nor UO_1825 (O_1825,N_17433,N_17545);
or UO_1826 (O_1826,N_17714,N_16908);
and UO_1827 (O_1827,N_18185,N_19996);
nor UO_1828 (O_1828,N_18558,N_16911);
nor UO_1829 (O_1829,N_16886,N_16794);
nor UO_1830 (O_1830,N_19905,N_16711);
nand UO_1831 (O_1831,N_17137,N_16841);
nand UO_1832 (O_1832,N_17557,N_19138);
nor UO_1833 (O_1833,N_19400,N_16725);
or UO_1834 (O_1834,N_16901,N_16830);
nor UO_1835 (O_1835,N_18077,N_16526);
or UO_1836 (O_1836,N_19910,N_19957);
nor UO_1837 (O_1837,N_19816,N_18214);
and UO_1838 (O_1838,N_17794,N_16560);
nand UO_1839 (O_1839,N_18627,N_16123);
nor UO_1840 (O_1840,N_17823,N_18545);
or UO_1841 (O_1841,N_16499,N_19696);
and UO_1842 (O_1842,N_18535,N_19340);
nor UO_1843 (O_1843,N_19545,N_16745);
nor UO_1844 (O_1844,N_16064,N_19426);
nor UO_1845 (O_1845,N_17293,N_17070);
or UO_1846 (O_1846,N_16611,N_16273);
nor UO_1847 (O_1847,N_17448,N_19383);
nor UO_1848 (O_1848,N_16051,N_16980);
nor UO_1849 (O_1849,N_17138,N_17571);
nand UO_1850 (O_1850,N_16801,N_19605);
nor UO_1851 (O_1851,N_19937,N_17620);
nand UO_1852 (O_1852,N_16978,N_18605);
or UO_1853 (O_1853,N_16928,N_19602);
or UO_1854 (O_1854,N_17235,N_17118);
or UO_1855 (O_1855,N_19960,N_16934);
and UO_1856 (O_1856,N_18868,N_18451);
and UO_1857 (O_1857,N_17577,N_17582);
and UO_1858 (O_1858,N_19408,N_16268);
and UO_1859 (O_1859,N_18805,N_17183);
or UO_1860 (O_1860,N_19728,N_16953);
nand UO_1861 (O_1861,N_16795,N_17750);
or UO_1862 (O_1862,N_17724,N_19311);
and UO_1863 (O_1863,N_17886,N_16783);
nand UO_1864 (O_1864,N_19793,N_19839);
nor UO_1865 (O_1865,N_16257,N_17980);
and UO_1866 (O_1866,N_19737,N_18439);
or UO_1867 (O_1867,N_16811,N_16929);
or UO_1868 (O_1868,N_19837,N_16286);
nor UO_1869 (O_1869,N_17143,N_18191);
and UO_1870 (O_1870,N_18552,N_16094);
nor UO_1871 (O_1871,N_18741,N_18107);
nor UO_1872 (O_1872,N_19169,N_18270);
nand UO_1873 (O_1873,N_19467,N_18170);
or UO_1874 (O_1874,N_18123,N_16965);
and UO_1875 (O_1875,N_18758,N_17933);
nand UO_1876 (O_1876,N_16344,N_17815);
or UO_1877 (O_1877,N_16226,N_18697);
nand UO_1878 (O_1878,N_19853,N_19112);
and UO_1879 (O_1879,N_16202,N_18005);
and UO_1880 (O_1880,N_16012,N_18378);
or UO_1881 (O_1881,N_16403,N_18744);
nor UO_1882 (O_1882,N_16337,N_17931);
nor UO_1883 (O_1883,N_19459,N_16769);
or UO_1884 (O_1884,N_16388,N_16169);
nor UO_1885 (O_1885,N_17196,N_19009);
nor UO_1886 (O_1886,N_19818,N_17626);
nand UO_1887 (O_1887,N_18119,N_16027);
and UO_1888 (O_1888,N_16621,N_17280);
and UO_1889 (O_1889,N_19182,N_17413);
nand UO_1890 (O_1890,N_19831,N_18904);
and UO_1891 (O_1891,N_16957,N_18138);
nand UO_1892 (O_1892,N_17292,N_18391);
and UO_1893 (O_1893,N_18333,N_19798);
or UO_1894 (O_1894,N_18178,N_19327);
nor UO_1895 (O_1895,N_19417,N_16579);
and UO_1896 (O_1896,N_19024,N_16072);
nor UO_1897 (O_1897,N_16310,N_18438);
nand UO_1898 (O_1898,N_18568,N_19388);
or UO_1899 (O_1899,N_16900,N_19105);
nand UO_1900 (O_1900,N_19175,N_18650);
nor UO_1901 (O_1901,N_16342,N_16695);
nand UO_1902 (O_1902,N_19592,N_19769);
nor UO_1903 (O_1903,N_16157,N_17796);
nor UO_1904 (O_1904,N_18976,N_17297);
or UO_1905 (O_1905,N_16154,N_19891);
nand UO_1906 (O_1906,N_19188,N_16590);
and UO_1907 (O_1907,N_16933,N_17155);
or UO_1908 (O_1908,N_17705,N_18081);
nand UO_1909 (O_1909,N_18569,N_18194);
or UO_1910 (O_1910,N_18377,N_17003);
nor UO_1911 (O_1911,N_16331,N_18820);
and UO_1912 (O_1912,N_16661,N_18702);
nand UO_1913 (O_1913,N_18125,N_16762);
nand UO_1914 (O_1914,N_16309,N_17165);
and UO_1915 (O_1915,N_17462,N_18035);
nor UO_1916 (O_1916,N_17770,N_19242);
nand UO_1917 (O_1917,N_19844,N_17688);
or UO_1918 (O_1918,N_18268,N_17642);
and UO_1919 (O_1919,N_19678,N_17084);
or UO_1920 (O_1920,N_17040,N_18953);
nor UO_1921 (O_1921,N_18475,N_16171);
or UO_1922 (O_1922,N_16237,N_18415);
nor UO_1923 (O_1923,N_16693,N_19489);
or UO_1924 (O_1924,N_18359,N_17879);
or UO_1925 (O_1925,N_19420,N_19547);
nand UO_1926 (O_1926,N_17051,N_17515);
and UO_1927 (O_1927,N_17692,N_19830);
nand UO_1928 (O_1928,N_19708,N_18933);
nor UO_1929 (O_1929,N_19474,N_19450);
and UO_1930 (O_1930,N_19504,N_17549);
nor UO_1931 (O_1931,N_19092,N_17579);
nor UO_1932 (O_1932,N_18085,N_19272);
nor UO_1933 (O_1933,N_18516,N_19908);
nand UO_1934 (O_1934,N_18583,N_19671);
nand UO_1935 (O_1935,N_17005,N_16489);
and UO_1936 (O_1936,N_17759,N_16470);
and UO_1937 (O_1937,N_19160,N_18942);
and UO_1938 (O_1938,N_19664,N_19345);
and UO_1939 (O_1939,N_17452,N_17135);
or UO_1940 (O_1940,N_19392,N_19829);
xnor UO_1941 (O_1941,N_19027,N_19285);
and UO_1942 (O_1942,N_16614,N_16359);
nor UO_1943 (O_1943,N_18966,N_17417);
and UO_1944 (O_1944,N_19794,N_17326);
or UO_1945 (O_1945,N_18811,N_19168);
nand UO_1946 (O_1946,N_18737,N_19023);
and UO_1947 (O_1947,N_19557,N_18122);
nand UO_1948 (O_1948,N_18768,N_18375);
or UO_1949 (O_1949,N_16111,N_18757);
nor UO_1950 (O_1950,N_18210,N_16684);
nand UO_1951 (O_1951,N_16617,N_17774);
and UO_1952 (O_1952,N_17656,N_18398);
or UO_1953 (O_1953,N_16305,N_17716);
or UO_1954 (O_1954,N_18704,N_16817);
or UO_1955 (O_1955,N_18127,N_19073);
nand UO_1956 (O_1956,N_19812,N_16942);
nor UO_1957 (O_1957,N_18855,N_17730);
xor UO_1958 (O_1958,N_19217,N_18262);
nor UO_1959 (O_1959,N_16587,N_18883);
or UO_1960 (O_1960,N_19570,N_16212);
nor UO_1961 (O_1961,N_17740,N_19756);
nand UO_1962 (O_1962,N_16797,N_18615);
nand UO_1963 (O_1963,N_16751,N_18488);
and UO_1964 (O_1964,N_19871,N_18562);
nand UO_1965 (O_1965,N_19103,N_19042);
nand UO_1966 (O_1966,N_17460,N_18743);
nand UO_1967 (O_1967,N_16097,N_16078);
nor UO_1968 (O_1968,N_17848,N_16085);
and UO_1969 (O_1969,N_19014,N_16606);
or UO_1970 (O_1970,N_17694,N_19860);
and UO_1971 (O_1971,N_18675,N_19353);
and UO_1972 (O_1972,N_17921,N_17217);
nor UO_1973 (O_1973,N_19606,N_16970);
nor UO_1974 (O_1974,N_18018,N_16334);
and UO_1975 (O_1975,N_18972,N_18973);
nor UO_1976 (O_1976,N_17616,N_17032);
nor UO_1977 (O_1977,N_16735,N_18218);
and UO_1978 (O_1978,N_19748,N_17928);
and UO_1979 (O_1979,N_16256,N_18477);
nand UO_1980 (O_1980,N_18269,N_18957);
or UO_1981 (O_1981,N_16807,N_16398);
or UO_1982 (O_1982,N_19026,N_17168);
nor UO_1983 (O_1983,N_17530,N_18371);
nand UO_1984 (O_1984,N_16081,N_18483);
or UO_1985 (O_1985,N_16748,N_19403);
nand UO_1986 (O_1986,N_16563,N_19364);
nor UO_1987 (O_1987,N_17994,N_16907);
and UO_1988 (O_1988,N_19020,N_16709);
nor UO_1989 (O_1989,N_19882,N_19768);
and UO_1990 (O_1990,N_17686,N_19722);
nand UO_1991 (O_1991,N_16086,N_18560);
nand UO_1992 (O_1992,N_19566,N_17004);
nand UO_1993 (O_1993,N_16071,N_18588);
or UO_1994 (O_1994,N_18128,N_16136);
nor UO_1995 (O_1995,N_19933,N_17228);
nor UO_1996 (O_1996,N_19350,N_17710);
nand UO_1997 (O_1997,N_18434,N_17628);
nor UO_1998 (O_1998,N_17733,N_19611);
or UO_1999 (O_1999,N_19351,N_19563);
and UO_2000 (O_2000,N_19903,N_16964);
nand UO_2001 (O_2001,N_17448,N_16056);
or UO_2002 (O_2002,N_19029,N_16322);
nor UO_2003 (O_2003,N_19638,N_17503);
nand UO_2004 (O_2004,N_17574,N_19482);
and UO_2005 (O_2005,N_18540,N_18214);
and UO_2006 (O_2006,N_19959,N_19837);
nor UO_2007 (O_2007,N_19163,N_19457);
nand UO_2008 (O_2008,N_19437,N_18087);
nor UO_2009 (O_2009,N_19064,N_16252);
nand UO_2010 (O_2010,N_19085,N_19665);
xor UO_2011 (O_2011,N_19665,N_19305);
nor UO_2012 (O_2012,N_19604,N_19859);
and UO_2013 (O_2013,N_17186,N_17472);
or UO_2014 (O_2014,N_16158,N_16647);
nor UO_2015 (O_2015,N_18140,N_17731);
nand UO_2016 (O_2016,N_19641,N_17092);
and UO_2017 (O_2017,N_16893,N_16172);
nor UO_2018 (O_2018,N_16582,N_16361);
and UO_2019 (O_2019,N_19154,N_16353);
or UO_2020 (O_2020,N_18937,N_16784);
or UO_2021 (O_2021,N_19793,N_18106);
nand UO_2022 (O_2022,N_18858,N_18677);
nor UO_2023 (O_2023,N_16679,N_18226);
nand UO_2024 (O_2024,N_18655,N_19343);
and UO_2025 (O_2025,N_16113,N_19507);
and UO_2026 (O_2026,N_18295,N_17941);
nor UO_2027 (O_2027,N_16472,N_16093);
and UO_2028 (O_2028,N_19864,N_18206);
or UO_2029 (O_2029,N_18083,N_16830);
nand UO_2030 (O_2030,N_16118,N_19066);
nand UO_2031 (O_2031,N_18902,N_17073);
nand UO_2032 (O_2032,N_17412,N_17890);
or UO_2033 (O_2033,N_18425,N_19762);
nor UO_2034 (O_2034,N_16268,N_17737);
nand UO_2035 (O_2035,N_16802,N_16583);
and UO_2036 (O_2036,N_18246,N_16061);
nand UO_2037 (O_2037,N_18924,N_19467);
or UO_2038 (O_2038,N_17137,N_19200);
and UO_2039 (O_2039,N_18279,N_18413);
xor UO_2040 (O_2040,N_16704,N_18517);
or UO_2041 (O_2041,N_17946,N_17365);
or UO_2042 (O_2042,N_19618,N_16228);
nand UO_2043 (O_2043,N_18309,N_16547);
nand UO_2044 (O_2044,N_19451,N_17097);
nor UO_2045 (O_2045,N_17906,N_19904);
or UO_2046 (O_2046,N_16139,N_18775);
nand UO_2047 (O_2047,N_18729,N_19986);
nor UO_2048 (O_2048,N_16168,N_17441);
and UO_2049 (O_2049,N_18068,N_19067);
nand UO_2050 (O_2050,N_16283,N_17907);
and UO_2051 (O_2051,N_19926,N_17306);
and UO_2052 (O_2052,N_18936,N_19893);
nand UO_2053 (O_2053,N_16973,N_17798);
and UO_2054 (O_2054,N_17478,N_17863);
and UO_2055 (O_2055,N_17292,N_18681);
or UO_2056 (O_2056,N_18358,N_18808);
nor UO_2057 (O_2057,N_16666,N_18172);
nand UO_2058 (O_2058,N_16702,N_19663);
nand UO_2059 (O_2059,N_18052,N_17074);
or UO_2060 (O_2060,N_19391,N_16734);
nand UO_2061 (O_2061,N_17723,N_18692);
xnor UO_2062 (O_2062,N_17444,N_17569);
nand UO_2063 (O_2063,N_16800,N_18695);
or UO_2064 (O_2064,N_18039,N_17425);
nand UO_2065 (O_2065,N_18104,N_18850);
or UO_2066 (O_2066,N_16769,N_18268);
nand UO_2067 (O_2067,N_16421,N_16118);
nand UO_2068 (O_2068,N_18325,N_17582);
nand UO_2069 (O_2069,N_18474,N_17280);
and UO_2070 (O_2070,N_16025,N_16110);
xor UO_2071 (O_2071,N_19745,N_16998);
or UO_2072 (O_2072,N_18294,N_19754);
nor UO_2073 (O_2073,N_17649,N_17529);
and UO_2074 (O_2074,N_17692,N_18950);
or UO_2075 (O_2075,N_17821,N_19936);
nor UO_2076 (O_2076,N_19192,N_18045);
and UO_2077 (O_2077,N_17451,N_17011);
nand UO_2078 (O_2078,N_17067,N_19424);
xor UO_2079 (O_2079,N_16314,N_19726);
or UO_2080 (O_2080,N_19084,N_19041);
nor UO_2081 (O_2081,N_16611,N_16297);
and UO_2082 (O_2082,N_16720,N_16803);
or UO_2083 (O_2083,N_19497,N_16836);
and UO_2084 (O_2084,N_16469,N_18566);
and UO_2085 (O_2085,N_16173,N_17568);
nand UO_2086 (O_2086,N_17219,N_19527);
nand UO_2087 (O_2087,N_19013,N_17837);
and UO_2088 (O_2088,N_16349,N_18055);
nand UO_2089 (O_2089,N_17511,N_19337);
or UO_2090 (O_2090,N_19702,N_16570);
nand UO_2091 (O_2091,N_19897,N_16607);
or UO_2092 (O_2092,N_19784,N_16164);
nand UO_2093 (O_2093,N_16296,N_18347);
nor UO_2094 (O_2094,N_18114,N_18463);
nand UO_2095 (O_2095,N_16955,N_18872);
nor UO_2096 (O_2096,N_17425,N_16910);
nor UO_2097 (O_2097,N_19594,N_16517);
and UO_2098 (O_2098,N_17577,N_19478);
or UO_2099 (O_2099,N_17368,N_18800);
xor UO_2100 (O_2100,N_19894,N_17729);
or UO_2101 (O_2101,N_16972,N_18211);
and UO_2102 (O_2102,N_19806,N_19360);
or UO_2103 (O_2103,N_18408,N_16324);
or UO_2104 (O_2104,N_19918,N_16607);
nand UO_2105 (O_2105,N_18694,N_18304);
or UO_2106 (O_2106,N_18487,N_19730);
and UO_2107 (O_2107,N_18647,N_18889);
nand UO_2108 (O_2108,N_19129,N_17579);
or UO_2109 (O_2109,N_17323,N_16696);
nor UO_2110 (O_2110,N_18518,N_17400);
and UO_2111 (O_2111,N_16055,N_16071);
and UO_2112 (O_2112,N_18233,N_19597);
nor UO_2113 (O_2113,N_19390,N_16539);
nor UO_2114 (O_2114,N_18859,N_17747);
and UO_2115 (O_2115,N_16326,N_16401);
nand UO_2116 (O_2116,N_17627,N_16893);
xor UO_2117 (O_2117,N_17221,N_16684);
xor UO_2118 (O_2118,N_17899,N_19517);
nor UO_2119 (O_2119,N_17076,N_19939);
nor UO_2120 (O_2120,N_17779,N_18329);
or UO_2121 (O_2121,N_16223,N_19522);
or UO_2122 (O_2122,N_19461,N_18330);
nor UO_2123 (O_2123,N_19821,N_19313);
or UO_2124 (O_2124,N_16906,N_16754);
or UO_2125 (O_2125,N_17009,N_16833);
nor UO_2126 (O_2126,N_16770,N_18618);
nor UO_2127 (O_2127,N_18286,N_16771);
nand UO_2128 (O_2128,N_17959,N_19314);
nor UO_2129 (O_2129,N_16807,N_17775);
nand UO_2130 (O_2130,N_18982,N_18930);
xor UO_2131 (O_2131,N_19060,N_19233);
nand UO_2132 (O_2132,N_17196,N_18842);
and UO_2133 (O_2133,N_19172,N_17614);
and UO_2134 (O_2134,N_16257,N_19217);
and UO_2135 (O_2135,N_19020,N_16045);
nor UO_2136 (O_2136,N_16906,N_19948);
xnor UO_2137 (O_2137,N_17648,N_19305);
nor UO_2138 (O_2138,N_16089,N_17741);
and UO_2139 (O_2139,N_17092,N_17934);
or UO_2140 (O_2140,N_19327,N_16322);
nand UO_2141 (O_2141,N_16839,N_18095);
or UO_2142 (O_2142,N_18914,N_19590);
or UO_2143 (O_2143,N_18470,N_16831);
xor UO_2144 (O_2144,N_16422,N_18393);
and UO_2145 (O_2145,N_16421,N_19261);
nand UO_2146 (O_2146,N_17930,N_18107);
nor UO_2147 (O_2147,N_19457,N_17739);
nor UO_2148 (O_2148,N_18973,N_18423);
nor UO_2149 (O_2149,N_19842,N_16780);
and UO_2150 (O_2150,N_17570,N_19426);
or UO_2151 (O_2151,N_18425,N_16680);
nor UO_2152 (O_2152,N_18967,N_16790);
nand UO_2153 (O_2153,N_16766,N_19242);
nor UO_2154 (O_2154,N_19212,N_18746);
and UO_2155 (O_2155,N_17963,N_19768);
nor UO_2156 (O_2156,N_18180,N_19775);
nand UO_2157 (O_2157,N_16259,N_19544);
nand UO_2158 (O_2158,N_19780,N_16264);
nand UO_2159 (O_2159,N_17670,N_18601);
and UO_2160 (O_2160,N_17286,N_19735);
nand UO_2161 (O_2161,N_18222,N_17068);
and UO_2162 (O_2162,N_17478,N_19358);
or UO_2163 (O_2163,N_17052,N_16727);
nand UO_2164 (O_2164,N_19297,N_17059);
or UO_2165 (O_2165,N_17718,N_19705);
nand UO_2166 (O_2166,N_19496,N_16515);
nor UO_2167 (O_2167,N_17021,N_17196);
nor UO_2168 (O_2168,N_16110,N_18952);
nor UO_2169 (O_2169,N_18276,N_17444);
and UO_2170 (O_2170,N_19203,N_19264);
nor UO_2171 (O_2171,N_16715,N_18679);
nor UO_2172 (O_2172,N_19323,N_19469);
and UO_2173 (O_2173,N_19567,N_18469);
or UO_2174 (O_2174,N_19558,N_19776);
nand UO_2175 (O_2175,N_19577,N_18426);
nor UO_2176 (O_2176,N_19030,N_17928);
nand UO_2177 (O_2177,N_19867,N_17813);
and UO_2178 (O_2178,N_19039,N_17910);
or UO_2179 (O_2179,N_16066,N_18125);
nor UO_2180 (O_2180,N_17127,N_17117);
nor UO_2181 (O_2181,N_18190,N_17726);
or UO_2182 (O_2182,N_16594,N_19083);
nand UO_2183 (O_2183,N_17071,N_18351);
nand UO_2184 (O_2184,N_19831,N_16658);
nor UO_2185 (O_2185,N_18283,N_16330);
or UO_2186 (O_2186,N_17295,N_18912);
nand UO_2187 (O_2187,N_18889,N_17179);
nor UO_2188 (O_2188,N_19340,N_18998);
nor UO_2189 (O_2189,N_18166,N_18841);
nor UO_2190 (O_2190,N_18510,N_16502);
nand UO_2191 (O_2191,N_19209,N_16594);
and UO_2192 (O_2192,N_19596,N_16603);
nand UO_2193 (O_2193,N_18567,N_16034);
nand UO_2194 (O_2194,N_17044,N_19319);
or UO_2195 (O_2195,N_19766,N_16383);
nor UO_2196 (O_2196,N_17097,N_17001);
nor UO_2197 (O_2197,N_16906,N_18899);
nand UO_2198 (O_2198,N_17237,N_16669);
or UO_2199 (O_2199,N_19531,N_16651);
or UO_2200 (O_2200,N_18443,N_16439);
nand UO_2201 (O_2201,N_18175,N_19171);
or UO_2202 (O_2202,N_17264,N_17068);
xor UO_2203 (O_2203,N_18093,N_16537);
and UO_2204 (O_2204,N_19698,N_19110);
nand UO_2205 (O_2205,N_19851,N_19320);
or UO_2206 (O_2206,N_18001,N_16730);
and UO_2207 (O_2207,N_18843,N_17894);
nand UO_2208 (O_2208,N_17405,N_19309);
nor UO_2209 (O_2209,N_17856,N_16588);
nor UO_2210 (O_2210,N_17160,N_18069);
nand UO_2211 (O_2211,N_19564,N_19073);
and UO_2212 (O_2212,N_19348,N_17940);
and UO_2213 (O_2213,N_16330,N_16416);
nor UO_2214 (O_2214,N_19040,N_18649);
and UO_2215 (O_2215,N_19805,N_16091);
nor UO_2216 (O_2216,N_18855,N_18595);
or UO_2217 (O_2217,N_19255,N_19263);
or UO_2218 (O_2218,N_17256,N_19343);
nor UO_2219 (O_2219,N_18860,N_18958);
and UO_2220 (O_2220,N_17083,N_18382);
nand UO_2221 (O_2221,N_17031,N_17013);
nor UO_2222 (O_2222,N_17375,N_16463);
or UO_2223 (O_2223,N_16986,N_19600);
nor UO_2224 (O_2224,N_16125,N_17641);
nand UO_2225 (O_2225,N_17693,N_17529);
nand UO_2226 (O_2226,N_18040,N_18655);
or UO_2227 (O_2227,N_16447,N_19216);
and UO_2228 (O_2228,N_19989,N_17620);
nand UO_2229 (O_2229,N_18522,N_19056);
nor UO_2230 (O_2230,N_16446,N_16135);
and UO_2231 (O_2231,N_16923,N_18078);
nand UO_2232 (O_2232,N_19671,N_16511);
nand UO_2233 (O_2233,N_16133,N_16316);
nor UO_2234 (O_2234,N_18010,N_16120);
nor UO_2235 (O_2235,N_16956,N_17885);
nand UO_2236 (O_2236,N_18205,N_16419);
nor UO_2237 (O_2237,N_16927,N_18503);
nand UO_2238 (O_2238,N_16982,N_16416);
nor UO_2239 (O_2239,N_18008,N_18414);
nor UO_2240 (O_2240,N_17087,N_16298);
and UO_2241 (O_2241,N_16596,N_19763);
nand UO_2242 (O_2242,N_18243,N_17315);
nor UO_2243 (O_2243,N_19835,N_17433);
and UO_2244 (O_2244,N_17505,N_16762);
nor UO_2245 (O_2245,N_17420,N_18215);
and UO_2246 (O_2246,N_17914,N_19873);
or UO_2247 (O_2247,N_16126,N_18383);
nand UO_2248 (O_2248,N_16404,N_17721);
or UO_2249 (O_2249,N_19746,N_19334);
nand UO_2250 (O_2250,N_19378,N_17503);
nor UO_2251 (O_2251,N_19221,N_18074);
and UO_2252 (O_2252,N_18633,N_17939);
nor UO_2253 (O_2253,N_18839,N_17910);
nand UO_2254 (O_2254,N_17423,N_16437);
xnor UO_2255 (O_2255,N_16145,N_17397);
or UO_2256 (O_2256,N_17922,N_18222);
nand UO_2257 (O_2257,N_18620,N_18175);
nor UO_2258 (O_2258,N_17136,N_19253);
and UO_2259 (O_2259,N_16895,N_16212);
nor UO_2260 (O_2260,N_19728,N_16658);
nor UO_2261 (O_2261,N_19222,N_19863);
or UO_2262 (O_2262,N_17905,N_17579);
nand UO_2263 (O_2263,N_18833,N_16054);
nand UO_2264 (O_2264,N_17832,N_18286);
nor UO_2265 (O_2265,N_19573,N_17687);
nand UO_2266 (O_2266,N_18674,N_17717);
and UO_2267 (O_2267,N_16304,N_16759);
and UO_2268 (O_2268,N_19205,N_19733);
or UO_2269 (O_2269,N_17630,N_18007);
and UO_2270 (O_2270,N_16587,N_18158);
nor UO_2271 (O_2271,N_16160,N_19708);
or UO_2272 (O_2272,N_16295,N_16725);
nand UO_2273 (O_2273,N_17092,N_19980);
nand UO_2274 (O_2274,N_18154,N_16421);
nand UO_2275 (O_2275,N_17626,N_19473);
nor UO_2276 (O_2276,N_18624,N_17993);
and UO_2277 (O_2277,N_16996,N_19666);
or UO_2278 (O_2278,N_18049,N_19947);
or UO_2279 (O_2279,N_18033,N_18438);
and UO_2280 (O_2280,N_18533,N_16900);
nor UO_2281 (O_2281,N_18506,N_19007);
and UO_2282 (O_2282,N_18484,N_16706);
nand UO_2283 (O_2283,N_19838,N_16489);
or UO_2284 (O_2284,N_17938,N_19656);
or UO_2285 (O_2285,N_19579,N_18421);
nand UO_2286 (O_2286,N_19052,N_16890);
or UO_2287 (O_2287,N_19443,N_17409);
nor UO_2288 (O_2288,N_17829,N_16608);
nand UO_2289 (O_2289,N_18444,N_17081);
and UO_2290 (O_2290,N_16466,N_16118);
or UO_2291 (O_2291,N_18398,N_16051);
nand UO_2292 (O_2292,N_17357,N_16291);
nor UO_2293 (O_2293,N_18081,N_19737);
nand UO_2294 (O_2294,N_17347,N_17485);
and UO_2295 (O_2295,N_19077,N_16809);
nor UO_2296 (O_2296,N_17654,N_16859);
or UO_2297 (O_2297,N_18923,N_19855);
nand UO_2298 (O_2298,N_19234,N_18834);
or UO_2299 (O_2299,N_19900,N_19337);
or UO_2300 (O_2300,N_17669,N_17719);
nor UO_2301 (O_2301,N_19450,N_16781);
and UO_2302 (O_2302,N_19002,N_19727);
nand UO_2303 (O_2303,N_16179,N_18289);
nand UO_2304 (O_2304,N_18441,N_18183);
or UO_2305 (O_2305,N_19577,N_16813);
and UO_2306 (O_2306,N_16509,N_18726);
and UO_2307 (O_2307,N_19019,N_18635);
nand UO_2308 (O_2308,N_17417,N_18179);
nor UO_2309 (O_2309,N_18383,N_18610);
and UO_2310 (O_2310,N_19134,N_16979);
nor UO_2311 (O_2311,N_17184,N_18901);
and UO_2312 (O_2312,N_16122,N_19452);
or UO_2313 (O_2313,N_19548,N_17225);
and UO_2314 (O_2314,N_17647,N_17440);
and UO_2315 (O_2315,N_17329,N_19046);
or UO_2316 (O_2316,N_17876,N_16371);
or UO_2317 (O_2317,N_16909,N_19087);
or UO_2318 (O_2318,N_19179,N_18321);
and UO_2319 (O_2319,N_17589,N_19494);
or UO_2320 (O_2320,N_17841,N_17474);
nor UO_2321 (O_2321,N_18689,N_16636);
nand UO_2322 (O_2322,N_17913,N_19877);
nand UO_2323 (O_2323,N_18690,N_16147);
nand UO_2324 (O_2324,N_18930,N_17413);
nor UO_2325 (O_2325,N_18433,N_16638);
or UO_2326 (O_2326,N_16147,N_18593);
and UO_2327 (O_2327,N_16295,N_17291);
nor UO_2328 (O_2328,N_17544,N_17071);
or UO_2329 (O_2329,N_17798,N_18575);
nand UO_2330 (O_2330,N_17341,N_17603);
nand UO_2331 (O_2331,N_19147,N_19242);
nor UO_2332 (O_2332,N_18574,N_19022);
and UO_2333 (O_2333,N_19952,N_17095);
nor UO_2334 (O_2334,N_18309,N_18447);
and UO_2335 (O_2335,N_19553,N_17345);
and UO_2336 (O_2336,N_19001,N_16707);
nor UO_2337 (O_2337,N_19045,N_18937);
and UO_2338 (O_2338,N_19087,N_19010);
or UO_2339 (O_2339,N_18605,N_18995);
or UO_2340 (O_2340,N_18698,N_16414);
and UO_2341 (O_2341,N_18506,N_18237);
and UO_2342 (O_2342,N_16711,N_19652);
nor UO_2343 (O_2343,N_17393,N_19945);
or UO_2344 (O_2344,N_18515,N_19636);
nand UO_2345 (O_2345,N_18553,N_18560);
or UO_2346 (O_2346,N_18533,N_17490);
and UO_2347 (O_2347,N_16112,N_19479);
or UO_2348 (O_2348,N_18482,N_17660);
nor UO_2349 (O_2349,N_16085,N_18333);
or UO_2350 (O_2350,N_18306,N_16161);
nor UO_2351 (O_2351,N_18796,N_19058);
nor UO_2352 (O_2352,N_16815,N_17224);
nand UO_2353 (O_2353,N_17374,N_17675);
nor UO_2354 (O_2354,N_17511,N_19811);
nor UO_2355 (O_2355,N_18177,N_17197);
nor UO_2356 (O_2356,N_19986,N_17929);
nor UO_2357 (O_2357,N_16002,N_19814);
and UO_2358 (O_2358,N_18248,N_19940);
and UO_2359 (O_2359,N_19245,N_18893);
nand UO_2360 (O_2360,N_19539,N_18440);
and UO_2361 (O_2361,N_16185,N_16267);
nand UO_2362 (O_2362,N_17286,N_19397);
or UO_2363 (O_2363,N_18954,N_16812);
and UO_2364 (O_2364,N_16105,N_17885);
nor UO_2365 (O_2365,N_18537,N_16780);
or UO_2366 (O_2366,N_18929,N_16769);
or UO_2367 (O_2367,N_16907,N_16331);
or UO_2368 (O_2368,N_19967,N_16919);
or UO_2369 (O_2369,N_16151,N_18860);
or UO_2370 (O_2370,N_19691,N_16436);
or UO_2371 (O_2371,N_19154,N_19415);
nand UO_2372 (O_2372,N_17517,N_17309);
and UO_2373 (O_2373,N_17871,N_17941);
and UO_2374 (O_2374,N_18433,N_18290);
nor UO_2375 (O_2375,N_19807,N_19628);
nor UO_2376 (O_2376,N_17931,N_17349);
nand UO_2377 (O_2377,N_17920,N_17740);
nor UO_2378 (O_2378,N_17585,N_16821);
or UO_2379 (O_2379,N_18873,N_16816);
and UO_2380 (O_2380,N_19054,N_18991);
or UO_2381 (O_2381,N_16774,N_16815);
or UO_2382 (O_2382,N_17914,N_18188);
and UO_2383 (O_2383,N_19824,N_19950);
and UO_2384 (O_2384,N_19773,N_17505);
nand UO_2385 (O_2385,N_17589,N_17776);
and UO_2386 (O_2386,N_19054,N_18393);
or UO_2387 (O_2387,N_19116,N_16082);
and UO_2388 (O_2388,N_16718,N_18301);
and UO_2389 (O_2389,N_17865,N_18983);
or UO_2390 (O_2390,N_18395,N_19293);
and UO_2391 (O_2391,N_18476,N_19330);
or UO_2392 (O_2392,N_19601,N_17930);
nor UO_2393 (O_2393,N_19248,N_19414);
or UO_2394 (O_2394,N_17308,N_18222);
nor UO_2395 (O_2395,N_19765,N_17558);
and UO_2396 (O_2396,N_19059,N_19249);
nand UO_2397 (O_2397,N_19615,N_18708);
nor UO_2398 (O_2398,N_18732,N_19897);
nor UO_2399 (O_2399,N_19016,N_18562);
nand UO_2400 (O_2400,N_18243,N_19558);
nor UO_2401 (O_2401,N_19315,N_19738);
nand UO_2402 (O_2402,N_18013,N_17406);
and UO_2403 (O_2403,N_16851,N_18603);
and UO_2404 (O_2404,N_16371,N_19629);
nor UO_2405 (O_2405,N_16369,N_17235);
nand UO_2406 (O_2406,N_19311,N_18881);
nor UO_2407 (O_2407,N_16628,N_18187);
nor UO_2408 (O_2408,N_19788,N_16832);
nand UO_2409 (O_2409,N_17630,N_16923);
nand UO_2410 (O_2410,N_18090,N_19902);
nor UO_2411 (O_2411,N_19377,N_19510);
nand UO_2412 (O_2412,N_18678,N_18077);
or UO_2413 (O_2413,N_17065,N_19460);
nand UO_2414 (O_2414,N_17754,N_17790);
nor UO_2415 (O_2415,N_19826,N_19521);
nor UO_2416 (O_2416,N_16295,N_17301);
or UO_2417 (O_2417,N_16437,N_19873);
nor UO_2418 (O_2418,N_16159,N_19659);
nand UO_2419 (O_2419,N_19583,N_17342);
and UO_2420 (O_2420,N_17700,N_16040);
and UO_2421 (O_2421,N_18484,N_19252);
nor UO_2422 (O_2422,N_16429,N_18194);
nor UO_2423 (O_2423,N_18042,N_19813);
or UO_2424 (O_2424,N_16530,N_18065);
nor UO_2425 (O_2425,N_16973,N_18593);
nand UO_2426 (O_2426,N_16755,N_18351);
or UO_2427 (O_2427,N_17436,N_17586);
nand UO_2428 (O_2428,N_19090,N_16975);
nand UO_2429 (O_2429,N_19324,N_17743);
or UO_2430 (O_2430,N_18139,N_19748);
or UO_2431 (O_2431,N_18914,N_18674);
nor UO_2432 (O_2432,N_16574,N_19651);
and UO_2433 (O_2433,N_19085,N_19229);
nor UO_2434 (O_2434,N_19241,N_19127);
nand UO_2435 (O_2435,N_19735,N_16698);
and UO_2436 (O_2436,N_18071,N_19070);
nor UO_2437 (O_2437,N_18151,N_19888);
and UO_2438 (O_2438,N_19146,N_19728);
nor UO_2439 (O_2439,N_16239,N_19585);
and UO_2440 (O_2440,N_18442,N_16867);
and UO_2441 (O_2441,N_18331,N_19664);
nand UO_2442 (O_2442,N_19563,N_16586);
or UO_2443 (O_2443,N_19649,N_16027);
and UO_2444 (O_2444,N_16291,N_17594);
nor UO_2445 (O_2445,N_18934,N_16844);
nor UO_2446 (O_2446,N_17204,N_19921);
or UO_2447 (O_2447,N_18636,N_19856);
and UO_2448 (O_2448,N_17720,N_16616);
and UO_2449 (O_2449,N_19598,N_18210);
nand UO_2450 (O_2450,N_16355,N_19005);
nand UO_2451 (O_2451,N_18041,N_18397);
or UO_2452 (O_2452,N_18605,N_16712);
nor UO_2453 (O_2453,N_19264,N_19811);
nor UO_2454 (O_2454,N_16813,N_17180);
nand UO_2455 (O_2455,N_18420,N_18673);
and UO_2456 (O_2456,N_19757,N_17665);
or UO_2457 (O_2457,N_16977,N_19470);
or UO_2458 (O_2458,N_16054,N_17540);
or UO_2459 (O_2459,N_17175,N_16232);
and UO_2460 (O_2460,N_16754,N_16008);
and UO_2461 (O_2461,N_18798,N_19503);
nor UO_2462 (O_2462,N_17458,N_16912);
and UO_2463 (O_2463,N_16808,N_16111);
nand UO_2464 (O_2464,N_17494,N_17714);
or UO_2465 (O_2465,N_18890,N_17594);
nand UO_2466 (O_2466,N_18428,N_19746);
and UO_2467 (O_2467,N_18986,N_19470);
and UO_2468 (O_2468,N_18139,N_18741);
or UO_2469 (O_2469,N_19094,N_16776);
nand UO_2470 (O_2470,N_18904,N_17649);
nor UO_2471 (O_2471,N_19498,N_16578);
nor UO_2472 (O_2472,N_18765,N_17719);
or UO_2473 (O_2473,N_19867,N_18657);
nand UO_2474 (O_2474,N_18165,N_18637);
xnor UO_2475 (O_2475,N_19863,N_18075);
nor UO_2476 (O_2476,N_17320,N_16566);
nand UO_2477 (O_2477,N_18868,N_16706);
or UO_2478 (O_2478,N_16788,N_19273);
or UO_2479 (O_2479,N_17467,N_19803);
nor UO_2480 (O_2480,N_16082,N_18224);
nand UO_2481 (O_2481,N_18469,N_16067);
and UO_2482 (O_2482,N_17562,N_17119);
or UO_2483 (O_2483,N_19959,N_16246);
and UO_2484 (O_2484,N_17957,N_16861);
and UO_2485 (O_2485,N_18864,N_16884);
nor UO_2486 (O_2486,N_19206,N_19214);
nor UO_2487 (O_2487,N_16415,N_16101);
xor UO_2488 (O_2488,N_16330,N_16785);
nand UO_2489 (O_2489,N_16411,N_18917);
or UO_2490 (O_2490,N_19203,N_19703);
nand UO_2491 (O_2491,N_17486,N_17684);
and UO_2492 (O_2492,N_16078,N_18482);
nand UO_2493 (O_2493,N_17394,N_16592);
nand UO_2494 (O_2494,N_16928,N_19167);
or UO_2495 (O_2495,N_18664,N_18715);
and UO_2496 (O_2496,N_19536,N_17022);
or UO_2497 (O_2497,N_18600,N_16464);
xor UO_2498 (O_2498,N_16652,N_19625);
and UO_2499 (O_2499,N_19926,N_17067);
endmodule