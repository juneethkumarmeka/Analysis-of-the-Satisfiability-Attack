module basic_750_5000_1000_10_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_23,In_299);
or U1 (N_1,In_589,In_391);
nand U2 (N_2,In_580,In_400);
or U3 (N_3,In_617,In_521);
nor U4 (N_4,In_574,In_9);
nand U5 (N_5,In_160,In_303);
and U6 (N_6,In_363,In_45);
nor U7 (N_7,In_470,In_564);
or U8 (N_8,In_118,In_138);
or U9 (N_9,In_727,In_502);
or U10 (N_10,In_595,In_596);
nor U11 (N_11,In_27,In_560);
nor U12 (N_12,In_29,In_104);
and U13 (N_13,In_707,In_642);
or U14 (N_14,In_384,In_656);
and U15 (N_15,In_427,In_612);
nand U16 (N_16,In_60,In_432);
nor U17 (N_17,In_183,In_336);
xnor U18 (N_18,In_33,In_377);
and U19 (N_19,In_148,In_629);
and U20 (N_20,In_155,In_307);
and U21 (N_21,In_90,In_451);
xnor U22 (N_22,In_353,In_214);
nand U23 (N_23,In_235,In_720);
and U24 (N_24,In_190,In_48);
xor U25 (N_25,In_181,In_714);
nor U26 (N_26,In_70,In_718);
nor U27 (N_27,In_539,In_211);
or U28 (N_28,In_593,In_298);
or U29 (N_29,In_58,In_217);
nand U30 (N_30,In_610,In_417);
nor U31 (N_31,In_227,In_263);
nand U32 (N_32,In_34,In_459);
or U33 (N_33,In_78,In_291);
nand U34 (N_34,In_609,In_339);
nor U35 (N_35,In_66,In_255);
and U36 (N_36,In_14,In_150);
nor U37 (N_37,In_397,In_650);
nor U38 (N_38,In_740,In_242);
or U39 (N_39,In_578,In_31);
nand U40 (N_40,In_5,In_477);
or U41 (N_41,In_172,In_346);
nor U42 (N_42,In_556,In_405);
nor U43 (N_43,In_409,In_97);
nor U44 (N_44,In_186,In_563);
nor U45 (N_45,In_110,In_337);
and U46 (N_46,In_329,In_107);
and U47 (N_47,In_476,In_261);
and U48 (N_48,In_39,In_387);
nor U49 (N_49,In_441,In_355);
nor U50 (N_50,In_527,In_260);
or U51 (N_51,In_666,In_591);
or U52 (N_52,In_370,In_334);
nand U53 (N_53,In_231,In_475);
nor U54 (N_54,In_598,In_233);
nor U55 (N_55,In_582,In_43);
or U56 (N_56,In_705,In_641);
and U57 (N_57,In_232,In_249);
xor U58 (N_58,In_361,In_471);
and U59 (N_59,In_736,In_505);
nor U60 (N_60,In_145,In_175);
or U61 (N_61,In_466,In_542);
or U62 (N_62,In_454,In_429);
nor U63 (N_63,In_635,In_710);
xnor U64 (N_64,In_219,In_238);
or U65 (N_65,In_621,In_32);
nor U66 (N_66,In_203,In_457);
and U67 (N_67,In_731,In_673);
nand U68 (N_68,In_220,In_706);
and U69 (N_69,In_597,In_108);
nor U70 (N_70,In_171,In_305);
nor U71 (N_71,In_91,In_488);
or U72 (N_72,In_47,In_732);
and U73 (N_73,In_557,In_366);
nand U74 (N_74,In_575,In_209);
nand U75 (N_75,In_1,In_453);
nand U76 (N_76,In_674,In_259);
and U77 (N_77,In_681,In_114);
and U78 (N_78,In_423,In_586);
and U79 (N_79,In_94,In_413);
nand U80 (N_80,In_695,In_742);
and U81 (N_81,In_716,In_501);
nand U82 (N_82,In_603,In_522);
nand U83 (N_83,In_380,In_498);
nand U84 (N_84,In_276,In_319);
nor U85 (N_85,In_98,In_274);
nand U86 (N_86,In_265,In_382);
and U87 (N_87,In_611,In_525);
or U88 (N_88,In_630,In_561);
and U89 (N_89,In_719,In_38);
nor U90 (N_90,In_665,In_661);
or U91 (N_91,In_179,In_210);
and U92 (N_92,In_65,In_101);
and U93 (N_93,In_270,In_395);
or U94 (N_94,In_544,In_469);
nand U95 (N_95,In_304,In_602);
nand U96 (N_96,In_317,In_663);
nor U97 (N_97,In_734,In_446);
and U98 (N_98,In_688,In_646);
nor U99 (N_99,In_80,In_606);
nand U100 (N_100,In_280,In_607);
or U101 (N_101,In_422,In_106);
and U102 (N_102,In_349,In_283);
or U103 (N_103,In_687,In_371);
nand U104 (N_104,In_576,In_394);
and U105 (N_105,In_416,In_415);
nor U106 (N_106,In_82,In_2);
nor U107 (N_107,In_581,In_37);
or U108 (N_108,In_320,In_121);
or U109 (N_109,In_748,In_123);
or U110 (N_110,In_500,In_335);
nand U111 (N_111,In_126,In_715);
and U112 (N_112,In_533,In_367);
nand U113 (N_113,In_301,In_89);
or U114 (N_114,In_306,In_484);
nor U115 (N_115,In_376,In_351);
nand U116 (N_116,In_52,In_153);
or U117 (N_117,In_701,In_11);
or U118 (N_118,In_96,In_450);
nand U119 (N_119,In_269,In_592);
nand U120 (N_120,In_573,In_133);
nor U121 (N_121,In_430,In_711);
or U122 (N_122,In_552,In_230);
nand U123 (N_123,In_61,In_166);
nand U124 (N_124,In_455,In_266);
nor U125 (N_125,In_467,In_638);
or U126 (N_126,In_691,In_653);
nand U127 (N_127,In_645,In_667);
xnor U128 (N_128,In_236,In_712);
nand U129 (N_129,In_657,In_508);
and U130 (N_130,In_253,In_187);
nand U131 (N_131,In_294,In_668);
nor U132 (N_132,In_496,In_4);
nand U133 (N_133,In_424,In_569);
or U134 (N_134,In_222,In_26);
and U135 (N_135,In_410,In_322);
nor U136 (N_136,In_130,In_683);
nor U137 (N_137,In_374,In_296);
nand U138 (N_138,In_141,In_509);
xor U139 (N_139,In_288,In_604);
xor U140 (N_140,In_461,In_435);
or U141 (N_141,In_401,In_315);
nor U142 (N_142,In_157,In_402);
and U143 (N_143,In_250,In_692);
and U144 (N_144,In_733,In_474);
and U145 (N_145,In_514,In_20);
and U146 (N_146,In_234,In_140);
nand U147 (N_147,In_614,In_343);
nand U148 (N_148,In_345,In_293);
nand U149 (N_149,In_690,In_633);
or U150 (N_150,In_749,In_318);
nand U151 (N_151,In_73,In_536);
or U152 (N_152,In_12,In_262);
and U153 (N_153,In_689,In_482);
and U154 (N_154,In_622,In_159);
nand U155 (N_155,In_543,In_511);
xor U156 (N_156,In_117,In_678);
nor U157 (N_157,In_42,In_601);
nand U158 (N_158,In_587,In_205);
nand U159 (N_159,In_243,In_88);
nand U160 (N_160,In_373,In_297);
nand U161 (N_161,In_347,In_137);
nor U162 (N_162,In_747,In_378);
or U163 (N_163,In_411,In_237);
and U164 (N_164,In_309,In_684);
nor U165 (N_165,In_745,In_340);
and U166 (N_166,In_41,In_652);
nand U167 (N_167,In_356,In_112);
nor U168 (N_168,In_228,In_443);
nor U169 (N_169,In_717,In_670);
nand U170 (N_170,In_333,In_81);
nand U171 (N_171,In_528,In_83);
nand U172 (N_172,In_448,In_134);
and U173 (N_173,In_702,In_693);
or U174 (N_174,In_440,In_169);
nand U175 (N_175,In_393,In_545);
or U176 (N_176,In_659,In_554);
nor U177 (N_177,In_344,In_464);
nor U178 (N_178,In_135,In_605);
and U179 (N_179,In_532,In_549);
xnor U180 (N_180,In_680,In_414);
xnor U181 (N_181,In_69,In_156);
or U182 (N_182,In_647,In_486);
nand U183 (N_183,In_77,In_462);
or U184 (N_184,In_178,In_103);
nand U185 (N_185,In_8,In_516);
nor U186 (N_186,In_512,In_627);
nor U187 (N_187,In_287,In_418);
and U188 (N_188,In_704,In_550);
nor U189 (N_189,In_531,In_698);
xor U190 (N_190,In_588,In_746);
nor U191 (N_191,In_127,In_568);
and U192 (N_192,In_245,In_634);
and U193 (N_193,In_28,In_24);
and U194 (N_194,In_649,In_201);
nand U195 (N_195,In_17,In_364);
and U196 (N_196,In_599,In_383);
or U197 (N_197,In_16,In_204);
or U198 (N_198,In_360,In_30);
or U199 (N_199,In_342,In_85);
or U200 (N_200,In_357,In_350);
and U201 (N_201,In_241,In_620);
nand U202 (N_202,In_485,In_163);
or U203 (N_203,In_285,In_679);
nor U204 (N_204,In_463,In_682);
nand U205 (N_205,In_664,In_338);
nor U206 (N_206,In_272,In_686);
nor U207 (N_207,In_628,In_308);
nand U208 (N_208,In_286,In_426);
or U209 (N_209,In_577,In_57);
nand U210 (N_210,In_566,In_392);
or U211 (N_211,In_654,In_200);
nand U212 (N_212,In_375,In_354);
and U213 (N_213,In_737,In_271);
xor U214 (N_214,In_473,In_626);
nand U215 (N_215,In_248,In_193);
nand U216 (N_216,In_481,In_225);
and U217 (N_217,In_267,In_128);
and U218 (N_218,In_321,In_313);
nor U219 (N_219,In_206,In_93);
or U220 (N_220,In_275,In_164);
nor U221 (N_221,In_672,In_412);
nor U222 (N_222,In_115,In_158);
nor U223 (N_223,In_18,In_503);
xor U224 (N_224,In_132,In_381);
or U225 (N_225,In_728,In_314);
nand U226 (N_226,In_709,In_102);
nand U227 (N_227,In_327,In_182);
nand U228 (N_228,In_144,In_15);
nor U229 (N_229,In_197,In_198);
or U230 (N_230,In_631,In_369);
nand U231 (N_231,In_289,In_660);
nand U232 (N_232,In_208,In_216);
or U233 (N_233,In_10,In_571);
nand U234 (N_234,In_420,In_0);
and U235 (N_235,In_725,In_438);
nor U236 (N_236,In_184,In_75);
nor U237 (N_237,In_724,In_729);
or U238 (N_238,In_215,In_331);
or U239 (N_239,In_460,In_221);
xor U240 (N_240,In_492,In_139);
or U241 (N_241,In_279,In_348);
or U242 (N_242,In_277,In_36);
or U243 (N_243,In_517,In_537);
nor U244 (N_244,In_559,In_252);
nor U245 (N_245,In_74,In_310);
or U246 (N_246,In_445,In_590);
and U247 (N_247,In_177,In_62);
xor U248 (N_248,In_493,In_49);
nor U249 (N_249,In_434,In_13);
nand U250 (N_250,In_64,In_616);
or U251 (N_251,In_311,In_192);
and U252 (N_252,In_379,In_146);
nor U253 (N_253,In_68,In_147);
nand U254 (N_254,In_312,In_708);
nor U255 (N_255,In_173,In_671);
or U256 (N_256,In_479,In_439);
or U257 (N_257,In_56,In_447);
nand U258 (N_258,In_555,In_365);
and U259 (N_259,In_726,In_565);
nand U260 (N_260,In_442,In_535);
or U261 (N_261,In_180,In_125);
nand U262 (N_262,In_76,In_399);
nor U263 (N_263,In_520,In_694);
nor U264 (N_264,In_185,In_515);
and U265 (N_265,In_324,In_491);
nor U266 (N_266,In_478,In_744);
nand U267 (N_267,In_669,In_558);
and U268 (N_268,In_195,In_456);
or U269 (N_269,In_300,In_239);
nor U270 (N_270,In_79,In_63);
or U271 (N_271,In_546,In_256);
xor U272 (N_272,In_741,In_613);
xor U273 (N_273,In_50,In_648);
nand U274 (N_274,In_67,In_675);
or U275 (N_275,In_273,In_189);
nor U276 (N_276,In_738,In_541);
xnor U277 (N_277,In_6,In_284);
nor U278 (N_278,In_168,In_735);
nor U279 (N_279,In_142,In_644);
and U280 (N_280,In_722,In_436);
nand U281 (N_281,In_406,In_325);
and U282 (N_282,In_676,In_510);
or U283 (N_283,In_584,In_99);
nor U284 (N_284,In_721,In_199);
or U285 (N_285,In_87,In_3);
or U286 (N_286,In_244,In_341);
and U287 (N_287,In_154,In_86);
nor U288 (N_288,In_444,In_703);
or U289 (N_289,In_408,In_119);
nor U290 (N_290,In_188,In_489);
nand U291 (N_291,In_389,In_40);
and U292 (N_292,In_562,In_174);
xor U293 (N_293,In_615,In_625);
or U294 (N_294,In_257,In_212);
or U295 (N_295,In_594,In_323);
nor U296 (N_296,In_251,In_696);
and U297 (N_297,In_518,In_385);
xnor U298 (N_298,In_7,In_585);
nand U299 (N_299,In_618,In_655);
nand U300 (N_300,In_55,In_643);
nand U301 (N_301,In_19,In_226);
or U302 (N_302,In_120,In_292);
or U303 (N_303,In_372,In_662);
nor U304 (N_304,In_472,In_92);
nor U305 (N_305,In_332,In_483);
nor U306 (N_306,In_290,In_538);
and U307 (N_307,In_35,In_328);
nand U308 (N_308,In_403,In_386);
xnor U309 (N_309,In_608,In_247);
or U310 (N_310,In_519,In_161);
nand U311 (N_311,In_224,In_529);
nand U312 (N_312,In_624,In_72);
nand U313 (N_313,In_143,In_111);
nor U314 (N_314,In_194,In_499);
nor U315 (N_315,In_524,In_513);
nand U316 (N_316,In_572,In_196);
nand U317 (N_317,In_637,In_419);
and U318 (N_318,In_95,In_109);
nand U319 (N_319,In_730,In_579);
and U320 (N_320,In_449,In_129);
nand U321 (N_321,In_362,In_390);
nor U322 (N_322,In_468,In_465);
nand U323 (N_323,In_743,In_480);
or U324 (N_324,In_636,In_431);
nand U325 (N_325,In_723,In_437);
and U326 (N_326,In_398,In_302);
nor U327 (N_327,In_122,In_358);
and U328 (N_328,In_21,In_428);
xor U329 (N_329,In_651,In_540);
or U330 (N_330,In_433,In_452);
nand U331 (N_331,In_697,In_116);
or U332 (N_332,In_100,In_25);
or U333 (N_333,In_639,In_551);
nand U334 (N_334,In_223,In_368);
and U335 (N_335,In_330,In_295);
nor U336 (N_336,In_167,In_113);
nand U337 (N_337,In_534,In_421);
xor U338 (N_338,In_553,In_53);
xnor U339 (N_339,In_425,In_526);
nor U340 (N_340,In_59,In_316);
and U341 (N_341,In_623,In_282);
nor U342 (N_342,In_264,In_523);
nor U343 (N_343,In_388,In_507);
and U344 (N_344,In_136,In_326);
nor U345 (N_345,In_497,In_51);
nand U346 (N_346,In_640,In_218);
or U347 (N_347,In_504,In_396);
xnor U348 (N_348,In_458,In_570);
and U349 (N_349,In_352,In_487);
nand U350 (N_350,In_54,In_152);
and U351 (N_351,In_162,In_567);
or U352 (N_352,In_739,In_191);
or U353 (N_353,In_149,In_165);
nand U354 (N_354,In_490,In_105);
nor U355 (N_355,In_700,In_22);
nor U356 (N_356,In_699,In_495);
nor U357 (N_357,In_685,In_407);
and U358 (N_358,In_202,In_268);
or U359 (N_359,In_207,In_254);
xor U360 (N_360,In_658,In_506);
nor U361 (N_361,In_548,In_619);
or U362 (N_362,In_713,In_213);
nor U363 (N_363,In_170,In_583);
or U364 (N_364,In_131,In_46);
nor U365 (N_365,In_44,In_677);
nand U366 (N_366,In_176,In_71);
nor U367 (N_367,In_151,In_278);
nor U368 (N_368,In_240,In_494);
xnor U369 (N_369,In_246,In_530);
xnor U370 (N_370,In_281,In_229);
and U371 (N_371,In_404,In_547);
xnor U372 (N_372,In_124,In_632);
xor U373 (N_373,In_258,In_84);
or U374 (N_374,In_359,In_600);
nor U375 (N_375,In_143,In_713);
or U376 (N_376,In_729,In_449);
and U377 (N_377,In_482,In_359);
nor U378 (N_378,In_106,In_403);
nand U379 (N_379,In_549,In_429);
nand U380 (N_380,In_344,In_425);
and U381 (N_381,In_538,In_472);
or U382 (N_382,In_637,In_225);
nand U383 (N_383,In_481,In_338);
nand U384 (N_384,In_292,In_724);
or U385 (N_385,In_452,In_418);
or U386 (N_386,In_735,In_623);
and U387 (N_387,In_684,In_612);
or U388 (N_388,In_251,In_727);
and U389 (N_389,In_286,In_360);
nand U390 (N_390,In_199,In_190);
nor U391 (N_391,In_440,In_35);
nand U392 (N_392,In_166,In_596);
or U393 (N_393,In_376,In_229);
nor U394 (N_394,In_67,In_94);
nand U395 (N_395,In_433,In_633);
or U396 (N_396,In_708,In_279);
and U397 (N_397,In_689,In_196);
nor U398 (N_398,In_647,In_63);
and U399 (N_399,In_213,In_62);
nor U400 (N_400,In_665,In_525);
and U401 (N_401,In_7,In_194);
nand U402 (N_402,In_619,In_425);
nand U403 (N_403,In_726,In_719);
or U404 (N_404,In_545,In_384);
or U405 (N_405,In_558,In_254);
and U406 (N_406,In_459,In_305);
xor U407 (N_407,In_70,In_0);
nand U408 (N_408,In_48,In_427);
and U409 (N_409,In_695,In_17);
nand U410 (N_410,In_369,In_596);
and U411 (N_411,In_112,In_560);
or U412 (N_412,In_44,In_247);
or U413 (N_413,In_133,In_723);
nor U414 (N_414,In_729,In_741);
and U415 (N_415,In_205,In_518);
nor U416 (N_416,In_745,In_512);
nor U417 (N_417,In_397,In_575);
nand U418 (N_418,In_659,In_56);
and U419 (N_419,In_260,In_69);
and U420 (N_420,In_171,In_14);
nor U421 (N_421,In_266,In_4);
xor U422 (N_422,In_188,In_237);
or U423 (N_423,In_410,In_440);
nand U424 (N_424,In_591,In_679);
nor U425 (N_425,In_621,In_6);
nand U426 (N_426,In_106,In_171);
or U427 (N_427,In_238,In_595);
nor U428 (N_428,In_738,In_250);
or U429 (N_429,In_477,In_400);
or U430 (N_430,In_157,In_240);
and U431 (N_431,In_280,In_302);
nand U432 (N_432,In_432,In_220);
nand U433 (N_433,In_33,In_284);
nor U434 (N_434,In_617,In_121);
or U435 (N_435,In_575,In_48);
and U436 (N_436,In_582,In_681);
or U437 (N_437,In_709,In_558);
xnor U438 (N_438,In_608,In_711);
nand U439 (N_439,In_407,In_388);
and U440 (N_440,In_362,In_554);
nor U441 (N_441,In_19,In_178);
and U442 (N_442,In_677,In_75);
nand U443 (N_443,In_601,In_708);
or U444 (N_444,In_721,In_71);
or U445 (N_445,In_412,In_425);
or U446 (N_446,In_250,In_526);
nand U447 (N_447,In_297,In_185);
nor U448 (N_448,In_14,In_3);
nand U449 (N_449,In_252,In_527);
or U450 (N_450,In_269,In_289);
nand U451 (N_451,In_298,In_746);
or U452 (N_452,In_516,In_60);
or U453 (N_453,In_460,In_563);
and U454 (N_454,In_333,In_140);
nor U455 (N_455,In_379,In_668);
nand U456 (N_456,In_239,In_743);
nor U457 (N_457,In_498,In_447);
nand U458 (N_458,In_135,In_569);
and U459 (N_459,In_419,In_350);
xnor U460 (N_460,In_15,In_25);
and U461 (N_461,In_484,In_274);
nor U462 (N_462,In_12,In_75);
and U463 (N_463,In_665,In_162);
nand U464 (N_464,In_430,In_243);
or U465 (N_465,In_248,In_654);
nand U466 (N_466,In_372,In_715);
or U467 (N_467,In_672,In_537);
nand U468 (N_468,In_331,In_643);
and U469 (N_469,In_74,In_701);
or U470 (N_470,In_324,In_457);
nor U471 (N_471,In_281,In_425);
xor U472 (N_472,In_466,In_232);
nor U473 (N_473,In_317,In_14);
xor U474 (N_474,In_280,In_241);
xnor U475 (N_475,In_656,In_293);
nand U476 (N_476,In_618,In_182);
nand U477 (N_477,In_282,In_97);
and U478 (N_478,In_252,In_712);
nor U479 (N_479,In_128,In_336);
xnor U480 (N_480,In_179,In_254);
or U481 (N_481,In_162,In_253);
and U482 (N_482,In_185,In_145);
xor U483 (N_483,In_108,In_427);
or U484 (N_484,In_465,In_683);
and U485 (N_485,In_124,In_319);
or U486 (N_486,In_381,In_729);
and U487 (N_487,In_112,In_358);
nor U488 (N_488,In_239,In_338);
and U489 (N_489,In_372,In_369);
nand U490 (N_490,In_405,In_547);
nor U491 (N_491,In_600,In_173);
nor U492 (N_492,In_275,In_548);
or U493 (N_493,In_660,In_528);
nor U494 (N_494,In_385,In_487);
and U495 (N_495,In_460,In_146);
and U496 (N_496,In_626,In_380);
nand U497 (N_497,In_145,In_371);
xnor U498 (N_498,In_459,In_484);
xor U499 (N_499,In_193,In_65);
and U500 (N_500,N_390,N_64);
or U501 (N_501,N_419,N_465);
or U502 (N_502,N_159,N_418);
or U503 (N_503,N_48,N_160);
or U504 (N_504,N_284,N_229);
nand U505 (N_505,N_446,N_110);
nand U506 (N_506,N_28,N_333);
nand U507 (N_507,N_234,N_275);
nor U508 (N_508,N_259,N_118);
xnor U509 (N_509,N_149,N_216);
and U510 (N_510,N_19,N_420);
or U511 (N_511,N_61,N_65);
or U512 (N_512,N_363,N_242);
nand U513 (N_513,N_290,N_417);
nor U514 (N_514,N_99,N_341);
nand U515 (N_515,N_354,N_493);
nand U516 (N_516,N_235,N_194);
and U517 (N_517,N_288,N_483);
and U518 (N_518,N_250,N_57);
nor U519 (N_519,N_185,N_466);
and U520 (N_520,N_166,N_31);
xnor U521 (N_521,N_252,N_477);
nand U522 (N_522,N_375,N_156);
or U523 (N_523,N_497,N_8);
or U524 (N_524,N_88,N_404);
and U525 (N_525,N_382,N_219);
or U526 (N_526,N_323,N_26);
nand U527 (N_527,N_260,N_475);
or U528 (N_528,N_123,N_415);
and U529 (N_529,N_189,N_262);
nand U530 (N_530,N_313,N_168);
and U531 (N_531,N_271,N_198);
nor U532 (N_532,N_264,N_277);
nand U533 (N_533,N_238,N_261);
and U534 (N_534,N_308,N_10);
and U535 (N_535,N_329,N_473);
nor U536 (N_536,N_312,N_398);
nor U537 (N_537,N_287,N_224);
or U538 (N_538,N_469,N_414);
nor U539 (N_539,N_315,N_208);
nor U540 (N_540,N_93,N_392);
nor U541 (N_541,N_474,N_41);
or U542 (N_542,N_139,N_309);
or U543 (N_543,N_131,N_267);
nor U544 (N_544,N_339,N_22);
xor U545 (N_545,N_396,N_217);
xnor U546 (N_546,N_338,N_316);
or U547 (N_547,N_448,N_306);
or U548 (N_548,N_92,N_12);
nor U549 (N_549,N_11,N_207);
nor U550 (N_550,N_162,N_321);
and U551 (N_551,N_154,N_257);
nor U552 (N_552,N_62,N_245);
and U553 (N_553,N_80,N_301);
xor U554 (N_554,N_244,N_40);
nand U555 (N_555,N_221,N_351);
nand U556 (N_556,N_322,N_455);
nor U557 (N_557,N_109,N_328);
or U558 (N_558,N_494,N_52);
or U559 (N_559,N_424,N_228);
xor U560 (N_560,N_176,N_412);
and U561 (N_561,N_326,N_478);
or U562 (N_562,N_370,N_56);
or U563 (N_563,N_201,N_492);
or U564 (N_564,N_425,N_128);
nand U565 (N_565,N_101,N_319);
or U566 (N_566,N_220,N_96);
or U567 (N_567,N_355,N_349);
or U568 (N_568,N_278,N_141);
nand U569 (N_569,N_268,N_479);
nor U570 (N_570,N_119,N_366);
nor U571 (N_571,N_318,N_68);
and U572 (N_572,N_361,N_37);
nand U573 (N_573,N_389,N_114);
and U574 (N_574,N_305,N_155);
and U575 (N_575,N_85,N_51);
or U576 (N_576,N_243,N_134);
xnor U577 (N_577,N_303,N_439);
or U578 (N_578,N_405,N_112);
nand U579 (N_579,N_387,N_472);
nor U580 (N_580,N_100,N_451);
xnor U581 (N_581,N_15,N_458);
xor U582 (N_582,N_274,N_350);
nand U583 (N_583,N_54,N_307);
or U584 (N_584,N_324,N_95);
and U585 (N_585,N_47,N_143);
and U586 (N_586,N_44,N_340);
or U587 (N_587,N_369,N_6);
nand U588 (N_588,N_77,N_342);
nor U589 (N_589,N_39,N_55);
nor U590 (N_590,N_4,N_280);
nor U591 (N_591,N_499,N_437);
nand U592 (N_592,N_222,N_188);
or U593 (N_593,N_391,N_358);
and U594 (N_594,N_460,N_202);
nand U595 (N_595,N_86,N_233);
nor U596 (N_596,N_468,N_276);
nand U597 (N_597,N_330,N_171);
nand U598 (N_598,N_124,N_152);
and U599 (N_599,N_317,N_447);
and U600 (N_600,N_18,N_476);
nor U601 (N_601,N_442,N_362);
or U602 (N_602,N_258,N_106);
and U603 (N_603,N_43,N_314);
nand U604 (N_604,N_334,N_163);
nor U605 (N_605,N_285,N_402);
nor U606 (N_606,N_140,N_78);
nand U607 (N_607,N_368,N_103);
or U608 (N_608,N_489,N_408);
or U609 (N_609,N_270,N_311);
or U610 (N_610,N_117,N_373);
nor U611 (N_611,N_122,N_429);
xnor U612 (N_612,N_2,N_331);
or U613 (N_613,N_50,N_133);
nand U614 (N_614,N_32,N_269);
or U615 (N_615,N_486,N_359);
nor U616 (N_616,N_121,N_304);
nand U617 (N_617,N_399,N_230);
nor U618 (N_618,N_147,N_191);
nor U619 (N_619,N_407,N_223);
and U620 (N_620,N_102,N_71);
and U621 (N_621,N_94,N_495);
nand U622 (N_622,N_81,N_403);
nor U623 (N_623,N_496,N_430);
nand U624 (N_624,N_192,N_169);
or U625 (N_625,N_246,N_416);
nor U626 (N_626,N_241,N_173);
xor U627 (N_627,N_218,N_428);
and U628 (N_628,N_248,N_33);
nor U629 (N_629,N_213,N_360);
and U630 (N_630,N_367,N_376);
nand U631 (N_631,N_127,N_423);
xor U632 (N_632,N_378,N_175);
and U633 (N_633,N_279,N_167);
xnor U634 (N_634,N_104,N_421);
and U635 (N_635,N_129,N_199);
xnor U636 (N_636,N_108,N_413);
and U637 (N_637,N_291,N_263);
nor U638 (N_638,N_209,N_247);
or U639 (N_639,N_178,N_254);
nand U640 (N_640,N_34,N_471);
nor U641 (N_641,N_197,N_181);
nor U642 (N_642,N_281,N_422);
nand U643 (N_643,N_299,N_27);
nand U644 (N_644,N_153,N_165);
nor U645 (N_645,N_137,N_225);
or U646 (N_646,N_464,N_381);
xor U647 (N_647,N_111,N_353);
nor U648 (N_648,N_75,N_98);
and U649 (N_649,N_325,N_142);
and U650 (N_650,N_174,N_84);
nor U651 (N_651,N_180,N_23);
or U652 (N_652,N_357,N_35);
xnor U653 (N_653,N_240,N_384);
nor U654 (N_654,N_498,N_431);
and U655 (N_655,N_16,N_292);
nor U656 (N_656,N_177,N_25);
or U657 (N_657,N_388,N_470);
or U658 (N_658,N_184,N_30);
xor U659 (N_659,N_226,N_148);
or U660 (N_660,N_371,N_186);
or U661 (N_661,N_249,N_3);
or U662 (N_662,N_14,N_255);
or U663 (N_663,N_193,N_42);
xnor U664 (N_664,N_345,N_426);
nor U665 (N_665,N_151,N_487);
or U666 (N_666,N_17,N_253);
xnor U667 (N_667,N_456,N_83);
nor U668 (N_668,N_344,N_294);
and U669 (N_669,N_132,N_73);
xor U670 (N_670,N_236,N_206);
and U671 (N_671,N_70,N_237);
nand U672 (N_672,N_195,N_449);
nor U673 (N_673,N_406,N_20);
nor U674 (N_674,N_365,N_239);
and U675 (N_675,N_214,N_190);
nor U676 (N_676,N_211,N_461);
and U677 (N_677,N_69,N_289);
and U678 (N_678,N_256,N_283);
or U679 (N_679,N_13,N_467);
nand U680 (N_680,N_66,N_432);
nor U681 (N_681,N_157,N_182);
nor U682 (N_682,N_462,N_136);
and U683 (N_683,N_296,N_302);
or U684 (N_684,N_266,N_463);
or U685 (N_685,N_29,N_282);
nand U686 (N_686,N_227,N_452);
and U687 (N_687,N_215,N_210);
and U688 (N_688,N_24,N_161);
or U689 (N_689,N_205,N_337);
nand U690 (N_690,N_297,N_273);
nor U691 (N_691,N_386,N_441);
and U692 (N_692,N_67,N_187);
xnor U693 (N_693,N_286,N_410);
xnor U694 (N_694,N_146,N_440);
and U695 (N_695,N_457,N_231);
nand U696 (N_696,N_58,N_395);
or U697 (N_697,N_265,N_481);
xor U698 (N_698,N_484,N_356);
and U699 (N_699,N_135,N_295);
xnor U700 (N_700,N_450,N_144);
or U701 (N_701,N_7,N_59);
nand U702 (N_702,N_401,N_126);
nand U703 (N_703,N_36,N_107);
nor U704 (N_704,N_374,N_380);
or U705 (N_705,N_411,N_364);
nand U706 (N_706,N_453,N_170);
nor U707 (N_707,N_179,N_443);
or U708 (N_708,N_183,N_120);
xor U709 (N_709,N_74,N_9);
and U710 (N_710,N_372,N_310);
and U711 (N_711,N_89,N_343);
nand U712 (N_712,N_158,N_138);
nand U713 (N_713,N_293,N_49);
or U714 (N_714,N_490,N_409);
nand U715 (N_715,N_485,N_79);
or U716 (N_716,N_196,N_346);
nand U717 (N_717,N_445,N_38);
nand U718 (N_718,N_438,N_393);
and U719 (N_719,N_383,N_125);
nor U720 (N_720,N_115,N_459);
or U721 (N_721,N_164,N_45);
nor U722 (N_722,N_336,N_145);
nor U723 (N_723,N_46,N_53);
and U724 (N_724,N_150,N_352);
and U725 (N_725,N_1,N_272);
nor U726 (N_726,N_397,N_480);
nor U727 (N_727,N_130,N_60);
nor U728 (N_728,N_200,N_204);
and U729 (N_729,N_5,N_444);
nor U730 (N_730,N_63,N_400);
nand U731 (N_731,N_379,N_113);
or U732 (N_732,N_72,N_348);
nor U733 (N_733,N_433,N_251);
or U734 (N_734,N_232,N_327);
and U735 (N_735,N_298,N_454);
or U736 (N_736,N_332,N_0);
or U737 (N_737,N_212,N_491);
nand U738 (N_738,N_91,N_436);
or U739 (N_739,N_377,N_347);
or U740 (N_740,N_335,N_434);
nand U741 (N_741,N_435,N_488);
nor U742 (N_742,N_482,N_300);
or U743 (N_743,N_87,N_82);
nand U744 (N_744,N_203,N_76);
nor U745 (N_745,N_97,N_320);
nor U746 (N_746,N_90,N_385);
nand U747 (N_747,N_21,N_394);
nand U748 (N_748,N_116,N_172);
and U749 (N_749,N_105,N_427);
and U750 (N_750,N_91,N_128);
and U751 (N_751,N_60,N_246);
or U752 (N_752,N_26,N_110);
or U753 (N_753,N_70,N_320);
nand U754 (N_754,N_365,N_398);
and U755 (N_755,N_112,N_116);
nor U756 (N_756,N_403,N_13);
or U757 (N_757,N_218,N_330);
and U758 (N_758,N_68,N_370);
xor U759 (N_759,N_154,N_385);
or U760 (N_760,N_140,N_478);
nor U761 (N_761,N_224,N_105);
nor U762 (N_762,N_119,N_65);
nor U763 (N_763,N_480,N_23);
nand U764 (N_764,N_487,N_53);
and U765 (N_765,N_97,N_134);
nand U766 (N_766,N_242,N_376);
or U767 (N_767,N_200,N_179);
nand U768 (N_768,N_251,N_293);
nor U769 (N_769,N_403,N_466);
or U770 (N_770,N_424,N_295);
or U771 (N_771,N_354,N_312);
nand U772 (N_772,N_390,N_332);
nand U773 (N_773,N_38,N_175);
nand U774 (N_774,N_327,N_169);
nor U775 (N_775,N_476,N_254);
nand U776 (N_776,N_363,N_285);
nand U777 (N_777,N_360,N_175);
and U778 (N_778,N_25,N_348);
and U779 (N_779,N_474,N_486);
nand U780 (N_780,N_321,N_456);
and U781 (N_781,N_139,N_236);
nand U782 (N_782,N_261,N_375);
or U783 (N_783,N_25,N_165);
nand U784 (N_784,N_202,N_424);
or U785 (N_785,N_268,N_47);
nand U786 (N_786,N_323,N_277);
and U787 (N_787,N_128,N_12);
or U788 (N_788,N_365,N_169);
and U789 (N_789,N_37,N_357);
nand U790 (N_790,N_212,N_381);
xor U791 (N_791,N_362,N_188);
nor U792 (N_792,N_32,N_346);
or U793 (N_793,N_85,N_184);
and U794 (N_794,N_131,N_362);
nand U795 (N_795,N_337,N_294);
nand U796 (N_796,N_102,N_54);
nor U797 (N_797,N_1,N_283);
xnor U798 (N_798,N_40,N_193);
nand U799 (N_799,N_81,N_13);
and U800 (N_800,N_244,N_468);
or U801 (N_801,N_20,N_25);
and U802 (N_802,N_10,N_331);
nand U803 (N_803,N_484,N_35);
and U804 (N_804,N_369,N_347);
or U805 (N_805,N_390,N_310);
nor U806 (N_806,N_41,N_462);
nor U807 (N_807,N_274,N_434);
nor U808 (N_808,N_324,N_371);
and U809 (N_809,N_191,N_354);
or U810 (N_810,N_347,N_92);
nor U811 (N_811,N_5,N_74);
or U812 (N_812,N_329,N_203);
nor U813 (N_813,N_158,N_163);
nand U814 (N_814,N_160,N_246);
or U815 (N_815,N_330,N_366);
and U816 (N_816,N_89,N_373);
nor U817 (N_817,N_145,N_282);
and U818 (N_818,N_424,N_169);
and U819 (N_819,N_76,N_237);
and U820 (N_820,N_130,N_76);
and U821 (N_821,N_22,N_273);
nand U822 (N_822,N_245,N_85);
or U823 (N_823,N_31,N_416);
xnor U824 (N_824,N_443,N_280);
nor U825 (N_825,N_476,N_235);
nor U826 (N_826,N_47,N_177);
and U827 (N_827,N_399,N_104);
nand U828 (N_828,N_344,N_2);
or U829 (N_829,N_173,N_397);
nor U830 (N_830,N_428,N_403);
and U831 (N_831,N_97,N_17);
xnor U832 (N_832,N_79,N_39);
nor U833 (N_833,N_298,N_396);
nor U834 (N_834,N_260,N_309);
or U835 (N_835,N_365,N_339);
nor U836 (N_836,N_185,N_332);
nor U837 (N_837,N_172,N_281);
nor U838 (N_838,N_366,N_317);
and U839 (N_839,N_408,N_45);
nand U840 (N_840,N_471,N_347);
or U841 (N_841,N_467,N_452);
nor U842 (N_842,N_26,N_479);
nor U843 (N_843,N_227,N_51);
nand U844 (N_844,N_195,N_179);
xnor U845 (N_845,N_334,N_217);
nand U846 (N_846,N_244,N_16);
nor U847 (N_847,N_216,N_175);
or U848 (N_848,N_395,N_423);
xor U849 (N_849,N_88,N_485);
xnor U850 (N_850,N_363,N_367);
nand U851 (N_851,N_408,N_248);
and U852 (N_852,N_72,N_324);
and U853 (N_853,N_193,N_428);
and U854 (N_854,N_421,N_15);
and U855 (N_855,N_78,N_336);
or U856 (N_856,N_41,N_179);
nand U857 (N_857,N_209,N_100);
nand U858 (N_858,N_121,N_265);
and U859 (N_859,N_450,N_168);
nor U860 (N_860,N_356,N_394);
xor U861 (N_861,N_392,N_75);
nor U862 (N_862,N_14,N_290);
and U863 (N_863,N_109,N_137);
nor U864 (N_864,N_336,N_483);
and U865 (N_865,N_399,N_312);
and U866 (N_866,N_221,N_433);
nor U867 (N_867,N_442,N_284);
and U868 (N_868,N_253,N_478);
and U869 (N_869,N_78,N_48);
or U870 (N_870,N_35,N_445);
nor U871 (N_871,N_186,N_221);
or U872 (N_872,N_380,N_195);
and U873 (N_873,N_178,N_176);
nand U874 (N_874,N_186,N_408);
and U875 (N_875,N_198,N_290);
nand U876 (N_876,N_145,N_122);
or U877 (N_877,N_470,N_183);
nor U878 (N_878,N_63,N_332);
nor U879 (N_879,N_230,N_268);
and U880 (N_880,N_54,N_257);
nand U881 (N_881,N_112,N_124);
and U882 (N_882,N_161,N_448);
and U883 (N_883,N_371,N_202);
nand U884 (N_884,N_4,N_381);
nand U885 (N_885,N_118,N_460);
nand U886 (N_886,N_380,N_100);
xnor U887 (N_887,N_486,N_72);
or U888 (N_888,N_333,N_137);
nand U889 (N_889,N_399,N_120);
or U890 (N_890,N_119,N_246);
or U891 (N_891,N_413,N_324);
nor U892 (N_892,N_345,N_171);
nor U893 (N_893,N_42,N_113);
xor U894 (N_894,N_436,N_447);
and U895 (N_895,N_155,N_85);
nor U896 (N_896,N_422,N_259);
nor U897 (N_897,N_147,N_233);
and U898 (N_898,N_198,N_326);
xnor U899 (N_899,N_447,N_28);
or U900 (N_900,N_367,N_53);
nor U901 (N_901,N_389,N_493);
or U902 (N_902,N_81,N_462);
nor U903 (N_903,N_54,N_232);
xnor U904 (N_904,N_307,N_200);
and U905 (N_905,N_196,N_114);
and U906 (N_906,N_37,N_294);
nand U907 (N_907,N_465,N_296);
or U908 (N_908,N_318,N_124);
and U909 (N_909,N_274,N_257);
and U910 (N_910,N_314,N_309);
nand U911 (N_911,N_427,N_64);
or U912 (N_912,N_465,N_33);
and U913 (N_913,N_453,N_294);
nand U914 (N_914,N_140,N_340);
nor U915 (N_915,N_129,N_73);
nand U916 (N_916,N_179,N_404);
and U917 (N_917,N_11,N_430);
nor U918 (N_918,N_142,N_347);
and U919 (N_919,N_354,N_132);
nor U920 (N_920,N_467,N_221);
and U921 (N_921,N_301,N_200);
nor U922 (N_922,N_4,N_205);
xor U923 (N_923,N_65,N_405);
nor U924 (N_924,N_187,N_289);
xnor U925 (N_925,N_124,N_39);
nand U926 (N_926,N_345,N_201);
nor U927 (N_927,N_329,N_72);
nand U928 (N_928,N_370,N_340);
xor U929 (N_929,N_106,N_189);
nor U930 (N_930,N_393,N_280);
or U931 (N_931,N_368,N_482);
nand U932 (N_932,N_462,N_157);
and U933 (N_933,N_285,N_44);
or U934 (N_934,N_365,N_424);
and U935 (N_935,N_172,N_205);
and U936 (N_936,N_67,N_481);
nand U937 (N_937,N_55,N_41);
nand U938 (N_938,N_10,N_75);
nor U939 (N_939,N_377,N_76);
and U940 (N_940,N_89,N_289);
or U941 (N_941,N_293,N_225);
xor U942 (N_942,N_294,N_48);
nor U943 (N_943,N_316,N_96);
or U944 (N_944,N_7,N_285);
and U945 (N_945,N_323,N_124);
and U946 (N_946,N_88,N_295);
nor U947 (N_947,N_63,N_100);
or U948 (N_948,N_497,N_238);
nand U949 (N_949,N_53,N_225);
nor U950 (N_950,N_223,N_21);
nor U951 (N_951,N_381,N_90);
or U952 (N_952,N_55,N_448);
or U953 (N_953,N_414,N_111);
nor U954 (N_954,N_121,N_319);
nand U955 (N_955,N_42,N_151);
and U956 (N_956,N_107,N_139);
nand U957 (N_957,N_405,N_135);
or U958 (N_958,N_361,N_29);
nor U959 (N_959,N_292,N_208);
nor U960 (N_960,N_353,N_150);
and U961 (N_961,N_388,N_366);
nand U962 (N_962,N_171,N_299);
or U963 (N_963,N_116,N_348);
or U964 (N_964,N_194,N_221);
nand U965 (N_965,N_347,N_499);
and U966 (N_966,N_0,N_59);
xnor U967 (N_967,N_14,N_316);
nor U968 (N_968,N_212,N_306);
and U969 (N_969,N_477,N_383);
nor U970 (N_970,N_21,N_456);
and U971 (N_971,N_440,N_168);
nand U972 (N_972,N_109,N_388);
nor U973 (N_973,N_134,N_470);
or U974 (N_974,N_239,N_166);
nor U975 (N_975,N_203,N_469);
or U976 (N_976,N_307,N_74);
or U977 (N_977,N_318,N_412);
and U978 (N_978,N_215,N_216);
and U979 (N_979,N_153,N_114);
nor U980 (N_980,N_220,N_400);
nand U981 (N_981,N_353,N_200);
or U982 (N_982,N_95,N_298);
or U983 (N_983,N_438,N_285);
nor U984 (N_984,N_378,N_62);
xnor U985 (N_985,N_245,N_449);
or U986 (N_986,N_261,N_307);
and U987 (N_987,N_424,N_82);
or U988 (N_988,N_412,N_253);
nand U989 (N_989,N_142,N_472);
nand U990 (N_990,N_189,N_405);
nand U991 (N_991,N_247,N_220);
nor U992 (N_992,N_131,N_51);
or U993 (N_993,N_447,N_356);
and U994 (N_994,N_139,N_353);
nor U995 (N_995,N_260,N_231);
nand U996 (N_996,N_325,N_427);
and U997 (N_997,N_487,N_450);
and U998 (N_998,N_429,N_15);
and U999 (N_999,N_320,N_256);
nor U1000 (N_1000,N_958,N_952);
nand U1001 (N_1001,N_734,N_939);
or U1002 (N_1002,N_873,N_797);
and U1003 (N_1003,N_747,N_905);
or U1004 (N_1004,N_779,N_940);
or U1005 (N_1005,N_613,N_578);
and U1006 (N_1006,N_677,N_833);
nor U1007 (N_1007,N_997,N_615);
xor U1008 (N_1008,N_549,N_519);
nand U1009 (N_1009,N_991,N_913);
xnor U1010 (N_1010,N_619,N_592);
nor U1011 (N_1011,N_612,N_564);
nand U1012 (N_1012,N_528,N_941);
and U1013 (N_1013,N_646,N_688);
nand U1014 (N_1014,N_978,N_740);
nor U1015 (N_1015,N_644,N_815);
and U1016 (N_1016,N_543,N_681);
or U1017 (N_1017,N_778,N_938);
nor U1018 (N_1018,N_785,N_822);
xnor U1019 (N_1019,N_558,N_553);
nor U1020 (N_1020,N_632,N_949);
and U1021 (N_1021,N_979,N_783);
and U1022 (N_1022,N_853,N_525);
nor U1023 (N_1023,N_561,N_529);
and U1024 (N_1024,N_977,N_879);
and U1025 (N_1025,N_934,N_864);
nand U1026 (N_1026,N_523,N_899);
and U1027 (N_1027,N_511,N_607);
and U1028 (N_1028,N_568,N_826);
nand U1029 (N_1029,N_507,N_774);
nand U1030 (N_1030,N_965,N_686);
and U1031 (N_1031,N_577,N_841);
nand U1032 (N_1032,N_936,N_522);
xor U1033 (N_1033,N_526,N_933);
and U1034 (N_1034,N_626,N_857);
nor U1035 (N_1035,N_699,N_521);
or U1036 (N_1036,N_673,N_658);
or U1037 (N_1037,N_791,N_571);
nand U1038 (N_1038,N_671,N_995);
or U1039 (N_1039,N_627,N_888);
nand U1040 (N_1040,N_756,N_987);
or U1041 (N_1041,N_884,N_892);
or U1042 (N_1042,N_618,N_812);
nor U1043 (N_1043,N_794,N_737);
nand U1044 (N_1044,N_817,N_844);
and U1045 (N_1045,N_945,N_551);
nand U1046 (N_1046,N_559,N_806);
or U1047 (N_1047,N_852,N_832);
and U1048 (N_1048,N_775,N_517);
or U1049 (N_1049,N_924,N_788);
xnor U1050 (N_1050,N_847,N_611);
nand U1051 (N_1051,N_849,N_850);
nor U1052 (N_1052,N_556,N_862);
nand U1053 (N_1053,N_895,N_754);
xnor U1054 (N_1054,N_750,N_777);
xnor U1055 (N_1055,N_620,N_982);
nand U1056 (N_1056,N_983,N_657);
and U1057 (N_1057,N_891,N_917);
or U1058 (N_1058,N_947,N_973);
nand U1059 (N_1059,N_880,N_769);
xnor U1060 (N_1060,N_859,N_856);
or U1061 (N_1061,N_565,N_836);
xnor U1062 (N_1062,N_961,N_547);
and U1063 (N_1063,N_825,N_820);
and U1064 (N_1064,N_953,N_903);
or U1065 (N_1065,N_690,N_871);
or U1066 (N_1066,N_911,N_759);
or U1067 (N_1067,N_683,N_799);
or U1068 (N_1068,N_972,N_868);
xnor U1069 (N_1069,N_649,N_638);
and U1070 (N_1070,N_996,N_976);
nand U1071 (N_1071,N_594,N_744);
and U1072 (N_1072,N_567,N_725);
nand U1073 (N_1073,N_893,N_942);
nor U1074 (N_1074,N_544,N_539);
and U1075 (N_1075,N_541,N_703);
or U1076 (N_1076,N_918,N_730);
nor U1077 (N_1077,N_610,N_957);
or U1078 (N_1078,N_697,N_768);
nand U1079 (N_1079,N_712,N_804);
and U1080 (N_1080,N_717,N_647);
xnor U1081 (N_1081,N_555,N_925);
nand U1082 (N_1082,N_763,N_998);
nand U1083 (N_1083,N_716,N_886);
and U1084 (N_1084,N_727,N_729);
nor U1085 (N_1085,N_574,N_513);
nor U1086 (N_1086,N_838,N_802);
nand U1087 (N_1087,N_732,N_524);
or U1088 (N_1088,N_660,N_629);
nand U1089 (N_1089,N_676,N_557);
nand U1090 (N_1090,N_731,N_509);
nor U1091 (N_1091,N_645,N_869);
or U1092 (N_1092,N_764,N_890);
nand U1093 (N_1093,N_948,N_811);
nand U1094 (N_1094,N_767,N_994);
or U1095 (N_1095,N_711,N_927);
or U1096 (N_1096,N_714,N_531);
and U1097 (N_1097,N_707,N_969);
or U1098 (N_1098,N_596,N_598);
nand U1099 (N_1099,N_861,N_602);
xnor U1100 (N_1100,N_765,N_622);
xor U1101 (N_1101,N_614,N_663);
xor U1102 (N_1102,N_661,N_692);
nand U1103 (N_1103,N_664,N_828);
nand U1104 (N_1104,N_776,N_789);
and U1105 (N_1105,N_784,N_700);
nand U1106 (N_1106,N_937,N_854);
nor U1107 (N_1107,N_781,N_746);
nand U1108 (N_1108,N_993,N_971);
and U1109 (N_1109,N_719,N_516);
or U1110 (N_1110,N_851,N_741);
or U1111 (N_1111,N_538,N_621);
xor U1112 (N_1112,N_989,N_751);
nand U1113 (N_1113,N_944,N_720);
nor U1114 (N_1114,N_867,N_588);
nand U1115 (N_1115,N_846,N_634);
xor U1116 (N_1116,N_668,N_882);
nand U1117 (N_1117,N_824,N_816);
nand U1118 (N_1118,N_883,N_562);
nor U1119 (N_1119,N_687,N_742);
nand U1120 (N_1120,N_738,N_837);
and U1121 (N_1121,N_827,N_748);
xnor U1122 (N_1122,N_921,N_582);
nor U1123 (N_1123,N_623,N_809);
or U1124 (N_1124,N_819,N_510);
nand U1125 (N_1125,N_653,N_518);
or U1126 (N_1126,N_520,N_585);
nand U1127 (N_1127,N_810,N_504);
nand U1128 (N_1128,N_662,N_902);
xnor U1129 (N_1129,N_943,N_967);
nor U1130 (N_1130,N_694,N_753);
or U1131 (N_1131,N_684,N_855);
nand U1132 (N_1132,N_984,N_915);
or U1133 (N_1133,N_569,N_752);
nand U1134 (N_1134,N_566,N_665);
xor U1135 (N_1135,N_723,N_900);
nand U1136 (N_1136,N_845,N_515);
and U1137 (N_1137,N_843,N_502);
or U1138 (N_1138,N_670,N_839);
and U1139 (N_1139,N_563,N_758);
or U1140 (N_1140,N_975,N_709);
and U1141 (N_1141,N_616,N_704);
nand U1142 (N_1142,N_587,N_534);
nor U1143 (N_1143,N_575,N_573);
nand U1144 (N_1144,N_930,N_887);
or U1145 (N_1145,N_666,N_985);
nor U1146 (N_1146,N_675,N_793);
or U1147 (N_1147,N_757,N_878);
or U1148 (N_1148,N_652,N_550);
and U1149 (N_1149,N_689,N_922);
or U1150 (N_1150,N_505,N_710);
nand U1151 (N_1151,N_964,N_698);
and U1152 (N_1152,N_705,N_894);
or U1153 (N_1153,N_637,N_795);
or U1154 (N_1154,N_735,N_914);
or U1155 (N_1155,N_678,N_858);
nand U1156 (N_1156,N_885,N_693);
or U1157 (N_1157,N_749,N_728);
and U1158 (N_1158,N_625,N_591);
or U1159 (N_1159,N_916,N_796);
and U1160 (N_1160,N_935,N_724);
xnor U1161 (N_1161,N_552,N_818);
nand U1162 (N_1162,N_980,N_907);
nand U1163 (N_1163,N_896,N_651);
nand U1164 (N_1164,N_990,N_981);
xnor U1165 (N_1165,N_722,N_954);
nor U1166 (N_1166,N_908,N_786);
and U1167 (N_1167,N_624,N_926);
and U1168 (N_1168,N_560,N_956);
nand U1169 (N_1169,N_805,N_875);
xnor U1170 (N_1170,N_766,N_963);
or U1171 (N_1171,N_733,N_514);
or U1172 (N_1172,N_576,N_955);
or U1173 (N_1173,N_606,N_608);
xor U1174 (N_1174,N_590,N_901);
nand U1175 (N_1175,N_770,N_848);
and U1176 (N_1176,N_881,N_530);
nor U1177 (N_1177,N_912,N_628);
nand U1178 (N_1178,N_701,N_721);
nand U1179 (N_1179,N_920,N_842);
or U1180 (N_1180,N_674,N_503);
nand U1181 (N_1181,N_762,N_792);
xor U1182 (N_1182,N_780,N_581);
xor U1183 (N_1183,N_572,N_589);
and U1184 (N_1184,N_960,N_506);
or U1185 (N_1185,N_597,N_772);
nor U1186 (N_1186,N_713,N_708);
or U1187 (N_1187,N_876,N_910);
nor U1188 (N_1188,N_546,N_702);
nor U1189 (N_1189,N_966,N_593);
and U1190 (N_1190,N_872,N_814);
or U1191 (N_1191,N_760,N_874);
nand U1192 (N_1192,N_715,N_527);
xor U1193 (N_1193,N_834,N_609);
nor U1194 (N_1194,N_648,N_898);
nor U1195 (N_1195,N_821,N_761);
nand U1196 (N_1196,N_743,N_974);
and U1197 (N_1197,N_928,N_840);
xnor U1198 (N_1198,N_535,N_823);
xnor U1199 (N_1199,N_669,N_736);
nand U1200 (N_1200,N_512,N_605);
and U1201 (N_1201,N_798,N_755);
nand U1202 (N_1202,N_642,N_641);
nor U1203 (N_1203,N_679,N_706);
or U1204 (N_1204,N_508,N_580);
and U1205 (N_1205,N_863,N_931);
and U1206 (N_1206,N_932,N_617);
nand U1207 (N_1207,N_680,N_542);
nand U1208 (N_1208,N_808,N_595);
xnor U1209 (N_1209,N_790,N_800);
and U1210 (N_1210,N_548,N_501);
nor U1211 (N_1211,N_829,N_691);
or U1212 (N_1212,N_787,N_570);
or U1213 (N_1213,N_654,N_537);
and U1214 (N_1214,N_601,N_959);
xnor U1215 (N_1215,N_659,N_636);
and U1216 (N_1216,N_682,N_919);
xnor U1217 (N_1217,N_771,N_532);
and U1218 (N_1218,N_831,N_865);
nor U1219 (N_1219,N_946,N_639);
nor U1220 (N_1220,N_860,N_726);
and U1221 (N_1221,N_745,N_635);
or U1222 (N_1222,N_667,N_603);
and U1223 (N_1223,N_500,N_718);
nor U1224 (N_1224,N_929,N_870);
or U1225 (N_1225,N_904,N_604);
nand U1226 (N_1226,N_579,N_889);
or U1227 (N_1227,N_672,N_813);
and U1228 (N_1228,N_968,N_962);
nand U1229 (N_1229,N_951,N_999);
or U1230 (N_1230,N_773,N_584);
nor U1231 (N_1231,N_631,N_643);
or U1232 (N_1232,N_782,N_803);
and U1233 (N_1233,N_897,N_540);
and U1234 (N_1234,N_650,N_630);
nand U1235 (N_1235,N_583,N_554);
and U1236 (N_1236,N_533,N_835);
or U1237 (N_1237,N_656,N_970);
nor U1238 (N_1238,N_640,N_633);
nor U1239 (N_1239,N_600,N_739);
and U1240 (N_1240,N_685,N_988);
nor U1241 (N_1241,N_696,N_909);
nand U1242 (N_1242,N_950,N_536);
nor U1243 (N_1243,N_992,N_695);
or U1244 (N_1244,N_586,N_599);
nor U1245 (N_1245,N_545,N_906);
nand U1246 (N_1246,N_923,N_986);
and U1247 (N_1247,N_807,N_830);
nand U1248 (N_1248,N_655,N_877);
and U1249 (N_1249,N_866,N_801);
and U1250 (N_1250,N_548,N_500);
and U1251 (N_1251,N_760,N_962);
or U1252 (N_1252,N_632,N_699);
nor U1253 (N_1253,N_652,N_947);
nor U1254 (N_1254,N_958,N_515);
nand U1255 (N_1255,N_929,N_857);
or U1256 (N_1256,N_890,N_671);
nor U1257 (N_1257,N_834,N_686);
or U1258 (N_1258,N_676,N_958);
xnor U1259 (N_1259,N_888,N_775);
nand U1260 (N_1260,N_517,N_982);
or U1261 (N_1261,N_845,N_542);
and U1262 (N_1262,N_978,N_767);
nand U1263 (N_1263,N_652,N_600);
nand U1264 (N_1264,N_894,N_844);
and U1265 (N_1265,N_803,N_603);
and U1266 (N_1266,N_628,N_769);
nand U1267 (N_1267,N_503,N_899);
nand U1268 (N_1268,N_563,N_588);
nand U1269 (N_1269,N_722,N_626);
nor U1270 (N_1270,N_828,N_721);
xnor U1271 (N_1271,N_965,N_982);
or U1272 (N_1272,N_592,N_975);
xnor U1273 (N_1273,N_815,N_637);
or U1274 (N_1274,N_631,N_634);
and U1275 (N_1275,N_680,N_670);
and U1276 (N_1276,N_514,N_511);
and U1277 (N_1277,N_599,N_697);
nor U1278 (N_1278,N_524,N_999);
nor U1279 (N_1279,N_668,N_923);
xor U1280 (N_1280,N_795,N_975);
xnor U1281 (N_1281,N_504,N_874);
nor U1282 (N_1282,N_719,N_752);
nand U1283 (N_1283,N_700,N_655);
or U1284 (N_1284,N_789,N_921);
nand U1285 (N_1285,N_615,N_974);
nand U1286 (N_1286,N_770,N_992);
nand U1287 (N_1287,N_598,N_545);
nand U1288 (N_1288,N_745,N_551);
or U1289 (N_1289,N_865,N_734);
or U1290 (N_1290,N_572,N_966);
nand U1291 (N_1291,N_932,N_866);
or U1292 (N_1292,N_563,N_771);
or U1293 (N_1293,N_677,N_930);
nor U1294 (N_1294,N_724,N_542);
nand U1295 (N_1295,N_772,N_580);
or U1296 (N_1296,N_674,N_976);
or U1297 (N_1297,N_578,N_574);
and U1298 (N_1298,N_751,N_603);
nor U1299 (N_1299,N_861,N_917);
nor U1300 (N_1300,N_551,N_627);
and U1301 (N_1301,N_985,N_944);
xor U1302 (N_1302,N_862,N_551);
nor U1303 (N_1303,N_625,N_674);
and U1304 (N_1304,N_833,N_648);
and U1305 (N_1305,N_796,N_961);
or U1306 (N_1306,N_686,N_784);
nand U1307 (N_1307,N_814,N_783);
or U1308 (N_1308,N_765,N_938);
or U1309 (N_1309,N_866,N_886);
and U1310 (N_1310,N_517,N_940);
or U1311 (N_1311,N_612,N_540);
or U1312 (N_1312,N_865,N_788);
nor U1313 (N_1313,N_836,N_541);
and U1314 (N_1314,N_691,N_819);
nor U1315 (N_1315,N_662,N_850);
and U1316 (N_1316,N_773,N_830);
and U1317 (N_1317,N_851,N_662);
nand U1318 (N_1318,N_705,N_781);
nand U1319 (N_1319,N_736,N_688);
nor U1320 (N_1320,N_817,N_519);
xnor U1321 (N_1321,N_694,N_816);
nor U1322 (N_1322,N_817,N_686);
nand U1323 (N_1323,N_652,N_993);
nand U1324 (N_1324,N_998,N_661);
and U1325 (N_1325,N_906,N_777);
xnor U1326 (N_1326,N_525,N_644);
nand U1327 (N_1327,N_643,N_573);
nand U1328 (N_1328,N_682,N_566);
nand U1329 (N_1329,N_769,N_522);
and U1330 (N_1330,N_598,N_975);
nand U1331 (N_1331,N_830,N_786);
or U1332 (N_1332,N_650,N_660);
nand U1333 (N_1333,N_581,N_909);
and U1334 (N_1334,N_942,N_618);
nand U1335 (N_1335,N_910,N_709);
or U1336 (N_1336,N_729,N_702);
xnor U1337 (N_1337,N_563,N_603);
or U1338 (N_1338,N_907,N_768);
nand U1339 (N_1339,N_734,N_600);
nand U1340 (N_1340,N_819,N_976);
and U1341 (N_1341,N_737,N_937);
nor U1342 (N_1342,N_644,N_583);
nor U1343 (N_1343,N_576,N_865);
and U1344 (N_1344,N_972,N_820);
or U1345 (N_1345,N_859,N_883);
and U1346 (N_1346,N_797,N_533);
or U1347 (N_1347,N_796,N_717);
and U1348 (N_1348,N_822,N_900);
and U1349 (N_1349,N_936,N_527);
nand U1350 (N_1350,N_511,N_705);
xor U1351 (N_1351,N_698,N_600);
nor U1352 (N_1352,N_874,N_803);
nor U1353 (N_1353,N_964,N_741);
xor U1354 (N_1354,N_813,N_808);
nor U1355 (N_1355,N_663,N_930);
and U1356 (N_1356,N_849,N_665);
xor U1357 (N_1357,N_993,N_848);
or U1358 (N_1358,N_569,N_505);
nand U1359 (N_1359,N_696,N_786);
and U1360 (N_1360,N_984,N_513);
or U1361 (N_1361,N_827,N_716);
nand U1362 (N_1362,N_647,N_662);
nand U1363 (N_1363,N_544,N_833);
xnor U1364 (N_1364,N_702,N_656);
or U1365 (N_1365,N_677,N_509);
nand U1366 (N_1366,N_623,N_833);
or U1367 (N_1367,N_852,N_630);
and U1368 (N_1368,N_976,N_763);
nand U1369 (N_1369,N_842,N_964);
or U1370 (N_1370,N_761,N_721);
or U1371 (N_1371,N_673,N_629);
or U1372 (N_1372,N_509,N_732);
or U1373 (N_1373,N_658,N_945);
nor U1374 (N_1374,N_818,N_609);
nand U1375 (N_1375,N_674,N_927);
or U1376 (N_1376,N_834,N_842);
nand U1377 (N_1377,N_957,N_797);
or U1378 (N_1378,N_850,N_756);
nand U1379 (N_1379,N_964,N_918);
or U1380 (N_1380,N_672,N_942);
nor U1381 (N_1381,N_761,N_957);
nor U1382 (N_1382,N_504,N_558);
or U1383 (N_1383,N_615,N_670);
or U1384 (N_1384,N_716,N_532);
nor U1385 (N_1385,N_786,N_845);
xor U1386 (N_1386,N_954,N_701);
or U1387 (N_1387,N_749,N_638);
or U1388 (N_1388,N_812,N_730);
nand U1389 (N_1389,N_975,N_819);
nor U1390 (N_1390,N_944,N_883);
xnor U1391 (N_1391,N_592,N_793);
nand U1392 (N_1392,N_954,N_689);
or U1393 (N_1393,N_987,N_886);
and U1394 (N_1394,N_810,N_523);
nand U1395 (N_1395,N_553,N_988);
and U1396 (N_1396,N_878,N_606);
nor U1397 (N_1397,N_562,N_773);
nor U1398 (N_1398,N_581,N_762);
nor U1399 (N_1399,N_575,N_563);
or U1400 (N_1400,N_979,N_983);
nor U1401 (N_1401,N_530,N_735);
or U1402 (N_1402,N_713,N_631);
or U1403 (N_1403,N_562,N_719);
and U1404 (N_1404,N_762,N_728);
and U1405 (N_1405,N_684,N_859);
or U1406 (N_1406,N_591,N_689);
nand U1407 (N_1407,N_907,N_571);
nand U1408 (N_1408,N_707,N_601);
or U1409 (N_1409,N_687,N_641);
nor U1410 (N_1410,N_739,N_737);
nor U1411 (N_1411,N_861,N_549);
nor U1412 (N_1412,N_991,N_529);
or U1413 (N_1413,N_525,N_574);
and U1414 (N_1414,N_633,N_973);
nor U1415 (N_1415,N_923,N_820);
or U1416 (N_1416,N_776,N_988);
nor U1417 (N_1417,N_652,N_532);
or U1418 (N_1418,N_801,N_544);
nand U1419 (N_1419,N_795,N_773);
or U1420 (N_1420,N_948,N_894);
xor U1421 (N_1421,N_946,N_542);
xor U1422 (N_1422,N_706,N_675);
nand U1423 (N_1423,N_750,N_781);
and U1424 (N_1424,N_702,N_500);
and U1425 (N_1425,N_657,N_929);
nor U1426 (N_1426,N_546,N_897);
or U1427 (N_1427,N_926,N_632);
nand U1428 (N_1428,N_566,N_737);
or U1429 (N_1429,N_808,N_682);
or U1430 (N_1430,N_897,N_651);
or U1431 (N_1431,N_603,N_627);
xor U1432 (N_1432,N_633,N_653);
and U1433 (N_1433,N_624,N_661);
and U1434 (N_1434,N_577,N_535);
or U1435 (N_1435,N_755,N_539);
nor U1436 (N_1436,N_953,N_677);
or U1437 (N_1437,N_654,N_684);
nand U1438 (N_1438,N_517,N_866);
nor U1439 (N_1439,N_632,N_626);
nand U1440 (N_1440,N_815,N_989);
and U1441 (N_1441,N_758,N_645);
nand U1442 (N_1442,N_892,N_829);
nand U1443 (N_1443,N_592,N_933);
nor U1444 (N_1444,N_685,N_830);
nor U1445 (N_1445,N_534,N_894);
nor U1446 (N_1446,N_782,N_945);
or U1447 (N_1447,N_739,N_890);
or U1448 (N_1448,N_762,N_724);
nand U1449 (N_1449,N_934,N_671);
and U1450 (N_1450,N_851,N_928);
nand U1451 (N_1451,N_623,N_887);
or U1452 (N_1452,N_846,N_732);
nor U1453 (N_1453,N_709,N_947);
xor U1454 (N_1454,N_974,N_859);
nor U1455 (N_1455,N_688,N_920);
or U1456 (N_1456,N_667,N_793);
nor U1457 (N_1457,N_918,N_819);
and U1458 (N_1458,N_655,N_878);
or U1459 (N_1459,N_869,N_745);
nor U1460 (N_1460,N_712,N_620);
nand U1461 (N_1461,N_795,N_663);
nand U1462 (N_1462,N_635,N_590);
nor U1463 (N_1463,N_937,N_553);
or U1464 (N_1464,N_929,N_555);
and U1465 (N_1465,N_660,N_949);
or U1466 (N_1466,N_808,N_901);
and U1467 (N_1467,N_869,N_651);
nand U1468 (N_1468,N_780,N_614);
or U1469 (N_1469,N_996,N_626);
and U1470 (N_1470,N_546,N_528);
or U1471 (N_1471,N_591,N_643);
nor U1472 (N_1472,N_605,N_759);
or U1473 (N_1473,N_777,N_945);
nand U1474 (N_1474,N_916,N_518);
or U1475 (N_1475,N_860,N_531);
nor U1476 (N_1476,N_906,N_766);
or U1477 (N_1477,N_606,N_928);
or U1478 (N_1478,N_695,N_932);
nor U1479 (N_1479,N_767,N_746);
and U1480 (N_1480,N_879,N_501);
and U1481 (N_1481,N_697,N_932);
and U1482 (N_1482,N_613,N_683);
or U1483 (N_1483,N_950,N_613);
nand U1484 (N_1484,N_679,N_661);
nor U1485 (N_1485,N_661,N_574);
nor U1486 (N_1486,N_523,N_826);
or U1487 (N_1487,N_584,N_760);
xnor U1488 (N_1488,N_600,N_602);
or U1489 (N_1489,N_576,N_879);
or U1490 (N_1490,N_663,N_548);
and U1491 (N_1491,N_701,N_953);
or U1492 (N_1492,N_671,N_596);
or U1493 (N_1493,N_548,N_978);
nor U1494 (N_1494,N_956,N_509);
and U1495 (N_1495,N_559,N_950);
xor U1496 (N_1496,N_834,N_936);
nand U1497 (N_1497,N_759,N_776);
nand U1498 (N_1498,N_729,N_671);
nand U1499 (N_1499,N_616,N_947);
nand U1500 (N_1500,N_1410,N_1027);
nand U1501 (N_1501,N_1316,N_1260);
and U1502 (N_1502,N_1416,N_1230);
nand U1503 (N_1503,N_1066,N_1268);
nor U1504 (N_1504,N_1065,N_1239);
nand U1505 (N_1505,N_1366,N_1157);
xor U1506 (N_1506,N_1156,N_1058);
and U1507 (N_1507,N_1294,N_1151);
or U1508 (N_1508,N_1097,N_1202);
nor U1509 (N_1509,N_1475,N_1322);
nand U1510 (N_1510,N_1024,N_1211);
and U1511 (N_1511,N_1125,N_1367);
nand U1512 (N_1512,N_1438,N_1080);
and U1513 (N_1513,N_1484,N_1148);
and U1514 (N_1514,N_1163,N_1033);
nand U1515 (N_1515,N_1489,N_1364);
nand U1516 (N_1516,N_1266,N_1324);
or U1517 (N_1517,N_1209,N_1473);
or U1518 (N_1518,N_1098,N_1405);
and U1519 (N_1519,N_1164,N_1096);
or U1520 (N_1520,N_1441,N_1281);
nand U1521 (N_1521,N_1348,N_1375);
nor U1522 (N_1522,N_1022,N_1210);
and U1523 (N_1523,N_1253,N_1422);
nor U1524 (N_1524,N_1259,N_1464);
nor U1525 (N_1525,N_1095,N_1196);
xnor U1526 (N_1526,N_1377,N_1166);
nand U1527 (N_1527,N_1143,N_1450);
nand U1528 (N_1528,N_1068,N_1251);
nand U1529 (N_1529,N_1458,N_1289);
nand U1530 (N_1530,N_1343,N_1406);
and U1531 (N_1531,N_1387,N_1398);
nand U1532 (N_1532,N_1413,N_1250);
and U1533 (N_1533,N_1409,N_1255);
or U1534 (N_1534,N_1257,N_1352);
and U1535 (N_1535,N_1477,N_1476);
and U1536 (N_1536,N_1036,N_1113);
or U1537 (N_1537,N_1331,N_1304);
or U1538 (N_1538,N_1178,N_1386);
or U1539 (N_1539,N_1168,N_1382);
or U1540 (N_1540,N_1445,N_1173);
or U1541 (N_1541,N_1019,N_1147);
or U1542 (N_1542,N_1174,N_1182);
and U1543 (N_1543,N_1213,N_1488);
and U1544 (N_1544,N_1146,N_1224);
nand U1545 (N_1545,N_1252,N_1160);
nand U1546 (N_1546,N_1053,N_1466);
or U1547 (N_1547,N_1002,N_1244);
nand U1548 (N_1548,N_1135,N_1045);
or U1549 (N_1549,N_1309,N_1431);
and U1550 (N_1550,N_1001,N_1329);
nor U1551 (N_1551,N_1059,N_1397);
nor U1552 (N_1552,N_1225,N_1028);
or U1553 (N_1553,N_1195,N_1403);
and U1554 (N_1554,N_1313,N_1305);
or U1555 (N_1555,N_1487,N_1060);
or U1556 (N_1556,N_1279,N_1256);
and U1557 (N_1557,N_1167,N_1470);
xnor U1558 (N_1558,N_1170,N_1054);
and U1559 (N_1559,N_1355,N_1443);
or U1560 (N_1560,N_1302,N_1049);
or U1561 (N_1561,N_1379,N_1123);
and U1562 (N_1562,N_1300,N_1128);
nand U1563 (N_1563,N_1333,N_1121);
and U1564 (N_1564,N_1064,N_1463);
nor U1565 (N_1565,N_1414,N_1342);
and U1566 (N_1566,N_1393,N_1437);
or U1567 (N_1567,N_1076,N_1479);
nand U1568 (N_1568,N_1424,N_1310);
xnor U1569 (N_1569,N_1104,N_1453);
xor U1570 (N_1570,N_1407,N_1181);
nand U1571 (N_1571,N_1234,N_1130);
and U1572 (N_1572,N_1044,N_1070);
and U1573 (N_1573,N_1042,N_1381);
and U1574 (N_1574,N_1419,N_1370);
and U1575 (N_1575,N_1353,N_1378);
nand U1576 (N_1576,N_1291,N_1275);
or U1577 (N_1577,N_1176,N_1385);
nor U1578 (N_1578,N_1103,N_1472);
nand U1579 (N_1579,N_1208,N_1047);
or U1580 (N_1580,N_1248,N_1442);
xor U1581 (N_1581,N_1184,N_1013);
nor U1582 (N_1582,N_1241,N_1344);
and U1583 (N_1583,N_1320,N_1117);
or U1584 (N_1584,N_1165,N_1292);
nor U1585 (N_1585,N_1391,N_1186);
nor U1586 (N_1586,N_1293,N_1051);
and U1587 (N_1587,N_1231,N_1287);
xnor U1588 (N_1588,N_1206,N_1242);
or U1589 (N_1589,N_1145,N_1220);
or U1590 (N_1590,N_1106,N_1152);
and U1591 (N_1591,N_1457,N_1420);
and U1592 (N_1592,N_1205,N_1188);
and U1593 (N_1593,N_1297,N_1086);
nor U1594 (N_1594,N_1035,N_1183);
and U1595 (N_1595,N_1325,N_1288);
or U1596 (N_1596,N_1428,N_1057);
and U1597 (N_1597,N_1228,N_1439);
nor U1598 (N_1598,N_1340,N_1417);
nor U1599 (N_1599,N_1101,N_1073);
or U1600 (N_1600,N_1011,N_1132);
nor U1601 (N_1601,N_1351,N_1021);
nor U1602 (N_1602,N_1043,N_1233);
nor U1603 (N_1603,N_1171,N_1223);
and U1604 (N_1604,N_1137,N_1278);
and U1605 (N_1605,N_1362,N_1298);
and U1606 (N_1606,N_1447,N_1238);
nor U1607 (N_1607,N_1193,N_1119);
and U1608 (N_1608,N_1478,N_1139);
xor U1609 (N_1609,N_1452,N_1109);
nor U1610 (N_1610,N_1199,N_1138);
and U1611 (N_1611,N_1454,N_1283);
or U1612 (N_1612,N_1107,N_1483);
or U1613 (N_1613,N_1460,N_1358);
and U1614 (N_1614,N_1299,N_1092);
and U1615 (N_1615,N_1020,N_1000);
or U1616 (N_1616,N_1034,N_1426);
and U1617 (N_1617,N_1079,N_1185);
nor U1618 (N_1618,N_1491,N_1069);
or U1619 (N_1619,N_1308,N_1154);
xnor U1620 (N_1620,N_1084,N_1236);
nor U1621 (N_1621,N_1235,N_1112);
nand U1622 (N_1622,N_1219,N_1081);
or U1623 (N_1623,N_1155,N_1025);
and U1624 (N_1624,N_1061,N_1161);
nand U1625 (N_1625,N_1448,N_1227);
and U1626 (N_1626,N_1421,N_1249);
nand U1627 (N_1627,N_1187,N_1031);
and U1628 (N_1628,N_1190,N_1203);
or U1629 (N_1629,N_1496,N_1306);
or U1630 (N_1630,N_1029,N_1356);
and U1631 (N_1631,N_1041,N_1087);
or U1632 (N_1632,N_1177,N_1232);
nand U1633 (N_1633,N_1380,N_1338);
nand U1634 (N_1634,N_1411,N_1039);
and U1635 (N_1635,N_1273,N_1335);
or U1636 (N_1636,N_1486,N_1179);
and U1637 (N_1637,N_1349,N_1032);
nor U1638 (N_1638,N_1245,N_1071);
or U1639 (N_1639,N_1090,N_1361);
and U1640 (N_1640,N_1451,N_1067);
or U1641 (N_1641,N_1471,N_1401);
and U1642 (N_1642,N_1493,N_1318);
or U1643 (N_1643,N_1094,N_1120);
nand U1644 (N_1644,N_1078,N_1446);
nor U1645 (N_1645,N_1267,N_1374);
nor U1646 (N_1646,N_1246,N_1400);
xor U1647 (N_1647,N_1144,N_1363);
or U1648 (N_1648,N_1074,N_1311);
nand U1649 (N_1649,N_1216,N_1383);
or U1650 (N_1650,N_1158,N_1023);
and U1651 (N_1651,N_1339,N_1394);
and U1652 (N_1652,N_1048,N_1371);
and U1653 (N_1653,N_1222,N_1492);
and U1654 (N_1654,N_1432,N_1296);
or U1655 (N_1655,N_1072,N_1347);
xnor U1656 (N_1656,N_1384,N_1323);
nand U1657 (N_1657,N_1360,N_1389);
nor U1658 (N_1658,N_1482,N_1425);
or U1659 (N_1659,N_1402,N_1328);
or U1660 (N_1660,N_1207,N_1388);
nand U1661 (N_1661,N_1142,N_1180);
nand U1662 (N_1662,N_1014,N_1277);
nand U1663 (N_1663,N_1373,N_1346);
nor U1664 (N_1664,N_1175,N_1435);
nor U1665 (N_1665,N_1404,N_1274);
or U1666 (N_1666,N_1429,N_1159);
nand U1667 (N_1667,N_1063,N_1494);
nand U1668 (N_1668,N_1110,N_1423);
nand U1669 (N_1669,N_1115,N_1485);
nor U1670 (N_1670,N_1026,N_1118);
or U1671 (N_1671,N_1007,N_1433);
and U1672 (N_1672,N_1499,N_1212);
and U1673 (N_1673,N_1136,N_1449);
and U1674 (N_1674,N_1010,N_1334);
nand U1675 (N_1675,N_1197,N_1262);
and U1676 (N_1676,N_1467,N_1462);
or U1677 (N_1677,N_1140,N_1200);
nand U1678 (N_1678,N_1469,N_1218);
and U1679 (N_1679,N_1189,N_1082);
nand U1680 (N_1680,N_1149,N_1495);
or U1681 (N_1681,N_1303,N_1263);
or U1682 (N_1682,N_1015,N_1427);
xor U1683 (N_1683,N_1192,N_1415);
xor U1684 (N_1684,N_1089,N_1396);
and U1685 (N_1685,N_1312,N_1099);
and U1686 (N_1686,N_1412,N_1271);
or U1687 (N_1687,N_1124,N_1392);
and U1688 (N_1688,N_1062,N_1172);
and U1689 (N_1689,N_1150,N_1436);
and U1690 (N_1690,N_1201,N_1075);
nor U1691 (N_1691,N_1016,N_1408);
nand U1692 (N_1692,N_1004,N_1226);
nor U1693 (N_1693,N_1102,N_1091);
and U1694 (N_1694,N_1088,N_1321);
or U1695 (N_1695,N_1214,N_1008);
or U1696 (N_1696,N_1134,N_1317);
nand U1697 (N_1697,N_1258,N_1085);
nand U1698 (N_1698,N_1127,N_1459);
nor U1699 (N_1699,N_1295,N_1114);
and U1700 (N_1700,N_1083,N_1272);
xnor U1701 (N_1701,N_1357,N_1005);
or U1702 (N_1702,N_1198,N_1133);
nor U1703 (N_1703,N_1399,N_1307);
or U1704 (N_1704,N_1395,N_1261);
and U1705 (N_1705,N_1116,N_1003);
or U1706 (N_1706,N_1490,N_1129);
or U1707 (N_1707,N_1037,N_1430);
nand U1708 (N_1708,N_1017,N_1055);
nand U1709 (N_1709,N_1350,N_1354);
and U1710 (N_1710,N_1265,N_1365);
and U1711 (N_1711,N_1341,N_1012);
nand U1712 (N_1712,N_1280,N_1286);
or U1713 (N_1713,N_1243,N_1284);
and U1714 (N_1714,N_1217,N_1314);
nand U1715 (N_1715,N_1481,N_1368);
nor U1716 (N_1716,N_1326,N_1056);
nor U1717 (N_1717,N_1369,N_1204);
nand U1718 (N_1718,N_1126,N_1315);
nand U1719 (N_1719,N_1319,N_1030);
xnor U1720 (N_1720,N_1169,N_1046);
and U1721 (N_1721,N_1221,N_1247);
nor U1722 (N_1722,N_1456,N_1131);
and U1723 (N_1723,N_1285,N_1497);
nor U1724 (N_1724,N_1093,N_1162);
nand U1725 (N_1725,N_1474,N_1077);
nor U1726 (N_1726,N_1465,N_1290);
xnor U1727 (N_1727,N_1038,N_1336);
and U1728 (N_1728,N_1359,N_1376);
nor U1729 (N_1729,N_1194,N_1468);
xor U1730 (N_1730,N_1372,N_1018);
and U1731 (N_1731,N_1330,N_1332);
and U1732 (N_1732,N_1282,N_1301);
nor U1733 (N_1733,N_1461,N_1006);
nor U1734 (N_1734,N_1440,N_1498);
nand U1735 (N_1735,N_1141,N_1418);
or U1736 (N_1736,N_1264,N_1480);
or U1737 (N_1737,N_1254,N_1111);
nor U1738 (N_1738,N_1229,N_1105);
xor U1739 (N_1739,N_1444,N_1237);
and U1740 (N_1740,N_1108,N_1345);
nand U1741 (N_1741,N_1276,N_1050);
or U1742 (N_1742,N_1327,N_1270);
or U1743 (N_1743,N_1040,N_1269);
nand U1744 (N_1744,N_1434,N_1052);
nor U1745 (N_1745,N_1240,N_1153);
or U1746 (N_1746,N_1215,N_1122);
nor U1747 (N_1747,N_1009,N_1337);
and U1748 (N_1748,N_1191,N_1390);
nand U1749 (N_1749,N_1100,N_1455);
and U1750 (N_1750,N_1126,N_1428);
nor U1751 (N_1751,N_1433,N_1340);
or U1752 (N_1752,N_1149,N_1033);
nand U1753 (N_1753,N_1452,N_1021);
nor U1754 (N_1754,N_1297,N_1410);
or U1755 (N_1755,N_1205,N_1460);
nand U1756 (N_1756,N_1106,N_1003);
or U1757 (N_1757,N_1013,N_1391);
xnor U1758 (N_1758,N_1223,N_1249);
xnor U1759 (N_1759,N_1097,N_1417);
or U1760 (N_1760,N_1444,N_1268);
nor U1761 (N_1761,N_1036,N_1214);
or U1762 (N_1762,N_1289,N_1339);
or U1763 (N_1763,N_1063,N_1077);
nor U1764 (N_1764,N_1211,N_1475);
nor U1765 (N_1765,N_1130,N_1387);
nor U1766 (N_1766,N_1147,N_1314);
nor U1767 (N_1767,N_1489,N_1356);
nor U1768 (N_1768,N_1230,N_1387);
nor U1769 (N_1769,N_1413,N_1213);
nor U1770 (N_1770,N_1318,N_1083);
or U1771 (N_1771,N_1042,N_1330);
and U1772 (N_1772,N_1162,N_1417);
xor U1773 (N_1773,N_1110,N_1123);
nor U1774 (N_1774,N_1355,N_1330);
nor U1775 (N_1775,N_1380,N_1353);
nor U1776 (N_1776,N_1283,N_1217);
and U1777 (N_1777,N_1287,N_1089);
and U1778 (N_1778,N_1184,N_1152);
nand U1779 (N_1779,N_1008,N_1495);
xnor U1780 (N_1780,N_1369,N_1335);
nor U1781 (N_1781,N_1044,N_1433);
nor U1782 (N_1782,N_1379,N_1388);
nor U1783 (N_1783,N_1219,N_1039);
nor U1784 (N_1784,N_1486,N_1359);
nand U1785 (N_1785,N_1199,N_1229);
nor U1786 (N_1786,N_1457,N_1402);
nand U1787 (N_1787,N_1484,N_1319);
or U1788 (N_1788,N_1455,N_1257);
or U1789 (N_1789,N_1351,N_1205);
and U1790 (N_1790,N_1374,N_1447);
xor U1791 (N_1791,N_1421,N_1255);
nand U1792 (N_1792,N_1354,N_1040);
xnor U1793 (N_1793,N_1398,N_1457);
and U1794 (N_1794,N_1410,N_1052);
or U1795 (N_1795,N_1368,N_1383);
nand U1796 (N_1796,N_1474,N_1338);
and U1797 (N_1797,N_1408,N_1214);
or U1798 (N_1798,N_1095,N_1493);
nand U1799 (N_1799,N_1105,N_1391);
nor U1800 (N_1800,N_1020,N_1306);
and U1801 (N_1801,N_1428,N_1249);
nand U1802 (N_1802,N_1171,N_1363);
nand U1803 (N_1803,N_1272,N_1389);
xnor U1804 (N_1804,N_1121,N_1141);
or U1805 (N_1805,N_1469,N_1343);
and U1806 (N_1806,N_1078,N_1289);
xor U1807 (N_1807,N_1408,N_1430);
or U1808 (N_1808,N_1016,N_1223);
or U1809 (N_1809,N_1036,N_1398);
and U1810 (N_1810,N_1387,N_1480);
nor U1811 (N_1811,N_1003,N_1143);
and U1812 (N_1812,N_1364,N_1453);
nand U1813 (N_1813,N_1159,N_1419);
and U1814 (N_1814,N_1319,N_1465);
xnor U1815 (N_1815,N_1261,N_1103);
nand U1816 (N_1816,N_1477,N_1013);
and U1817 (N_1817,N_1244,N_1321);
and U1818 (N_1818,N_1388,N_1265);
nand U1819 (N_1819,N_1425,N_1451);
or U1820 (N_1820,N_1392,N_1237);
nand U1821 (N_1821,N_1222,N_1345);
nor U1822 (N_1822,N_1483,N_1217);
nand U1823 (N_1823,N_1448,N_1023);
or U1824 (N_1824,N_1293,N_1283);
and U1825 (N_1825,N_1117,N_1255);
and U1826 (N_1826,N_1074,N_1130);
nor U1827 (N_1827,N_1008,N_1446);
nand U1828 (N_1828,N_1190,N_1309);
nor U1829 (N_1829,N_1396,N_1235);
nand U1830 (N_1830,N_1164,N_1288);
and U1831 (N_1831,N_1177,N_1015);
or U1832 (N_1832,N_1029,N_1033);
nand U1833 (N_1833,N_1229,N_1489);
or U1834 (N_1834,N_1132,N_1317);
nor U1835 (N_1835,N_1144,N_1221);
or U1836 (N_1836,N_1444,N_1031);
nor U1837 (N_1837,N_1318,N_1195);
or U1838 (N_1838,N_1354,N_1083);
or U1839 (N_1839,N_1332,N_1227);
or U1840 (N_1840,N_1141,N_1435);
nor U1841 (N_1841,N_1338,N_1218);
xnor U1842 (N_1842,N_1473,N_1449);
nand U1843 (N_1843,N_1238,N_1212);
nor U1844 (N_1844,N_1356,N_1252);
and U1845 (N_1845,N_1380,N_1357);
or U1846 (N_1846,N_1272,N_1448);
or U1847 (N_1847,N_1274,N_1289);
or U1848 (N_1848,N_1332,N_1451);
and U1849 (N_1849,N_1409,N_1232);
nand U1850 (N_1850,N_1150,N_1393);
nand U1851 (N_1851,N_1188,N_1313);
or U1852 (N_1852,N_1408,N_1241);
and U1853 (N_1853,N_1206,N_1155);
or U1854 (N_1854,N_1107,N_1333);
nor U1855 (N_1855,N_1188,N_1307);
nand U1856 (N_1856,N_1174,N_1381);
nor U1857 (N_1857,N_1014,N_1251);
or U1858 (N_1858,N_1035,N_1097);
nor U1859 (N_1859,N_1069,N_1103);
and U1860 (N_1860,N_1219,N_1445);
or U1861 (N_1861,N_1482,N_1411);
or U1862 (N_1862,N_1329,N_1425);
and U1863 (N_1863,N_1016,N_1395);
nand U1864 (N_1864,N_1188,N_1165);
xor U1865 (N_1865,N_1205,N_1415);
nand U1866 (N_1866,N_1466,N_1335);
xnor U1867 (N_1867,N_1176,N_1488);
nand U1868 (N_1868,N_1024,N_1317);
nor U1869 (N_1869,N_1438,N_1062);
or U1870 (N_1870,N_1157,N_1236);
or U1871 (N_1871,N_1177,N_1359);
or U1872 (N_1872,N_1071,N_1037);
nand U1873 (N_1873,N_1204,N_1352);
and U1874 (N_1874,N_1417,N_1051);
and U1875 (N_1875,N_1144,N_1464);
or U1876 (N_1876,N_1320,N_1274);
nor U1877 (N_1877,N_1153,N_1486);
nand U1878 (N_1878,N_1457,N_1060);
or U1879 (N_1879,N_1252,N_1321);
nor U1880 (N_1880,N_1064,N_1090);
nor U1881 (N_1881,N_1309,N_1033);
or U1882 (N_1882,N_1036,N_1017);
or U1883 (N_1883,N_1341,N_1109);
and U1884 (N_1884,N_1365,N_1493);
nand U1885 (N_1885,N_1050,N_1113);
nand U1886 (N_1886,N_1148,N_1252);
nor U1887 (N_1887,N_1033,N_1379);
and U1888 (N_1888,N_1022,N_1190);
nand U1889 (N_1889,N_1134,N_1090);
and U1890 (N_1890,N_1047,N_1076);
nor U1891 (N_1891,N_1459,N_1093);
or U1892 (N_1892,N_1134,N_1398);
or U1893 (N_1893,N_1232,N_1234);
or U1894 (N_1894,N_1303,N_1408);
xor U1895 (N_1895,N_1470,N_1161);
nand U1896 (N_1896,N_1316,N_1303);
nor U1897 (N_1897,N_1037,N_1062);
nand U1898 (N_1898,N_1345,N_1429);
nor U1899 (N_1899,N_1418,N_1223);
or U1900 (N_1900,N_1092,N_1161);
and U1901 (N_1901,N_1381,N_1346);
nor U1902 (N_1902,N_1459,N_1068);
nor U1903 (N_1903,N_1251,N_1231);
nand U1904 (N_1904,N_1006,N_1237);
or U1905 (N_1905,N_1161,N_1397);
or U1906 (N_1906,N_1433,N_1220);
or U1907 (N_1907,N_1364,N_1347);
and U1908 (N_1908,N_1215,N_1177);
nand U1909 (N_1909,N_1087,N_1145);
nor U1910 (N_1910,N_1195,N_1442);
and U1911 (N_1911,N_1311,N_1293);
and U1912 (N_1912,N_1267,N_1006);
nand U1913 (N_1913,N_1428,N_1402);
and U1914 (N_1914,N_1031,N_1177);
nand U1915 (N_1915,N_1209,N_1208);
nand U1916 (N_1916,N_1266,N_1382);
or U1917 (N_1917,N_1034,N_1368);
or U1918 (N_1918,N_1190,N_1068);
and U1919 (N_1919,N_1168,N_1046);
nor U1920 (N_1920,N_1257,N_1058);
and U1921 (N_1921,N_1033,N_1165);
and U1922 (N_1922,N_1066,N_1449);
and U1923 (N_1923,N_1053,N_1325);
nor U1924 (N_1924,N_1071,N_1032);
or U1925 (N_1925,N_1279,N_1266);
or U1926 (N_1926,N_1319,N_1441);
nor U1927 (N_1927,N_1129,N_1020);
and U1928 (N_1928,N_1264,N_1420);
or U1929 (N_1929,N_1192,N_1060);
and U1930 (N_1930,N_1171,N_1434);
and U1931 (N_1931,N_1451,N_1471);
nor U1932 (N_1932,N_1130,N_1344);
nor U1933 (N_1933,N_1333,N_1411);
and U1934 (N_1934,N_1010,N_1003);
xor U1935 (N_1935,N_1095,N_1417);
nor U1936 (N_1936,N_1004,N_1314);
and U1937 (N_1937,N_1321,N_1462);
nor U1938 (N_1938,N_1472,N_1098);
nand U1939 (N_1939,N_1090,N_1066);
nand U1940 (N_1940,N_1133,N_1149);
nand U1941 (N_1941,N_1126,N_1452);
nand U1942 (N_1942,N_1011,N_1033);
xnor U1943 (N_1943,N_1482,N_1380);
and U1944 (N_1944,N_1364,N_1323);
and U1945 (N_1945,N_1353,N_1146);
nor U1946 (N_1946,N_1498,N_1054);
nand U1947 (N_1947,N_1127,N_1085);
nor U1948 (N_1948,N_1233,N_1290);
nand U1949 (N_1949,N_1310,N_1078);
or U1950 (N_1950,N_1189,N_1325);
nor U1951 (N_1951,N_1482,N_1325);
or U1952 (N_1952,N_1275,N_1170);
nand U1953 (N_1953,N_1325,N_1024);
and U1954 (N_1954,N_1235,N_1160);
nor U1955 (N_1955,N_1322,N_1218);
nor U1956 (N_1956,N_1455,N_1439);
nand U1957 (N_1957,N_1232,N_1221);
xor U1958 (N_1958,N_1216,N_1189);
and U1959 (N_1959,N_1115,N_1321);
and U1960 (N_1960,N_1477,N_1168);
nand U1961 (N_1961,N_1386,N_1468);
nand U1962 (N_1962,N_1414,N_1170);
nand U1963 (N_1963,N_1099,N_1479);
and U1964 (N_1964,N_1390,N_1203);
nand U1965 (N_1965,N_1033,N_1030);
and U1966 (N_1966,N_1328,N_1199);
or U1967 (N_1967,N_1050,N_1070);
nand U1968 (N_1968,N_1286,N_1093);
and U1969 (N_1969,N_1168,N_1164);
nand U1970 (N_1970,N_1036,N_1361);
or U1971 (N_1971,N_1240,N_1497);
and U1972 (N_1972,N_1464,N_1447);
or U1973 (N_1973,N_1058,N_1401);
and U1974 (N_1974,N_1133,N_1472);
and U1975 (N_1975,N_1392,N_1181);
or U1976 (N_1976,N_1149,N_1360);
and U1977 (N_1977,N_1133,N_1002);
and U1978 (N_1978,N_1446,N_1341);
nand U1979 (N_1979,N_1195,N_1186);
nor U1980 (N_1980,N_1163,N_1077);
nand U1981 (N_1981,N_1442,N_1283);
and U1982 (N_1982,N_1423,N_1351);
nand U1983 (N_1983,N_1252,N_1443);
or U1984 (N_1984,N_1254,N_1394);
and U1985 (N_1985,N_1404,N_1446);
nand U1986 (N_1986,N_1219,N_1494);
and U1987 (N_1987,N_1013,N_1490);
nor U1988 (N_1988,N_1435,N_1261);
nand U1989 (N_1989,N_1305,N_1137);
nor U1990 (N_1990,N_1032,N_1174);
nand U1991 (N_1991,N_1202,N_1267);
xor U1992 (N_1992,N_1211,N_1347);
nor U1993 (N_1993,N_1385,N_1482);
and U1994 (N_1994,N_1112,N_1363);
nand U1995 (N_1995,N_1311,N_1384);
or U1996 (N_1996,N_1365,N_1394);
nand U1997 (N_1997,N_1015,N_1145);
nor U1998 (N_1998,N_1386,N_1484);
and U1999 (N_1999,N_1291,N_1085);
nor U2000 (N_2000,N_1554,N_1536);
xor U2001 (N_2001,N_1849,N_1697);
and U2002 (N_2002,N_1622,N_1659);
nand U2003 (N_2003,N_1821,N_1918);
nand U2004 (N_2004,N_1983,N_1970);
nand U2005 (N_2005,N_1759,N_1567);
nand U2006 (N_2006,N_1840,N_1606);
xor U2007 (N_2007,N_1894,N_1757);
or U2008 (N_2008,N_1820,N_1559);
nor U2009 (N_2009,N_1708,N_1786);
nand U2010 (N_2010,N_1674,N_1873);
and U2011 (N_2011,N_1898,N_1914);
and U2012 (N_2012,N_1778,N_1928);
nand U2013 (N_2013,N_1616,N_1777);
nor U2014 (N_2014,N_1959,N_1602);
nor U2015 (N_2015,N_1828,N_1792);
or U2016 (N_2016,N_1515,N_1767);
or U2017 (N_2017,N_1871,N_1860);
and U2018 (N_2018,N_1818,N_1895);
and U2019 (N_2019,N_1858,N_1637);
nand U2020 (N_2020,N_1965,N_1938);
or U2021 (N_2021,N_1884,N_1856);
or U2022 (N_2022,N_1885,N_1916);
and U2023 (N_2023,N_1874,N_1621);
nor U2024 (N_2024,N_1800,N_1580);
or U2025 (N_2025,N_1682,N_1592);
xor U2026 (N_2026,N_1508,N_1953);
or U2027 (N_2027,N_1794,N_1814);
nor U2028 (N_2028,N_1958,N_1688);
nand U2029 (N_2029,N_1500,N_1903);
nand U2030 (N_2030,N_1556,N_1825);
and U2031 (N_2031,N_1913,N_1925);
nor U2032 (N_2032,N_1547,N_1891);
nand U2033 (N_2033,N_1996,N_1607);
nor U2034 (N_2034,N_1990,N_1579);
and U2035 (N_2035,N_1775,N_1549);
nor U2036 (N_2036,N_1839,N_1670);
or U2037 (N_2037,N_1807,N_1521);
nor U2038 (N_2038,N_1577,N_1736);
and U2039 (N_2039,N_1655,N_1717);
or U2040 (N_2040,N_1641,N_1713);
or U2041 (N_2041,N_1528,N_1940);
nand U2042 (N_2042,N_1980,N_1529);
or U2043 (N_2043,N_1752,N_1747);
nor U2044 (N_2044,N_1975,N_1861);
xnor U2045 (N_2045,N_1564,N_1583);
nand U2046 (N_2046,N_1982,N_1572);
nand U2047 (N_2047,N_1544,N_1608);
and U2048 (N_2048,N_1543,N_1626);
or U2049 (N_2049,N_1684,N_1919);
and U2050 (N_2050,N_1598,N_1756);
and U2051 (N_2051,N_1739,N_1628);
or U2052 (N_2052,N_1838,N_1941);
or U2053 (N_2053,N_1636,N_1877);
nand U2054 (N_2054,N_1563,N_1710);
nor U2055 (N_2055,N_1788,N_1900);
nand U2056 (N_2056,N_1888,N_1907);
nand U2057 (N_2057,N_1934,N_1876);
and U2058 (N_2058,N_1805,N_1780);
nor U2059 (N_2059,N_1935,N_1504);
xor U2060 (N_2060,N_1687,N_1582);
and U2061 (N_2061,N_1712,N_1514);
nor U2062 (N_2062,N_1615,N_1526);
and U2063 (N_2063,N_1978,N_1661);
nand U2064 (N_2064,N_1944,N_1748);
and U2065 (N_2065,N_1664,N_1618);
or U2066 (N_2066,N_1964,N_1816);
nand U2067 (N_2067,N_1764,N_1966);
and U2068 (N_2068,N_1784,N_1981);
and U2069 (N_2069,N_1799,N_1848);
nand U2070 (N_2070,N_1960,N_1623);
or U2071 (N_2071,N_1501,N_1823);
nor U2072 (N_2072,N_1709,N_1802);
or U2073 (N_2073,N_1597,N_1984);
nor U2074 (N_2074,N_1705,N_1942);
or U2075 (N_2075,N_1589,N_1902);
nand U2076 (N_2076,N_1893,N_1973);
nor U2077 (N_2077,N_1590,N_1692);
and U2078 (N_2078,N_1988,N_1926);
and U2079 (N_2079,N_1812,N_1698);
and U2080 (N_2080,N_1864,N_1969);
or U2081 (N_2081,N_1985,N_1790);
or U2082 (N_2082,N_1968,N_1663);
or U2083 (N_2083,N_1963,N_1831);
nor U2084 (N_2084,N_1773,N_1796);
or U2085 (N_2085,N_1976,N_1594);
and U2086 (N_2086,N_1974,N_1545);
or U2087 (N_2087,N_1870,N_1803);
nand U2088 (N_2088,N_1678,N_1555);
nand U2089 (N_2089,N_1505,N_1511);
or U2090 (N_2090,N_1746,N_1774);
and U2091 (N_2091,N_1855,N_1931);
nor U2092 (N_2092,N_1844,N_1811);
nor U2093 (N_2093,N_1890,N_1630);
nor U2094 (N_2094,N_1993,N_1904);
nand U2095 (N_2095,N_1610,N_1720);
and U2096 (N_2096,N_1769,N_1977);
or U2097 (N_2097,N_1881,N_1806);
and U2098 (N_2098,N_1875,N_1677);
or U2099 (N_2099,N_1765,N_1771);
nand U2100 (N_2100,N_1612,N_1634);
and U2101 (N_2101,N_1826,N_1967);
xor U2102 (N_2102,N_1892,N_1866);
nand U2103 (N_2103,N_1952,N_1955);
nand U2104 (N_2104,N_1599,N_1561);
nand U2105 (N_2105,N_1865,N_1723);
nor U2106 (N_2106,N_1879,N_1728);
nand U2107 (N_2107,N_1666,N_1851);
and U2108 (N_2108,N_1961,N_1569);
nor U2109 (N_2109,N_1742,N_1939);
nor U2110 (N_2110,N_1937,N_1842);
or U2111 (N_2111,N_1933,N_1603);
or U2112 (N_2112,N_1915,N_1945);
and U2113 (N_2113,N_1815,N_1729);
nor U2114 (N_2114,N_1843,N_1776);
nor U2115 (N_2115,N_1857,N_1750);
or U2116 (N_2116,N_1715,N_1558);
nand U2117 (N_2117,N_1732,N_1546);
and U2118 (N_2118,N_1585,N_1568);
nand U2119 (N_2119,N_1633,N_1600);
nand U2120 (N_2120,N_1629,N_1791);
or U2121 (N_2121,N_1910,N_1617);
nand U2122 (N_2122,N_1760,N_1658);
nand U2123 (N_2123,N_1927,N_1524);
or U2124 (N_2124,N_1645,N_1689);
or U2125 (N_2125,N_1754,N_1932);
or U2126 (N_2126,N_1995,N_1954);
or U2127 (N_2127,N_1669,N_1749);
nand U2128 (N_2128,N_1518,N_1531);
or U2129 (N_2129,N_1758,N_1810);
or U2130 (N_2130,N_1699,N_1520);
nand U2131 (N_2131,N_1835,N_1638);
and U2132 (N_2132,N_1516,N_1650);
nand U2133 (N_2133,N_1575,N_1847);
and U2134 (N_2134,N_1644,N_1987);
and U2135 (N_2135,N_1829,N_1539);
nand U2136 (N_2136,N_1726,N_1643);
and U2137 (N_2137,N_1672,N_1667);
or U2138 (N_2138,N_1783,N_1523);
and U2139 (N_2139,N_1946,N_1782);
or U2140 (N_2140,N_1586,N_1971);
xnor U2141 (N_2141,N_1869,N_1862);
and U2142 (N_2142,N_1624,N_1513);
nor U2143 (N_2143,N_1766,N_1763);
or U2144 (N_2144,N_1772,N_1921);
and U2145 (N_2145,N_1951,N_1830);
nand U2146 (N_2146,N_1647,N_1882);
and U2147 (N_2147,N_1787,N_1552);
or U2148 (N_2148,N_1679,N_1741);
and U2149 (N_2149,N_1761,N_1581);
nor U2150 (N_2150,N_1734,N_1770);
nand U2151 (N_2151,N_1700,N_1639);
nor U2152 (N_2152,N_1542,N_1956);
nor U2153 (N_2153,N_1817,N_1999);
or U2154 (N_2154,N_1906,N_1917);
and U2155 (N_2155,N_1745,N_1834);
nand U2156 (N_2156,N_1571,N_1837);
or U2157 (N_2157,N_1943,N_1897);
nor U2158 (N_2158,N_1753,N_1541);
nand U2159 (N_2159,N_1537,N_1789);
nand U2160 (N_2160,N_1525,N_1886);
nand U2161 (N_2161,N_1948,N_1722);
nand U2162 (N_2162,N_1642,N_1804);
nand U2163 (N_2163,N_1872,N_1595);
xnor U2164 (N_2164,N_1868,N_1587);
nor U2165 (N_2165,N_1795,N_1922);
and U2166 (N_2166,N_1992,N_1880);
or U2167 (N_2167,N_1593,N_1727);
nand U2168 (N_2168,N_1744,N_1517);
or U2169 (N_2169,N_1681,N_1668);
or U2170 (N_2170,N_1704,N_1702);
and U2171 (N_2171,N_1706,N_1614);
or U2172 (N_2172,N_1649,N_1716);
or U2173 (N_2173,N_1801,N_1781);
and U2174 (N_2174,N_1994,N_1991);
nor U2175 (N_2175,N_1797,N_1652);
nor U2176 (N_2176,N_1680,N_1566);
and U2177 (N_2177,N_1863,N_1920);
nor U2178 (N_2178,N_1665,N_1620);
or U2179 (N_2179,N_1519,N_1768);
nand U2180 (N_2180,N_1905,N_1574);
nor U2181 (N_2181,N_1535,N_1853);
or U2182 (N_2182,N_1588,N_1711);
nor U2183 (N_2183,N_1813,N_1532);
nand U2184 (N_2184,N_1733,N_1793);
nand U2185 (N_2185,N_1625,N_1507);
and U2186 (N_2186,N_1671,N_1675);
and U2187 (N_2187,N_1998,N_1836);
nor U2188 (N_2188,N_1950,N_1512);
or U2189 (N_2189,N_1653,N_1755);
or U2190 (N_2190,N_1506,N_1632);
nand U2191 (N_2191,N_1845,N_1827);
or U2192 (N_2192,N_1701,N_1657);
nor U2193 (N_2193,N_1724,N_1735);
nor U2194 (N_2194,N_1929,N_1751);
or U2195 (N_2195,N_1613,N_1596);
nor U2196 (N_2196,N_1693,N_1949);
nor U2197 (N_2197,N_1550,N_1605);
nor U2198 (N_2198,N_1627,N_1901);
nand U2199 (N_2199,N_1832,N_1957);
or U2200 (N_2200,N_1997,N_1648);
nand U2201 (N_2201,N_1924,N_1762);
nor U2202 (N_2202,N_1565,N_1779);
and U2203 (N_2203,N_1591,N_1730);
and U2204 (N_2204,N_1846,N_1573);
or U2205 (N_2205,N_1850,N_1611);
and U2206 (N_2206,N_1721,N_1527);
or U2207 (N_2207,N_1899,N_1911);
and U2208 (N_2208,N_1930,N_1578);
xor U2209 (N_2209,N_1609,N_1534);
xnor U2210 (N_2210,N_1740,N_1551);
nor U2211 (N_2211,N_1651,N_1576);
nand U2212 (N_2212,N_1635,N_1824);
and U2213 (N_2213,N_1841,N_1533);
xnor U2214 (N_2214,N_1540,N_1503);
nand U2215 (N_2215,N_1833,N_1695);
xor U2216 (N_2216,N_1947,N_1662);
or U2217 (N_2217,N_1557,N_1601);
nor U2218 (N_2218,N_1936,N_1676);
or U2219 (N_2219,N_1619,N_1719);
nor U2220 (N_2220,N_1972,N_1731);
or U2221 (N_2221,N_1703,N_1867);
xnor U2222 (N_2222,N_1553,N_1854);
and U2223 (N_2223,N_1883,N_1819);
or U2224 (N_2224,N_1989,N_1646);
nor U2225 (N_2225,N_1584,N_1570);
or U2226 (N_2226,N_1604,N_1798);
nor U2227 (N_2227,N_1538,N_1562);
nand U2228 (N_2228,N_1889,N_1690);
or U2229 (N_2229,N_1691,N_1707);
nand U2230 (N_2230,N_1522,N_1631);
xnor U2231 (N_2231,N_1923,N_1696);
xor U2232 (N_2232,N_1822,N_1912);
nor U2233 (N_2233,N_1640,N_1530);
nand U2234 (N_2234,N_1852,N_1986);
nor U2235 (N_2235,N_1808,N_1785);
and U2236 (N_2236,N_1502,N_1683);
nand U2237 (N_2237,N_1673,N_1908);
nand U2238 (N_2238,N_1685,N_1896);
or U2239 (N_2239,N_1887,N_1694);
and U2240 (N_2240,N_1979,N_1743);
or U2241 (N_2241,N_1510,N_1859);
nor U2242 (N_2242,N_1686,N_1660);
nand U2243 (N_2243,N_1548,N_1909);
nor U2244 (N_2244,N_1718,N_1878);
and U2245 (N_2245,N_1714,N_1809);
xor U2246 (N_2246,N_1560,N_1509);
or U2247 (N_2247,N_1725,N_1654);
nand U2248 (N_2248,N_1656,N_1962);
or U2249 (N_2249,N_1738,N_1737);
nor U2250 (N_2250,N_1510,N_1621);
nor U2251 (N_2251,N_1935,N_1523);
nand U2252 (N_2252,N_1581,N_1856);
nand U2253 (N_2253,N_1544,N_1995);
or U2254 (N_2254,N_1777,N_1697);
or U2255 (N_2255,N_1799,N_1631);
nand U2256 (N_2256,N_1736,N_1603);
nand U2257 (N_2257,N_1542,N_1813);
xnor U2258 (N_2258,N_1643,N_1796);
xnor U2259 (N_2259,N_1807,N_1841);
nor U2260 (N_2260,N_1780,N_1865);
nor U2261 (N_2261,N_1767,N_1556);
nor U2262 (N_2262,N_1642,N_1751);
nand U2263 (N_2263,N_1805,N_1928);
nor U2264 (N_2264,N_1763,N_1586);
nor U2265 (N_2265,N_1697,N_1871);
nor U2266 (N_2266,N_1801,N_1684);
xor U2267 (N_2267,N_1617,N_1647);
or U2268 (N_2268,N_1803,N_1534);
nor U2269 (N_2269,N_1540,N_1700);
nand U2270 (N_2270,N_1670,N_1925);
nand U2271 (N_2271,N_1789,N_1894);
and U2272 (N_2272,N_1573,N_1641);
or U2273 (N_2273,N_1823,N_1930);
and U2274 (N_2274,N_1951,N_1725);
or U2275 (N_2275,N_1961,N_1544);
nor U2276 (N_2276,N_1673,N_1800);
and U2277 (N_2277,N_1681,N_1737);
nand U2278 (N_2278,N_1806,N_1679);
nand U2279 (N_2279,N_1799,N_1808);
and U2280 (N_2280,N_1749,N_1724);
nor U2281 (N_2281,N_1827,N_1652);
nand U2282 (N_2282,N_1592,N_1736);
xor U2283 (N_2283,N_1623,N_1729);
or U2284 (N_2284,N_1546,N_1729);
nor U2285 (N_2285,N_1721,N_1551);
or U2286 (N_2286,N_1798,N_1739);
or U2287 (N_2287,N_1570,N_1822);
xor U2288 (N_2288,N_1500,N_1522);
and U2289 (N_2289,N_1511,N_1886);
nand U2290 (N_2290,N_1675,N_1772);
and U2291 (N_2291,N_1887,N_1904);
nor U2292 (N_2292,N_1582,N_1789);
and U2293 (N_2293,N_1702,N_1968);
nor U2294 (N_2294,N_1525,N_1616);
and U2295 (N_2295,N_1641,N_1754);
nor U2296 (N_2296,N_1776,N_1971);
nand U2297 (N_2297,N_1838,N_1574);
xnor U2298 (N_2298,N_1845,N_1885);
nor U2299 (N_2299,N_1922,N_1545);
nor U2300 (N_2300,N_1820,N_1599);
nor U2301 (N_2301,N_1914,N_1729);
or U2302 (N_2302,N_1684,N_1941);
xnor U2303 (N_2303,N_1748,N_1803);
and U2304 (N_2304,N_1769,N_1803);
nand U2305 (N_2305,N_1592,N_1767);
nor U2306 (N_2306,N_1776,N_1648);
nand U2307 (N_2307,N_1507,N_1877);
nand U2308 (N_2308,N_1845,N_1551);
and U2309 (N_2309,N_1816,N_1952);
and U2310 (N_2310,N_1543,N_1518);
xnor U2311 (N_2311,N_1912,N_1735);
nor U2312 (N_2312,N_1885,N_1922);
and U2313 (N_2313,N_1913,N_1627);
nand U2314 (N_2314,N_1622,N_1897);
and U2315 (N_2315,N_1724,N_1527);
xnor U2316 (N_2316,N_1531,N_1709);
nor U2317 (N_2317,N_1762,N_1841);
nor U2318 (N_2318,N_1774,N_1685);
or U2319 (N_2319,N_1598,N_1993);
or U2320 (N_2320,N_1628,N_1560);
and U2321 (N_2321,N_1826,N_1806);
nand U2322 (N_2322,N_1593,N_1535);
nand U2323 (N_2323,N_1539,N_1555);
nor U2324 (N_2324,N_1712,N_1721);
xor U2325 (N_2325,N_1913,N_1769);
or U2326 (N_2326,N_1506,N_1979);
nor U2327 (N_2327,N_1506,N_1983);
nand U2328 (N_2328,N_1647,N_1795);
nand U2329 (N_2329,N_1718,N_1804);
nor U2330 (N_2330,N_1725,N_1849);
and U2331 (N_2331,N_1546,N_1731);
and U2332 (N_2332,N_1784,N_1527);
and U2333 (N_2333,N_1825,N_1813);
or U2334 (N_2334,N_1636,N_1901);
nand U2335 (N_2335,N_1539,N_1759);
or U2336 (N_2336,N_1508,N_1844);
nor U2337 (N_2337,N_1764,N_1601);
nand U2338 (N_2338,N_1992,N_1546);
or U2339 (N_2339,N_1630,N_1621);
xnor U2340 (N_2340,N_1600,N_1970);
and U2341 (N_2341,N_1897,N_1929);
xor U2342 (N_2342,N_1616,N_1747);
nand U2343 (N_2343,N_1979,N_1634);
nor U2344 (N_2344,N_1576,N_1503);
and U2345 (N_2345,N_1596,N_1969);
xor U2346 (N_2346,N_1535,N_1814);
and U2347 (N_2347,N_1609,N_1928);
or U2348 (N_2348,N_1546,N_1660);
and U2349 (N_2349,N_1902,N_1849);
and U2350 (N_2350,N_1653,N_1790);
and U2351 (N_2351,N_1669,N_1787);
or U2352 (N_2352,N_1744,N_1995);
nand U2353 (N_2353,N_1693,N_1745);
and U2354 (N_2354,N_1713,N_1658);
xor U2355 (N_2355,N_1904,N_1558);
and U2356 (N_2356,N_1863,N_1712);
nand U2357 (N_2357,N_1813,N_1500);
and U2358 (N_2358,N_1691,N_1638);
or U2359 (N_2359,N_1939,N_1722);
and U2360 (N_2360,N_1837,N_1626);
or U2361 (N_2361,N_1920,N_1739);
nand U2362 (N_2362,N_1541,N_1729);
or U2363 (N_2363,N_1947,N_1878);
nand U2364 (N_2364,N_1808,N_1575);
and U2365 (N_2365,N_1540,N_1736);
nand U2366 (N_2366,N_1663,N_1884);
and U2367 (N_2367,N_1702,N_1537);
nor U2368 (N_2368,N_1585,N_1678);
or U2369 (N_2369,N_1558,N_1759);
nor U2370 (N_2370,N_1706,N_1738);
and U2371 (N_2371,N_1563,N_1513);
or U2372 (N_2372,N_1794,N_1832);
or U2373 (N_2373,N_1521,N_1769);
and U2374 (N_2374,N_1781,N_1870);
or U2375 (N_2375,N_1664,N_1923);
nor U2376 (N_2376,N_1676,N_1680);
nand U2377 (N_2377,N_1720,N_1966);
nor U2378 (N_2378,N_1753,N_1773);
xor U2379 (N_2379,N_1905,N_1636);
nand U2380 (N_2380,N_1595,N_1870);
nand U2381 (N_2381,N_1786,N_1534);
xnor U2382 (N_2382,N_1791,N_1807);
nand U2383 (N_2383,N_1940,N_1599);
xor U2384 (N_2384,N_1934,N_1758);
and U2385 (N_2385,N_1945,N_1659);
or U2386 (N_2386,N_1527,N_1931);
or U2387 (N_2387,N_1732,N_1513);
or U2388 (N_2388,N_1547,N_1623);
or U2389 (N_2389,N_1635,N_1900);
xor U2390 (N_2390,N_1800,N_1820);
and U2391 (N_2391,N_1853,N_1988);
and U2392 (N_2392,N_1875,N_1652);
nor U2393 (N_2393,N_1956,N_1927);
xnor U2394 (N_2394,N_1853,N_1837);
and U2395 (N_2395,N_1839,N_1647);
and U2396 (N_2396,N_1871,N_1870);
xnor U2397 (N_2397,N_1674,N_1571);
nor U2398 (N_2398,N_1802,N_1874);
or U2399 (N_2399,N_1961,N_1935);
nand U2400 (N_2400,N_1817,N_1721);
nor U2401 (N_2401,N_1684,N_1630);
or U2402 (N_2402,N_1697,N_1863);
and U2403 (N_2403,N_1822,N_1886);
and U2404 (N_2404,N_1941,N_1544);
nand U2405 (N_2405,N_1906,N_1732);
nor U2406 (N_2406,N_1815,N_1919);
or U2407 (N_2407,N_1532,N_1730);
xor U2408 (N_2408,N_1694,N_1843);
nand U2409 (N_2409,N_1897,N_1700);
or U2410 (N_2410,N_1910,N_1689);
or U2411 (N_2411,N_1886,N_1798);
or U2412 (N_2412,N_1868,N_1814);
nor U2413 (N_2413,N_1517,N_1533);
nand U2414 (N_2414,N_1508,N_1952);
and U2415 (N_2415,N_1878,N_1615);
nand U2416 (N_2416,N_1802,N_1527);
xor U2417 (N_2417,N_1890,N_1942);
xor U2418 (N_2418,N_1789,N_1549);
nor U2419 (N_2419,N_1711,N_1838);
nor U2420 (N_2420,N_1635,N_1925);
nor U2421 (N_2421,N_1563,N_1524);
and U2422 (N_2422,N_1951,N_1509);
and U2423 (N_2423,N_1542,N_1567);
nand U2424 (N_2424,N_1993,N_1840);
or U2425 (N_2425,N_1949,N_1663);
nand U2426 (N_2426,N_1786,N_1624);
nor U2427 (N_2427,N_1773,N_1648);
nor U2428 (N_2428,N_1736,N_1621);
and U2429 (N_2429,N_1524,N_1747);
nor U2430 (N_2430,N_1615,N_1875);
and U2431 (N_2431,N_1569,N_1738);
and U2432 (N_2432,N_1748,N_1723);
xnor U2433 (N_2433,N_1644,N_1740);
nand U2434 (N_2434,N_1762,N_1821);
or U2435 (N_2435,N_1889,N_1740);
nor U2436 (N_2436,N_1654,N_1952);
or U2437 (N_2437,N_1917,N_1897);
nor U2438 (N_2438,N_1804,N_1570);
nand U2439 (N_2439,N_1647,N_1935);
nand U2440 (N_2440,N_1501,N_1667);
nand U2441 (N_2441,N_1592,N_1982);
or U2442 (N_2442,N_1665,N_1577);
and U2443 (N_2443,N_1719,N_1927);
and U2444 (N_2444,N_1686,N_1602);
or U2445 (N_2445,N_1591,N_1802);
and U2446 (N_2446,N_1807,N_1753);
and U2447 (N_2447,N_1775,N_1843);
or U2448 (N_2448,N_1991,N_1885);
nand U2449 (N_2449,N_1885,N_1626);
or U2450 (N_2450,N_1889,N_1733);
or U2451 (N_2451,N_1575,N_1617);
xnor U2452 (N_2452,N_1584,N_1732);
nand U2453 (N_2453,N_1829,N_1713);
and U2454 (N_2454,N_1545,N_1527);
nand U2455 (N_2455,N_1712,N_1885);
nor U2456 (N_2456,N_1712,N_1602);
nor U2457 (N_2457,N_1539,N_1899);
nor U2458 (N_2458,N_1638,N_1623);
or U2459 (N_2459,N_1587,N_1734);
and U2460 (N_2460,N_1786,N_1655);
or U2461 (N_2461,N_1549,N_1726);
xnor U2462 (N_2462,N_1636,N_1610);
or U2463 (N_2463,N_1965,N_1701);
nor U2464 (N_2464,N_1887,N_1597);
and U2465 (N_2465,N_1685,N_1730);
and U2466 (N_2466,N_1644,N_1695);
and U2467 (N_2467,N_1591,N_1611);
or U2468 (N_2468,N_1643,N_1879);
or U2469 (N_2469,N_1528,N_1514);
xnor U2470 (N_2470,N_1698,N_1644);
and U2471 (N_2471,N_1927,N_1680);
or U2472 (N_2472,N_1710,N_1653);
and U2473 (N_2473,N_1784,N_1877);
nor U2474 (N_2474,N_1674,N_1744);
nand U2475 (N_2475,N_1633,N_1754);
nand U2476 (N_2476,N_1937,N_1984);
nand U2477 (N_2477,N_1640,N_1658);
nor U2478 (N_2478,N_1654,N_1740);
nor U2479 (N_2479,N_1726,N_1622);
nand U2480 (N_2480,N_1527,N_1637);
and U2481 (N_2481,N_1785,N_1739);
and U2482 (N_2482,N_1524,N_1764);
nand U2483 (N_2483,N_1773,N_1794);
and U2484 (N_2484,N_1637,N_1937);
or U2485 (N_2485,N_1604,N_1948);
nand U2486 (N_2486,N_1926,N_1709);
nand U2487 (N_2487,N_1953,N_1749);
and U2488 (N_2488,N_1689,N_1952);
nand U2489 (N_2489,N_1822,N_1897);
nand U2490 (N_2490,N_1781,N_1831);
and U2491 (N_2491,N_1742,N_1573);
and U2492 (N_2492,N_1857,N_1801);
nor U2493 (N_2493,N_1513,N_1610);
nand U2494 (N_2494,N_1857,N_1842);
nor U2495 (N_2495,N_1985,N_1965);
nand U2496 (N_2496,N_1650,N_1904);
nor U2497 (N_2497,N_1739,N_1679);
nand U2498 (N_2498,N_1968,N_1532);
and U2499 (N_2499,N_1957,N_1995);
and U2500 (N_2500,N_2487,N_2267);
and U2501 (N_2501,N_2416,N_2360);
and U2502 (N_2502,N_2430,N_2139);
nor U2503 (N_2503,N_2488,N_2050);
xnor U2504 (N_2504,N_2034,N_2148);
nor U2505 (N_2505,N_2038,N_2471);
xnor U2506 (N_2506,N_2068,N_2373);
and U2507 (N_2507,N_2400,N_2223);
nand U2508 (N_2508,N_2270,N_2285);
nor U2509 (N_2509,N_2458,N_2411);
or U2510 (N_2510,N_2449,N_2394);
or U2511 (N_2511,N_2186,N_2396);
nor U2512 (N_2512,N_2438,N_2194);
and U2513 (N_2513,N_2330,N_2136);
nor U2514 (N_2514,N_2296,N_2078);
and U2515 (N_2515,N_2132,N_2174);
xnor U2516 (N_2516,N_2257,N_2066);
or U2517 (N_2517,N_2406,N_2221);
and U2518 (N_2518,N_2474,N_2156);
nor U2519 (N_2519,N_2260,N_2439);
nor U2520 (N_2520,N_2003,N_2345);
xnor U2521 (N_2521,N_2173,N_2448);
xnor U2522 (N_2522,N_2399,N_2486);
nand U2523 (N_2523,N_2307,N_2379);
nand U2524 (N_2524,N_2249,N_2142);
nor U2525 (N_2525,N_2404,N_2189);
nor U2526 (N_2526,N_2427,N_2370);
nand U2527 (N_2527,N_2405,N_2178);
nor U2528 (N_2528,N_2278,N_2299);
nor U2529 (N_2529,N_2141,N_2305);
or U2530 (N_2530,N_2137,N_2262);
nand U2531 (N_2531,N_2089,N_2140);
and U2532 (N_2532,N_2105,N_2030);
and U2533 (N_2533,N_2154,N_2101);
and U2534 (N_2534,N_2375,N_2339);
nand U2535 (N_2535,N_2205,N_2244);
nor U2536 (N_2536,N_2341,N_2079);
nand U2537 (N_2537,N_2494,N_2317);
or U2538 (N_2538,N_2426,N_2331);
or U2539 (N_2539,N_2199,N_2028);
and U2540 (N_2540,N_2462,N_2453);
or U2541 (N_2541,N_2049,N_2364);
and U2542 (N_2542,N_2151,N_2145);
nor U2543 (N_2543,N_2445,N_2304);
nand U2544 (N_2544,N_2150,N_2232);
and U2545 (N_2545,N_2401,N_2010);
or U2546 (N_2546,N_2366,N_2460);
xnor U2547 (N_2547,N_2433,N_2209);
nand U2548 (N_2548,N_2193,N_2253);
or U2549 (N_2549,N_2006,N_2246);
nor U2550 (N_2550,N_2286,N_2423);
or U2551 (N_2551,N_2091,N_2340);
nand U2552 (N_2552,N_2429,N_2387);
and U2553 (N_2553,N_2316,N_2302);
nor U2554 (N_2554,N_2033,N_2061);
nand U2555 (N_2555,N_2212,N_2022);
and U2556 (N_2556,N_2226,N_2032);
nand U2557 (N_2557,N_2467,N_2385);
xnor U2558 (N_2558,N_2171,N_2300);
xor U2559 (N_2559,N_2265,N_2256);
and U2560 (N_2560,N_2046,N_2388);
nand U2561 (N_2561,N_2273,N_2224);
nand U2562 (N_2562,N_2198,N_2029);
and U2563 (N_2563,N_2037,N_2197);
or U2564 (N_2564,N_2104,N_2422);
and U2565 (N_2565,N_2052,N_2452);
and U2566 (N_2566,N_2324,N_2362);
or U2567 (N_2567,N_2475,N_2359);
or U2568 (N_2568,N_2319,N_2441);
or U2569 (N_2569,N_2268,N_2227);
or U2570 (N_2570,N_2352,N_2073);
and U2571 (N_2571,N_2229,N_2255);
nand U2572 (N_2572,N_2167,N_2208);
or U2573 (N_2573,N_2081,N_2131);
or U2574 (N_2574,N_2347,N_2496);
nand U2575 (N_2575,N_2060,N_2200);
xnor U2576 (N_2576,N_2009,N_2125);
and U2577 (N_2577,N_2220,N_2014);
nor U2578 (N_2578,N_2292,N_2111);
nand U2579 (N_2579,N_2211,N_2418);
nor U2580 (N_2580,N_2251,N_2088);
nor U2581 (N_2581,N_2040,N_2202);
nor U2582 (N_2582,N_2110,N_2196);
or U2583 (N_2583,N_2086,N_2469);
or U2584 (N_2584,N_2397,N_2204);
nand U2585 (N_2585,N_2381,N_2044);
and U2586 (N_2586,N_2412,N_2436);
nor U2587 (N_2587,N_2019,N_2447);
nor U2588 (N_2588,N_2077,N_2280);
xor U2589 (N_2589,N_2376,N_2369);
xor U2590 (N_2590,N_2041,N_2365);
nand U2591 (N_2591,N_2311,N_2410);
nand U2592 (N_2592,N_2297,N_2228);
or U2593 (N_2593,N_2168,N_2463);
and U2594 (N_2594,N_2398,N_2002);
nor U2595 (N_2595,N_2084,N_2259);
xor U2596 (N_2596,N_2323,N_2218);
nand U2597 (N_2597,N_2337,N_2456);
nand U2598 (N_2598,N_2057,N_2306);
nand U2599 (N_2599,N_2461,N_2000);
xor U2600 (N_2600,N_2358,N_2415);
xor U2601 (N_2601,N_2020,N_2138);
nor U2602 (N_2602,N_2015,N_2035);
and U2603 (N_2603,N_2217,N_2016);
or U2604 (N_2604,N_2389,N_2266);
nand U2605 (N_2605,N_2318,N_2153);
nand U2606 (N_2606,N_2333,N_2238);
or U2607 (N_2607,N_2314,N_2087);
nor U2608 (N_2608,N_2025,N_2085);
or U2609 (N_2609,N_2069,N_2272);
and U2610 (N_2610,N_2126,N_2393);
nor U2611 (N_2611,N_2384,N_2011);
nor U2612 (N_2612,N_2294,N_2036);
nor U2613 (N_2613,N_2207,N_2083);
or U2614 (N_2614,N_2313,N_2236);
or U2615 (N_2615,N_2017,N_2166);
nand U2616 (N_2616,N_2464,N_2160);
or U2617 (N_2617,N_2013,N_2308);
nand U2618 (N_2618,N_2417,N_2161);
nand U2619 (N_2619,N_2372,N_2233);
or U2620 (N_2620,N_2071,N_2203);
and U2621 (N_2621,N_2130,N_2230);
nand U2622 (N_2622,N_2301,N_2484);
nor U2623 (N_2623,N_2325,N_2004);
xnor U2624 (N_2624,N_2216,N_2225);
nand U2625 (N_2625,N_2390,N_2261);
nand U2626 (N_2626,N_2332,N_2348);
nor U2627 (N_2627,N_2413,N_2492);
or U2628 (N_2628,N_2144,N_2134);
or U2629 (N_2629,N_2334,N_2328);
nor U2630 (N_2630,N_2112,N_2100);
or U2631 (N_2631,N_2149,N_2420);
and U2632 (N_2632,N_2027,N_2195);
or U2633 (N_2633,N_2491,N_2407);
xnor U2634 (N_2634,N_2187,N_2129);
nand U2635 (N_2635,N_2382,N_2241);
and U2636 (N_2636,N_2170,N_2054);
nor U2637 (N_2637,N_2001,N_2283);
nor U2638 (N_2638,N_2498,N_2021);
nor U2639 (N_2639,N_2113,N_2277);
nor U2640 (N_2640,N_2152,N_2219);
nand U2641 (N_2641,N_2455,N_2062);
nand U2642 (N_2642,N_2143,N_2175);
nand U2643 (N_2643,N_2063,N_2479);
nand U2644 (N_2644,N_2440,N_2076);
or U2645 (N_2645,N_2124,N_2179);
nor U2646 (N_2646,N_2431,N_2248);
or U2647 (N_2647,N_2135,N_2499);
or U2648 (N_2648,N_2048,N_2192);
nor U2649 (N_2649,N_2095,N_2329);
or U2650 (N_2650,N_2258,N_2284);
and U2651 (N_2651,N_2099,N_2293);
nor U2652 (N_2652,N_2481,N_2031);
nor U2653 (N_2653,N_2184,N_2287);
or U2654 (N_2654,N_2242,N_2008);
or U2655 (N_2655,N_2155,N_2109);
or U2656 (N_2656,N_2428,N_2018);
nand U2657 (N_2657,N_2082,N_2443);
and U2658 (N_2658,N_2042,N_2237);
nor U2659 (N_2659,N_2094,N_2056);
and U2660 (N_2660,N_2096,N_2005);
and U2661 (N_2661,N_2213,N_2451);
and U2662 (N_2662,N_2424,N_2162);
nand U2663 (N_2663,N_2327,N_2465);
or U2664 (N_2664,N_2103,N_2190);
or U2665 (N_2665,N_2122,N_2177);
or U2666 (N_2666,N_2210,N_2480);
nor U2667 (N_2667,N_2403,N_2444);
or U2668 (N_2668,N_2419,N_2466);
nor U2669 (N_2669,N_2146,N_2367);
or U2670 (N_2670,N_2392,N_2408);
nand U2671 (N_2671,N_2092,N_2493);
nor U2672 (N_2672,N_2435,N_2371);
nand U2673 (N_2673,N_2402,N_2395);
or U2674 (N_2674,N_2201,N_2495);
nand U2675 (N_2675,N_2039,N_2275);
nand U2676 (N_2676,N_2107,N_2102);
nand U2677 (N_2677,N_2374,N_2473);
or U2678 (N_2678,N_2108,N_2391);
or U2679 (N_2679,N_2239,N_2222);
nor U2680 (N_2680,N_2043,N_2181);
or U2681 (N_2681,N_2377,N_2240);
or U2682 (N_2682,N_2414,N_2432);
xnor U2683 (N_2683,N_2361,N_2214);
or U2684 (N_2684,N_2354,N_2070);
xor U2685 (N_2685,N_2117,N_2353);
nand U2686 (N_2686,N_2123,N_2380);
nand U2687 (N_2687,N_2065,N_2234);
nor U2688 (N_2688,N_2356,N_2497);
or U2689 (N_2689,N_2472,N_2064);
nor U2690 (N_2690,N_2342,N_2243);
nor U2691 (N_2691,N_2271,N_2483);
nand U2692 (N_2692,N_2279,N_2349);
or U2693 (N_2693,N_2059,N_2386);
nand U2694 (N_2694,N_2183,N_2119);
and U2695 (N_2695,N_2485,N_2383);
nor U2696 (N_2696,N_2343,N_2072);
and U2697 (N_2697,N_2090,N_2158);
nand U2698 (N_2698,N_2098,N_2315);
or U2699 (N_2699,N_2409,N_2350);
nor U2700 (N_2700,N_2074,N_2450);
nand U2701 (N_2701,N_2164,N_2312);
xnor U2702 (N_2702,N_2442,N_2169);
nor U2703 (N_2703,N_2106,N_2476);
nand U2704 (N_2704,N_2254,N_2295);
xor U2705 (N_2705,N_2276,N_2310);
or U2706 (N_2706,N_2326,N_2097);
or U2707 (N_2707,N_2288,N_2180);
or U2708 (N_2708,N_2176,N_2128);
or U2709 (N_2709,N_2289,N_2378);
nor U2710 (N_2710,N_2490,N_2172);
nand U2711 (N_2711,N_2459,N_2264);
or U2712 (N_2712,N_2421,N_2437);
nor U2713 (N_2713,N_2336,N_2454);
and U2714 (N_2714,N_2206,N_2351);
nor U2715 (N_2715,N_2185,N_2163);
or U2716 (N_2716,N_2457,N_2231);
or U2717 (N_2717,N_2290,N_2026);
nand U2718 (N_2718,N_2274,N_2120);
or U2719 (N_2719,N_2075,N_2355);
or U2720 (N_2720,N_2053,N_2055);
nor U2721 (N_2721,N_2127,N_2115);
and U2722 (N_2722,N_2045,N_2188);
nand U2723 (N_2723,N_2470,N_2252);
and U2724 (N_2724,N_2215,N_2446);
nor U2725 (N_2725,N_2058,N_2247);
nand U2726 (N_2726,N_2309,N_2478);
nor U2727 (N_2727,N_2335,N_2133);
nand U2728 (N_2728,N_2489,N_2344);
nor U2729 (N_2729,N_2118,N_2282);
nand U2730 (N_2730,N_2250,N_2191);
nand U2731 (N_2731,N_2322,N_2114);
nand U2732 (N_2732,N_2093,N_2165);
or U2733 (N_2733,N_2007,N_2303);
nand U2734 (N_2734,N_2346,N_2338);
nand U2735 (N_2735,N_2263,N_2482);
and U2736 (N_2736,N_2051,N_2269);
nor U2737 (N_2737,N_2320,N_2024);
xor U2738 (N_2738,N_2477,N_2368);
nand U2739 (N_2739,N_2235,N_2425);
nand U2740 (N_2740,N_2157,N_2357);
xnor U2741 (N_2741,N_2281,N_2468);
and U2742 (N_2742,N_2147,N_2245);
nor U2743 (N_2743,N_2159,N_2023);
or U2744 (N_2744,N_2080,N_2012);
or U2745 (N_2745,N_2298,N_2121);
xnor U2746 (N_2746,N_2434,N_2321);
nand U2747 (N_2747,N_2067,N_2291);
and U2748 (N_2748,N_2116,N_2182);
nand U2749 (N_2749,N_2047,N_2363);
nor U2750 (N_2750,N_2294,N_2404);
nand U2751 (N_2751,N_2476,N_2492);
nand U2752 (N_2752,N_2457,N_2304);
nand U2753 (N_2753,N_2051,N_2330);
nand U2754 (N_2754,N_2445,N_2421);
nand U2755 (N_2755,N_2154,N_2458);
nor U2756 (N_2756,N_2412,N_2344);
nand U2757 (N_2757,N_2445,N_2280);
xnor U2758 (N_2758,N_2277,N_2049);
and U2759 (N_2759,N_2436,N_2176);
or U2760 (N_2760,N_2322,N_2312);
xnor U2761 (N_2761,N_2180,N_2462);
nand U2762 (N_2762,N_2245,N_2205);
or U2763 (N_2763,N_2450,N_2219);
nor U2764 (N_2764,N_2112,N_2446);
or U2765 (N_2765,N_2287,N_2356);
nor U2766 (N_2766,N_2300,N_2057);
or U2767 (N_2767,N_2306,N_2125);
xor U2768 (N_2768,N_2392,N_2128);
or U2769 (N_2769,N_2481,N_2174);
or U2770 (N_2770,N_2239,N_2137);
or U2771 (N_2771,N_2322,N_2158);
nor U2772 (N_2772,N_2300,N_2424);
nor U2773 (N_2773,N_2003,N_2039);
nand U2774 (N_2774,N_2068,N_2263);
nor U2775 (N_2775,N_2019,N_2416);
or U2776 (N_2776,N_2096,N_2394);
nand U2777 (N_2777,N_2160,N_2426);
xor U2778 (N_2778,N_2406,N_2113);
xor U2779 (N_2779,N_2316,N_2359);
nor U2780 (N_2780,N_2237,N_2226);
and U2781 (N_2781,N_2327,N_2295);
nor U2782 (N_2782,N_2116,N_2430);
or U2783 (N_2783,N_2120,N_2171);
and U2784 (N_2784,N_2008,N_2498);
nand U2785 (N_2785,N_2000,N_2305);
or U2786 (N_2786,N_2455,N_2160);
or U2787 (N_2787,N_2383,N_2083);
and U2788 (N_2788,N_2177,N_2286);
nand U2789 (N_2789,N_2468,N_2246);
xnor U2790 (N_2790,N_2407,N_2115);
or U2791 (N_2791,N_2310,N_2115);
nor U2792 (N_2792,N_2090,N_2023);
nand U2793 (N_2793,N_2036,N_2185);
nand U2794 (N_2794,N_2015,N_2308);
and U2795 (N_2795,N_2032,N_2262);
or U2796 (N_2796,N_2286,N_2295);
or U2797 (N_2797,N_2231,N_2332);
nor U2798 (N_2798,N_2461,N_2393);
and U2799 (N_2799,N_2288,N_2257);
xnor U2800 (N_2800,N_2101,N_2434);
or U2801 (N_2801,N_2001,N_2432);
nor U2802 (N_2802,N_2280,N_2099);
nor U2803 (N_2803,N_2064,N_2440);
or U2804 (N_2804,N_2149,N_2476);
and U2805 (N_2805,N_2279,N_2094);
and U2806 (N_2806,N_2270,N_2002);
nor U2807 (N_2807,N_2254,N_2343);
and U2808 (N_2808,N_2146,N_2424);
or U2809 (N_2809,N_2440,N_2495);
nand U2810 (N_2810,N_2072,N_2176);
or U2811 (N_2811,N_2019,N_2267);
and U2812 (N_2812,N_2391,N_2066);
and U2813 (N_2813,N_2404,N_2119);
or U2814 (N_2814,N_2162,N_2499);
nand U2815 (N_2815,N_2309,N_2268);
or U2816 (N_2816,N_2398,N_2174);
or U2817 (N_2817,N_2030,N_2342);
or U2818 (N_2818,N_2123,N_2477);
nand U2819 (N_2819,N_2402,N_2213);
and U2820 (N_2820,N_2463,N_2277);
or U2821 (N_2821,N_2496,N_2236);
xnor U2822 (N_2822,N_2317,N_2459);
nand U2823 (N_2823,N_2187,N_2285);
and U2824 (N_2824,N_2269,N_2183);
nand U2825 (N_2825,N_2109,N_2231);
or U2826 (N_2826,N_2014,N_2194);
or U2827 (N_2827,N_2264,N_2158);
nand U2828 (N_2828,N_2162,N_2418);
and U2829 (N_2829,N_2426,N_2306);
or U2830 (N_2830,N_2211,N_2054);
nand U2831 (N_2831,N_2174,N_2218);
nand U2832 (N_2832,N_2491,N_2250);
or U2833 (N_2833,N_2010,N_2079);
or U2834 (N_2834,N_2239,N_2037);
nor U2835 (N_2835,N_2158,N_2292);
or U2836 (N_2836,N_2269,N_2250);
and U2837 (N_2837,N_2232,N_2126);
xor U2838 (N_2838,N_2200,N_2122);
or U2839 (N_2839,N_2002,N_2066);
and U2840 (N_2840,N_2461,N_2339);
and U2841 (N_2841,N_2064,N_2211);
and U2842 (N_2842,N_2388,N_2240);
and U2843 (N_2843,N_2093,N_2340);
nor U2844 (N_2844,N_2134,N_2156);
or U2845 (N_2845,N_2184,N_2039);
or U2846 (N_2846,N_2189,N_2149);
nand U2847 (N_2847,N_2000,N_2392);
nor U2848 (N_2848,N_2322,N_2398);
nor U2849 (N_2849,N_2451,N_2162);
nand U2850 (N_2850,N_2385,N_2378);
and U2851 (N_2851,N_2312,N_2031);
nor U2852 (N_2852,N_2166,N_2154);
or U2853 (N_2853,N_2300,N_2058);
xor U2854 (N_2854,N_2124,N_2115);
nand U2855 (N_2855,N_2105,N_2180);
or U2856 (N_2856,N_2220,N_2110);
nand U2857 (N_2857,N_2421,N_2054);
xor U2858 (N_2858,N_2079,N_2264);
and U2859 (N_2859,N_2266,N_2169);
or U2860 (N_2860,N_2168,N_2330);
nor U2861 (N_2861,N_2163,N_2385);
or U2862 (N_2862,N_2060,N_2251);
and U2863 (N_2863,N_2325,N_2032);
or U2864 (N_2864,N_2210,N_2329);
or U2865 (N_2865,N_2003,N_2463);
and U2866 (N_2866,N_2136,N_2400);
nand U2867 (N_2867,N_2271,N_2415);
and U2868 (N_2868,N_2444,N_2484);
and U2869 (N_2869,N_2396,N_2015);
nor U2870 (N_2870,N_2094,N_2271);
or U2871 (N_2871,N_2311,N_2412);
nor U2872 (N_2872,N_2149,N_2265);
nor U2873 (N_2873,N_2332,N_2171);
or U2874 (N_2874,N_2255,N_2481);
nand U2875 (N_2875,N_2272,N_2314);
nand U2876 (N_2876,N_2493,N_2347);
nand U2877 (N_2877,N_2459,N_2434);
nand U2878 (N_2878,N_2496,N_2101);
or U2879 (N_2879,N_2365,N_2484);
nand U2880 (N_2880,N_2190,N_2220);
nand U2881 (N_2881,N_2478,N_2357);
or U2882 (N_2882,N_2200,N_2058);
nor U2883 (N_2883,N_2009,N_2105);
or U2884 (N_2884,N_2465,N_2382);
nand U2885 (N_2885,N_2203,N_2322);
nor U2886 (N_2886,N_2394,N_2003);
and U2887 (N_2887,N_2117,N_2149);
nor U2888 (N_2888,N_2425,N_2250);
nand U2889 (N_2889,N_2484,N_2336);
nor U2890 (N_2890,N_2171,N_2282);
nor U2891 (N_2891,N_2425,N_2147);
nand U2892 (N_2892,N_2392,N_2493);
and U2893 (N_2893,N_2399,N_2122);
nand U2894 (N_2894,N_2378,N_2035);
or U2895 (N_2895,N_2424,N_2438);
or U2896 (N_2896,N_2077,N_2127);
nor U2897 (N_2897,N_2112,N_2236);
nand U2898 (N_2898,N_2000,N_2226);
and U2899 (N_2899,N_2474,N_2236);
and U2900 (N_2900,N_2123,N_2009);
nand U2901 (N_2901,N_2155,N_2395);
nor U2902 (N_2902,N_2350,N_2005);
or U2903 (N_2903,N_2382,N_2391);
nand U2904 (N_2904,N_2249,N_2462);
or U2905 (N_2905,N_2251,N_2156);
and U2906 (N_2906,N_2283,N_2480);
nand U2907 (N_2907,N_2306,N_2025);
and U2908 (N_2908,N_2384,N_2425);
or U2909 (N_2909,N_2081,N_2458);
and U2910 (N_2910,N_2253,N_2405);
xor U2911 (N_2911,N_2266,N_2074);
xnor U2912 (N_2912,N_2076,N_2124);
xnor U2913 (N_2913,N_2109,N_2306);
and U2914 (N_2914,N_2244,N_2070);
or U2915 (N_2915,N_2044,N_2159);
xnor U2916 (N_2916,N_2497,N_2372);
nand U2917 (N_2917,N_2216,N_2002);
nor U2918 (N_2918,N_2371,N_2450);
nand U2919 (N_2919,N_2077,N_2439);
nand U2920 (N_2920,N_2418,N_2273);
or U2921 (N_2921,N_2326,N_2220);
nand U2922 (N_2922,N_2307,N_2328);
xnor U2923 (N_2923,N_2005,N_2264);
and U2924 (N_2924,N_2083,N_2248);
or U2925 (N_2925,N_2016,N_2436);
and U2926 (N_2926,N_2090,N_2054);
nand U2927 (N_2927,N_2100,N_2246);
nand U2928 (N_2928,N_2401,N_2096);
xnor U2929 (N_2929,N_2417,N_2338);
or U2930 (N_2930,N_2460,N_2327);
nand U2931 (N_2931,N_2284,N_2397);
nor U2932 (N_2932,N_2461,N_2204);
nand U2933 (N_2933,N_2051,N_2066);
nand U2934 (N_2934,N_2468,N_2043);
and U2935 (N_2935,N_2322,N_2281);
nor U2936 (N_2936,N_2312,N_2027);
nand U2937 (N_2937,N_2423,N_2427);
xor U2938 (N_2938,N_2086,N_2249);
nor U2939 (N_2939,N_2109,N_2455);
nor U2940 (N_2940,N_2292,N_2424);
nor U2941 (N_2941,N_2498,N_2424);
and U2942 (N_2942,N_2022,N_2175);
nand U2943 (N_2943,N_2291,N_2302);
nand U2944 (N_2944,N_2351,N_2109);
or U2945 (N_2945,N_2002,N_2277);
or U2946 (N_2946,N_2118,N_2009);
nor U2947 (N_2947,N_2111,N_2201);
or U2948 (N_2948,N_2081,N_2097);
and U2949 (N_2949,N_2475,N_2393);
and U2950 (N_2950,N_2258,N_2319);
nand U2951 (N_2951,N_2321,N_2260);
or U2952 (N_2952,N_2066,N_2026);
or U2953 (N_2953,N_2351,N_2213);
nand U2954 (N_2954,N_2060,N_2459);
or U2955 (N_2955,N_2482,N_2309);
nor U2956 (N_2956,N_2400,N_2211);
nor U2957 (N_2957,N_2177,N_2328);
nand U2958 (N_2958,N_2160,N_2407);
nor U2959 (N_2959,N_2213,N_2179);
nor U2960 (N_2960,N_2083,N_2202);
nand U2961 (N_2961,N_2089,N_2189);
or U2962 (N_2962,N_2399,N_2379);
or U2963 (N_2963,N_2351,N_2080);
nor U2964 (N_2964,N_2141,N_2354);
and U2965 (N_2965,N_2347,N_2263);
or U2966 (N_2966,N_2233,N_2456);
and U2967 (N_2967,N_2068,N_2257);
or U2968 (N_2968,N_2407,N_2075);
nor U2969 (N_2969,N_2357,N_2426);
and U2970 (N_2970,N_2290,N_2031);
and U2971 (N_2971,N_2418,N_2332);
nand U2972 (N_2972,N_2196,N_2431);
and U2973 (N_2973,N_2076,N_2386);
and U2974 (N_2974,N_2081,N_2407);
and U2975 (N_2975,N_2174,N_2065);
or U2976 (N_2976,N_2031,N_2327);
xor U2977 (N_2977,N_2000,N_2056);
or U2978 (N_2978,N_2032,N_2346);
nand U2979 (N_2979,N_2471,N_2496);
and U2980 (N_2980,N_2121,N_2490);
and U2981 (N_2981,N_2297,N_2255);
and U2982 (N_2982,N_2174,N_2489);
and U2983 (N_2983,N_2485,N_2126);
or U2984 (N_2984,N_2374,N_2447);
xnor U2985 (N_2985,N_2451,N_2459);
xor U2986 (N_2986,N_2270,N_2075);
xor U2987 (N_2987,N_2127,N_2308);
nor U2988 (N_2988,N_2286,N_2317);
nand U2989 (N_2989,N_2100,N_2319);
nand U2990 (N_2990,N_2014,N_2400);
or U2991 (N_2991,N_2306,N_2213);
nor U2992 (N_2992,N_2329,N_2498);
or U2993 (N_2993,N_2243,N_2141);
nor U2994 (N_2994,N_2079,N_2001);
and U2995 (N_2995,N_2117,N_2187);
nand U2996 (N_2996,N_2456,N_2384);
nor U2997 (N_2997,N_2340,N_2259);
xor U2998 (N_2998,N_2073,N_2007);
and U2999 (N_2999,N_2076,N_2409);
or U3000 (N_3000,N_2673,N_2884);
nor U3001 (N_3001,N_2568,N_2923);
nand U3002 (N_3002,N_2723,N_2877);
xnor U3003 (N_3003,N_2599,N_2852);
nor U3004 (N_3004,N_2827,N_2839);
and U3005 (N_3005,N_2646,N_2627);
nand U3006 (N_3006,N_2843,N_2714);
and U3007 (N_3007,N_2631,N_2793);
nor U3008 (N_3008,N_2851,N_2887);
or U3009 (N_3009,N_2737,N_2639);
and U3010 (N_3010,N_2593,N_2792);
nor U3011 (N_3011,N_2751,N_2986);
nor U3012 (N_3012,N_2623,N_2881);
or U3013 (N_3013,N_2721,N_2542);
nand U3014 (N_3014,N_2904,N_2768);
and U3015 (N_3015,N_2720,N_2590);
nand U3016 (N_3016,N_2836,N_2759);
or U3017 (N_3017,N_2841,N_2628);
and U3018 (N_3018,N_2809,N_2529);
nand U3019 (N_3019,N_2562,N_2971);
nand U3020 (N_3020,N_2619,N_2592);
xnor U3021 (N_3021,N_2826,N_2758);
nand U3022 (N_3022,N_2535,N_2557);
or U3023 (N_3023,N_2519,N_2561);
and U3024 (N_3024,N_2832,N_2840);
nor U3025 (N_3025,N_2794,N_2596);
nor U3026 (N_3026,N_2928,N_2833);
and U3027 (N_3027,N_2776,N_2766);
nor U3028 (N_3028,N_2615,N_2888);
and U3029 (N_3029,N_2658,N_2732);
nand U3030 (N_3030,N_2802,N_2985);
and U3031 (N_3031,N_2508,N_2518);
or U3032 (N_3032,N_2604,N_2964);
nor U3033 (N_3033,N_2527,N_2886);
and U3034 (N_3034,N_2609,N_2689);
nand U3035 (N_3035,N_2944,N_2653);
and U3036 (N_3036,N_2989,N_2883);
or U3037 (N_3037,N_2539,N_2976);
nand U3038 (N_3038,N_2830,N_2581);
nor U3039 (N_3039,N_2805,N_2716);
nand U3040 (N_3040,N_2774,N_2893);
and U3041 (N_3041,N_2761,N_2548);
or U3042 (N_3042,N_2540,N_2547);
or U3043 (N_3043,N_2650,N_2878);
nor U3044 (N_3044,N_2586,N_2645);
or U3045 (N_3045,N_2949,N_2808);
xnor U3046 (N_3046,N_2507,N_2820);
nand U3047 (N_3047,N_2762,N_2734);
nor U3048 (N_3048,N_2783,N_2867);
nor U3049 (N_3049,N_2828,N_2853);
nor U3050 (N_3050,N_2857,N_2670);
and U3051 (N_3051,N_2974,N_2598);
xor U3052 (N_3052,N_2665,N_2757);
or U3053 (N_3053,N_2513,N_2861);
nand U3054 (N_3054,N_2688,N_2991);
or U3055 (N_3055,N_2937,N_2743);
nor U3056 (N_3056,N_2501,N_2709);
and U3057 (N_3057,N_2552,N_2848);
xnor U3058 (N_3058,N_2966,N_2775);
nand U3059 (N_3059,N_2522,N_2636);
or U3060 (N_3060,N_2907,N_2580);
or U3061 (N_3061,N_2876,N_2678);
nor U3062 (N_3062,N_2778,N_2591);
nor U3063 (N_3063,N_2902,N_2973);
and U3064 (N_3064,N_2536,N_2555);
nand U3065 (N_3065,N_2697,N_2772);
nand U3066 (N_3066,N_2831,N_2917);
nand U3067 (N_3067,N_2717,N_2703);
nor U3068 (N_3068,N_2891,N_2858);
nor U3069 (N_3069,N_2895,N_2629);
and U3070 (N_3070,N_2728,N_2649);
nand U3071 (N_3071,N_2582,N_2938);
and U3072 (N_3072,N_2834,N_2677);
nand U3073 (N_3073,N_2968,N_2722);
nand U3074 (N_3074,N_2784,N_2998);
nand U3075 (N_3075,N_2651,N_2683);
or U3076 (N_3076,N_2630,N_2686);
nor U3077 (N_3077,N_2691,N_2660);
or U3078 (N_3078,N_2789,N_2909);
xnor U3079 (N_3079,N_2936,N_2959);
or U3080 (N_3080,N_2578,N_2659);
nand U3081 (N_3081,N_2892,N_2738);
nor U3082 (N_3082,N_2781,N_2569);
nor U3083 (N_3083,N_2556,N_2756);
or U3084 (N_3084,N_2845,N_2875);
or U3085 (N_3085,N_2829,N_2754);
or U3086 (N_3086,N_2896,N_2600);
or U3087 (N_3087,N_2503,N_2963);
nor U3088 (N_3088,N_2584,N_2786);
xnor U3089 (N_3089,N_2915,N_2779);
nor U3090 (N_3090,N_2559,N_2900);
or U3091 (N_3091,N_2725,N_2795);
and U3092 (N_3092,N_2687,N_2702);
nor U3093 (N_3093,N_2641,N_2988);
nor U3094 (N_3094,N_2864,N_2745);
or U3095 (N_3095,N_2564,N_2602);
or U3096 (N_3096,N_2999,N_2940);
nand U3097 (N_3097,N_2773,N_2572);
and U3098 (N_3098,N_2606,N_2618);
nand U3099 (N_3099,N_2685,N_2695);
xnor U3100 (N_3100,N_2777,N_2983);
nor U3101 (N_3101,N_2594,N_2967);
or U3102 (N_3102,N_2588,N_2718);
and U3103 (N_3103,N_2755,N_2610);
xnor U3104 (N_3104,N_2538,N_2731);
nor U3105 (N_3105,N_2908,N_2837);
nor U3106 (N_3106,N_2696,N_2987);
and U3107 (N_3107,N_2595,N_2662);
nand U3108 (N_3108,N_2932,N_2943);
xor U3109 (N_3109,N_2934,N_2939);
and U3110 (N_3110,N_2873,N_2632);
nand U3111 (N_3111,N_2626,N_2872);
or U3112 (N_3112,N_2769,N_2933);
nor U3113 (N_3113,N_2981,N_2544);
or U3114 (N_3114,N_2742,N_2929);
or U3115 (N_3115,N_2563,N_2972);
nand U3116 (N_3116,N_2996,N_2969);
or U3117 (N_3117,N_2978,N_2553);
or U3118 (N_3118,N_2710,N_2741);
xnor U3119 (N_3119,N_2617,N_2819);
or U3120 (N_3120,N_2707,N_2679);
and U3121 (N_3121,N_2713,N_2704);
or U3122 (N_3122,N_2511,N_2791);
xor U3123 (N_3123,N_2847,N_2856);
nor U3124 (N_3124,N_2672,N_2577);
and U3125 (N_3125,N_2790,N_2894);
and U3126 (N_3126,N_2960,N_2882);
and U3127 (N_3127,N_2705,N_2825);
or U3128 (N_3128,N_2782,N_2621);
nand U3129 (N_3129,N_2748,N_2620);
nand U3130 (N_3130,N_2854,N_2997);
or U3131 (N_3131,N_2541,N_2865);
xor U3132 (N_3132,N_2648,N_2637);
nand U3133 (N_3133,N_2597,N_2505);
or U3134 (N_3134,N_2700,N_2545);
and U3135 (N_3135,N_2885,N_2694);
and U3136 (N_3136,N_2680,N_2913);
and U3137 (N_3137,N_2862,N_2583);
nor U3138 (N_3138,N_2706,N_2798);
or U3139 (N_3139,N_2500,N_2765);
nor U3140 (N_3140,N_2666,N_2749);
or U3141 (N_3141,N_2947,N_2824);
or U3142 (N_3142,N_2954,N_2815);
and U3143 (N_3143,N_2567,N_2855);
nor U3144 (N_3144,N_2879,N_2638);
nand U3145 (N_3145,N_2952,N_2990);
or U3146 (N_3146,N_2961,N_2711);
nor U3147 (N_3147,N_2520,N_2953);
and U3148 (N_3148,N_2912,N_2570);
nor U3149 (N_3149,N_2925,N_2640);
nor U3150 (N_3150,N_2514,N_2753);
or U3151 (N_3151,N_2526,N_2549);
nand U3152 (N_3152,N_2510,N_2589);
and U3153 (N_3153,N_2530,N_2760);
nand U3154 (N_3154,N_2931,N_2803);
nand U3155 (N_3155,N_2554,N_2616);
and U3156 (N_3156,N_2930,N_2977);
or U3157 (N_3157,N_2980,N_2740);
nor U3158 (N_3158,N_2780,N_2681);
nor U3159 (N_3159,N_2668,N_2729);
and U3160 (N_3160,N_2945,N_2537);
nand U3161 (N_3161,N_2838,N_2633);
or U3162 (N_3162,N_2655,N_2560);
and U3163 (N_3163,N_2574,N_2771);
or U3164 (N_3164,N_2935,N_2512);
nand U3165 (N_3165,N_2763,N_2899);
nor U3166 (N_3166,N_2652,N_2962);
nor U3167 (N_3167,N_2533,N_2579);
nand U3168 (N_3168,N_2796,N_2657);
nor U3169 (N_3169,N_2920,N_2799);
nand U3170 (N_3170,N_2642,N_2995);
and U3171 (N_3171,N_2515,N_2752);
and U3172 (N_3172,N_2903,N_2587);
or U3173 (N_3173,N_2676,N_2941);
and U3174 (N_3174,N_2647,N_2788);
and U3175 (N_3175,N_2558,N_2750);
or U3176 (N_3176,N_2951,N_2914);
or U3177 (N_3177,N_2661,N_2524);
or U3178 (N_3178,N_2571,N_2992);
nor U3179 (N_3179,N_2576,N_2921);
or U3180 (N_3180,N_2504,N_2984);
nand U3181 (N_3181,N_2622,N_2625);
nor U3182 (N_3182,N_2746,N_2897);
or U3183 (N_3183,N_2898,N_2835);
nor U3184 (N_3184,N_2575,N_2546);
nor U3185 (N_3185,N_2849,N_2927);
or U3186 (N_3186,N_2733,N_2603);
nor U3187 (N_3187,N_2674,N_2712);
xnor U3188 (N_3188,N_2684,N_2979);
nor U3189 (N_3189,N_2955,N_2889);
or U3190 (N_3190,N_2624,N_2611);
and U3191 (N_3191,N_2810,N_2656);
or U3192 (N_3192,N_2525,N_2534);
and U3193 (N_3193,N_2502,N_2654);
and U3194 (N_3194,N_2911,N_2550);
or U3195 (N_3195,N_2787,N_2664);
or U3196 (N_3196,N_2715,N_2817);
nor U3197 (N_3197,N_2764,N_2735);
and U3198 (N_3198,N_2675,N_2880);
and U3199 (N_3199,N_2724,N_2601);
nand U3200 (N_3200,N_2926,N_2747);
nand U3201 (N_3201,N_2607,N_2958);
xnor U3202 (N_3202,N_2859,N_2821);
and U3203 (N_3203,N_2922,N_2605);
xor U3204 (N_3204,N_2906,N_2918);
nand U3205 (N_3205,N_2634,N_2823);
nor U3206 (N_3206,N_2736,N_2608);
nor U3207 (N_3207,N_2744,N_2946);
nand U3208 (N_3208,N_2956,N_2890);
nor U3209 (N_3209,N_2813,N_2950);
and U3210 (N_3210,N_2871,N_2874);
nor U3211 (N_3211,N_2585,N_2994);
nand U3212 (N_3212,N_2682,N_2663);
and U3213 (N_3213,N_2516,N_2785);
and U3214 (N_3214,N_2869,N_2818);
and U3215 (N_3215,N_2669,N_2730);
and U3216 (N_3216,N_2806,N_2726);
nand U3217 (N_3217,N_2532,N_2612);
nand U3218 (N_3218,N_2844,N_2509);
nand U3219 (N_3219,N_2506,N_2901);
or U3220 (N_3220,N_2643,N_2671);
or U3221 (N_3221,N_2708,N_2957);
and U3222 (N_3222,N_2531,N_2905);
or U3223 (N_3223,N_2812,N_2767);
nor U3224 (N_3224,N_2868,N_2846);
or U3225 (N_3225,N_2910,N_2667);
or U3226 (N_3226,N_2565,N_2517);
xor U3227 (N_3227,N_2699,N_2644);
and U3228 (N_3228,N_2528,N_2635);
nand U3229 (N_3229,N_2942,N_2692);
xor U3230 (N_3230,N_2770,N_2523);
or U3231 (N_3231,N_2919,N_2811);
or U3232 (N_3232,N_2814,N_2727);
and U3233 (N_3233,N_2863,N_2521);
xnor U3234 (N_3234,N_2804,N_2816);
and U3235 (N_3235,N_2719,N_2698);
xor U3236 (N_3236,N_2739,N_2860);
nor U3237 (N_3237,N_2690,N_2551);
and U3238 (N_3238,N_2800,N_2797);
or U3239 (N_3239,N_2870,N_2982);
and U3240 (N_3240,N_2573,N_2993);
and U3241 (N_3241,N_2693,N_2822);
or U3242 (N_3242,N_2613,N_2801);
nor U3243 (N_3243,N_2807,N_2948);
or U3244 (N_3244,N_2850,N_2543);
nor U3245 (N_3245,N_2965,N_2916);
nand U3246 (N_3246,N_2866,N_2975);
xor U3247 (N_3247,N_2566,N_2970);
and U3248 (N_3248,N_2842,N_2924);
nand U3249 (N_3249,N_2614,N_2701);
or U3250 (N_3250,N_2616,N_2712);
and U3251 (N_3251,N_2928,N_2832);
xnor U3252 (N_3252,N_2970,N_2792);
nor U3253 (N_3253,N_2995,N_2579);
or U3254 (N_3254,N_2795,N_2679);
and U3255 (N_3255,N_2523,N_2659);
nor U3256 (N_3256,N_2614,N_2772);
nand U3257 (N_3257,N_2534,N_2896);
nand U3258 (N_3258,N_2862,N_2513);
and U3259 (N_3259,N_2885,N_2634);
and U3260 (N_3260,N_2793,N_2996);
and U3261 (N_3261,N_2756,N_2731);
and U3262 (N_3262,N_2506,N_2680);
and U3263 (N_3263,N_2559,N_2996);
nand U3264 (N_3264,N_2758,N_2959);
and U3265 (N_3265,N_2920,N_2697);
nor U3266 (N_3266,N_2842,N_2665);
xnor U3267 (N_3267,N_2911,N_2530);
and U3268 (N_3268,N_2875,N_2871);
xnor U3269 (N_3269,N_2556,N_2506);
and U3270 (N_3270,N_2535,N_2623);
nor U3271 (N_3271,N_2778,N_2575);
nor U3272 (N_3272,N_2908,N_2670);
and U3273 (N_3273,N_2762,N_2813);
or U3274 (N_3274,N_2832,N_2966);
and U3275 (N_3275,N_2612,N_2570);
nor U3276 (N_3276,N_2584,N_2575);
nand U3277 (N_3277,N_2759,N_2823);
or U3278 (N_3278,N_2831,N_2879);
and U3279 (N_3279,N_2579,N_2921);
and U3280 (N_3280,N_2556,N_2619);
nor U3281 (N_3281,N_2624,N_2971);
and U3282 (N_3282,N_2716,N_2963);
nor U3283 (N_3283,N_2588,N_2990);
or U3284 (N_3284,N_2549,N_2624);
nor U3285 (N_3285,N_2836,N_2597);
xor U3286 (N_3286,N_2853,N_2749);
xor U3287 (N_3287,N_2562,N_2660);
nand U3288 (N_3288,N_2666,N_2844);
nand U3289 (N_3289,N_2709,N_2865);
and U3290 (N_3290,N_2831,N_2779);
or U3291 (N_3291,N_2810,N_2552);
or U3292 (N_3292,N_2664,N_2500);
or U3293 (N_3293,N_2945,N_2562);
or U3294 (N_3294,N_2882,N_2916);
nor U3295 (N_3295,N_2886,N_2767);
xnor U3296 (N_3296,N_2779,N_2962);
and U3297 (N_3297,N_2674,N_2937);
or U3298 (N_3298,N_2532,N_2662);
and U3299 (N_3299,N_2547,N_2952);
nand U3300 (N_3300,N_2957,N_2941);
and U3301 (N_3301,N_2626,N_2822);
or U3302 (N_3302,N_2954,N_2799);
or U3303 (N_3303,N_2998,N_2780);
and U3304 (N_3304,N_2951,N_2857);
nor U3305 (N_3305,N_2715,N_2874);
and U3306 (N_3306,N_2902,N_2986);
or U3307 (N_3307,N_2852,N_2628);
or U3308 (N_3308,N_2700,N_2659);
or U3309 (N_3309,N_2763,N_2971);
or U3310 (N_3310,N_2844,N_2757);
nand U3311 (N_3311,N_2565,N_2842);
nor U3312 (N_3312,N_2601,N_2800);
nand U3313 (N_3313,N_2686,N_2813);
nand U3314 (N_3314,N_2553,N_2997);
or U3315 (N_3315,N_2724,N_2964);
or U3316 (N_3316,N_2862,N_2894);
and U3317 (N_3317,N_2691,N_2672);
nor U3318 (N_3318,N_2542,N_2924);
xnor U3319 (N_3319,N_2902,N_2680);
and U3320 (N_3320,N_2864,N_2711);
xnor U3321 (N_3321,N_2943,N_2887);
or U3322 (N_3322,N_2716,N_2966);
and U3323 (N_3323,N_2857,N_2559);
or U3324 (N_3324,N_2598,N_2779);
xnor U3325 (N_3325,N_2708,N_2784);
or U3326 (N_3326,N_2849,N_2794);
nor U3327 (N_3327,N_2830,N_2669);
nor U3328 (N_3328,N_2539,N_2780);
nand U3329 (N_3329,N_2714,N_2688);
and U3330 (N_3330,N_2672,N_2915);
nor U3331 (N_3331,N_2916,N_2881);
or U3332 (N_3332,N_2898,N_2604);
or U3333 (N_3333,N_2957,N_2880);
nand U3334 (N_3334,N_2999,N_2806);
and U3335 (N_3335,N_2909,N_2557);
nand U3336 (N_3336,N_2878,N_2584);
and U3337 (N_3337,N_2840,N_2773);
xor U3338 (N_3338,N_2617,N_2980);
or U3339 (N_3339,N_2670,N_2931);
nor U3340 (N_3340,N_2929,N_2729);
and U3341 (N_3341,N_2543,N_2984);
nand U3342 (N_3342,N_2692,N_2603);
and U3343 (N_3343,N_2609,N_2592);
and U3344 (N_3344,N_2998,N_2760);
nor U3345 (N_3345,N_2605,N_2844);
nor U3346 (N_3346,N_2562,N_2731);
or U3347 (N_3347,N_2743,N_2985);
nand U3348 (N_3348,N_2624,N_2601);
nand U3349 (N_3349,N_2785,N_2649);
or U3350 (N_3350,N_2782,N_2582);
nand U3351 (N_3351,N_2980,N_2863);
nor U3352 (N_3352,N_2880,N_2711);
and U3353 (N_3353,N_2733,N_2753);
nor U3354 (N_3354,N_2511,N_2644);
or U3355 (N_3355,N_2820,N_2557);
or U3356 (N_3356,N_2849,N_2798);
xnor U3357 (N_3357,N_2724,N_2665);
and U3358 (N_3358,N_2624,N_2597);
nor U3359 (N_3359,N_2509,N_2763);
nor U3360 (N_3360,N_2722,N_2980);
and U3361 (N_3361,N_2993,N_2997);
xnor U3362 (N_3362,N_2902,N_2514);
nor U3363 (N_3363,N_2583,N_2861);
nand U3364 (N_3364,N_2579,N_2554);
nor U3365 (N_3365,N_2581,N_2689);
nand U3366 (N_3366,N_2953,N_2870);
nor U3367 (N_3367,N_2901,N_2830);
or U3368 (N_3368,N_2969,N_2984);
and U3369 (N_3369,N_2760,N_2666);
nand U3370 (N_3370,N_2924,N_2729);
and U3371 (N_3371,N_2933,N_2650);
nand U3372 (N_3372,N_2528,N_2813);
and U3373 (N_3373,N_2690,N_2974);
nand U3374 (N_3374,N_2584,N_2892);
or U3375 (N_3375,N_2937,N_2681);
or U3376 (N_3376,N_2524,N_2539);
xor U3377 (N_3377,N_2890,N_2609);
xor U3378 (N_3378,N_2552,N_2633);
and U3379 (N_3379,N_2826,N_2590);
nand U3380 (N_3380,N_2592,N_2837);
or U3381 (N_3381,N_2716,N_2745);
nand U3382 (N_3382,N_2571,N_2608);
or U3383 (N_3383,N_2885,N_2510);
and U3384 (N_3384,N_2887,N_2643);
and U3385 (N_3385,N_2870,N_2521);
nand U3386 (N_3386,N_2575,N_2932);
and U3387 (N_3387,N_2972,N_2796);
and U3388 (N_3388,N_2869,N_2692);
or U3389 (N_3389,N_2972,N_2737);
xor U3390 (N_3390,N_2714,N_2674);
or U3391 (N_3391,N_2692,N_2827);
xor U3392 (N_3392,N_2583,N_2957);
or U3393 (N_3393,N_2538,N_2754);
or U3394 (N_3394,N_2977,N_2809);
and U3395 (N_3395,N_2873,N_2974);
xor U3396 (N_3396,N_2711,N_2823);
or U3397 (N_3397,N_2741,N_2541);
xor U3398 (N_3398,N_2940,N_2542);
nor U3399 (N_3399,N_2998,N_2882);
nor U3400 (N_3400,N_2934,N_2574);
and U3401 (N_3401,N_2697,N_2959);
or U3402 (N_3402,N_2735,N_2641);
and U3403 (N_3403,N_2812,N_2561);
nor U3404 (N_3404,N_2789,N_2829);
or U3405 (N_3405,N_2906,N_2820);
nand U3406 (N_3406,N_2535,N_2548);
or U3407 (N_3407,N_2868,N_2831);
and U3408 (N_3408,N_2742,N_2861);
xor U3409 (N_3409,N_2804,N_2701);
nor U3410 (N_3410,N_2881,N_2622);
xnor U3411 (N_3411,N_2709,N_2716);
nor U3412 (N_3412,N_2957,N_2714);
or U3413 (N_3413,N_2936,N_2729);
nand U3414 (N_3414,N_2573,N_2985);
nand U3415 (N_3415,N_2974,N_2594);
and U3416 (N_3416,N_2642,N_2885);
and U3417 (N_3417,N_2667,N_2536);
nand U3418 (N_3418,N_2760,N_2845);
and U3419 (N_3419,N_2731,N_2863);
nor U3420 (N_3420,N_2947,N_2694);
or U3421 (N_3421,N_2512,N_2971);
nand U3422 (N_3422,N_2919,N_2760);
xor U3423 (N_3423,N_2578,N_2880);
xnor U3424 (N_3424,N_2683,N_2761);
nor U3425 (N_3425,N_2554,N_2503);
and U3426 (N_3426,N_2527,N_2524);
or U3427 (N_3427,N_2825,N_2845);
nor U3428 (N_3428,N_2713,N_2905);
nand U3429 (N_3429,N_2828,N_2725);
nand U3430 (N_3430,N_2623,N_2536);
or U3431 (N_3431,N_2937,N_2860);
nand U3432 (N_3432,N_2558,N_2963);
nor U3433 (N_3433,N_2961,N_2819);
and U3434 (N_3434,N_2961,N_2911);
nor U3435 (N_3435,N_2674,N_2556);
or U3436 (N_3436,N_2873,N_2890);
nand U3437 (N_3437,N_2681,N_2711);
or U3438 (N_3438,N_2723,N_2608);
nor U3439 (N_3439,N_2855,N_2558);
or U3440 (N_3440,N_2749,N_2628);
nor U3441 (N_3441,N_2992,N_2948);
nand U3442 (N_3442,N_2947,N_2720);
nor U3443 (N_3443,N_2842,N_2836);
and U3444 (N_3444,N_2930,N_2554);
and U3445 (N_3445,N_2773,N_2644);
nand U3446 (N_3446,N_2724,N_2993);
and U3447 (N_3447,N_2967,N_2819);
nor U3448 (N_3448,N_2574,N_2926);
nor U3449 (N_3449,N_2871,N_2598);
nor U3450 (N_3450,N_2503,N_2656);
nand U3451 (N_3451,N_2775,N_2769);
or U3452 (N_3452,N_2762,N_2602);
nand U3453 (N_3453,N_2704,N_2920);
and U3454 (N_3454,N_2575,N_2807);
or U3455 (N_3455,N_2546,N_2909);
or U3456 (N_3456,N_2824,N_2805);
and U3457 (N_3457,N_2522,N_2934);
xnor U3458 (N_3458,N_2503,N_2722);
and U3459 (N_3459,N_2589,N_2970);
or U3460 (N_3460,N_2799,N_2988);
nand U3461 (N_3461,N_2748,N_2749);
nor U3462 (N_3462,N_2856,N_2813);
nor U3463 (N_3463,N_2708,N_2959);
or U3464 (N_3464,N_2954,N_2674);
and U3465 (N_3465,N_2674,N_2928);
xor U3466 (N_3466,N_2577,N_2653);
or U3467 (N_3467,N_2932,N_2667);
nor U3468 (N_3468,N_2727,N_2798);
nor U3469 (N_3469,N_2616,N_2532);
or U3470 (N_3470,N_2523,N_2686);
nand U3471 (N_3471,N_2534,N_2883);
and U3472 (N_3472,N_2519,N_2875);
nand U3473 (N_3473,N_2636,N_2798);
or U3474 (N_3474,N_2991,N_2596);
or U3475 (N_3475,N_2746,N_2703);
and U3476 (N_3476,N_2545,N_2739);
nor U3477 (N_3477,N_2921,N_2843);
xor U3478 (N_3478,N_2753,N_2810);
and U3479 (N_3479,N_2510,N_2887);
xnor U3480 (N_3480,N_2959,N_2644);
xor U3481 (N_3481,N_2869,N_2512);
nand U3482 (N_3482,N_2667,N_2637);
nand U3483 (N_3483,N_2538,N_2869);
and U3484 (N_3484,N_2939,N_2844);
and U3485 (N_3485,N_2712,N_2879);
nand U3486 (N_3486,N_2805,N_2792);
nand U3487 (N_3487,N_2919,N_2579);
nor U3488 (N_3488,N_2586,N_2944);
and U3489 (N_3489,N_2546,N_2813);
and U3490 (N_3490,N_2743,N_2877);
nor U3491 (N_3491,N_2677,N_2867);
nand U3492 (N_3492,N_2973,N_2541);
nand U3493 (N_3493,N_2507,N_2780);
nor U3494 (N_3494,N_2533,N_2510);
or U3495 (N_3495,N_2686,N_2765);
or U3496 (N_3496,N_2939,N_2668);
and U3497 (N_3497,N_2743,N_2856);
or U3498 (N_3498,N_2717,N_2689);
nand U3499 (N_3499,N_2724,N_2712);
and U3500 (N_3500,N_3146,N_3335);
nor U3501 (N_3501,N_3121,N_3408);
nand U3502 (N_3502,N_3482,N_3226);
and U3503 (N_3503,N_3297,N_3163);
or U3504 (N_3504,N_3131,N_3143);
nor U3505 (N_3505,N_3476,N_3398);
xor U3506 (N_3506,N_3463,N_3273);
and U3507 (N_3507,N_3489,N_3011);
nor U3508 (N_3508,N_3350,N_3475);
or U3509 (N_3509,N_3327,N_3422);
xnor U3510 (N_3510,N_3303,N_3008);
nor U3511 (N_3511,N_3015,N_3212);
nand U3512 (N_3512,N_3188,N_3043);
xnor U3513 (N_3513,N_3107,N_3116);
xor U3514 (N_3514,N_3112,N_3404);
nand U3515 (N_3515,N_3492,N_3364);
and U3516 (N_3516,N_3256,N_3374);
and U3517 (N_3517,N_3018,N_3400);
and U3518 (N_3518,N_3448,N_3021);
nor U3519 (N_3519,N_3344,N_3378);
nand U3520 (N_3520,N_3328,N_3318);
or U3521 (N_3521,N_3170,N_3167);
and U3522 (N_3522,N_3373,N_3034);
nor U3523 (N_3523,N_3098,N_3391);
and U3524 (N_3524,N_3093,N_3109);
nor U3525 (N_3525,N_3030,N_3035);
and U3526 (N_3526,N_3345,N_3294);
and U3527 (N_3527,N_3007,N_3236);
nor U3528 (N_3528,N_3359,N_3083);
nor U3529 (N_3529,N_3300,N_3355);
nor U3530 (N_3530,N_3057,N_3401);
or U3531 (N_3531,N_3331,N_3249);
or U3532 (N_3532,N_3101,N_3321);
or U3533 (N_3533,N_3380,N_3044);
nand U3534 (N_3534,N_3117,N_3495);
xor U3535 (N_3535,N_3037,N_3186);
nor U3536 (N_3536,N_3177,N_3435);
or U3537 (N_3537,N_3175,N_3198);
nand U3538 (N_3538,N_3136,N_3356);
or U3539 (N_3539,N_3078,N_3111);
or U3540 (N_3540,N_3323,N_3258);
and U3541 (N_3541,N_3394,N_3058);
or U3542 (N_3542,N_3081,N_3001);
or U3543 (N_3543,N_3106,N_3076);
and U3544 (N_3544,N_3269,N_3029);
and U3545 (N_3545,N_3077,N_3144);
or U3546 (N_3546,N_3329,N_3499);
nor U3547 (N_3547,N_3241,N_3099);
and U3548 (N_3548,N_3465,N_3082);
xor U3549 (N_3549,N_3484,N_3016);
and U3550 (N_3550,N_3187,N_3341);
xor U3551 (N_3551,N_3485,N_3085);
or U3552 (N_3552,N_3494,N_3147);
or U3553 (N_3553,N_3181,N_3261);
and U3554 (N_3554,N_3122,N_3279);
nor U3555 (N_3555,N_3061,N_3075);
and U3556 (N_3556,N_3429,N_3458);
nand U3557 (N_3557,N_3063,N_3202);
or U3558 (N_3558,N_3245,N_3421);
or U3559 (N_3559,N_3173,N_3383);
and U3560 (N_3560,N_3259,N_3480);
or U3561 (N_3561,N_3488,N_3237);
nand U3562 (N_3562,N_3191,N_3453);
nor U3563 (N_3563,N_3119,N_3326);
nor U3564 (N_3564,N_3340,N_3159);
nand U3565 (N_3565,N_3151,N_3419);
nor U3566 (N_3566,N_3068,N_3434);
and U3567 (N_3567,N_3090,N_3314);
or U3568 (N_3568,N_3417,N_3062);
and U3569 (N_3569,N_3005,N_3403);
nand U3570 (N_3570,N_3246,N_3054);
and U3571 (N_3571,N_3330,N_3320);
or U3572 (N_3572,N_3006,N_3218);
or U3573 (N_3573,N_3456,N_3095);
nand U3574 (N_3574,N_3120,N_3051);
xnor U3575 (N_3575,N_3277,N_3036);
or U3576 (N_3576,N_3288,N_3406);
nor U3577 (N_3577,N_3221,N_3071);
nand U3578 (N_3578,N_3020,N_3092);
or U3579 (N_3579,N_3307,N_3490);
nand U3580 (N_3580,N_3225,N_3268);
nand U3581 (N_3581,N_3309,N_3405);
nand U3582 (N_3582,N_3185,N_3128);
or U3583 (N_3583,N_3299,N_3487);
nor U3584 (N_3584,N_3275,N_3274);
or U3585 (N_3585,N_3442,N_3156);
or U3586 (N_3586,N_3497,N_3293);
or U3587 (N_3587,N_3334,N_3467);
and U3588 (N_3588,N_3336,N_3368);
nor U3589 (N_3589,N_3301,N_3390);
or U3590 (N_3590,N_3420,N_3289);
nand U3591 (N_3591,N_3457,N_3140);
or U3592 (N_3592,N_3281,N_3280);
nor U3593 (N_3593,N_3347,N_3209);
nand U3594 (N_3594,N_3250,N_3089);
and U3595 (N_3595,N_3074,N_3471);
and U3596 (N_3596,N_3462,N_3257);
and U3597 (N_3597,N_3348,N_3284);
xor U3598 (N_3598,N_3166,N_3211);
nor U3599 (N_3599,N_3362,N_3047);
nor U3600 (N_3600,N_3079,N_3325);
and U3601 (N_3601,N_3113,N_3477);
nor U3602 (N_3602,N_3133,N_3402);
nand U3603 (N_3603,N_3148,N_3324);
or U3604 (N_3604,N_3255,N_3000);
or U3605 (N_3605,N_3445,N_3152);
nand U3606 (N_3606,N_3266,N_3153);
nand U3607 (N_3607,N_3239,N_3118);
nor U3608 (N_3608,N_3426,N_3038);
nor U3609 (N_3609,N_3385,N_3206);
and U3610 (N_3610,N_3014,N_3103);
nor U3611 (N_3611,N_3424,N_3413);
and U3612 (N_3612,N_3127,N_3418);
and U3613 (N_3613,N_3407,N_3428);
and U3614 (N_3614,N_3179,N_3194);
nand U3615 (N_3615,N_3392,N_3260);
or U3616 (N_3616,N_3027,N_3414);
or U3617 (N_3617,N_3028,N_3222);
or U3618 (N_3618,N_3282,N_3278);
or U3619 (N_3619,N_3010,N_3454);
nand U3620 (N_3620,N_3161,N_3322);
nand U3621 (N_3621,N_3009,N_3064);
nand U3622 (N_3622,N_3339,N_3104);
or U3623 (N_3623,N_3395,N_3039);
and U3624 (N_3624,N_3270,N_3097);
and U3625 (N_3625,N_3411,N_3253);
and U3626 (N_3626,N_3486,N_3283);
or U3627 (N_3627,N_3470,N_3204);
or U3628 (N_3628,N_3369,N_3017);
nor U3629 (N_3629,N_3313,N_3180);
and U3630 (N_3630,N_3498,N_3139);
nor U3631 (N_3631,N_3142,N_3479);
and U3632 (N_3632,N_3022,N_3168);
or U3633 (N_3633,N_3472,N_3088);
nand U3634 (N_3634,N_3172,N_3041);
nor U3635 (N_3635,N_3137,N_3271);
and U3636 (N_3636,N_3304,N_3254);
nand U3637 (N_3637,N_3365,N_3376);
nor U3638 (N_3638,N_3114,N_3134);
or U3639 (N_3639,N_3354,N_3003);
and U3640 (N_3640,N_3023,N_3178);
nand U3641 (N_3641,N_3232,N_3375);
and U3642 (N_3642,N_3048,N_3311);
nand U3643 (N_3643,N_3425,N_3229);
or U3644 (N_3644,N_3205,N_3182);
nor U3645 (N_3645,N_3295,N_3440);
nor U3646 (N_3646,N_3124,N_3013);
nand U3647 (N_3647,N_3491,N_3149);
or U3648 (N_3648,N_3308,N_3252);
or U3649 (N_3649,N_3358,N_3032);
or U3650 (N_3650,N_3130,N_3216);
and U3651 (N_3651,N_3203,N_3310);
nand U3652 (N_3652,N_3438,N_3220);
nand U3653 (N_3653,N_3416,N_3040);
nand U3654 (N_3654,N_3315,N_3070);
and U3655 (N_3655,N_3357,N_3223);
nand U3656 (N_3656,N_3195,N_3102);
and U3657 (N_3657,N_3481,N_3306);
or U3658 (N_3658,N_3285,N_3371);
nand U3659 (N_3659,N_3265,N_3312);
nor U3660 (N_3660,N_3343,N_3444);
nand U3661 (N_3661,N_3069,N_3110);
nand U3662 (N_3662,N_3351,N_3353);
nor U3663 (N_3663,N_3410,N_3100);
or U3664 (N_3664,N_3230,N_3461);
xnor U3665 (N_3665,N_3189,N_3138);
or U3666 (N_3666,N_3412,N_3105);
and U3667 (N_3667,N_3091,N_3056);
nand U3668 (N_3668,N_3415,N_3427);
and U3669 (N_3669,N_3352,N_3165);
nor U3670 (N_3670,N_3393,N_3046);
and U3671 (N_3671,N_3349,N_3086);
or U3672 (N_3672,N_3446,N_3478);
and U3673 (N_3673,N_3384,N_3377);
nand U3674 (N_3674,N_3233,N_3200);
nand U3675 (N_3675,N_3342,N_3267);
nor U3676 (N_3676,N_3240,N_3024);
or U3677 (N_3677,N_3060,N_3319);
nand U3678 (N_3678,N_3238,N_3396);
and U3679 (N_3679,N_3108,N_3433);
and U3680 (N_3680,N_3154,N_3192);
nand U3681 (N_3681,N_3333,N_3447);
or U3682 (N_3682,N_3251,N_3316);
or U3683 (N_3683,N_3449,N_3235);
nand U3684 (N_3684,N_3367,N_3432);
nor U3685 (N_3685,N_3399,N_3468);
and U3686 (N_3686,N_3437,N_3087);
xnor U3687 (N_3687,N_3452,N_3224);
xnor U3688 (N_3688,N_3066,N_3228);
and U3689 (N_3689,N_3055,N_3065);
and U3690 (N_3690,N_3171,N_3460);
or U3691 (N_3691,N_3217,N_3025);
nand U3692 (N_3692,N_3459,N_3372);
xor U3693 (N_3693,N_3387,N_3272);
nor U3694 (N_3694,N_3451,N_3298);
and U3695 (N_3695,N_3244,N_3389);
or U3696 (N_3696,N_3286,N_3231);
nor U3697 (N_3697,N_3002,N_3409);
nor U3698 (N_3698,N_3439,N_3431);
nand U3699 (N_3699,N_3450,N_3196);
nand U3700 (N_3700,N_3164,N_3469);
nand U3701 (N_3701,N_3262,N_3346);
nor U3702 (N_3702,N_3363,N_3123);
nor U3703 (N_3703,N_3243,N_3248);
nand U3704 (N_3704,N_3292,N_3466);
or U3705 (N_3705,N_3126,N_3464);
and U3706 (N_3706,N_3215,N_3474);
nand U3707 (N_3707,N_3263,N_3094);
and U3708 (N_3708,N_3073,N_3162);
nand U3709 (N_3709,N_3042,N_3199);
and U3710 (N_3710,N_3157,N_3052);
nor U3711 (N_3711,N_3207,N_3338);
and U3712 (N_3712,N_3496,N_3072);
nand U3713 (N_3713,N_3059,N_3115);
nand U3714 (N_3714,N_3141,N_3155);
nor U3715 (N_3715,N_3135,N_3381);
nand U3716 (N_3716,N_3067,N_3049);
or U3717 (N_3717,N_3158,N_3483);
nor U3718 (N_3718,N_3305,N_3388);
nor U3719 (N_3719,N_3302,N_3264);
and U3720 (N_3720,N_3019,N_3096);
and U3721 (N_3721,N_3493,N_3004);
and U3722 (N_3722,N_3183,N_3361);
or U3723 (N_3723,N_3296,N_3053);
nand U3724 (N_3724,N_3234,N_3360);
or U3725 (N_3725,N_3012,N_3382);
and U3726 (N_3726,N_3208,N_3227);
and U3727 (N_3727,N_3190,N_3337);
nand U3728 (N_3728,N_3287,N_3430);
or U3729 (N_3729,N_3379,N_3366);
and U3730 (N_3730,N_3050,N_3080);
or U3731 (N_3731,N_3291,N_3370);
or U3732 (N_3732,N_3441,N_3033);
nand U3733 (N_3733,N_3276,N_3201);
and U3734 (N_3734,N_3386,N_3184);
nand U3735 (N_3735,N_3045,N_3423);
and U3736 (N_3736,N_3031,N_3242);
nand U3737 (N_3737,N_3473,N_3397);
xnor U3738 (N_3738,N_3193,N_3290);
nor U3739 (N_3739,N_3214,N_3455);
and U3740 (N_3740,N_3084,N_3317);
or U3741 (N_3741,N_3125,N_3197);
nand U3742 (N_3742,N_3210,N_3150);
xor U3743 (N_3743,N_3132,N_3160);
and U3744 (N_3744,N_3174,N_3145);
nand U3745 (N_3745,N_3176,N_3247);
or U3746 (N_3746,N_3169,N_3026);
nand U3747 (N_3747,N_3443,N_3332);
or U3748 (N_3748,N_3219,N_3213);
nand U3749 (N_3749,N_3436,N_3129);
and U3750 (N_3750,N_3278,N_3106);
or U3751 (N_3751,N_3474,N_3399);
nor U3752 (N_3752,N_3354,N_3217);
nor U3753 (N_3753,N_3213,N_3288);
or U3754 (N_3754,N_3163,N_3340);
nor U3755 (N_3755,N_3195,N_3368);
and U3756 (N_3756,N_3203,N_3416);
nor U3757 (N_3757,N_3308,N_3131);
nor U3758 (N_3758,N_3300,N_3001);
or U3759 (N_3759,N_3172,N_3295);
xor U3760 (N_3760,N_3119,N_3040);
and U3761 (N_3761,N_3346,N_3172);
or U3762 (N_3762,N_3099,N_3180);
and U3763 (N_3763,N_3380,N_3365);
and U3764 (N_3764,N_3016,N_3320);
nor U3765 (N_3765,N_3343,N_3249);
or U3766 (N_3766,N_3016,N_3414);
and U3767 (N_3767,N_3060,N_3351);
xnor U3768 (N_3768,N_3314,N_3281);
xor U3769 (N_3769,N_3026,N_3098);
and U3770 (N_3770,N_3287,N_3375);
and U3771 (N_3771,N_3050,N_3093);
nor U3772 (N_3772,N_3071,N_3064);
and U3773 (N_3773,N_3355,N_3107);
and U3774 (N_3774,N_3265,N_3301);
and U3775 (N_3775,N_3335,N_3427);
xor U3776 (N_3776,N_3253,N_3049);
or U3777 (N_3777,N_3032,N_3304);
xnor U3778 (N_3778,N_3351,N_3475);
or U3779 (N_3779,N_3221,N_3477);
and U3780 (N_3780,N_3048,N_3103);
nand U3781 (N_3781,N_3266,N_3326);
or U3782 (N_3782,N_3445,N_3267);
or U3783 (N_3783,N_3144,N_3135);
nand U3784 (N_3784,N_3102,N_3327);
nand U3785 (N_3785,N_3443,N_3064);
and U3786 (N_3786,N_3324,N_3300);
nand U3787 (N_3787,N_3299,N_3495);
and U3788 (N_3788,N_3265,N_3213);
or U3789 (N_3789,N_3281,N_3427);
or U3790 (N_3790,N_3041,N_3267);
or U3791 (N_3791,N_3050,N_3236);
nand U3792 (N_3792,N_3077,N_3266);
or U3793 (N_3793,N_3110,N_3219);
nand U3794 (N_3794,N_3060,N_3085);
and U3795 (N_3795,N_3479,N_3237);
nand U3796 (N_3796,N_3356,N_3451);
nor U3797 (N_3797,N_3434,N_3318);
or U3798 (N_3798,N_3432,N_3167);
or U3799 (N_3799,N_3451,N_3184);
xnor U3800 (N_3800,N_3049,N_3262);
nor U3801 (N_3801,N_3321,N_3459);
and U3802 (N_3802,N_3169,N_3159);
and U3803 (N_3803,N_3133,N_3398);
xnor U3804 (N_3804,N_3085,N_3224);
or U3805 (N_3805,N_3228,N_3346);
nand U3806 (N_3806,N_3246,N_3142);
or U3807 (N_3807,N_3258,N_3294);
and U3808 (N_3808,N_3175,N_3156);
xnor U3809 (N_3809,N_3023,N_3255);
xnor U3810 (N_3810,N_3372,N_3473);
or U3811 (N_3811,N_3032,N_3145);
and U3812 (N_3812,N_3238,N_3315);
and U3813 (N_3813,N_3022,N_3103);
nor U3814 (N_3814,N_3453,N_3187);
xor U3815 (N_3815,N_3193,N_3437);
nor U3816 (N_3816,N_3213,N_3089);
and U3817 (N_3817,N_3186,N_3406);
or U3818 (N_3818,N_3090,N_3440);
and U3819 (N_3819,N_3297,N_3275);
or U3820 (N_3820,N_3271,N_3286);
nand U3821 (N_3821,N_3267,N_3215);
and U3822 (N_3822,N_3380,N_3228);
nand U3823 (N_3823,N_3383,N_3118);
nand U3824 (N_3824,N_3341,N_3029);
nor U3825 (N_3825,N_3227,N_3119);
xor U3826 (N_3826,N_3373,N_3129);
xor U3827 (N_3827,N_3086,N_3339);
nand U3828 (N_3828,N_3032,N_3399);
xnor U3829 (N_3829,N_3240,N_3089);
or U3830 (N_3830,N_3226,N_3224);
nand U3831 (N_3831,N_3058,N_3169);
nand U3832 (N_3832,N_3176,N_3236);
nand U3833 (N_3833,N_3194,N_3221);
nand U3834 (N_3834,N_3015,N_3401);
nand U3835 (N_3835,N_3382,N_3299);
and U3836 (N_3836,N_3059,N_3437);
xor U3837 (N_3837,N_3258,N_3297);
nand U3838 (N_3838,N_3251,N_3204);
or U3839 (N_3839,N_3494,N_3190);
or U3840 (N_3840,N_3104,N_3493);
nand U3841 (N_3841,N_3061,N_3188);
nor U3842 (N_3842,N_3080,N_3411);
or U3843 (N_3843,N_3035,N_3452);
xnor U3844 (N_3844,N_3226,N_3360);
nand U3845 (N_3845,N_3428,N_3130);
xnor U3846 (N_3846,N_3204,N_3295);
or U3847 (N_3847,N_3486,N_3358);
xor U3848 (N_3848,N_3453,N_3149);
nor U3849 (N_3849,N_3142,N_3375);
nor U3850 (N_3850,N_3119,N_3373);
nand U3851 (N_3851,N_3145,N_3463);
and U3852 (N_3852,N_3254,N_3037);
and U3853 (N_3853,N_3296,N_3380);
and U3854 (N_3854,N_3038,N_3307);
and U3855 (N_3855,N_3413,N_3475);
xnor U3856 (N_3856,N_3108,N_3370);
or U3857 (N_3857,N_3305,N_3325);
or U3858 (N_3858,N_3425,N_3423);
or U3859 (N_3859,N_3095,N_3336);
and U3860 (N_3860,N_3432,N_3163);
or U3861 (N_3861,N_3103,N_3387);
or U3862 (N_3862,N_3455,N_3176);
or U3863 (N_3863,N_3160,N_3419);
and U3864 (N_3864,N_3468,N_3050);
nand U3865 (N_3865,N_3337,N_3046);
nor U3866 (N_3866,N_3144,N_3032);
nor U3867 (N_3867,N_3437,N_3078);
nand U3868 (N_3868,N_3308,N_3223);
xor U3869 (N_3869,N_3223,N_3210);
or U3870 (N_3870,N_3424,N_3243);
or U3871 (N_3871,N_3195,N_3340);
nor U3872 (N_3872,N_3247,N_3439);
nand U3873 (N_3873,N_3485,N_3039);
nor U3874 (N_3874,N_3465,N_3230);
and U3875 (N_3875,N_3104,N_3465);
and U3876 (N_3876,N_3360,N_3103);
nor U3877 (N_3877,N_3379,N_3188);
nand U3878 (N_3878,N_3395,N_3427);
nand U3879 (N_3879,N_3148,N_3406);
nand U3880 (N_3880,N_3262,N_3193);
or U3881 (N_3881,N_3210,N_3176);
or U3882 (N_3882,N_3000,N_3310);
nor U3883 (N_3883,N_3077,N_3091);
nand U3884 (N_3884,N_3091,N_3335);
nor U3885 (N_3885,N_3085,N_3427);
nor U3886 (N_3886,N_3326,N_3221);
or U3887 (N_3887,N_3378,N_3234);
nand U3888 (N_3888,N_3166,N_3105);
or U3889 (N_3889,N_3323,N_3385);
nand U3890 (N_3890,N_3439,N_3146);
or U3891 (N_3891,N_3115,N_3252);
or U3892 (N_3892,N_3277,N_3490);
nor U3893 (N_3893,N_3059,N_3281);
and U3894 (N_3894,N_3323,N_3371);
and U3895 (N_3895,N_3409,N_3191);
nand U3896 (N_3896,N_3014,N_3297);
nand U3897 (N_3897,N_3481,N_3342);
and U3898 (N_3898,N_3214,N_3481);
and U3899 (N_3899,N_3074,N_3270);
nor U3900 (N_3900,N_3052,N_3355);
nand U3901 (N_3901,N_3465,N_3353);
nand U3902 (N_3902,N_3085,N_3120);
xnor U3903 (N_3903,N_3094,N_3078);
nor U3904 (N_3904,N_3175,N_3478);
and U3905 (N_3905,N_3172,N_3370);
nand U3906 (N_3906,N_3384,N_3425);
nor U3907 (N_3907,N_3004,N_3345);
or U3908 (N_3908,N_3472,N_3361);
nor U3909 (N_3909,N_3274,N_3204);
nand U3910 (N_3910,N_3240,N_3343);
nor U3911 (N_3911,N_3298,N_3348);
xor U3912 (N_3912,N_3457,N_3084);
and U3913 (N_3913,N_3489,N_3423);
nand U3914 (N_3914,N_3324,N_3111);
nand U3915 (N_3915,N_3151,N_3003);
and U3916 (N_3916,N_3273,N_3304);
and U3917 (N_3917,N_3476,N_3040);
or U3918 (N_3918,N_3149,N_3221);
xnor U3919 (N_3919,N_3261,N_3152);
and U3920 (N_3920,N_3057,N_3325);
xnor U3921 (N_3921,N_3328,N_3032);
or U3922 (N_3922,N_3397,N_3436);
nand U3923 (N_3923,N_3139,N_3017);
or U3924 (N_3924,N_3418,N_3410);
and U3925 (N_3925,N_3136,N_3076);
and U3926 (N_3926,N_3103,N_3347);
xor U3927 (N_3927,N_3279,N_3002);
nor U3928 (N_3928,N_3339,N_3297);
nor U3929 (N_3929,N_3369,N_3498);
nand U3930 (N_3930,N_3049,N_3375);
or U3931 (N_3931,N_3442,N_3166);
and U3932 (N_3932,N_3468,N_3466);
xnor U3933 (N_3933,N_3360,N_3352);
nand U3934 (N_3934,N_3030,N_3302);
nor U3935 (N_3935,N_3013,N_3087);
nor U3936 (N_3936,N_3164,N_3341);
nor U3937 (N_3937,N_3009,N_3037);
nand U3938 (N_3938,N_3301,N_3476);
nor U3939 (N_3939,N_3202,N_3352);
and U3940 (N_3940,N_3121,N_3458);
or U3941 (N_3941,N_3036,N_3108);
nand U3942 (N_3942,N_3292,N_3021);
nor U3943 (N_3943,N_3041,N_3409);
nand U3944 (N_3944,N_3271,N_3069);
and U3945 (N_3945,N_3091,N_3203);
and U3946 (N_3946,N_3036,N_3084);
or U3947 (N_3947,N_3131,N_3067);
or U3948 (N_3948,N_3327,N_3333);
nor U3949 (N_3949,N_3472,N_3111);
and U3950 (N_3950,N_3351,N_3287);
or U3951 (N_3951,N_3287,N_3443);
nand U3952 (N_3952,N_3249,N_3018);
and U3953 (N_3953,N_3404,N_3011);
or U3954 (N_3954,N_3468,N_3436);
nor U3955 (N_3955,N_3146,N_3180);
and U3956 (N_3956,N_3276,N_3384);
xor U3957 (N_3957,N_3425,N_3354);
or U3958 (N_3958,N_3005,N_3481);
or U3959 (N_3959,N_3040,N_3375);
and U3960 (N_3960,N_3445,N_3393);
nor U3961 (N_3961,N_3178,N_3198);
or U3962 (N_3962,N_3200,N_3499);
and U3963 (N_3963,N_3371,N_3028);
xor U3964 (N_3964,N_3053,N_3109);
nor U3965 (N_3965,N_3052,N_3361);
or U3966 (N_3966,N_3392,N_3412);
nor U3967 (N_3967,N_3046,N_3049);
or U3968 (N_3968,N_3204,N_3208);
and U3969 (N_3969,N_3456,N_3168);
and U3970 (N_3970,N_3291,N_3299);
nor U3971 (N_3971,N_3488,N_3044);
nor U3972 (N_3972,N_3170,N_3358);
xnor U3973 (N_3973,N_3091,N_3155);
xnor U3974 (N_3974,N_3057,N_3495);
nor U3975 (N_3975,N_3167,N_3239);
nor U3976 (N_3976,N_3275,N_3040);
nor U3977 (N_3977,N_3191,N_3291);
or U3978 (N_3978,N_3264,N_3246);
nor U3979 (N_3979,N_3358,N_3221);
or U3980 (N_3980,N_3487,N_3377);
nor U3981 (N_3981,N_3424,N_3096);
and U3982 (N_3982,N_3059,N_3400);
xnor U3983 (N_3983,N_3060,N_3382);
nand U3984 (N_3984,N_3336,N_3443);
nand U3985 (N_3985,N_3316,N_3312);
nand U3986 (N_3986,N_3374,N_3467);
nand U3987 (N_3987,N_3210,N_3309);
and U3988 (N_3988,N_3422,N_3128);
xor U3989 (N_3989,N_3154,N_3243);
or U3990 (N_3990,N_3013,N_3169);
nand U3991 (N_3991,N_3089,N_3448);
or U3992 (N_3992,N_3237,N_3310);
and U3993 (N_3993,N_3470,N_3085);
nand U3994 (N_3994,N_3471,N_3172);
and U3995 (N_3995,N_3007,N_3375);
nand U3996 (N_3996,N_3309,N_3372);
xnor U3997 (N_3997,N_3281,N_3283);
or U3998 (N_3998,N_3152,N_3312);
nor U3999 (N_3999,N_3475,N_3054);
xnor U4000 (N_4000,N_3696,N_3855);
nor U4001 (N_4001,N_3642,N_3879);
nor U4002 (N_4002,N_3638,N_3953);
nor U4003 (N_4003,N_3903,N_3687);
nand U4004 (N_4004,N_3780,N_3663);
or U4005 (N_4005,N_3977,N_3555);
and U4006 (N_4006,N_3521,N_3991);
nor U4007 (N_4007,N_3618,N_3765);
or U4008 (N_4008,N_3827,N_3681);
nand U4009 (N_4009,N_3536,N_3677);
nor U4010 (N_4010,N_3829,N_3598);
and U4011 (N_4011,N_3649,N_3510);
and U4012 (N_4012,N_3632,N_3878);
and U4013 (N_4013,N_3816,N_3695);
and U4014 (N_4014,N_3810,N_3584);
xnor U4015 (N_4015,N_3509,N_3538);
and U4016 (N_4016,N_3885,N_3843);
or U4017 (N_4017,N_3704,N_3819);
nor U4018 (N_4018,N_3852,N_3660);
and U4019 (N_4019,N_3934,N_3769);
and U4020 (N_4020,N_3662,N_3782);
and U4021 (N_4021,N_3808,N_3725);
nand U4022 (N_4022,N_3506,N_3888);
xnor U4023 (N_4023,N_3954,N_3964);
xor U4024 (N_4024,N_3791,N_3668);
nand U4025 (N_4025,N_3925,N_3548);
nand U4026 (N_4026,N_3607,N_3856);
nand U4027 (N_4027,N_3570,N_3661);
and U4028 (N_4028,N_3535,N_3796);
nor U4029 (N_4029,N_3659,N_3970);
nand U4030 (N_4030,N_3624,N_3591);
nor U4031 (N_4031,N_3701,N_3545);
or U4032 (N_4032,N_3542,N_3576);
or U4033 (N_4033,N_3636,N_3669);
nor U4034 (N_4034,N_3914,N_3945);
and U4035 (N_4035,N_3919,N_3958);
nor U4036 (N_4036,N_3795,N_3920);
nor U4037 (N_4037,N_3771,N_3844);
and U4038 (N_4038,N_3626,N_3528);
nand U4039 (N_4039,N_3941,N_3880);
nand U4040 (N_4040,N_3889,N_3788);
nand U4041 (N_4041,N_3899,N_3520);
xnor U4042 (N_4042,N_3666,N_3806);
nand U4043 (N_4043,N_3875,N_3841);
xnor U4044 (N_4044,N_3730,N_3755);
nor U4045 (N_4045,N_3680,N_3734);
or U4046 (N_4046,N_3742,N_3840);
and U4047 (N_4047,N_3686,N_3505);
nand U4048 (N_4048,N_3747,N_3698);
and U4049 (N_4049,N_3532,N_3592);
and U4050 (N_4050,N_3785,N_3824);
or U4051 (N_4051,N_3679,N_3751);
nor U4052 (N_4052,N_3574,N_3719);
and U4053 (N_4053,N_3857,N_3552);
or U4054 (N_4054,N_3781,N_3616);
nand U4055 (N_4055,N_3717,N_3603);
nand U4056 (N_4056,N_3718,N_3709);
and U4057 (N_4057,N_3842,N_3646);
and U4058 (N_4058,N_3516,N_3942);
or U4059 (N_4059,N_3502,N_3514);
xnor U4060 (N_4060,N_3926,N_3960);
nor U4061 (N_4061,N_3931,N_3873);
or U4062 (N_4062,N_3923,N_3994);
xor U4063 (N_4063,N_3947,N_3815);
nor U4064 (N_4064,N_3537,N_3943);
xor U4065 (N_4065,N_3645,N_3764);
and U4066 (N_4066,N_3956,N_3614);
xnor U4067 (N_4067,N_3658,N_3861);
nand U4068 (N_4068,N_3775,N_3854);
nand U4069 (N_4069,N_3590,N_3809);
nand U4070 (N_4070,N_3665,N_3524);
or U4071 (N_4071,N_3541,N_3507);
nand U4072 (N_4072,N_3863,N_3884);
nand U4073 (N_4073,N_3901,N_3556);
nor U4074 (N_4074,N_3655,N_3729);
nor U4075 (N_4075,N_3776,N_3896);
nor U4076 (N_4076,N_3594,N_3741);
or U4077 (N_4077,N_3948,N_3969);
or U4078 (N_4078,N_3817,N_3721);
nand U4079 (N_4079,N_3876,N_3579);
nor U4080 (N_4080,N_3886,N_3830);
nor U4081 (N_4081,N_3581,N_3911);
and U4082 (N_4082,N_3800,N_3732);
or U4083 (N_4083,N_3531,N_3743);
and U4084 (N_4084,N_3568,N_3892);
nor U4085 (N_4085,N_3707,N_3625);
xnor U4086 (N_4086,N_3980,N_3508);
nand U4087 (N_4087,N_3727,N_3897);
nor U4088 (N_4088,N_3550,N_3768);
and U4089 (N_4089,N_3848,N_3786);
nand U4090 (N_4090,N_3986,N_3564);
and U4091 (N_4091,N_3601,N_3975);
or U4092 (N_4092,N_3998,N_3647);
xnor U4093 (N_4093,N_3544,N_3546);
nor U4094 (N_4094,N_3633,N_3569);
and U4095 (N_4095,N_3613,N_3551);
or U4096 (N_4096,N_3756,N_3676);
nor U4097 (N_4097,N_3936,N_3959);
nor U4098 (N_4098,N_3804,N_3835);
xor U4099 (N_4099,N_3723,N_3833);
and U4100 (N_4100,N_3987,N_3634);
nand U4101 (N_4101,N_3602,N_3553);
or U4102 (N_4102,N_3990,N_3600);
nand U4103 (N_4103,N_3525,N_3907);
nand U4104 (N_4104,N_3716,N_3682);
and U4105 (N_4105,N_3563,N_3512);
or U4106 (N_4106,N_3823,N_3963);
or U4107 (N_4107,N_3706,N_3916);
and U4108 (N_4108,N_3818,N_3891);
nand U4109 (N_4109,N_3801,N_3710);
nor U4110 (N_4110,N_3978,N_3935);
and U4111 (N_4111,N_3872,N_3587);
nor U4112 (N_4112,N_3639,N_3859);
and U4113 (N_4113,N_3641,N_3828);
or U4114 (N_4114,N_3597,N_3648);
nand U4115 (N_4115,N_3714,N_3814);
nand U4116 (N_4116,N_3517,N_3928);
and U4117 (N_4117,N_3985,N_3692);
and U4118 (N_4118,N_3612,N_3789);
and U4119 (N_4119,N_3684,N_3893);
and U4120 (N_4120,N_3733,N_3699);
nand U4121 (N_4121,N_3922,N_3866);
nand U4122 (N_4122,N_3713,N_3522);
or U4123 (N_4123,N_3562,N_3822);
nor U4124 (N_4124,N_3534,N_3939);
and U4125 (N_4125,N_3580,N_3573);
nand U4126 (N_4126,N_3883,N_3983);
and U4127 (N_4127,N_3627,N_3981);
nor U4128 (N_4128,N_3762,N_3858);
nor U4129 (N_4129,N_3500,N_3740);
nand U4130 (N_4130,N_3974,N_3831);
and U4131 (N_4131,N_3637,N_3606);
nor U4132 (N_4132,N_3685,N_3812);
and U4133 (N_4133,N_3595,N_3558);
nand U4134 (N_4134,N_3797,N_3838);
and U4135 (N_4135,N_3862,N_3644);
nand U4136 (N_4136,N_3811,N_3973);
and U4137 (N_4137,N_3937,N_3547);
nor U4138 (N_4138,N_3825,N_3993);
nor U4139 (N_4139,N_3772,N_3674);
or U4140 (N_4140,N_3820,N_3821);
and U4141 (N_4141,N_3582,N_3615);
and U4142 (N_4142,N_3846,N_3657);
or U4143 (N_4143,N_3715,N_3708);
nand U4144 (N_4144,N_3799,N_3955);
or U4145 (N_4145,N_3807,N_3503);
nand U4146 (N_4146,N_3930,N_3794);
or U4147 (N_4147,N_3826,N_3868);
nor U4148 (N_4148,N_3513,N_3559);
nand U4149 (N_4149,N_3654,N_3611);
xnor U4150 (N_4150,N_3619,N_3881);
or U4151 (N_4151,N_3577,N_3608);
and U4152 (N_4152,N_3766,N_3770);
xnor U4153 (N_4153,N_3629,N_3750);
xor U4154 (N_4154,N_3957,N_3999);
and U4155 (N_4155,N_3773,N_3691);
or U4156 (N_4156,N_3683,N_3620);
nor U4157 (N_4157,N_3643,N_3927);
nor U4158 (N_4158,N_3705,N_3805);
nor U4159 (N_4159,N_3748,N_3908);
and U4160 (N_4160,N_3651,N_3752);
or U4161 (N_4161,N_3539,N_3790);
nor U4162 (N_4162,N_3971,N_3952);
or U4163 (N_4163,N_3519,N_3864);
nor U4164 (N_4164,N_3837,N_3917);
and U4165 (N_4165,N_3774,N_3929);
xnor U4166 (N_4166,N_3898,N_3951);
and U4167 (N_4167,N_3921,N_3874);
or U4168 (N_4168,N_3554,N_3787);
and U4169 (N_4169,N_3754,N_3966);
and U4170 (N_4170,N_3967,N_3915);
and U4171 (N_4171,N_3575,N_3736);
nand U4172 (N_4172,N_3778,N_3972);
or U4173 (N_4173,N_3869,N_3895);
nor U4174 (N_4174,N_3913,N_3739);
nor U4175 (N_4175,N_3832,N_3653);
xnor U4176 (N_4176,N_3995,N_3757);
and U4177 (N_4177,N_3759,N_3902);
and U4178 (N_4178,N_3912,N_3567);
nor U4179 (N_4179,N_3882,N_3946);
nand U4180 (N_4180,N_3758,N_3847);
xnor U4181 (N_4181,N_3924,N_3753);
nand U4182 (N_4182,N_3932,N_3851);
and U4183 (N_4183,N_3617,N_3760);
or U4184 (N_4184,N_3565,N_3802);
nand U4185 (N_4185,N_3693,N_3652);
and U4186 (N_4186,N_3867,N_3989);
nand U4187 (N_4187,N_3673,N_3877);
xnor U4188 (N_4188,N_3529,N_3839);
nor U4189 (N_4189,N_3511,N_3560);
nand U4190 (N_4190,N_3585,N_3557);
or U4191 (N_4191,N_3656,N_3792);
xor U4192 (N_4192,N_3783,N_3853);
nor U4193 (N_4193,N_3890,N_3870);
nand U4194 (N_4194,N_3860,N_3672);
nor U4195 (N_4195,N_3635,N_3593);
xor U4196 (N_4196,N_3530,N_3578);
xor U4197 (N_4197,N_3744,N_3533);
or U4198 (N_4198,N_3523,N_3605);
nor U4199 (N_4199,N_3737,N_3933);
nand U4200 (N_4200,N_3887,N_3767);
or U4201 (N_4201,N_3982,N_3678);
nand U4202 (N_4202,N_3992,N_3621);
nand U4203 (N_4203,N_3849,N_3588);
and U4204 (N_4204,N_3738,N_3749);
nor U4205 (N_4205,N_3798,N_3720);
and U4206 (N_4206,N_3664,N_3640);
and U4207 (N_4207,N_3979,N_3905);
nand U4208 (N_4208,N_3604,N_3813);
or U4209 (N_4209,N_3962,N_3894);
and U4210 (N_4210,N_3845,N_3630);
nor U4211 (N_4211,N_3540,N_3865);
or U4212 (N_4212,N_3728,N_3900);
xor U4213 (N_4213,N_3735,N_3566);
and U4214 (N_4214,N_3918,N_3834);
nor U4215 (N_4215,N_3504,N_3910);
nor U4216 (N_4216,N_3631,N_3984);
nand U4217 (N_4217,N_3694,N_3961);
or U4218 (N_4218,N_3724,N_3777);
or U4219 (N_4219,N_3988,N_3561);
nor U4220 (N_4220,N_3596,N_3609);
or U4221 (N_4221,N_3622,N_3906);
nor U4222 (N_4222,N_3836,N_3722);
and U4223 (N_4223,N_3518,N_3700);
nor U4224 (N_4224,N_3549,N_3589);
nor U4225 (N_4225,N_3731,N_3586);
nand U4226 (N_4226,N_3940,N_3583);
nand U4227 (N_4227,N_3976,N_3965);
nor U4228 (N_4228,N_3697,N_3793);
xnor U4229 (N_4229,N_3726,N_3689);
and U4230 (N_4230,N_3904,N_3850);
xor U4231 (N_4231,N_3670,N_3690);
nand U4232 (N_4232,N_3871,N_3628);
nor U4233 (N_4233,N_3688,N_3599);
nor U4234 (N_4234,N_3711,N_3944);
nand U4235 (N_4235,N_3909,N_3543);
and U4236 (N_4236,N_3996,N_3997);
or U4237 (N_4237,N_3675,N_3950);
nand U4238 (N_4238,N_3526,N_3779);
and U4239 (N_4239,N_3968,N_3938);
xnor U4240 (N_4240,N_3527,N_3623);
xor U4241 (N_4241,N_3610,N_3949);
or U4242 (N_4242,N_3572,N_3571);
or U4243 (N_4243,N_3515,N_3763);
and U4244 (N_4244,N_3671,N_3784);
nor U4245 (N_4245,N_3501,N_3702);
and U4246 (N_4246,N_3803,N_3650);
nand U4247 (N_4247,N_3761,N_3667);
and U4248 (N_4248,N_3746,N_3745);
and U4249 (N_4249,N_3703,N_3712);
and U4250 (N_4250,N_3579,N_3747);
or U4251 (N_4251,N_3589,N_3762);
nand U4252 (N_4252,N_3632,N_3927);
or U4253 (N_4253,N_3688,N_3674);
xor U4254 (N_4254,N_3537,N_3646);
nand U4255 (N_4255,N_3692,N_3606);
nand U4256 (N_4256,N_3505,N_3597);
and U4257 (N_4257,N_3802,N_3702);
nor U4258 (N_4258,N_3984,N_3828);
xor U4259 (N_4259,N_3907,N_3667);
nand U4260 (N_4260,N_3945,N_3580);
and U4261 (N_4261,N_3734,N_3584);
nor U4262 (N_4262,N_3909,N_3953);
and U4263 (N_4263,N_3998,N_3595);
nor U4264 (N_4264,N_3696,N_3852);
nor U4265 (N_4265,N_3879,N_3902);
nor U4266 (N_4266,N_3772,N_3900);
or U4267 (N_4267,N_3530,N_3550);
nor U4268 (N_4268,N_3760,N_3628);
or U4269 (N_4269,N_3606,N_3665);
or U4270 (N_4270,N_3922,N_3576);
and U4271 (N_4271,N_3986,N_3604);
nand U4272 (N_4272,N_3952,N_3616);
and U4273 (N_4273,N_3935,N_3681);
nor U4274 (N_4274,N_3645,N_3906);
xnor U4275 (N_4275,N_3513,N_3535);
and U4276 (N_4276,N_3890,N_3902);
nor U4277 (N_4277,N_3776,N_3804);
or U4278 (N_4278,N_3709,N_3952);
and U4279 (N_4279,N_3945,N_3736);
nor U4280 (N_4280,N_3620,N_3623);
nor U4281 (N_4281,N_3769,N_3847);
or U4282 (N_4282,N_3827,N_3651);
nand U4283 (N_4283,N_3604,N_3893);
or U4284 (N_4284,N_3792,N_3619);
nor U4285 (N_4285,N_3662,N_3920);
nand U4286 (N_4286,N_3863,N_3580);
nor U4287 (N_4287,N_3834,N_3657);
or U4288 (N_4288,N_3834,N_3660);
or U4289 (N_4289,N_3626,N_3603);
xor U4290 (N_4290,N_3614,N_3903);
or U4291 (N_4291,N_3856,N_3584);
nand U4292 (N_4292,N_3621,N_3903);
and U4293 (N_4293,N_3980,N_3725);
or U4294 (N_4294,N_3506,N_3783);
nand U4295 (N_4295,N_3557,N_3822);
nand U4296 (N_4296,N_3942,N_3976);
nand U4297 (N_4297,N_3960,N_3614);
nand U4298 (N_4298,N_3665,N_3899);
xnor U4299 (N_4299,N_3873,N_3990);
or U4300 (N_4300,N_3554,N_3840);
nor U4301 (N_4301,N_3671,N_3812);
nor U4302 (N_4302,N_3500,N_3651);
nand U4303 (N_4303,N_3781,N_3787);
nor U4304 (N_4304,N_3527,N_3692);
or U4305 (N_4305,N_3786,N_3887);
nand U4306 (N_4306,N_3966,N_3777);
or U4307 (N_4307,N_3842,N_3708);
or U4308 (N_4308,N_3766,N_3721);
or U4309 (N_4309,N_3587,N_3605);
nand U4310 (N_4310,N_3927,N_3727);
nor U4311 (N_4311,N_3715,N_3772);
or U4312 (N_4312,N_3950,N_3960);
and U4313 (N_4313,N_3671,N_3624);
and U4314 (N_4314,N_3959,N_3608);
xor U4315 (N_4315,N_3829,N_3611);
nand U4316 (N_4316,N_3821,N_3782);
nand U4317 (N_4317,N_3588,N_3793);
and U4318 (N_4318,N_3525,N_3831);
or U4319 (N_4319,N_3660,N_3939);
nor U4320 (N_4320,N_3552,N_3541);
or U4321 (N_4321,N_3774,N_3865);
nand U4322 (N_4322,N_3708,N_3750);
or U4323 (N_4323,N_3550,N_3874);
or U4324 (N_4324,N_3846,N_3826);
nor U4325 (N_4325,N_3978,N_3912);
nand U4326 (N_4326,N_3572,N_3965);
or U4327 (N_4327,N_3861,N_3511);
and U4328 (N_4328,N_3696,N_3721);
and U4329 (N_4329,N_3631,N_3642);
nor U4330 (N_4330,N_3877,N_3830);
and U4331 (N_4331,N_3898,N_3857);
and U4332 (N_4332,N_3739,N_3798);
or U4333 (N_4333,N_3987,N_3915);
nor U4334 (N_4334,N_3804,N_3716);
nor U4335 (N_4335,N_3983,N_3605);
and U4336 (N_4336,N_3500,N_3875);
and U4337 (N_4337,N_3737,N_3729);
nand U4338 (N_4338,N_3727,N_3780);
nand U4339 (N_4339,N_3952,N_3969);
nor U4340 (N_4340,N_3817,N_3672);
nand U4341 (N_4341,N_3711,N_3931);
and U4342 (N_4342,N_3893,N_3735);
nand U4343 (N_4343,N_3939,N_3686);
xor U4344 (N_4344,N_3548,N_3621);
nand U4345 (N_4345,N_3640,N_3993);
and U4346 (N_4346,N_3983,N_3919);
nand U4347 (N_4347,N_3906,N_3866);
nor U4348 (N_4348,N_3818,N_3895);
nor U4349 (N_4349,N_3735,N_3800);
or U4350 (N_4350,N_3671,N_3838);
nor U4351 (N_4351,N_3517,N_3597);
nand U4352 (N_4352,N_3817,N_3614);
nand U4353 (N_4353,N_3993,N_3525);
nor U4354 (N_4354,N_3916,N_3763);
nor U4355 (N_4355,N_3644,N_3682);
and U4356 (N_4356,N_3880,N_3663);
or U4357 (N_4357,N_3513,N_3871);
nand U4358 (N_4358,N_3985,N_3723);
and U4359 (N_4359,N_3775,N_3823);
or U4360 (N_4360,N_3808,N_3611);
nor U4361 (N_4361,N_3975,N_3646);
or U4362 (N_4362,N_3786,N_3811);
and U4363 (N_4363,N_3661,N_3911);
and U4364 (N_4364,N_3638,N_3787);
and U4365 (N_4365,N_3718,N_3810);
nor U4366 (N_4366,N_3563,N_3664);
nand U4367 (N_4367,N_3721,N_3504);
nor U4368 (N_4368,N_3610,N_3700);
and U4369 (N_4369,N_3639,N_3895);
and U4370 (N_4370,N_3893,N_3673);
nand U4371 (N_4371,N_3970,N_3717);
or U4372 (N_4372,N_3616,N_3752);
xor U4373 (N_4373,N_3905,N_3692);
nand U4374 (N_4374,N_3674,N_3904);
nor U4375 (N_4375,N_3726,N_3810);
and U4376 (N_4376,N_3637,N_3856);
and U4377 (N_4377,N_3527,N_3877);
nor U4378 (N_4378,N_3585,N_3728);
and U4379 (N_4379,N_3920,N_3700);
and U4380 (N_4380,N_3750,N_3522);
or U4381 (N_4381,N_3906,N_3730);
nor U4382 (N_4382,N_3806,N_3690);
nor U4383 (N_4383,N_3900,N_3501);
xor U4384 (N_4384,N_3645,N_3926);
or U4385 (N_4385,N_3654,N_3644);
and U4386 (N_4386,N_3928,N_3516);
nand U4387 (N_4387,N_3535,N_3559);
nor U4388 (N_4388,N_3998,N_3722);
nand U4389 (N_4389,N_3903,N_3818);
or U4390 (N_4390,N_3984,N_3807);
nor U4391 (N_4391,N_3997,N_3759);
nor U4392 (N_4392,N_3597,N_3547);
xnor U4393 (N_4393,N_3661,N_3874);
nor U4394 (N_4394,N_3846,N_3939);
nand U4395 (N_4395,N_3971,N_3593);
or U4396 (N_4396,N_3849,N_3535);
nand U4397 (N_4397,N_3816,N_3595);
nand U4398 (N_4398,N_3737,N_3685);
and U4399 (N_4399,N_3983,N_3917);
or U4400 (N_4400,N_3979,N_3523);
nand U4401 (N_4401,N_3700,N_3880);
nand U4402 (N_4402,N_3930,N_3671);
xor U4403 (N_4403,N_3717,N_3978);
nand U4404 (N_4404,N_3526,N_3919);
nor U4405 (N_4405,N_3946,N_3901);
xnor U4406 (N_4406,N_3891,N_3678);
and U4407 (N_4407,N_3916,N_3905);
nor U4408 (N_4408,N_3996,N_3753);
nor U4409 (N_4409,N_3523,N_3865);
xnor U4410 (N_4410,N_3537,N_3761);
and U4411 (N_4411,N_3942,N_3537);
nand U4412 (N_4412,N_3682,N_3925);
xnor U4413 (N_4413,N_3927,N_3779);
and U4414 (N_4414,N_3557,N_3728);
and U4415 (N_4415,N_3932,N_3762);
nand U4416 (N_4416,N_3735,N_3814);
nand U4417 (N_4417,N_3814,N_3598);
and U4418 (N_4418,N_3663,N_3904);
nor U4419 (N_4419,N_3984,N_3650);
nand U4420 (N_4420,N_3939,N_3584);
or U4421 (N_4421,N_3689,N_3965);
nor U4422 (N_4422,N_3849,N_3799);
and U4423 (N_4423,N_3954,N_3753);
nor U4424 (N_4424,N_3575,N_3953);
nor U4425 (N_4425,N_3688,N_3691);
xor U4426 (N_4426,N_3988,N_3599);
nand U4427 (N_4427,N_3701,N_3581);
or U4428 (N_4428,N_3637,N_3645);
nor U4429 (N_4429,N_3797,N_3613);
nand U4430 (N_4430,N_3578,N_3675);
nand U4431 (N_4431,N_3547,N_3924);
xor U4432 (N_4432,N_3862,N_3899);
and U4433 (N_4433,N_3797,N_3992);
or U4434 (N_4434,N_3594,N_3792);
and U4435 (N_4435,N_3904,N_3846);
and U4436 (N_4436,N_3787,N_3894);
nor U4437 (N_4437,N_3594,N_3790);
nand U4438 (N_4438,N_3969,N_3752);
or U4439 (N_4439,N_3851,N_3597);
or U4440 (N_4440,N_3718,N_3629);
nor U4441 (N_4441,N_3900,N_3907);
and U4442 (N_4442,N_3960,N_3602);
xnor U4443 (N_4443,N_3793,N_3907);
xnor U4444 (N_4444,N_3518,N_3699);
xor U4445 (N_4445,N_3937,N_3817);
nand U4446 (N_4446,N_3983,N_3937);
or U4447 (N_4447,N_3710,N_3742);
xnor U4448 (N_4448,N_3617,N_3856);
xor U4449 (N_4449,N_3512,N_3597);
or U4450 (N_4450,N_3750,N_3731);
or U4451 (N_4451,N_3938,N_3703);
nor U4452 (N_4452,N_3669,N_3961);
nand U4453 (N_4453,N_3974,N_3765);
nand U4454 (N_4454,N_3993,N_3580);
and U4455 (N_4455,N_3813,N_3859);
or U4456 (N_4456,N_3943,N_3647);
or U4457 (N_4457,N_3912,N_3509);
nand U4458 (N_4458,N_3760,N_3898);
or U4459 (N_4459,N_3855,N_3939);
nand U4460 (N_4460,N_3564,N_3864);
xnor U4461 (N_4461,N_3845,N_3708);
nand U4462 (N_4462,N_3643,N_3565);
nand U4463 (N_4463,N_3807,N_3803);
nand U4464 (N_4464,N_3901,N_3700);
and U4465 (N_4465,N_3793,N_3806);
nand U4466 (N_4466,N_3838,N_3983);
and U4467 (N_4467,N_3735,N_3671);
or U4468 (N_4468,N_3697,N_3698);
nor U4469 (N_4469,N_3844,N_3669);
nand U4470 (N_4470,N_3996,N_3649);
nor U4471 (N_4471,N_3950,N_3933);
or U4472 (N_4472,N_3862,N_3548);
nor U4473 (N_4473,N_3665,N_3891);
xor U4474 (N_4474,N_3766,N_3724);
and U4475 (N_4475,N_3945,N_3560);
and U4476 (N_4476,N_3606,N_3851);
nor U4477 (N_4477,N_3535,N_3913);
nor U4478 (N_4478,N_3976,N_3986);
and U4479 (N_4479,N_3812,N_3609);
nand U4480 (N_4480,N_3751,N_3942);
and U4481 (N_4481,N_3945,N_3944);
or U4482 (N_4482,N_3850,N_3967);
nor U4483 (N_4483,N_3948,N_3644);
or U4484 (N_4484,N_3894,N_3651);
and U4485 (N_4485,N_3961,N_3800);
and U4486 (N_4486,N_3910,N_3791);
nand U4487 (N_4487,N_3558,N_3682);
or U4488 (N_4488,N_3770,N_3719);
xor U4489 (N_4489,N_3665,N_3601);
nor U4490 (N_4490,N_3895,N_3796);
nor U4491 (N_4491,N_3635,N_3795);
nor U4492 (N_4492,N_3888,N_3960);
nor U4493 (N_4493,N_3648,N_3946);
xnor U4494 (N_4494,N_3652,N_3962);
or U4495 (N_4495,N_3562,N_3759);
and U4496 (N_4496,N_3528,N_3610);
nand U4497 (N_4497,N_3711,N_3998);
nor U4498 (N_4498,N_3925,N_3999);
nand U4499 (N_4499,N_3593,N_3579);
nor U4500 (N_4500,N_4084,N_4362);
xor U4501 (N_4501,N_4267,N_4283);
or U4502 (N_4502,N_4399,N_4341);
and U4503 (N_4503,N_4478,N_4214);
and U4504 (N_4504,N_4481,N_4237);
or U4505 (N_4505,N_4291,N_4077);
nor U4506 (N_4506,N_4152,N_4236);
nand U4507 (N_4507,N_4171,N_4038);
and U4508 (N_4508,N_4022,N_4133);
nand U4509 (N_4509,N_4434,N_4095);
or U4510 (N_4510,N_4012,N_4272);
nor U4511 (N_4511,N_4223,N_4053);
nor U4512 (N_4512,N_4484,N_4170);
nor U4513 (N_4513,N_4311,N_4342);
or U4514 (N_4514,N_4492,N_4121);
or U4515 (N_4515,N_4308,N_4381);
or U4516 (N_4516,N_4245,N_4301);
and U4517 (N_4517,N_4396,N_4195);
xor U4518 (N_4518,N_4213,N_4243);
nor U4519 (N_4519,N_4219,N_4003);
nor U4520 (N_4520,N_4450,N_4444);
or U4521 (N_4521,N_4394,N_4234);
or U4522 (N_4522,N_4360,N_4462);
nand U4523 (N_4523,N_4007,N_4324);
nor U4524 (N_4524,N_4108,N_4011);
and U4525 (N_4525,N_4157,N_4140);
and U4526 (N_4526,N_4310,N_4355);
and U4527 (N_4527,N_4040,N_4432);
nor U4528 (N_4528,N_4368,N_4338);
or U4529 (N_4529,N_4065,N_4281);
and U4530 (N_4530,N_4202,N_4044);
xnor U4531 (N_4531,N_4015,N_4403);
or U4532 (N_4532,N_4296,N_4114);
xor U4533 (N_4533,N_4454,N_4318);
nand U4534 (N_4534,N_4079,N_4106);
nor U4535 (N_4535,N_4261,N_4174);
nor U4536 (N_4536,N_4321,N_4176);
nor U4537 (N_4537,N_4257,N_4104);
nand U4538 (N_4538,N_4485,N_4410);
nor U4539 (N_4539,N_4442,N_4193);
xor U4540 (N_4540,N_4378,N_4329);
and U4541 (N_4541,N_4000,N_4169);
nand U4542 (N_4542,N_4465,N_4071);
nand U4543 (N_4543,N_4070,N_4479);
xnor U4544 (N_4544,N_4109,N_4483);
or U4545 (N_4545,N_4134,N_4043);
nor U4546 (N_4546,N_4069,N_4282);
nor U4547 (N_4547,N_4495,N_4313);
nand U4548 (N_4548,N_4178,N_4029);
or U4549 (N_4549,N_4499,N_4209);
and U4550 (N_4550,N_4182,N_4306);
xnor U4551 (N_4551,N_4027,N_4112);
and U4552 (N_4552,N_4383,N_4331);
or U4553 (N_4553,N_4074,N_4404);
nand U4554 (N_4554,N_4340,N_4167);
xor U4555 (N_4555,N_4420,N_4183);
xnor U4556 (N_4556,N_4008,N_4446);
xnor U4557 (N_4557,N_4392,N_4142);
nand U4558 (N_4558,N_4376,N_4299);
xor U4559 (N_4559,N_4421,N_4231);
nand U4560 (N_4560,N_4486,N_4302);
xnor U4561 (N_4561,N_4312,N_4241);
nand U4562 (N_4562,N_4041,N_4339);
and U4563 (N_4563,N_4405,N_4344);
or U4564 (N_4564,N_4482,N_4039);
or U4565 (N_4565,N_4144,N_4131);
nand U4566 (N_4566,N_4349,N_4107);
and U4567 (N_4567,N_4045,N_4292);
nor U4568 (N_4568,N_4210,N_4058);
nand U4569 (N_4569,N_4150,N_4332);
or U4570 (N_4570,N_4147,N_4162);
or U4571 (N_4571,N_4297,N_4286);
nand U4572 (N_4572,N_4409,N_4232);
nor U4573 (N_4573,N_4244,N_4087);
and U4574 (N_4574,N_4093,N_4060);
and U4575 (N_4575,N_4334,N_4161);
nand U4576 (N_4576,N_4494,N_4250);
and U4577 (N_4577,N_4304,N_4320);
and U4578 (N_4578,N_4326,N_4088);
or U4579 (N_4579,N_4290,N_4135);
xor U4580 (N_4580,N_4389,N_4227);
or U4581 (N_4581,N_4363,N_4051);
and U4582 (N_4582,N_4422,N_4464);
nand U4583 (N_4583,N_4033,N_4366);
nand U4584 (N_4584,N_4215,N_4443);
or U4585 (N_4585,N_4004,N_4371);
and U4586 (N_4586,N_4273,N_4120);
nand U4587 (N_4587,N_4110,N_4279);
and U4588 (N_4588,N_4092,N_4258);
xor U4589 (N_4589,N_4449,N_4159);
or U4590 (N_4590,N_4248,N_4055);
nand U4591 (N_4591,N_4487,N_4179);
nor U4592 (N_4592,N_4374,N_4445);
and U4593 (N_4593,N_4190,N_4315);
nand U4594 (N_4594,N_4316,N_4327);
nor U4595 (N_4595,N_4275,N_4201);
and U4596 (N_4596,N_4163,N_4205);
or U4597 (N_4597,N_4325,N_4252);
or U4598 (N_4598,N_4437,N_4006);
xnor U4599 (N_4599,N_4390,N_4056);
nor U4600 (N_4600,N_4351,N_4280);
and U4601 (N_4601,N_4352,N_4030);
and U4602 (N_4602,N_4274,N_4278);
nand U4603 (N_4603,N_4059,N_4222);
and U4604 (N_4604,N_4328,N_4477);
and U4605 (N_4605,N_4211,N_4253);
or U4606 (N_4606,N_4300,N_4016);
and U4607 (N_4607,N_4469,N_4401);
or U4608 (N_4608,N_4141,N_4269);
nand U4609 (N_4609,N_4001,N_4361);
and U4610 (N_4610,N_4345,N_4406);
nand U4611 (N_4611,N_4013,N_4184);
nand U4612 (N_4612,N_4028,N_4375);
or U4613 (N_4613,N_4259,N_4117);
nand U4614 (N_4614,N_4335,N_4149);
nand U4615 (N_4615,N_4382,N_4224);
or U4616 (N_4616,N_4357,N_4132);
nand U4617 (N_4617,N_4010,N_4398);
nor U4618 (N_4618,N_4451,N_4367);
xnor U4619 (N_4619,N_4026,N_4113);
and U4620 (N_4620,N_4452,N_4350);
and U4621 (N_4621,N_4294,N_4271);
and U4622 (N_4622,N_4025,N_4090);
and U4623 (N_4623,N_4393,N_4139);
nand U4624 (N_4624,N_4124,N_4458);
xnor U4625 (N_4625,N_4086,N_4433);
nor U4626 (N_4626,N_4032,N_4081);
xnor U4627 (N_4627,N_4066,N_4154);
or U4628 (N_4628,N_4118,N_4097);
nor U4629 (N_4629,N_4192,N_4457);
nor U4630 (N_4630,N_4125,N_4158);
xor U4631 (N_4631,N_4031,N_4206);
nand U4632 (N_4632,N_4387,N_4343);
nor U4633 (N_4633,N_4220,N_4212);
and U4634 (N_4634,N_4050,N_4194);
and U4635 (N_4635,N_4242,N_4166);
or U4636 (N_4636,N_4230,N_4129);
or U4637 (N_4637,N_4436,N_4122);
nor U4638 (N_4638,N_4100,N_4412);
or U4639 (N_4639,N_4415,N_4498);
and U4640 (N_4640,N_4238,N_4063);
nand U4641 (N_4641,N_4068,N_4018);
xor U4642 (N_4642,N_4263,N_4397);
nand U4643 (N_4643,N_4064,N_4151);
xor U4644 (N_4644,N_4333,N_4395);
nor U4645 (N_4645,N_4293,N_4438);
nand U4646 (N_4646,N_4094,N_4285);
nor U4647 (N_4647,N_4468,N_4021);
and U4648 (N_4648,N_4189,N_4160);
or U4649 (N_4649,N_4049,N_4091);
and U4650 (N_4650,N_4270,N_4148);
nor U4651 (N_4651,N_4076,N_4372);
or U4652 (N_4652,N_4407,N_4384);
and U4653 (N_4653,N_4284,N_4348);
nor U4654 (N_4654,N_4082,N_4491);
nor U4655 (N_4655,N_4359,N_4448);
and U4656 (N_4656,N_4254,N_4233);
and U4657 (N_4657,N_4369,N_4196);
xnor U4658 (N_4658,N_4089,N_4489);
or U4659 (N_4659,N_4020,N_4146);
nor U4660 (N_4660,N_4370,N_4391);
nand U4661 (N_4661,N_4240,N_4052);
nor U4662 (N_4662,N_4036,N_4187);
xnor U4663 (N_4663,N_4400,N_4102);
nand U4664 (N_4664,N_4046,N_4017);
xor U4665 (N_4665,N_4085,N_4019);
or U4666 (N_4666,N_4456,N_4365);
and U4667 (N_4667,N_4143,N_4256);
nand U4668 (N_4668,N_4098,N_4266);
nor U4669 (N_4669,N_4164,N_4439);
nor U4670 (N_4670,N_4153,N_4411);
nor U4671 (N_4671,N_4062,N_4042);
nor U4672 (N_4672,N_4037,N_4061);
and U4673 (N_4673,N_4474,N_4265);
nor U4674 (N_4674,N_4425,N_4221);
and U4675 (N_4675,N_4002,N_4471);
nand U4676 (N_4676,N_4466,N_4358);
nor U4677 (N_4677,N_4101,N_4228);
nand U4678 (N_4678,N_4145,N_4418);
xor U4679 (N_4679,N_4175,N_4111);
nand U4680 (N_4680,N_4128,N_4277);
nand U4681 (N_4681,N_4009,N_4419);
and U4682 (N_4682,N_4435,N_4298);
and U4683 (N_4683,N_4386,N_4305);
nor U4684 (N_4684,N_4136,N_4460);
nand U4685 (N_4685,N_4138,N_4226);
nor U4686 (N_4686,N_4441,N_4322);
or U4687 (N_4687,N_4126,N_4303);
nand U4688 (N_4688,N_4289,N_4105);
nand U4689 (N_4689,N_4057,N_4216);
nor U4690 (N_4690,N_4005,N_4455);
or U4691 (N_4691,N_4480,N_4496);
xor U4692 (N_4692,N_4309,N_4307);
and U4693 (N_4693,N_4354,N_4264);
and U4694 (N_4694,N_4488,N_4472);
nor U4695 (N_4695,N_4229,N_4078);
and U4696 (N_4696,N_4048,N_4225);
or U4697 (N_4697,N_4218,N_4447);
and U4698 (N_4698,N_4180,N_4346);
xnor U4699 (N_4699,N_4119,N_4430);
or U4700 (N_4700,N_4424,N_4072);
xor U4701 (N_4701,N_4127,N_4380);
and U4702 (N_4702,N_4373,N_4385);
and U4703 (N_4703,N_4168,N_4185);
and U4704 (N_4704,N_4073,N_4199);
or U4705 (N_4705,N_4249,N_4423);
and U4706 (N_4706,N_4251,N_4083);
and U4707 (N_4707,N_4208,N_4497);
or U4708 (N_4708,N_4356,N_4200);
or U4709 (N_4709,N_4188,N_4276);
nand U4710 (N_4710,N_4463,N_4337);
nor U4711 (N_4711,N_4247,N_4155);
nor U4712 (N_4712,N_4156,N_4217);
nor U4713 (N_4713,N_4130,N_4408);
and U4714 (N_4714,N_4476,N_4467);
or U4715 (N_4715,N_4414,N_4388);
and U4716 (N_4716,N_4426,N_4014);
nand U4717 (N_4717,N_4440,N_4428);
xor U4718 (N_4718,N_4416,N_4123);
or U4719 (N_4719,N_4314,N_4235);
or U4720 (N_4720,N_4493,N_4490);
and U4721 (N_4721,N_4172,N_4475);
nor U4722 (N_4722,N_4287,N_4103);
or U4723 (N_4723,N_4075,N_4198);
or U4724 (N_4724,N_4186,N_4431);
or U4725 (N_4725,N_4067,N_4402);
and U4726 (N_4726,N_4379,N_4099);
nor U4727 (N_4727,N_4096,N_4080);
nand U4728 (N_4728,N_4288,N_4255);
nor U4729 (N_4729,N_4262,N_4024);
nand U4730 (N_4730,N_4364,N_4260);
and U4731 (N_4731,N_4239,N_4417);
nor U4732 (N_4732,N_4181,N_4177);
xor U4733 (N_4733,N_4377,N_4246);
or U4734 (N_4734,N_4427,N_4023);
and U4735 (N_4735,N_4034,N_4115);
or U4736 (N_4736,N_4459,N_4165);
nand U4737 (N_4737,N_4035,N_4295);
and U4738 (N_4738,N_4353,N_4336);
nand U4739 (N_4739,N_4470,N_4054);
or U4740 (N_4740,N_4203,N_4268);
and U4741 (N_4741,N_4317,N_4116);
nor U4742 (N_4742,N_4330,N_4319);
nor U4743 (N_4743,N_4191,N_4429);
nand U4744 (N_4744,N_4453,N_4197);
or U4745 (N_4745,N_4207,N_4473);
and U4746 (N_4746,N_4047,N_4413);
or U4747 (N_4747,N_4204,N_4173);
nor U4748 (N_4748,N_4323,N_4461);
nor U4749 (N_4749,N_4347,N_4137);
xor U4750 (N_4750,N_4156,N_4454);
nand U4751 (N_4751,N_4077,N_4380);
nor U4752 (N_4752,N_4130,N_4145);
nor U4753 (N_4753,N_4243,N_4138);
nor U4754 (N_4754,N_4376,N_4050);
and U4755 (N_4755,N_4447,N_4202);
nand U4756 (N_4756,N_4191,N_4005);
and U4757 (N_4757,N_4174,N_4429);
nor U4758 (N_4758,N_4438,N_4066);
nor U4759 (N_4759,N_4075,N_4217);
xor U4760 (N_4760,N_4006,N_4163);
nor U4761 (N_4761,N_4008,N_4332);
nand U4762 (N_4762,N_4116,N_4070);
and U4763 (N_4763,N_4401,N_4162);
nor U4764 (N_4764,N_4068,N_4008);
nand U4765 (N_4765,N_4065,N_4375);
or U4766 (N_4766,N_4216,N_4334);
or U4767 (N_4767,N_4262,N_4260);
and U4768 (N_4768,N_4493,N_4212);
nor U4769 (N_4769,N_4436,N_4124);
nand U4770 (N_4770,N_4108,N_4331);
and U4771 (N_4771,N_4138,N_4051);
nand U4772 (N_4772,N_4390,N_4170);
or U4773 (N_4773,N_4324,N_4155);
nand U4774 (N_4774,N_4277,N_4039);
xor U4775 (N_4775,N_4214,N_4049);
or U4776 (N_4776,N_4141,N_4389);
xnor U4777 (N_4777,N_4224,N_4229);
xor U4778 (N_4778,N_4007,N_4155);
xor U4779 (N_4779,N_4272,N_4240);
nor U4780 (N_4780,N_4028,N_4100);
or U4781 (N_4781,N_4184,N_4454);
nor U4782 (N_4782,N_4192,N_4088);
or U4783 (N_4783,N_4035,N_4165);
and U4784 (N_4784,N_4188,N_4441);
nor U4785 (N_4785,N_4244,N_4290);
xor U4786 (N_4786,N_4065,N_4360);
nand U4787 (N_4787,N_4302,N_4329);
xnor U4788 (N_4788,N_4188,N_4388);
and U4789 (N_4789,N_4410,N_4173);
nand U4790 (N_4790,N_4357,N_4432);
nor U4791 (N_4791,N_4442,N_4360);
and U4792 (N_4792,N_4094,N_4095);
nand U4793 (N_4793,N_4304,N_4471);
and U4794 (N_4794,N_4052,N_4291);
or U4795 (N_4795,N_4086,N_4379);
and U4796 (N_4796,N_4446,N_4360);
xnor U4797 (N_4797,N_4485,N_4000);
or U4798 (N_4798,N_4214,N_4339);
or U4799 (N_4799,N_4110,N_4010);
and U4800 (N_4800,N_4416,N_4200);
or U4801 (N_4801,N_4301,N_4401);
or U4802 (N_4802,N_4130,N_4373);
nor U4803 (N_4803,N_4495,N_4113);
and U4804 (N_4804,N_4420,N_4029);
nor U4805 (N_4805,N_4129,N_4443);
and U4806 (N_4806,N_4200,N_4097);
nand U4807 (N_4807,N_4272,N_4232);
or U4808 (N_4808,N_4086,N_4217);
and U4809 (N_4809,N_4001,N_4392);
xnor U4810 (N_4810,N_4251,N_4250);
nand U4811 (N_4811,N_4377,N_4482);
nand U4812 (N_4812,N_4113,N_4069);
nand U4813 (N_4813,N_4161,N_4117);
nor U4814 (N_4814,N_4113,N_4432);
nor U4815 (N_4815,N_4257,N_4364);
and U4816 (N_4816,N_4465,N_4079);
or U4817 (N_4817,N_4218,N_4023);
and U4818 (N_4818,N_4059,N_4140);
nand U4819 (N_4819,N_4316,N_4317);
and U4820 (N_4820,N_4087,N_4151);
nor U4821 (N_4821,N_4380,N_4157);
and U4822 (N_4822,N_4466,N_4372);
nor U4823 (N_4823,N_4297,N_4063);
and U4824 (N_4824,N_4125,N_4396);
nand U4825 (N_4825,N_4038,N_4137);
nand U4826 (N_4826,N_4002,N_4164);
or U4827 (N_4827,N_4117,N_4080);
nor U4828 (N_4828,N_4031,N_4171);
and U4829 (N_4829,N_4060,N_4180);
and U4830 (N_4830,N_4138,N_4027);
or U4831 (N_4831,N_4154,N_4013);
nor U4832 (N_4832,N_4472,N_4058);
nand U4833 (N_4833,N_4040,N_4108);
or U4834 (N_4834,N_4413,N_4361);
nand U4835 (N_4835,N_4411,N_4489);
nor U4836 (N_4836,N_4313,N_4316);
or U4837 (N_4837,N_4133,N_4083);
nand U4838 (N_4838,N_4210,N_4321);
nor U4839 (N_4839,N_4225,N_4142);
nand U4840 (N_4840,N_4344,N_4039);
xnor U4841 (N_4841,N_4226,N_4233);
or U4842 (N_4842,N_4037,N_4409);
or U4843 (N_4843,N_4422,N_4037);
and U4844 (N_4844,N_4380,N_4322);
nor U4845 (N_4845,N_4097,N_4145);
nor U4846 (N_4846,N_4473,N_4105);
xor U4847 (N_4847,N_4241,N_4494);
nand U4848 (N_4848,N_4473,N_4369);
and U4849 (N_4849,N_4150,N_4136);
nor U4850 (N_4850,N_4343,N_4473);
nand U4851 (N_4851,N_4009,N_4308);
nor U4852 (N_4852,N_4442,N_4296);
or U4853 (N_4853,N_4230,N_4499);
nor U4854 (N_4854,N_4151,N_4083);
nor U4855 (N_4855,N_4102,N_4433);
or U4856 (N_4856,N_4177,N_4252);
and U4857 (N_4857,N_4329,N_4373);
xor U4858 (N_4858,N_4023,N_4060);
xnor U4859 (N_4859,N_4462,N_4249);
or U4860 (N_4860,N_4306,N_4269);
or U4861 (N_4861,N_4091,N_4106);
and U4862 (N_4862,N_4277,N_4191);
nand U4863 (N_4863,N_4055,N_4221);
or U4864 (N_4864,N_4229,N_4186);
nand U4865 (N_4865,N_4237,N_4495);
and U4866 (N_4866,N_4442,N_4358);
and U4867 (N_4867,N_4078,N_4362);
and U4868 (N_4868,N_4036,N_4242);
or U4869 (N_4869,N_4263,N_4276);
and U4870 (N_4870,N_4427,N_4456);
and U4871 (N_4871,N_4241,N_4131);
nor U4872 (N_4872,N_4009,N_4185);
nand U4873 (N_4873,N_4176,N_4363);
nand U4874 (N_4874,N_4343,N_4261);
and U4875 (N_4875,N_4095,N_4212);
nand U4876 (N_4876,N_4162,N_4326);
and U4877 (N_4877,N_4339,N_4383);
or U4878 (N_4878,N_4223,N_4335);
nand U4879 (N_4879,N_4124,N_4128);
nand U4880 (N_4880,N_4246,N_4139);
or U4881 (N_4881,N_4053,N_4092);
nand U4882 (N_4882,N_4173,N_4217);
and U4883 (N_4883,N_4151,N_4347);
or U4884 (N_4884,N_4319,N_4376);
nor U4885 (N_4885,N_4499,N_4264);
or U4886 (N_4886,N_4375,N_4166);
and U4887 (N_4887,N_4437,N_4250);
nand U4888 (N_4888,N_4386,N_4181);
nand U4889 (N_4889,N_4404,N_4203);
nand U4890 (N_4890,N_4067,N_4396);
nand U4891 (N_4891,N_4483,N_4116);
nand U4892 (N_4892,N_4437,N_4471);
nand U4893 (N_4893,N_4419,N_4347);
nand U4894 (N_4894,N_4492,N_4306);
or U4895 (N_4895,N_4030,N_4487);
or U4896 (N_4896,N_4140,N_4008);
and U4897 (N_4897,N_4144,N_4346);
nor U4898 (N_4898,N_4338,N_4442);
nand U4899 (N_4899,N_4032,N_4481);
xor U4900 (N_4900,N_4256,N_4213);
nand U4901 (N_4901,N_4370,N_4166);
nor U4902 (N_4902,N_4205,N_4074);
or U4903 (N_4903,N_4055,N_4222);
or U4904 (N_4904,N_4299,N_4026);
nand U4905 (N_4905,N_4003,N_4425);
nor U4906 (N_4906,N_4118,N_4321);
and U4907 (N_4907,N_4359,N_4060);
nand U4908 (N_4908,N_4222,N_4402);
nand U4909 (N_4909,N_4281,N_4012);
and U4910 (N_4910,N_4170,N_4497);
and U4911 (N_4911,N_4036,N_4190);
nor U4912 (N_4912,N_4491,N_4075);
or U4913 (N_4913,N_4302,N_4356);
nor U4914 (N_4914,N_4462,N_4046);
nand U4915 (N_4915,N_4278,N_4280);
nor U4916 (N_4916,N_4486,N_4455);
nor U4917 (N_4917,N_4002,N_4378);
nor U4918 (N_4918,N_4240,N_4027);
or U4919 (N_4919,N_4051,N_4040);
nor U4920 (N_4920,N_4001,N_4245);
or U4921 (N_4921,N_4424,N_4202);
or U4922 (N_4922,N_4161,N_4210);
xnor U4923 (N_4923,N_4206,N_4466);
nor U4924 (N_4924,N_4170,N_4291);
nor U4925 (N_4925,N_4128,N_4223);
nand U4926 (N_4926,N_4289,N_4139);
and U4927 (N_4927,N_4299,N_4384);
and U4928 (N_4928,N_4476,N_4149);
nor U4929 (N_4929,N_4446,N_4017);
nand U4930 (N_4930,N_4424,N_4043);
nand U4931 (N_4931,N_4418,N_4036);
nand U4932 (N_4932,N_4413,N_4348);
and U4933 (N_4933,N_4341,N_4283);
xor U4934 (N_4934,N_4145,N_4163);
nor U4935 (N_4935,N_4114,N_4027);
nand U4936 (N_4936,N_4102,N_4427);
and U4937 (N_4937,N_4100,N_4273);
or U4938 (N_4938,N_4266,N_4116);
nor U4939 (N_4939,N_4076,N_4226);
or U4940 (N_4940,N_4441,N_4315);
nor U4941 (N_4941,N_4102,N_4037);
and U4942 (N_4942,N_4303,N_4493);
xnor U4943 (N_4943,N_4101,N_4028);
nand U4944 (N_4944,N_4091,N_4325);
nor U4945 (N_4945,N_4156,N_4475);
or U4946 (N_4946,N_4151,N_4411);
nand U4947 (N_4947,N_4334,N_4069);
xnor U4948 (N_4948,N_4070,N_4034);
nand U4949 (N_4949,N_4391,N_4300);
xor U4950 (N_4950,N_4341,N_4094);
nand U4951 (N_4951,N_4494,N_4435);
and U4952 (N_4952,N_4202,N_4144);
nand U4953 (N_4953,N_4410,N_4494);
and U4954 (N_4954,N_4335,N_4251);
or U4955 (N_4955,N_4350,N_4025);
xnor U4956 (N_4956,N_4054,N_4223);
and U4957 (N_4957,N_4071,N_4306);
or U4958 (N_4958,N_4239,N_4071);
nand U4959 (N_4959,N_4309,N_4389);
and U4960 (N_4960,N_4056,N_4376);
or U4961 (N_4961,N_4403,N_4021);
and U4962 (N_4962,N_4142,N_4341);
or U4963 (N_4963,N_4385,N_4038);
nand U4964 (N_4964,N_4359,N_4424);
nor U4965 (N_4965,N_4209,N_4435);
or U4966 (N_4966,N_4405,N_4099);
and U4967 (N_4967,N_4299,N_4438);
or U4968 (N_4968,N_4000,N_4158);
or U4969 (N_4969,N_4090,N_4063);
and U4970 (N_4970,N_4173,N_4287);
and U4971 (N_4971,N_4112,N_4163);
nor U4972 (N_4972,N_4076,N_4310);
nand U4973 (N_4973,N_4243,N_4460);
nand U4974 (N_4974,N_4045,N_4036);
nor U4975 (N_4975,N_4035,N_4237);
or U4976 (N_4976,N_4381,N_4320);
nor U4977 (N_4977,N_4004,N_4434);
nor U4978 (N_4978,N_4094,N_4464);
nor U4979 (N_4979,N_4241,N_4034);
nand U4980 (N_4980,N_4104,N_4347);
nor U4981 (N_4981,N_4392,N_4367);
nor U4982 (N_4982,N_4347,N_4427);
or U4983 (N_4983,N_4282,N_4122);
nor U4984 (N_4984,N_4048,N_4168);
or U4985 (N_4985,N_4267,N_4171);
and U4986 (N_4986,N_4311,N_4037);
nor U4987 (N_4987,N_4259,N_4288);
nand U4988 (N_4988,N_4062,N_4428);
and U4989 (N_4989,N_4367,N_4313);
and U4990 (N_4990,N_4490,N_4244);
and U4991 (N_4991,N_4390,N_4208);
and U4992 (N_4992,N_4384,N_4007);
nor U4993 (N_4993,N_4088,N_4047);
or U4994 (N_4994,N_4494,N_4014);
nor U4995 (N_4995,N_4172,N_4054);
and U4996 (N_4996,N_4256,N_4458);
nand U4997 (N_4997,N_4218,N_4132);
or U4998 (N_4998,N_4411,N_4237);
or U4999 (N_4999,N_4202,N_4198);
and UO_0 (O_0,N_4607,N_4587);
nor UO_1 (O_1,N_4955,N_4851);
nand UO_2 (O_2,N_4641,N_4591);
nor UO_3 (O_3,N_4692,N_4502);
nand UO_4 (O_4,N_4725,N_4678);
nor UO_5 (O_5,N_4662,N_4980);
nor UO_6 (O_6,N_4584,N_4648);
xnor UO_7 (O_7,N_4860,N_4884);
or UO_8 (O_8,N_4543,N_4828);
and UO_9 (O_9,N_4650,N_4913);
nor UO_10 (O_10,N_4962,N_4726);
xor UO_11 (O_11,N_4682,N_4701);
or UO_12 (O_12,N_4970,N_4529);
nand UO_13 (O_13,N_4659,N_4912);
and UO_14 (O_14,N_4891,N_4803);
nor UO_15 (O_15,N_4842,N_4723);
nand UO_16 (O_16,N_4578,N_4753);
nand UO_17 (O_17,N_4612,N_4854);
and UO_18 (O_18,N_4611,N_4558);
and UO_19 (O_19,N_4791,N_4879);
nor UO_20 (O_20,N_4592,N_4594);
nand UO_21 (O_21,N_4646,N_4972);
or UO_22 (O_22,N_4976,N_4874);
nor UO_23 (O_23,N_4640,N_4695);
and UO_24 (O_24,N_4812,N_4769);
and UO_25 (O_25,N_4570,N_4835);
nor UO_26 (O_26,N_4947,N_4602);
nor UO_27 (O_27,N_4889,N_4520);
or UO_28 (O_28,N_4523,N_4622);
nor UO_29 (O_29,N_4738,N_4559);
or UO_30 (O_30,N_4525,N_4804);
or UO_31 (O_31,N_4674,N_4939);
nor UO_32 (O_32,N_4600,N_4623);
nor UO_33 (O_33,N_4831,N_4948);
or UO_34 (O_34,N_4876,N_4554);
nor UO_35 (O_35,N_4784,N_4596);
or UO_36 (O_36,N_4586,N_4973);
or UO_37 (O_37,N_4673,N_4810);
nor UO_38 (O_38,N_4500,N_4820);
and UO_39 (O_39,N_4763,N_4661);
and UO_40 (O_40,N_4652,N_4569);
nand UO_41 (O_41,N_4895,N_4902);
and UO_42 (O_42,N_4671,N_4690);
or UO_43 (O_43,N_4909,N_4907);
nor UO_44 (O_44,N_4518,N_4667);
nand UO_45 (O_45,N_4867,N_4811);
and UO_46 (O_46,N_4880,N_4953);
or UO_47 (O_47,N_4670,N_4802);
nand UO_48 (O_48,N_4786,N_4821);
nor UO_49 (O_49,N_4762,N_4657);
nor UO_50 (O_50,N_4778,N_4750);
or UO_51 (O_51,N_4537,N_4732);
and UO_52 (O_52,N_4741,N_4615);
nor UO_53 (O_53,N_4633,N_4631);
nor UO_54 (O_54,N_4644,N_4969);
nor UO_55 (O_55,N_4524,N_4903);
nand UO_56 (O_56,N_4833,N_4509);
nor UO_57 (O_57,N_4745,N_4512);
nor UO_58 (O_58,N_4510,N_4798);
and UO_59 (O_59,N_4647,N_4736);
nor UO_60 (O_60,N_4562,N_4789);
nand UO_61 (O_61,N_4504,N_4885);
and UO_62 (O_62,N_4551,N_4838);
or UO_63 (O_63,N_4629,N_4944);
nand UO_64 (O_64,N_4931,N_4950);
nand UO_65 (O_65,N_4904,N_4681);
or UO_66 (O_66,N_4527,N_4740);
and UO_67 (O_67,N_4758,N_4914);
nand UO_68 (O_68,N_4966,N_4548);
and UO_69 (O_69,N_4850,N_4634);
and UO_70 (O_70,N_4579,N_4768);
nand UO_71 (O_71,N_4731,N_4937);
nand UO_72 (O_72,N_4691,N_4795);
nor UO_73 (O_73,N_4557,N_4935);
nand UO_74 (O_74,N_4781,N_4744);
nand UO_75 (O_75,N_4882,N_4997);
and UO_76 (O_76,N_4981,N_4721);
nor UO_77 (O_77,N_4555,N_4775);
and UO_78 (O_78,N_4624,N_4837);
and UO_79 (O_79,N_4883,N_4794);
nor UO_80 (O_80,N_4963,N_4720);
or UO_81 (O_81,N_4968,N_4601);
or UO_82 (O_82,N_4800,N_4603);
nor UO_83 (O_83,N_4893,N_4638);
nand UO_84 (O_84,N_4897,N_4971);
nor UO_85 (O_85,N_4806,N_4565);
nor UO_86 (O_86,N_4545,N_4534);
and UO_87 (O_87,N_4730,N_4958);
nor UO_88 (O_88,N_4544,N_4906);
nor UO_89 (O_89,N_4696,N_4830);
and UO_90 (O_90,N_4700,N_4877);
or UO_91 (O_91,N_4748,N_4561);
and UO_92 (O_92,N_4892,N_4776);
nor UO_93 (O_93,N_4853,N_4869);
nor UO_94 (O_94,N_4908,N_4668);
nand UO_95 (O_95,N_4552,N_4605);
or UO_96 (O_96,N_4943,N_4761);
and UO_97 (O_97,N_4777,N_4826);
nand UO_98 (O_98,N_4714,N_4549);
or UO_99 (O_99,N_4697,N_4566);
and UO_100 (O_100,N_4809,N_4577);
nor UO_101 (O_101,N_4526,N_4949);
or UO_102 (O_102,N_4653,N_4597);
or UO_103 (O_103,N_4746,N_4834);
and UO_104 (O_104,N_4711,N_4856);
nor UO_105 (O_105,N_4922,N_4737);
or UO_106 (O_106,N_4530,N_4941);
nand UO_107 (O_107,N_4986,N_4954);
or UO_108 (O_108,N_4799,N_4749);
nand UO_109 (O_109,N_4604,N_4772);
or UO_110 (O_110,N_4698,N_4735);
or UO_111 (O_111,N_4628,N_4616);
nand UO_112 (O_112,N_4642,N_4664);
nand UO_113 (O_113,N_4679,N_4663);
and UO_114 (O_114,N_4796,N_4887);
and UO_115 (O_115,N_4705,N_4766);
or UO_116 (O_116,N_4733,N_4547);
nand UO_117 (O_117,N_4627,N_4507);
or UO_118 (O_118,N_4606,N_4747);
xnor UO_119 (O_119,N_4693,N_4621);
nor UO_120 (O_120,N_4875,N_4888);
and UO_121 (O_121,N_4576,N_4996);
nor UO_122 (O_122,N_4703,N_4739);
and UO_123 (O_123,N_4654,N_4538);
and UO_124 (O_124,N_4780,N_4734);
nand UO_125 (O_125,N_4774,N_4991);
or UO_126 (O_126,N_4901,N_4580);
and UO_127 (O_127,N_4508,N_4614);
or UO_128 (O_128,N_4506,N_4709);
nand UO_129 (O_129,N_4643,N_4568);
nand UO_130 (O_130,N_4719,N_4801);
or UO_131 (O_131,N_4755,N_4896);
and UO_132 (O_132,N_4560,N_4505);
nand UO_133 (O_133,N_4932,N_4832);
or UO_134 (O_134,N_4983,N_4930);
and UO_135 (O_135,N_4940,N_4936);
nand UO_136 (O_136,N_4609,N_4511);
or UO_137 (O_137,N_4751,N_4864);
xor UO_138 (O_138,N_4994,N_4848);
nand UO_139 (O_139,N_4637,N_4998);
nor UO_140 (O_140,N_4857,N_4952);
nand UO_141 (O_141,N_4951,N_4843);
nand UO_142 (O_142,N_4919,N_4742);
and UO_143 (O_143,N_4649,N_4503);
nand UO_144 (O_144,N_4704,N_4546);
and UO_145 (O_145,N_4844,N_4722);
and UO_146 (O_146,N_4898,N_4900);
or UO_147 (O_147,N_4535,N_4757);
nor UO_148 (O_148,N_4689,N_4626);
or UO_149 (O_149,N_4686,N_4756);
nor UO_150 (O_150,N_4975,N_4598);
or UO_151 (O_151,N_4694,N_4849);
and UO_152 (O_152,N_4599,N_4839);
nor UO_153 (O_153,N_4574,N_4993);
nor UO_154 (O_154,N_4760,N_4571);
and UO_155 (O_155,N_4868,N_4590);
xor UO_156 (O_156,N_4706,N_4639);
and UO_157 (O_157,N_4808,N_4878);
and UO_158 (O_158,N_4871,N_4620);
and UO_159 (O_159,N_4564,N_4672);
nor UO_160 (O_160,N_4585,N_4788);
and UO_161 (O_161,N_4684,N_4595);
nand UO_162 (O_162,N_4528,N_4729);
and UO_163 (O_163,N_4905,N_4790);
nand UO_164 (O_164,N_4881,N_4934);
nand UO_165 (O_165,N_4517,N_4918);
nor UO_166 (O_166,N_4677,N_4645);
xnor UO_167 (O_167,N_4823,N_4836);
and UO_168 (O_168,N_4924,N_4656);
xnor UO_169 (O_169,N_4979,N_4593);
nor UO_170 (O_170,N_4818,N_4707);
nand UO_171 (O_171,N_4921,N_4974);
nand UO_172 (O_172,N_4522,N_4541);
and UO_173 (O_173,N_4859,N_4608);
or UO_174 (O_174,N_4533,N_4945);
nand UO_175 (O_175,N_4959,N_4956);
nor UO_176 (O_176,N_4999,N_4539);
and UO_177 (O_177,N_4687,N_4819);
nand UO_178 (O_178,N_4754,N_4967);
or UO_179 (O_179,N_4816,N_4925);
nor UO_180 (O_180,N_4787,N_4960);
or UO_181 (O_181,N_4770,N_4872);
and UO_182 (O_182,N_4567,N_4635);
nor UO_183 (O_183,N_4824,N_4515);
or UO_184 (O_184,N_4660,N_4521);
and UO_185 (O_185,N_4655,N_4588);
and UO_186 (O_186,N_4531,N_4792);
xnor UO_187 (O_187,N_4752,N_4702);
or UO_188 (O_188,N_4542,N_4610);
and UO_189 (O_189,N_4676,N_4782);
nand UO_190 (O_190,N_4669,N_4990);
nor UO_191 (O_191,N_4536,N_4890);
nand UO_192 (O_192,N_4814,N_4910);
or UO_193 (O_193,N_4718,N_4845);
nand UO_194 (O_194,N_4710,N_4942);
or UO_195 (O_195,N_4688,N_4516);
nor UO_196 (O_196,N_4743,N_4783);
nor UO_197 (O_197,N_4501,N_4613);
nor UO_198 (O_198,N_4625,N_4765);
nor UO_199 (O_199,N_4556,N_4861);
nor UO_200 (O_200,N_4866,N_4822);
and UO_201 (O_201,N_4727,N_4513);
xor UO_202 (O_202,N_4575,N_4840);
nand UO_203 (O_203,N_4989,N_4965);
or UO_204 (O_204,N_4573,N_4618);
or UO_205 (O_205,N_4827,N_4855);
nor UO_206 (O_206,N_4916,N_4617);
nor UO_207 (O_207,N_4886,N_4665);
and UO_208 (O_208,N_4699,N_4933);
nand UO_209 (O_209,N_4728,N_4841);
or UO_210 (O_210,N_4926,N_4563);
nand UO_211 (O_211,N_4865,N_4708);
or UO_212 (O_212,N_4817,N_4675);
nand UO_213 (O_213,N_4685,N_4977);
nand UO_214 (O_214,N_4873,N_4713);
and UO_215 (O_215,N_4961,N_4995);
nor UO_216 (O_216,N_4658,N_4987);
and UO_217 (O_217,N_4847,N_4858);
and UO_218 (O_218,N_4852,N_4813);
xnor UO_219 (O_219,N_4785,N_4797);
nand UO_220 (O_220,N_4982,N_4553);
xor UO_221 (O_221,N_4992,N_4519);
nand UO_222 (O_222,N_4724,N_4771);
nand UO_223 (O_223,N_4815,N_4805);
or UO_224 (O_224,N_4985,N_4572);
and UO_225 (O_225,N_4957,N_4915);
and UO_226 (O_226,N_4532,N_4589);
and UO_227 (O_227,N_4680,N_4759);
or UO_228 (O_228,N_4550,N_4581);
and UO_229 (O_229,N_4964,N_4863);
nand UO_230 (O_230,N_4583,N_4793);
and UO_231 (O_231,N_4946,N_4988);
or UO_232 (O_232,N_4911,N_4923);
and UO_233 (O_233,N_4764,N_4683);
or UO_234 (O_234,N_4929,N_4927);
nand UO_235 (O_235,N_4846,N_4899);
or UO_236 (O_236,N_4540,N_4807);
nand UO_237 (O_237,N_4712,N_4632);
nand UO_238 (O_238,N_4630,N_4779);
or UO_239 (O_239,N_4717,N_4984);
and UO_240 (O_240,N_4716,N_4773);
nor UO_241 (O_241,N_4894,N_4651);
nand UO_242 (O_242,N_4514,N_4825);
nand UO_243 (O_243,N_4619,N_4666);
and UO_244 (O_244,N_4715,N_4917);
nor UO_245 (O_245,N_4636,N_4862);
nor UO_246 (O_246,N_4582,N_4978);
and UO_247 (O_247,N_4938,N_4829);
nand UO_248 (O_248,N_4920,N_4767);
and UO_249 (O_249,N_4870,N_4928);
and UO_250 (O_250,N_4566,N_4526);
and UO_251 (O_251,N_4979,N_4824);
nor UO_252 (O_252,N_4571,N_4857);
nand UO_253 (O_253,N_4665,N_4951);
and UO_254 (O_254,N_4947,N_4820);
nor UO_255 (O_255,N_4550,N_4871);
xnor UO_256 (O_256,N_4758,N_4682);
nand UO_257 (O_257,N_4947,N_4816);
nand UO_258 (O_258,N_4798,N_4630);
or UO_259 (O_259,N_4951,N_4713);
nand UO_260 (O_260,N_4660,N_4921);
or UO_261 (O_261,N_4709,N_4628);
nor UO_262 (O_262,N_4925,N_4948);
or UO_263 (O_263,N_4537,N_4705);
nand UO_264 (O_264,N_4755,N_4839);
and UO_265 (O_265,N_4507,N_4905);
and UO_266 (O_266,N_4987,N_4814);
and UO_267 (O_267,N_4972,N_4853);
or UO_268 (O_268,N_4702,N_4701);
nand UO_269 (O_269,N_4780,N_4794);
or UO_270 (O_270,N_4527,N_4713);
nand UO_271 (O_271,N_4761,N_4570);
or UO_272 (O_272,N_4713,N_4798);
and UO_273 (O_273,N_4592,N_4647);
nand UO_274 (O_274,N_4933,N_4845);
or UO_275 (O_275,N_4822,N_4681);
xor UO_276 (O_276,N_4623,N_4526);
nand UO_277 (O_277,N_4563,N_4654);
and UO_278 (O_278,N_4714,N_4667);
nand UO_279 (O_279,N_4794,N_4515);
nand UO_280 (O_280,N_4719,N_4667);
or UO_281 (O_281,N_4665,N_4772);
and UO_282 (O_282,N_4848,N_4720);
nand UO_283 (O_283,N_4820,N_4894);
and UO_284 (O_284,N_4776,N_4666);
nor UO_285 (O_285,N_4735,N_4590);
nor UO_286 (O_286,N_4896,N_4537);
or UO_287 (O_287,N_4827,N_4530);
and UO_288 (O_288,N_4947,N_4624);
nand UO_289 (O_289,N_4516,N_4744);
or UO_290 (O_290,N_4525,N_4884);
nand UO_291 (O_291,N_4874,N_4692);
nand UO_292 (O_292,N_4817,N_4608);
and UO_293 (O_293,N_4969,N_4819);
or UO_294 (O_294,N_4819,N_4539);
and UO_295 (O_295,N_4709,N_4646);
nand UO_296 (O_296,N_4673,N_4681);
nand UO_297 (O_297,N_4569,N_4679);
xor UO_298 (O_298,N_4998,N_4635);
nor UO_299 (O_299,N_4887,N_4761);
and UO_300 (O_300,N_4658,N_4528);
or UO_301 (O_301,N_4768,N_4690);
nand UO_302 (O_302,N_4709,N_4536);
nand UO_303 (O_303,N_4769,N_4807);
xor UO_304 (O_304,N_4685,N_4624);
nand UO_305 (O_305,N_4527,N_4646);
and UO_306 (O_306,N_4864,N_4883);
or UO_307 (O_307,N_4674,N_4858);
or UO_308 (O_308,N_4598,N_4753);
and UO_309 (O_309,N_4662,N_4893);
xnor UO_310 (O_310,N_4971,N_4936);
and UO_311 (O_311,N_4932,N_4786);
or UO_312 (O_312,N_4762,N_4504);
and UO_313 (O_313,N_4776,N_4850);
nand UO_314 (O_314,N_4511,N_4984);
nor UO_315 (O_315,N_4772,N_4819);
and UO_316 (O_316,N_4652,N_4949);
nor UO_317 (O_317,N_4757,N_4628);
or UO_318 (O_318,N_4687,N_4694);
nand UO_319 (O_319,N_4507,N_4845);
nor UO_320 (O_320,N_4955,N_4801);
or UO_321 (O_321,N_4944,N_4746);
xor UO_322 (O_322,N_4826,N_4522);
nor UO_323 (O_323,N_4831,N_4818);
or UO_324 (O_324,N_4843,N_4984);
or UO_325 (O_325,N_4701,N_4699);
xor UO_326 (O_326,N_4617,N_4966);
and UO_327 (O_327,N_4736,N_4561);
nor UO_328 (O_328,N_4550,N_4877);
nor UO_329 (O_329,N_4957,N_4657);
nand UO_330 (O_330,N_4709,N_4606);
nand UO_331 (O_331,N_4524,N_4811);
or UO_332 (O_332,N_4992,N_4725);
or UO_333 (O_333,N_4620,N_4779);
nor UO_334 (O_334,N_4507,N_4919);
nand UO_335 (O_335,N_4974,N_4600);
nand UO_336 (O_336,N_4568,N_4585);
or UO_337 (O_337,N_4834,N_4813);
or UO_338 (O_338,N_4774,N_4876);
and UO_339 (O_339,N_4641,N_4556);
nand UO_340 (O_340,N_4811,N_4827);
nand UO_341 (O_341,N_4586,N_4648);
xnor UO_342 (O_342,N_4568,N_4939);
and UO_343 (O_343,N_4856,N_4789);
nand UO_344 (O_344,N_4738,N_4995);
nor UO_345 (O_345,N_4514,N_4838);
nand UO_346 (O_346,N_4601,N_4829);
or UO_347 (O_347,N_4937,N_4630);
or UO_348 (O_348,N_4751,N_4898);
and UO_349 (O_349,N_4823,N_4966);
nor UO_350 (O_350,N_4595,N_4970);
nor UO_351 (O_351,N_4597,N_4580);
nand UO_352 (O_352,N_4522,N_4639);
and UO_353 (O_353,N_4894,N_4728);
nand UO_354 (O_354,N_4869,N_4803);
and UO_355 (O_355,N_4603,N_4929);
or UO_356 (O_356,N_4907,N_4798);
or UO_357 (O_357,N_4730,N_4799);
xor UO_358 (O_358,N_4946,N_4612);
nor UO_359 (O_359,N_4937,N_4844);
nor UO_360 (O_360,N_4715,N_4963);
and UO_361 (O_361,N_4501,N_4917);
and UO_362 (O_362,N_4854,N_4666);
and UO_363 (O_363,N_4778,N_4672);
and UO_364 (O_364,N_4899,N_4964);
or UO_365 (O_365,N_4923,N_4641);
nor UO_366 (O_366,N_4696,N_4575);
nor UO_367 (O_367,N_4991,N_4542);
or UO_368 (O_368,N_4547,N_4707);
and UO_369 (O_369,N_4672,N_4675);
xnor UO_370 (O_370,N_4671,N_4541);
xnor UO_371 (O_371,N_4888,N_4953);
nand UO_372 (O_372,N_4521,N_4766);
nand UO_373 (O_373,N_4948,N_4507);
and UO_374 (O_374,N_4799,N_4664);
and UO_375 (O_375,N_4625,N_4939);
xor UO_376 (O_376,N_4742,N_4752);
or UO_377 (O_377,N_4827,N_4879);
and UO_378 (O_378,N_4547,N_4873);
nand UO_379 (O_379,N_4544,N_4521);
or UO_380 (O_380,N_4821,N_4992);
or UO_381 (O_381,N_4828,N_4957);
or UO_382 (O_382,N_4618,N_4543);
nand UO_383 (O_383,N_4819,N_4868);
and UO_384 (O_384,N_4816,N_4524);
or UO_385 (O_385,N_4682,N_4634);
and UO_386 (O_386,N_4695,N_4592);
nor UO_387 (O_387,N_4594,N_4865);
nor UO_388 (O_388,N_4718,N_4628);
xor UO_389 (O_389,N_4654,N_4921);
nand UO_390 (O_390,N_4640,N_4560);
xor UO_391 (O_391,N_4547,N_4569);
nand UO_392 (O_392,N_4994,N_4619);
nand UO_393 (O_393,N_4538,N_4655);
or UO_394 (O_394,N_4610,N_4695);
nand UO_395 (O_395,N_4534,N_4558);
or UO_396 (O_396,N_4811,N_4673);
xor UO_397 (O_397,N_4820,N_4773);
nand UO_398 (O_398,N_4583,N_4670);
nor UO_399 (O_399,N_4749,N_4741);
nand UO_400 (O_400,N_4604,N_4941);
and UO_401 (O_401,N_4607,N_4706);
xor UO_402 (O_402,N_4725,N_4600);
xnor UO_403 (O_403,N_4902,N_4710);
nand UO_404 (O_404,N_4626,N_4633);
or UO_405 (O_405,N_4970,N_4513);
and UO_406 (O_406,N_4851,N_4623);
nand UO_407 (O_407,N_4661,N_4879);
xnor UO_408 (O_408,N_4794,N_4874);
or UO_409 (O_409,N_4786,N_4889);
nor UO_410 (O_410,N_4528,N_4801);
and UO_411 (O_411,N_4808,N_4748);
nand UO_412 (O_412,N_4557,N_4764);
xnor UO_413 (O_413,N_4885,N_4852);
nand UO_414 (O_414,N_4935,N_4840);
and UO_415 (O_415,N_4789,N_4555);
or UO_416 (O_416,N_4887,N_4999);
and UO_417 (O_417,N_4512,N_4709);
or UO_418 (O_418,N_4937,N_4995);
or UO_419 (O_419,N_4725,N_4988);
nor UO_420 (O_420,N_4710,N_4682);
xor UO_421 (O_421,N_4708,N_4717);
or UO_422 (O_422,N_4845,N_4833);
and UO_423 (O_423,N_4584,N_4757);
or UO_424 (O_424,N_4812,N_4868);
xnor UO_425 (O_425,N_4725,N_4656);
nand UO_426 (O_426,N_4734,N_4641);
nor UO_427 (O_427,N_4552,N_4507);
nand UO_428 (O_428,N_4600,N_4873);
nor UO_429 (O_429,N_4593,N_4850);
and UO_430 (O_430,N_4701,N_4921);
and UO_431 (O_431,N_4944,N_4770);
or UO_432 (O_432,N_4870,N_4680);
nand UO_433 (O_433,N_4589,N_4565);
and UO_434 (O_434,N_4644,N_4666);
nand UO_435 (O_435,N_4730,N_4966);
nand UO_436 (O_436,N_4504,N_4694);
nand UO_437 (O_437,N_4899,N_4588);
nor UO_438 (O_438,N_4555,N_4605);
xor UO_439 (O_439,N_4510,N_4533);
nand UO_440 (O_440,N_4950,N_4514);
xor UO_441 (O_441,N_4659,N_4681);
nor UO_442 (O_442,N_4707,N_4819);
xnor UO_443 (O_443,N_4745,N_4958);
xor UO_444 (O_444,N_4678,N_4772);
nor UO_445 (O_445,N_4684,N_4752);
nand UO_446 (O_446,N_4910,N_4903);
or UO_447 (O_447,N_4569,N_4772);
nand UO_448 (O_448,N_4642,N_4867);
and UO_449 (O_449,N_4574,N_4567);
or UO_450 (O_450,N_4653,N_4997);
and UO_451 (O_451,N_4620,N_4903);
nand UO_452 (O_452,N_4702,N_4686);
nand UO_453 (O_453,N_4538,N_4556);
or UO_454 (O_454,N_4603,N_4921);
nand UO_455 (O_455,N_4644,N_4865);
and UO_456 (O_456,N_4967,N_4811);
xnor UO_457 (O_457,N_4954,N_4877);
and UO_458 (O_458,N_4706,N_4728);
nor UO_459 (O_459,N_4829,N_4503);
nor UO_460 (O_460,N_4659,N_4515);
xor UO_461 (O_461,N_4945,N_4794);
nand UO_462 (O_462,N_4734,N_4825);
or UO_463 (O_463,N_4949,N_4968);
nor UO_464 (O_464,N_4520,N_4711);
nor UO_465 (O_465,N_4790,N_4965);
nor UO_466 (O_466,N_4783,N_4821);
nand UO_467 (O_467,N_4963,N_4880);
xor UO_468 (O_468,N_4943,N_4869);
and UO_469 (O_469,N_4597,N_4983);
and UO_470 (O_470,N_4767,N_4593);
nand UO_471 (O_471,N_4565,N_4845);
nor UO_472 (O_472,N_4881,N_4595);
and UO_473 (O_473,N_4668,N_4856);
xnor UO_474 (O_474,N_4622,N_4842);
nand UO_475 (O_475,N_4647,N_4955);
or UO_476 (O_476,N_4793,N_4977);
nor UO_477 (O_477,N_4735,N_4522);
nand UO_478 (O_478,N_4590,N_4944);
xor UO_479 (O_479,N_4779,N_4532);
xnor UO_480 (O_480,N_4777,N_4859);
and UO_481 (O_481,N_4899,N_4993);
or UO_482 (O_482,N_4723,N_4638);
and UO_483 (O_483,N_4865,N_4608);
and UO_484 (O_484,N_4953,N_4759);
and UO_485 (O_485,N_4696,N_4545);
nand UO_486 (O_486,N_4918,N_4981);
xor UO_487 (O_487,N_4503,N_4736);
and UO_488 (O_488,N_4874,N_4576);
or UO_489 (O_489,N_4853,N_4639);
or UO_490 (O_490,N_4954,N_4876);
and UO_491 (O_491,N_4531,N_4808);
nor UO_492 (O_492,N_4771,N_4855);
xor UO_493 (O_493,N_4916,N_4607);
or UO_494 (O_494,N_4909,N_4866);
and UO_495 (O_495,N_4569,N_4692);
nor UO_496 (O_496,N_4502,N_4750);
nor UO_497 (O_497,N_4836,N_4955);
or UO_498 (O_498,N_4874,N_4606);
nor UO_499 (O_499,N_4644,N_4935);
nand UO_500 (O_500,N_4528,N_4526);
nand UO_501 (O_501,N_4557,N_4531);
and UO_502 (O_502,N_4568,N_4686);
or UO_503 (O_503,N_4941,N_4646);
xnor UO_504 (O_504,N_4815,N_4922);
or UO_505 (O_505,N_4822,N_4873);
nand UO_506 (O_506,N_4835,N_4899);
nand UO_507 (O_507,N_4774,N_4890);
and UO_508 (O_508,N_4841,N_4685);
nor UO_509 (O_509,N_4683,N_4969);
and UO_510 (O_510,N_4780,N_4634);
and UO_511 (O_511,N_4553,N_4742);
or UO_512 (O_512,N_4962,N_4634);
nand UO_513 (O_513,N_4575,N_4614);
or UO_514 (O_514,N_4519,N_4545);
nor UO_515 (O_515,N_4861,N_4597);
or UO_516 (O_516,N_4851,N_4942);
nand UO_517 (O_517,N_4937,N_4607);
xor UO_518 (O_518,N_4931,N_4648);
xor UO_519 (O_519,N_4722,N_4850);
nor UO_520 (O_520,N_4553,N_4513);
xnor UO_521 (O_521,N_4771,N_4895);
xnor UO_522 (O_522,N_4989,N_4948);
nand UO_523 (O_523,N_4751,N_4736);
xnor UO_524 (O_524,N_4771,N_4870);
or UO_525 (O_525,N_4549,N_4631);
or UO_526 (O_526,N_4613,N_4776);
or UO_527 (O_527,N_4513,N_4902);
or UO_528 (O_528,N_4630,N_4994);
nor UO_529 (O_529,N_4861,N_4969);
or UO_530 (O_530,N_4523,N_4890);
and UO_531 (O_531,N_4652,N_4782);
nand UO_532 (O_532,N_4596,N_4666);
or UO_533 (O_533,N_4958,N_4924);
nor UO_534 (O_534,N_4913,N_4756);
or UO_535 (O_535,N_4931,N_4658);
and UO_536 (O_536,N_4971,N_4756);
and UO_537 (O_537,N_4646,N_4626);
and UO_538 (O_538,N_4677,N_4675);
xor UO_539 (O_539,N_4873,N_4580);
nor UO_540 (O_540,N_4811,N_4966);
or UO_541 (O_541,N_4915,N_4862);
nand UO_542 (O_542,N_4706,N_4545);
and UO_543 (O_543,N_4949,N_4820);
nand UO_544 (O_544,N_4579,N_4731);
nor UO_545 (O_545,N_4626,N_4844);
nor UO_546 (O_546,N_4717,N_4519);
or UO_547 (O_547,N_4643,N_4775);
and UO_548 (O_548,N_4516,N_4842);
xor UO_549 (O_549,N_4649,N_4816);
or UO_550 (O_550,N_4521,N_4819);
or UO_551 (O_551,N_4821,N_4955);
or UO_552 (O_552,N_4752,N_4647);
nand UO_553 (O_553,N_4921,N_4764);
nor UO_554 (O_554,N_4612,N_4593);
xnor UO_555 (O_555,N_4867,N_4511);
or UO_556 (O_556,N_4573,N_4617);
and UO_557 (O_557,N_4509,N_4692);
and UO_558 (O_558,N_4773,N_4863);
and UO_559 (O_559,N_4984,N_4510);
nor UO_560 (O_560,N_4815,N_4655);
nor UO_561 (O_561,N_4882,N_4731);
nand UO_562 (O_562,N_4843,N_4639);
nor UO_563 (O_563,N_4859,N_4872);
and UO_564 (O_564,N_4596,N_4505);
nand UO_565 (O_565,N_4714,N_4605);
or UO_566 (O_566,N_4682,N_4640);
xnor UO_567 (O_567,N_4592,N_4994);
nand UO_568 (O_568,N_4589,N_4677);
nor UO_569 (O_569,N_4915,N_4821);
nor UO_570 (O_570,N_4651,N_4647);
nand UO_571 (O_571,N_4592,N_4645);
or UO_572 (O_572,N_4513,N_4893);
xor UO_573 (O_573,N_4514,N_4739);
and UO_574 (O_574,N_4602,N_4684);
and UO_575 (O_575,N_4625,N_4592);
nor UO_576 (O_576,N_4631,N_4552);
and UO_577 (O_577,N_4819,N_4660);
and UO_578 (O_578,N_4709,N_4568);
or UO_579 (O_579,N_4709,N_4885);
or UO_580 (O_580,N_4878,N_4510);
nor UO_581 (O_581,N_4538,N_4815);
nand UO_582 (O_582,N_4774,N_4547);
and UO_583 (O_583,N_4538,N_4553);
nor UO_584 (O_584,N_4989,N_4870);
nand UO_585 (O_585,N_4933,N_4510);
nand UO_586 (O_586,N_4503,N_4885);
and UO_587 (O_587,N_4949,N_4839);
nand UO_588 (O_588,N_4875,N_4514);
xnor UO_589 (O_589,N_4644,N_4955);
and UO_590 (O_590,N_4779,N_4819);
or UO_591 (O_591,N_4828,N_4670);
nand UO_592 (O_592,N_4633,N_4539);
or UO_593 (O_593,N_4854,N_4641);
nor UO_594 (O_594,N_4753,N_4687);
nor UO_595 (O_595,N_4835,N_4987);
nor UO_596 (O_596,N_4743,N_4841);
and UO_597 (O_597,N_4521,N_4902);
or UO_598 (O_598,N_4625,N_4578);
nand UO_599 (O_599,N_4845,N_4731);
nand UO_600 (O_600,N_4922,N_4659);
nand UO_601 (O_601,N_4910,N_4630);
xor UO_602 (O_602,N_4971,N_4828);
nor UO_603 (O_603,N_4676,N_4958);
or UO_604 (O_604,N_4943,N_4828);
nand UO_605 (O_605,N_4516,N_4733);
or UO_606 (O_606,N_4533,N_4631);
nor UO_607 (O_607,N_4573,N_4994);
or UO_608 (O_608,N_4948,N_4915);
and UO_609 (O_609,N_4969,N_4597);
and UO_610 (O_610,N_4639,N_4928);
nor UO_611 (O_611,N_4604,N_4576);
or UO_612 (O_612,N_4785,N_4948);
or UO_613 (O_613,N_4511,N_4910);
or UO_614 (O_614,N_4911,N_4687);
nand UO_615 (O_615,N_4885,N_4871);
xor UO_616 (O_616,N_4918,N_4899);
xnor UO_617 (O_617,N_4785,N_4665);
nor UO_618 (O_618,N_4652,N_4506);
nor UO_619 (O_619,N_4899,N_4661);
xor UO_620 (O_620,N_4909,N_4791);
xor UO_621 (O_621,N_4958,N_4686);
xor UO_622 (O_622,N_4846,N_4831);
and UO_623 (O_623,N_4707,N_4532);
and UO_624 (O_624,N_4522,N_4872);
nor UO_625 (O_625,N_4536,N_4981);
nor UO_626 (O_626,N_4620,N_4984);
nor UO_627 (O_627,N_4688,N_4784);
and UO_628 (O_628,N_4709,N_4951);
nand UO_629 (O_629,N_4643,N_4707);
nand UO_630 (O_630,N_4524,N_4924);
and UO_631 (O_631,N_4500,N_4907);
xor UO_632 (O_632,N_4727,N_4716);
or UO_633 (O_633,N_4968,N_4621);
or UO_634 (O_634,N_4993,N_4926);
nand UO_635 (O_635,N_4649,N_4625);
nand UO_636 (O_636,N_4736,N_4724);
xnor UO_637 (O_637,N_4989,N_4835);
and UO_638 (O_638,N_4515,N_4954);
nand UO_639 (O_639,N_4615,N_4538);
xor UO_640 (O_640,N_4892,N_4829);
nand UO_641 (O_641,N_4518,N_4745);
nor UO_642 (O_642,N_4509,N_4845);
nand UO_643 (O_643,N_4608,N_4535);
and UO_644 (O_644,N_4535,N_4761);
nand UO_645 (O_645,N_4572,N_4920);
nor UO_646 (O_646,N_4754,N_4713);
nor UO_647 (O_647,N_4831,N_4508);
and UO_648 (O_648,N_4819,N_4810);
and UO_649 (O_649,N_4939,N_4599);
or UO_650 (O_650,N_4926,N_4923);
and UO_651 (O_651,N_4933,N_4772);
and UO_652 (O_652,N_4863,N_4708);
nor UO_653 (O_653,N_4794,N_4720);
and UO_654 (O_654,N_4742,N_4687);
nand UO_655 (O_655,N_4587,N_4848);
nor UO_656 (O_656,N_4788,N_4759);
and UO_657 (O_657,N_4928,N_4692);
nand UO_658 (O_658,N_4982,N_4549);
or UO_659 (O_659,N_4760,N_4917);
and UO_660 (O_660,N_4689,N_4870);
xnor UO_661 (O_661,N_4879,N_4695);
xor UO_662 (O_662,N_4846,N_4756);
or UO_663 (O_663,N_4523,N_4512);
or UO_664 (O_664,N_4635,N_4738);
nor UO_665 (O_665,N_4738,N_4579);
or UO_666 (O_666,N_4549,N_4869);
xor UO_667 (O_667,N_4947,N_4560);
xnor UO_668 (O_668,N_4555,N_4858);
or UO_669 (O_669,N_4614,N_4649);
and UO_670 (O_670,N_4868,N_4976);
xnor UO_671 (O_671,N_4754,N_4987);
and UO_672 (O_672,N_4963,N_4713);
xor UO_673 (O_673,N_4652,N_4651);
xor UO_674 (O_674,N_4785,N_4853);
and UO_675 (O_675,N_4811,N_4648);
or UO_676 (O_676,N_4935,N_4526);
nor UO_677 (O_677,N_4658,N_4950);
or UO_678 (O_678,N_4620,N_4891);
and UO_679 (O_679,N_4757,N_4967);
nand UO_680 (O_680,N_4591,N_4931);
or UO_681 (O_681,N_4766,N_4780);
and UO_682 (O_682,N_4522,N_4772);
nand UO_683 (O_683,N_4765,N_4855);
nand UO_684 (O_684,N_4881,N_4726);
nand UO_685 (O_685,N_4966,N_4775);
xor UO_686 (O_686,N_4819,N_4704);
nor UO_687 (O_687,N_4934,N_4820);
and UO_688 (O_688,N_4627,N_4570);
nor UO_689 (O_689,N_4966,N_4843);
nand UO_690 (O_690,N_4637,N_4661);
and UO_691 (O_691,N_4804,N_4594);
or UO_692 (O_692,N_4686,N_4874);
nor UO_693 (O_693,N_4921,N_4536);
nor UO_694 (O_694,N_4708,N_4778);
nor UO_695 (O_695,N_4590,N_4759);
nand UO_696 (O_696,N_4510,N_4731);
nor UO_697 (O_697,N_4865,N_4998);
or UO_698 (O_698,N_4627,N_4775);
or UO_699 (O_699,N_4784,N_4685);
and UO_700 (O_700,N_4677,N_4718);
nor UO_701 (O_701,N_4566,N_4807);
xnor UO_702 (O_702,N_4786,N_4654);
nand UO_703 (O_703,N_4891,N_4556);
nor UO_704 (O_704,N_4517,N_4740);
xor UO_705 (O_705,N_4560,N_4681);
and UO_706 (O_706,N_4860,N_4618);
xor UO_707 (O_707,N_4714,N_4785);
nand UO_708 (O_708,N_4739,N_4590);
and UO_709 (O_709,N_4504,N_4828);
nor UO_710 (O_710,N_4580,N_4727);
nor UO_711 (O_711,N_4819,N_4813);
nand UO_712 (O_712,N_4545,N_4828);
nor UO_713 (O_713,N_4616,N_4567);
or UO_714 (O_714,N_4564,N_4616);
xor UO_715 (O_715,N_4785,N_4968);
nor UO_716 (O_716,N_4562,N_4935);
and UO_717 (O_717,N_4749,N_4586);
nor UO_718 (O_718,N_4978,N_4608);
and UO_719 (O_719,N_4524,N_4933);
nand UO_720 (O_720,N_4975,N_4970);
and UO_721 (O_721,N_4583,N_4741);
nand UO_722 (O_722,N_4841,N_4688);
xor UO_723 (O_723,N_4702,N_4602);
xor UO_724 (O_724,N_4914,N_4728);
nor UO_725 (O_725,N_4574,N_4720);
or UO_726 (O_726,N_4973,N_4563);
xor UO_727 (O_727,N_4578,N_4778);
nor UO_728 (O_728,N_4749,N_4903);
or UO_729 (O_729,N_4690,N_4691);
nand UO_730 (O_730,N_4659,N_4899);
nand UO_731 (O_731,N_4889,N_4948);
xnor UO_732 (O_732,N_4901,N_4519);
nand UO_733 (O_733,N_4931,N_4763);
xor UO_734 (O_734,N_4948,N_4861);
nand UO_735 (O_735,N_4818,N_4734);
or UO_736 (O_736,N_4598,N_4947);
and UO_737 (O_737,N_4961,N_4868);
and UO_738 (O_738,N_4898,N_4881);
nor UO_739 (O_739,N_4562,N_4503);
or UO_740 (O_740,N_4592,N_4895);
nand UO_741 (O_741,N_4686,N_4993);
nand UO_742 (O_742,N_4667,N_4552);
and UO_743 (O_743,N_4708,N_4775);
or UO_744 (O_744,N_4904,N_4825);
or UO_745 (O_745,N_4883,N_4778);
and UO_746 (O_746,N_4762,N_4816);
nand UO_747 (O_747,N_4896,N_4549);
nor UO_748 (O_748,N_4967,N_4924);
nand UO_749 (O_749,N_4640,N_4768);
or UO_750 (O_750,N_4531,N_4784);
nor UO_751 (O_751,N_4642,N_4893);
and UO_752 (O_752,N_4643,N_4617);
nand UO_753 (O_753,N_4623,N_4751);
nand UO_754 (O_754,N_4964,N_4898);
or UO_755 (O_755,N_4977,N_4864);
and UO_756 (O_756,N_4847,N_4542);
nand UO_757 (O_757,N_4561,N_4622);
and UO_758 (O_758,N_4832,N_4870);
and UO_759 (O_759,N_4871,N_4648);
or UO_760 (O_760,N_4787,N_4648);
and UO_761 (O_761,N_4583,N_4517);
or UO_762 (O_762,N_4530,N_4899);
nor UO_763 (O_763,N_4647,N_4948);
nand UO_764 (O_764,N_4632,N_4627);
nor UO_765 (O_765,N_4509,N_4670);
nand UO_766 (O_766,N_4821,N_4591);
or UO_767 (O_767,N_4577,N_4597);
nand UO_768 (O_768,N_4893,N_4835);
nor UO_769 (O_769,N_4502,N_4677);
and UO_770 (O_770,N_4822,N_4511);
and UO_771 (O_771,N_4942,N_4707);
nor UO_772 (O_772,N_4538,N_4676);
nor UO_773 (O_773,N_4811,N_4952);
nand UO_774 (O_774,N_4738,N_4602);
nand UO_775 (O_775,N_4559,N_4976);
or UO_776 (O_776,N_4981,N_4895);
nand UO_777 (O_777,N_4560,N_4729);
nand UO_778 (O_778,N_4717,N_4638);
or UO_779 (O_779,N_4683,N_4991);
or UO_780 (O_780,N_4576,N_4896);
nor UO_781 (O_781,N_4690,N_4589);
xor UO_782 (O_782,N_4857,N_4909);
and UO_783 (O_783,N_4719,N_4752);
and UO_784 (O_784,N_4751,N_4717);
nor UO_785 (O_785,N_4627,N_4689);
nand UO_786 (O_786,N_4594,N_4668);
nand UO_787 (O_787,N_4693,N_4903);
nor UO_788 (O_788,N_4793,N_4633);
and UO_789 (O_789,N_4679,N_4868);
nor UO_790 (O_790,N_4622,N_4611);
and UO_791 (O_791,N_4796,N_4805);
nand UO_792 (O_792,N_4800,N_4850);
or UO_793 (O_793,N_4812,N_4502);
nor UO_794 (O_794,N_4685,N_4753);
and UO_795 (O_795,N_4852,N_4986);
xnor UO_796 (O_796,N_4706,N_4669);
nor UO_797 (O_797,N_4986,N_4864);
or UO_798 (O_798,N_4721,N_4685);
nand UO_799 (O_799,N_4885,N_4679);
and UO_800 (O_800,N_4524,N_4870);
or UO_801 (O_801,N_4703,N_4871);
and UO_802 (O_802,N_4660,N_4833);
and UO_803 (O_803,N_4669,N_4547);
or UO_804 (O_804,N_4676,N_4716);
nand UO_805 (O_805,N_4778,N_4853);
nor UO_806 (O_806,N_4820,N_4841);
nor UO_807 (O_807,N_4806,N_4967);
and UO_808 (O_808,N_4633,N_4813);
or UO_809 (O_809,N_4875,N_4615);
or UO_810 (O_810,N_4646,N_4618);
nor UO_811 (O_811,N_4520,N_4535);
xor UO_812 (O_812,N_4854,N_4662);
xor UO_813 (O_813,N_4561,N_4870);
and UO_814 (O_814,N_4697,N_4832);
and UO_815 (O_815,N_4814,N_4935);
nor UO_816 (O_816,N_4882,N_4857);
or UO_817 (O_817,N_4966,N_4551);
nor UO_818 (O_818,N_4702,N_4817);
xnor UO_819 (O_819,N_4602,N_4509);
nand UO_820 (O_820,N_4884,N_4811);
or UO_821 (O_821,N_4926,N_4610);
and UO_822 (O_822,N_4557,N_4822);
and UO_823 (O_823,N_4640,N_4508);
or UO_824 (O_824,N_4508,N_4950);
nor UO_825 (O_825,N_4562,N_4724);
or UO_826 (O_826,N_4688,N_4584);
nand UO_827 (O_827,N_4872,N_4676);
and UO_828 (O_828,N_4604,N_4558);
xnor UO_829 (O_829,N_4990,N_4832);
nor UO_830 (O_830,N_4787,N_4541);
or UO_831 (O_831,N_4657,N_4950);
nand UO_832 (O_832,N_4793,N_4993);
nand UO_833 (O_833,N_4931,N_4770);
or UO_834 (O_834,N_4538,N_4502);
and UO_835 (O_835,N_4791,N_4651);
nand UO_836 (O_836,N_4634,N_4590);
nor UO_837 (O_837,N_4500,N_4610);
nor UO_838 (O_838,N_4568,N_4586);
xnor UO_839 (O_839,N_4905,N_4587);
and UO_840 (O_840,N_4573,N_4953);
and UO_841 (O_841,N_4773,N_4894);
nor UO_842 (O_842,N_4695,N_4722);
nand UO_843 (O_843,N_4611,N_4707);
or UO_844 (O_844,N_4825,N_4596);
nand UO_845 (O_845,N_4923,N_4906);
or UO_846 (O_846,N_4558,N_4768);
or UO_847 (O_847,N_4666,N_4807);
nand UO_848 (O_848,N_4858,N_4532);
nand UO_849 (O_849,N_4864,N_4506);
and UO_850 (O_850,N_4871,N_4812);
xnor UO_851 (O_851,N_4941,N_4700);
or UO_852 (O_852,N_4672,N_4513);
nor UO_853 (O_853,N_4865,N_4899);
xor UO_854 (O_854,N_4956,N_4749);
nand UO_855 (O_855,N_4881,N_4812);
nand UO_856 (O_856,N_4601,N_4970);
nand UO_857 (O_857,N_4903,N_4606);
xor UO_858 (O_858,N_4591,N_4592);
or UO_859 (O_859,N_4762,N_4785);
nand UO_860 (O_860,N_4782,N_4889);
nor UO_861 (O_861,N_4712,N_4734);
nand UO_862 (O_862,N_4680,N_4622);
or UO_863 (O_863,N_4803,N_4737);
nor UO_864 (O_864,N_4861,N_4889);
nor UO_865 (O_865,N_4829,N_4995);
and UO_866 (O_866,N_4764,N_4752);
nand UO_867 (O_867,N_4679,N_4634);
xnor UO_868 (O_868,N_4633,N_4745);
and UO_869 (O_869,N_4663,N_4810);
or UO_870 (O_870,N_4830,N_4755);
nand UO_871 (O_871,N_4842,N_4600);
nor UO_872 (O_872,N_4947,N_4650);
nand UO_873 (O_873,N_4669,N_4716);
and UO_874 (O_874,N_4867,N_4876);
nand UO_875 (O_875,N_4651,N_4629);
nand UO_876 (O_876,N_4506,N_4936);
xnor UO_877 (O_877,N_4777,N_4603);
nor UO_878 (O_878,N_4530,N_4888);
nand UO_879 (O_879,N_4830,N_4961);
and UO_880 (O_880,N_4759,N_4520);
and UO_881 (O_881,N_4990,N_4603);
and UO_882 (O_882,N_4729,N_4566);
nand UO_883 (O_883,N_4910,N_4663);
or UO_884 (O_884,N_4527,N_4884);
and UO_885 (O_885,N_4990,N_4907);
and UO_886 (O_886,N_4959,N_4523);
or UO_887 (O_887,N_4830,N_4728);
nor UO_888 (O_888,N_4901,N_4637);
nor UO_889 (O_889,N_4516,N_4545);
and UO_890 (O_890,N_4807,N_4943);
or UO_891 (O_891,N_4562,N_4510);
nand UO_892 (O_892,N_4725,N_4518);
nand UO_893 (O_893,N_4710,N_4925);
or UO_894 (O_894,N_4641,N_4547);
and UO_895 (O_895,N_4874,N_4634);
nand UO_896 (O_896,N_4920,N_4907);
or UO_897 (O_897,N_4550,N_4583);
and UO_898 (O_898,N_4738,N_4778);
nand UO_899 (O_899,N_4727,N_4625);
nor UO_900 (O_900,N_4779,N_4650);
nor UO_901 (O_901,N_4960,N_4888);
and UO_902 (O_902,N_4597,N_4816);
or UO_903 (O_903,N_4708,N_4813);
nand UO_904 (O_904,N_4866,N_4948);
xnor UO_905 (O_905,N_4864,N_4828);
nand UO_906 (O_906,N_4717,N_4526);
and UO_907 (O_907,N_4600,N_4990);
and UO_908 (O_908,N_4706,N_4585);
xnor UO_909 (O_909,N_4941,N_4918);
xnor UO_910 (O_910,N_4980,N_4603);
nor UO_911 (O_911,N_4532,N_4754);
xor UO_912 (O_912,N_4674,N_4848);
nor UO_913 (O_913,N_4983,N_4871);
and UO_914 (O_914,N_4613,N_4515);
or UO_915 (O_915,N_4625,N_4679);
xor UO_916 (O_916,N_4850,N_4654);
and UO_917 (O_917,N_4760,N_4825);
nor UO_918 (O_918,N_4583,N_4904);
and UO_919 (O_919,N_4640,N_4903);
nand UO_920 (O_920,N_4952,N_4704);
or UO_921 (O_921,N_4992,N_4887);
xor UO_922 (O_922,N_4706,N_4533);
nor UO_923 (O_923,N_4555,N_4704);
xnor UO_924 (O_924,N_4828,N_4771);
and UO_925 (O_925,N_4931,N_4978);
nand UO_926 (O_926,N_4913,N_4618);
nor UO_927 (O_927,N_4793,N_4567);
nor UO_928 (O_928,N_4967,N_4560);
and UO_929 (O_929,N_4932,N_4908);
nand UO_930 (O_930,N_4504,N_4733);
nand UO_931 (O_931,N_4689,N_4820);
nand UO_932 (O_932,N_4813,N_4963);
and UO_933 (O_933,N_4913,N_4958);
and UO_934 (O_934,N_4590,N_4609);
nand UO_935 (O_935,N_4816,N_4848);
or UO_936 (O_936,N_4584,N_4645);
or UO_937 (O_937,N_4729,N_4888);
nor UO_938 (O_938,N_4606,N_4654);
nand UO_939 (O_939,N_4806,N_4534);
xnor UO_940 (O_940,N_4956,N_4538);
and UO_941 (O_941,N_4884,N_4990);
nor UO_942 (O_942,N_4615,N_4568);
nor UO_943 (O_943,N_4665,N_4807);
xnor UO_944 (O_944,N_4987,N_4747);
and UO_945 (O_945,N_4707,N_4647);
nor UO_946 (O_946,N_4551,N_4533);
nand UO_947 (O_947,N_4998,N_4913);
nor UO_948 (O_948,N_4823,N_4783);
nand UO_949 (O_949,N_4671,N_4775);
or UO_950 (O_950,N_4886,N_4920);
or UO_951 (O_951,N_4959,N_4563);
or UO_952 (O_952,N_4997,N_4664);
nand UO_953 (O_953,N_4935,N_4839);
xnor UO_954 (O_954,N_4678,N_4544);
or UO_955 (O_955,N_4593,N_4566);
or UO_956 (O_956,N_4854,N_4593);
nor UO_957 (O_957,N_4595,N_4559);
and UO_958 (O_958,N_4779,N_4550);
nand UO_959 (O_959,N_4973,N_4630);
and UO_960 (O_960,N_4717,N_4929);
or UO_961 (O_961,N_4520,N_4522);
nor UO_962 (O_962,N_4620,N_4625);
and UO_963 (O_963,N_4685,N_4567);
or UO_964 (O_964,N_4973,N_4891);
and UO_965 (O_965,N_4712,N_4762);
nor UO_966 (O_966,N_4710,N_4708);
or UO_967 (O_967,N_4947,N_4710);
and UO_968 (O_968,N_4591,N_4827);
nand UO_969 (O_969,N_4896,N_4810);
or UO_970 (O_970,N_4755,N_4597);
and UO_971 (O_971,N_4529,N_4857);
and UO_972 (O_972,N_4671,N_4621);
or UO_973 (O_973,N_4947,N_4866);
nand UO_974 (O_974,N_4833,N_4873);
and UO_975 (O_975,N_4897,N_4718);
nand UO_976 (O_976,N_4504,N_4674);
and UO_977 (O_977,N_4849,N_4961);
and UO_978 (O_978,N_4778,N_4861);
nor UO_979 (O_979,N_4832,N_4534);
nand UO_980 (O_980,N_4916,N_4806);
and UO_981 (O_981,N_4755,N_4835);
and UO_982 (O_982,N_4577,N_4887);
nor UO_983 (O_983,N_4552,N_4633);
or UO_984 (O_984,N_4749,N_4999);
xor UO_985 (O_985,N_4581,N_4969);
nor UO_986 (O_986,N_4847,N_4885);
xor UO_987 (O_987,N_4544,N_4848);
and UO_988 (O_988,N_4812,N_4623);
or UO_989 (O_989,N_4936,N_4518);
and UO_990 (O_990,N_4898,N_4610);
and UO_991 (O_991,N_4811,N_4681);
nand UO_992 (O_992,N_4999,N_4885);
or UO_993 (O_993,N_4692,N_4879);
nand UO_994 (O_994,N_4866,N_4845);
nor UO_995 (O_995,N_4542,N_4570);
xnor UO_996 (O_996,N_4878,N_4642);
or UO_997 (O_997,N_4791,N_4579);
nand UO_998 (O_998,N_4796,N_4579);
nand UO_999 (O_999,N_4930,N_4797);
endmodule