module basic_500_3000_500_60_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_425,In_172);
nand U1 (N_1,In_493,In_161);
and U2 (N_2,In_96,In_317);
nand U3 (N_3,In_227,In_176);
and U4 (N_4,In_271,In_0);
nor U5 (N_5,In_115,In_222);
or U6 (N_6,In_43,In_343);
xor U7 (N_7,In_132,In_488);
or U8 (N_8,In_275,In_373);
xnor U9 (N_9,In_146,In_205);
nand U10 (N_10,In_203,In_72);
and U11 (N_11,In_1,In_30);
xor U12 (N_12,In_434,In_218);
xnor U13 (N_13,In_260,In_293);
and U14 (N_14,In_264,In_420);
nand U15 (N_15,In_394,In_285);
xnor U16 (N_16,In_333,In_177);
nand U17 (N_17,In_261,In_40);
nor U18 (N_18,In_269,In_313);
nand U19 (N_19,In_456,In_376);
nand U20 (N_20,In_395,In_138);
nand U21 (N_21,In_492,In_358);
nor U22 (N_22,In_85,In_254);
xor U23 (N_23,In_344,In_296);
nor U24 (N_24,In_153,In_372);
nor U25 (N_25,In_482,In_291);
nand U26 (N_26,In_249,In_448);
xnor U27 (N_27,In_332,In_457);
or U28 (N_28,In_320,In_143);
and U29 (N_29,In_472,In_196);
xnor U30 (N_30,In_364,In_474);
nand U31 (N_31,In_360,In_89);
nor U32 (N_32,In_449,In_315);
nor U33 (N_33,In_441,In_237);
or U34 (N_34,In_169,In_232);
and U35 (N_35,In_215,In_209);
nor U36 (N_36,In_246,In_4);
and U37 (N_37,In_487,In_286);
nor U38 (N_38,In_170,In_74);
xor U39 (N_39,In_413,In_7);
and U40 (N_40,In_159,In_411);
nor U41 (N_41,In_499,In_188);
nor U42 (N_42,In_314,In_450);
and U43 (N_43,In_212,In_114);
xnor U44 (N_44,In_124,In_155);
xnor U45 (N_45,In_479,In_219);
nand U46 (N_46,In_186,In_464);
nor U47 (N_47,In_105,In_113);
nand U48 (N_48,In_335,In_135);
and U49 (N_49,In_3,In_173);
and U50 (N_50,In_2,In_381);
and U51 (N_51,In_147,In_13);
nor U52 (N_52,In_483,In_243);
or U53 (N_53,In_91,In_162);
nand U54 (N_54,In_348,In_255);
nand U55 (N_55,In_42,In_330);
nand U56 (N_56,In_489,In_9);
xnor U57 (N_57,In_240,In_357);
nand U58 (N_58,In_192,In_412);
nand U59 (N_59,In_301,In_356);
or U60 (N_60,N_48,In_340);
or U61 (N_61,In_148,In_415);
or U62 (N_62,In_495,N_42);
nand U63 (N_63,In_111,In_213);
nand U64 (N_64,In_104,In_62);
and U65 (N_65,In_36,In_128);
and U66 (N_66,In_157,In_382);
or U67 (N_67,In_10,In_447);
and U68 (N_68,In_87,In_353);
nand U69 (N_69,In_48,In_436);
xor U70 (N_70,In_14,In_79);
nor U71 (N_71,In_295,In_136);
xor U72 (N_72,In_389,N_26);
nor U73 (N_73,In_459,In_362);
xnor U74 (N_74,In_365,In_83);
xor U75 (N_75,In_6,In_103);
xor U76 (N_76,In_429,In_211);
and U77 (N_77,In_262,In_354);
and U78 (N_78,In_478,In_366);
xor U79 (N_79,N_16,In_476);
xor U80 (N_80,In_331,In_280);
or U81 (N_81,In_34,In_51);
xor U82 (N_82,In_184,N_44);
nor U83 (N_83,In_398,In_99);
or U84 (N_84,In_50,N_6);
or U85 (N_85,In_20,In_145);
and U86 (N_86,In_187,In_416);
and U87 (N_87,In_207,In_175);
or U88 (N_88,In_134,In_17);
xnor U89 (N_89,In_225,In_116);
or U90 (N_90,In_279,In_29);
or U91 (N_91,In_133,In_309);
nor U92 (N_92,In_297,In_310);
nand U93 (N_93,In_403,In_463);
xor U94 (N_94,In_126,In_235);
or U95 (N_95,In_433,In_258);
or U96 (N_96,In_350,N_38);
and U97 (N_97,In_257,In_108);
nor U98 (N_98,In_191,N_35);
nand U99 (N_99,In_67,N_43);
and U100 (N_100,In_181,In_253);
nand U101 (N_101,In_82,N_18);
or U102 (N_102,In_345,In_438);
nand U103 (N_103,N_0,In_458);
and U104 (N_104,In_149,In_106);
or U105 (N_105,In_117,In_454);
or U106 (N_106,N_20,In_204);
and U107 (N_107,In_210,N_7);
or U108 (N_108,N_81,In_351);
xor U109 (N_109,In_361,In_468);
nand U110 (N_110,In_251,N_29);
and U111 (N_111,In_77,In_303);
nor U112 (N_112,In_432,In_470);
xnor U113 (N_113,In_379,In_247);
or U114 (N_114,In_273,In_63);
and U115 (N_115,In_337,In_221);
nand U116 (N_116,In_21,N_85);
nand U117 (N_117,In_431,In_405);
nor U118 (N_118,In_54,In_206);
or U119 (N_119,In_274,In_102);
or U120 (N_120,In_202,In_76);
nor U121 (N_121,N_36,N_9);
or U122 (N_122,In_75,In_22);
or U123 (N_123,N_90,In_152);
or U124 (N_124,N_28,In_28);
or U125 (N_125,N_14,In_460);
xor U126 (N_126,In_109,In_107);
or U127 (N_127,In_27,In_88);
nor U128 (N_128,N_25,In_110);
nand U129 (N_129,In_178,N_70);
nand U130 (N_130,In_370,In_305);
nor U131 (N_131,In_461,In_248);
nor U132 (N_132,N_32,In_266);
or U133 (N_133,In_90,N_65);
xor U134 (N_134,In_197,In_371);
or U135 (N_135,In_312,In_400);
or U136 (N_136,N_47,In_122);
nand U137 (N_137,In_236,N_99);
and U138 (N_138,In_341,N_97);
or U139 (N_139,N_76,In_220);
nand U140 (N_140,In_497,In_195);
nand U141 (N_141,In_231,In_426);
xor U142 (N_142,In_46,In_70);
and U143 (N_143,In_328,In_24);
and U144 (N_144,In_25,In_56);
nand U145 (N_145,In_59,In_491);
and U146 (N_146,In_435,In_302);
nor U147 (N_147,In_445,In_452);
or U148 (N_148,In_224,In_140);
nand U149 (N_149,In_244,In_352);
xnor U150 (N_150,N_24,N_73);
nand U151 (N_151,In_334,N_39);
and U152 (N_152,In_383,N_10);
nand U153 (N_153,N_143,N_134);
and U154 (N_154,In_39,N_112);
xnor U155 (N_155,In_198,N_147);
xnor U156 (N_156,In_327,N_116);
nand U157 (N_157,In_38,In_120);
xor U158 (N_158,In_73,In_130);
nor U159 (N_159,In_217,In_384);
and U160 (N_160,In_60,N_105);
and U161 (N_161,N_144,In_481);
nor U162 (N_162,In_339,N_67);
nand U163 (N_163,In_101,In_57);
nand U164 (N_164,N_40,In_137);
xor U165 (N_165,In_439,In_119);
nor U166 (N_166,N_66,In_131);
nand U167 (N_167,N_57,In_473);
xnor U168 (N_168,N_132,In_467);
xor U169 (N_169,In_5,In_256);
nand U170 (N_170,In_167,In_388);
and U171 (N_171,In_375,In_123);
nor U172 (N_172,In_234,In_223);
xnor U173 (N_173,N_82,N_108);
or U174 (N_174,In_252,In_486);
and U175 (N_175,In_377,N_115);
and U176 (N_176,N_119,In_11);
or U177 (N_177,In_55,In_469);
and U178 (N_178,In_18,In_462);
nor U179 (N_179,In_319,In_430);
nor U180 (N_180,N_58,N_109);
xnor U181 (N_181,In_23,In_378);
or U182 (N_182,In_214,In_282);
nor U183 (N_183,In_325,N_117);
xnor U184 (N_184,N_3,In_239);
and U185 (N_185,In_277,In_406);
nor U186 (N_186,N_96,N_93);
xor U187 (N_187,In_408,N_52);
nor U188 (N_188,In_444,In_369);
and U189 (N_189,In_386,In_485);
xor U190 (N_190,In_242,N_17);
and U191 (N_191,In_283,In_97);
nor U192 (N_192,N_142,N_104);
xnor U193 (N_193,In_190,In_100);
nand U194 (N_194,In_94,In_342);
xnor U195 (N_195,In_47,In_98);
nand U196 (N_196,In_141,In_194);
or U197 (N_197,In_31,In_78);
or U198 (N_198,In_49,In_471);
nand U199 (N_199,In_71,In_19);
xnor U200 (N_200,N_8,In_455);
xor U201 (N_201,N_15,N_41);
and U202 (N_202,In_26,N_50);
nand U203 (N_203,In_477,N_191);
nor U204 (N_204,In_427,In_68);
nor U205 (N_205,In_396,N_118);
nor U206 (N_206,N_12,N_155);
nand U207 (N_207,N_107,In_346);
nor U208 (N_208,N_184,In_81);
and U209 (N_209,N_188,In_387);
or U210 (N_210,In_156,N_2);
nand U211 (N_211,In_401,N_71);
or U212 (N_212,In_267,N_37);
or U213 (N_213,In_144,In_93);
nand U214 (N_214,N_179,N_163);
nand U215 (N_215,N_21,N_131);
nor U216 (N_216,N_94,N_124);
xnor U217 (N_217,In_428,N_56);
nor U218 (N_218,N_169,N_168);
nand U219 (N_219,In_245,N_197);
and U220 (N_220,N_149,N_154);
xor U221 (N_221,In_53,In_259);
nor U222 (N_222,N_140,In_69);
nor U223 (N_223,In_58,N_100);
and U224 (N_224,N_4,In_16);
and U225 (N_225,N_87,In_12);
and U226 (N_226,In_407,In_45);
nor U227 (N_227,In_287,In_185);
or U228 (N_228,In_419,In_437);
xor U229 (N_229,N_174,In_380);
and U230 (N_230,N_139,N_181);
nand U231 (N_231,N_183,N_171);
and U232 (N_232,N_49,In_289);
nand U233 (N_233,In_174,In_480);
nor U234 (N_234,In_183,N_120);
and U235 (N_235,N_146,In_451);
nand U236 (N_236,N_68,N_113);
xnor U237 (N_237,In_453,In_32);
nor U238 (N_238,In_440,N_150);
nor U239 (N_239,N_78,N_159);
or U240 (N_240,In_306,In_86);
and U241 (N_241,N_126,In_446);
xor U242 (N_242,N_122,In_397);
nand U243 (N_243,In_33,In_150);
and U244 (N_244,N_27,N_114);
or U245 (N_245,In_201,N_92);
xor U246 (N_246,In_84,N_111);
or U247 (N_247,N_106,N_138);
nor U248 (N_248,In_180,In_368);
xor U249 (N_249,In_199,N_130);
or U250 (N_250,N_239,In_300);
or U251 (N_251,In_179,N_95);
nor U252 (N_252,N_246,N_137);
xnor U253 (N_253,In_484,N_190);
or U254 (N_254,N_243,N_125);
and U255 (N_255,In_298,N_77);
nand U256 (N_256,N_121,In_238);
nand U257 (N_257,N_211,N_54);
xor U258 (N_258,N_152,N_164);
nand U259 (N_259,N_238,N_135);
or U260 (N_260,In_321,N_222);
nor U261 (N_261,N_194,N_170);
xor U262 (N_262,In_250,N_213);
xor U263 (N_263,N_11,N_178);
and U264 (N_264,In_41,N_46);
nor U265 (N_265,N_34,In_349);
and U266 (N_266,In_304,N_196);
and U267 (N_267,In_182,N_208);
nand U268 (N_268,In_490,N_217);
nor U269 (N_269,In_158,N_200);
xnor U270 (N_270,N_53,In_465);
nand U271 (N_271,In_391,N_102);
nand U272 (N_272,In_265,In_127);
xor U273 (N_273,In_399,In_374);
xnor U274 (N_274,N_221,N_167);
xnor U275 (N_275,In_318,N_242);
nand U276 (N_276,In_61,N_226);
or U277 (N_277,In_44,In_121);
nand U278 (N_278,N_72,N_199);
nand U279 (N_279,In_423,In_166);
xor U280 (N_280,N_153,N_51);
xor U281 (N_281,In_311,N_205);
nand U282 (N_282,In_494,N_210);
xor U283 (N_283,N_173,N_22);
or U284 (N_284,N_63,In_95);
and U285 (N_285,N_248,In_226);
and U286 (N_286,N_193,In_336);
xor U287 (N_287,In_118,N_236);
xnor U288 (N_288,N_215,In_263);
xnor U289 (N_289,In_64,In_208);
and U290 (N_290,In_324,In_417);
nand U291 (N_291,In_270,In_363);
and U292 (N_292,N_23,In_466);
or U293 (N_293,In_288,N_192);
and U294 (N_294,In_307,N_198);
or U295 (N_295,In_475,N_45);
xnor U296 (N_296,In_410,In_329);
or U297 (N_297,N_176,In_385);
or U298 (N_298,N_133,In_163);
nand U299 (N_299,N_158,In_402);
or U300 (N_300,In_422,N_202);
nor U301 (N_301,In_294,N_275);
or U302 (N_302,In_355,In_316);
or U303 (N_303,N_261,N_281);
nand U304 (N_304,N_148,N_185);
xnor U305 (N_305,N_253,In_367);
xnor U306 (N_306,N_75,In_404);
xnor U307 (N_307,In_200,N_264);
and U308 (N_308,In_165,N_214);
or U309 (N_309,N_295,N_278);
and U310 (N_310,N_228,In_35);
nor U311 (N_311,N_235,N_299);
nand U312 (N_312,N_55,N_273);
or U313 (N_313,N_98,In_359);
or U314 (N_314,N_216,N_33);
xnor U315 (N_315,N_282,N_288);
nand U316 (N_316,N_127,N_31);
xor U317 (N_317,In_92,N_234);
or U318 (N_318,In_414,In_151);
and U319 (N_319,In_322,N_260);
and U320 (N_320,N_101,N_250);
and U321 (N_321,N_180,In_66);
and U322 (N_322,In_125,N_145);
or U323 (N_323,N_269,N_224);
xor U324 (N_324,N_209,N_60);
nand U325 (N_325,In_233,N_290);
nor U326 (N_326,N_247,In_216);
and U327 (N_327,N_177,In_442);
nand U328 (N_328,In_281,N_91);
xor U329 (N_329,N_136,In_290);
nor U330 (N_330,N_219,N_284);
and U331 (N_331,In_229,In_154);
and U332 (N_332,In_299,N_258);
nor U333 (N_333,N_285,In_65);
and U334 (N_334,N_128,In_347);
or U335 (N_335,N_187,N_13);
and U336 (N_336,N_161,N_298);
nand U337 (N_337,N_289,N_103);
and U338 (N_338,In_37,N_61);
xor U339 (N_339,N_283,In_112);
nand U340 (N_340,N_123,N_277);
and U341 (N_341,N_59,In_160);
or U342 (N_342,N_156,In_272);
nor U343 (N_343,In_284,N_79);
and U344 (N_344,N_244,N_255);
xnor U345 (N_345,N_160,In_142);
xor U346 (N_346,N_263,In_393);
and U347 (N_347,N_241,N_141);
and U348 (N_348,N_64,In_139);
and U349 (N_349,N_229,In_171);
nand U350 (N_350,N_347,N_339);
or U351 (N_351,N_320,N_296);
and U352 (N_352,N_83,N_251);
and U353 (N_353,In_228,N_330);
nor U354 (N_354,N_319,In_421);
nor U355 (N_355,N_341,N_175);
nand U356 (N_356,N_1,In_168);
nor U357 (N_357,In_326,N_338);
nand U358 (N_358,N_30,In_424);
nand U359 (N_359,N_337,N_300);
or U360 (N_360,N_322,In_80);
or U361 (N_361,N_309,N_332);
nand U362 (N_362,N_280,N_343);
xnor U363 (N_363,In_323,N_306);
or U364 (N_364,In_308,In_129);
nor U365 (N_365,N_203,N_333);
nand U366 (N_366,N_157,N_349);
nand U367 (N_367,N_318,In_52);
nor U368 (N_368,N_272,N_312);
or U369 (N_369,N_227,N_19);
or U370 (N_370,N_256,N_297);
nor U371 (N_371,N_329,In_443);
nor U372 (N_372,N_310,N_189);
and U373 (N_373,N_88,N_336);
or U374 (N_374,In_276,N_317);
nor U375 (N_375,N_232,N_328);
nor U376 (N_376,N_311,N_86);
nand U377 (N_377,N_302,N_321);
and U378 (N_378,N_207,N_334);
or U379 (N_379,N_265,In_278);
xor U380 (N_380,N_270,N_195);
and U381 (N_381,N_315,N_324);
or U382 (N_382,N_292,N_276);
or U383 (N_383,N_266,N_162);
or U384 (N_384,N_182,In_8);
or U385 (N_385,N_231,N_331);
nand U386 (N_386,N_69,N_335);
nand U387 (N_387,N_294,N_305);
xor U388 (N_388,In_418,N_346);
xnor U389 (N_389,N_74,N_5);
or U390 (N_390,N_342,In_392);
nand U391 (N_391,N_268,N_165);
nor U392 (N_392,N_344,N_172);
nor U393 (N_393,N_204,In_390);
or U394 (N_394,In_409,N_225);
xnor U395 (N_395,N_286,N_257);
nor U396 (N_396,N_304,N_327);
nand U397 (N_397,N_262,N_240);
nand U398 (N_398,N_237,N_223);
nor U399 (N_399,In_189,N_316);
or U400 (N_400,N_274,N_397);
and U401 (N_401,N_303,N_387);
nand U402 (N_402,In_268,N_353);
xor U403 (N_403,N_259,N_357);
xor U404 (N_404,N_366,N_389);
or U405 (N_405,N_84,N_291);
nand U406 (N_406,N_355,N_206);
and U407 (N_407,N_386,N_313);
and U408 (N_408,N_381,N_369);
and U409 (N_409,N_380,N_372);
or U410 (N_410,In_193,N_359);
nand U411 (N_411,N_249,N_352);
nor U412 (N_412,N_377,N_340);
and U413 (N_413,N_233,N_186);
nor U414 (N_414,N_391,N_218);
or U415 (N_415,N_271,N_368);
or U416 (N_416,N_129,N_252);
or U417 (N_417,N_379,N_314);
and U418 (N_418,N_395,N_308);
nand U419 (N_419,N_361,N_398);
or U420 (N_420,N_358,In_15);
xor U421 (N_421,N_399,N_375);
nor U422 (N_422,N_393,N_370);
and U423 (N_423,N_362,N_287);
nor U424 (N_424,N_350,N_388);
nor U425 (N_425,N_371,N_356);
xor U426 (N_426,N_374,N_323);
xnor U427 (N_427,N_62,N_326);
xnor U428 (N_428,N_293,In_230);
or U429 (N_429,N_384,N_220);
and U430 (N_430,N_363,In_241);
xor U431 (N_431,In_496,N_80);
nor U432 (N_432,N_301,N_279);
or U433 (N_433,N_382,N_151);
and U434 (N_434,N_230,N_385);
or U435 (N_435,In_292,N_325);
or U436 (N_436,N_354,In_498);
and U437 (N_437,N_390,N_392);
nand U438 (N_438,N_254,N_245);
or U439 (N_439,N_166,N_376);
nand U440 (N_440,N_396,N_351);
nand U441 (N_441,N_383,N_267);
and U442 (N_442,N_360,N_364);
or U443 (N_443,N_110,N_348);
nand U444 (N_444,N_212,N_394);
xor U445 (N_445,N_89,N_365);
xnor U446 (N_446,N_373,N_345);
nand U447 (N_447,In_338,N_307);
nand U448 (N_448,In_164,N_378);
and U449 (N_449,N_367,N_201);
xnor U450 (N_450,N_432,N_410);
nand U451 (N_451,N_443,N_431);
and U452 (N_452,N_414,N_400);
and U453 (N_453,N_407,N_418);
xor U454 (N_454,N_424,N_411);
xor U455 (N_455,N_403,N_436);
and U456 (N_456,N_415,N_420);
xnor U457 (N_457,N_438,N_427);
and U458 (N_458,N_401,N_413);
xnor U459 (N_459,N_434,N_445);
xnor U460 (N_460,N_439,N_406);
nand U461 (N_461,N_409,N_448);
xnor U462 (N_462,N_442,N_402);
or U463 (N_463,N_423,N_444);
or U464 (N_464,N_428,N_422);
or U465 (N_465,N_447,N_404);
nand U466 (N_466,N_419,N_425);
or U467 (N_467,N_412,N_430);
xor U468 (N_468,N_421,N_446);
nor U469 (N_469,N_440,N_449);
nand U470 (N_470,N_426,N_429);
xor U471 (N_471,N_417,N_441);
nand U472 (N_472,N_437,N_433);
or U473 (N_473,N_405,N_435);
xor U474 (N_474,N_416,N_408);
nand U475 (N_475,N_438,N_413);
nor U476 (N_476,N_433,N_415);
or U477 (N_477,N_403,N_443);
nor U478 (N_478,N_424,N_441);
or U479 (N_479,N_438,N_416);
and U480 (N_480,N_434,N_439);
nand U481 (N_481,N_435,N_428);
nor U482 (N_482,N_420,N_406);
xor U483 (N_483,N_447,N_402);
and U484 (N_484,N_445,N_443);
nor U485 (N_485,N_415,N_424);
or U486 (N_486,N_408,N_443);
nor U487 (N_487,N_447,N_448);
nand U488 (N_488,N_413,N_429);
and U489 (N_489,N_448,N_426);
xnor U490 (N_490,N_404,N_414);
xnor U491 (N_491,N_426,N_411);
or U492 (N_492,N_431,N_410);
or U493 (N_493,N_413,N_404);
nor U494 (N_494,N_430,N_447);
and U495 (N_495,N_401,N_410);
or U496 (N_496,N_437,N_413);
nor U497 (N_497,N_444,N_414);
nand U498 (N_498,N_428,N_423);
xor U499 (N_499,N_445,N_406);
or U500 (N_500,N_486,N_468);
and U501 (N_501,N_463,N_479);
or U502 (N_502,N_453,N_461);
nor U503 (N_503,N_492,N_466);
nor U504 (N_504,N_496,N_476);
and U505 (N_505,N_458,N_481);
or U506 (N_506,N_467,N_459);
xnor U507 (N_507,N_457,N_471);
and U508 (N_508,N_482,N_480);
xor U509 (N_509,N_499,N_487);
and U510 (N_510,N_491,N_490);
nand U511 (N_511,N_483,N_474);
xnor U512 (N_512,N_475,N_460);
or U513 (N_513,N_452,N_456);
or U514 (N_514,N_473,N_497);
xnor U515 (N_515,N_493,N_455);
and U516 (N_516,N_450,N_489);
nor U517 (N_517,N_498,N_472);
xnor U518 (N_518,N_477,N_462);
or U519 (N_519,N_454,N_451);
nor U520 (N_520,N_470,N_465);
and U521 (N_521,N_469,N_464);
or U522 (N_522,N_485,N_484);
and U523 (N_523,N_494,N_478);
nor U524 (N_524,N_495,N_488);
nand U525 (N_525,N_488,N_451);
xnor U526 (N_526,N_484,N_475);
xor U527 (N_527,N_471,N_455);
nor U528 (N_528,N_464,N_473);
nor U529 (N_529,N_477,N_456);
nor U530 (N_530,N_459,N_499);
xnor U531 (N_531,N_485,N_492);
nand U532 (N_532,N_451,N_453);
xnor U533 (N_533,N_465,N_462);
and U534 (N_534,N_489,N_483);
xor U535 (N_535,N_452,N_499);
nor U536 (N_536,N_491,N_466);
xor U537 (N_537,N_460,N_450);
or U538 (N_538,N_457,N_476);
xnor U539 (N_539,N_472,N_481);
nand U540 (N_540,N_496,N_456);
nor U541 (N_541,N_467,N_466);
and U542 (N_542,N_488,N_497);
and U543 (N_543,N_488,N_466);
nand U544 (N_544,N_464,N_466);
xor U545 (N_545,N_486,N_499);
nor U546 (N_546,N_452,N_477);
xor U547 (N_547,N_494,N_477);
nor U548 (N_548,N_465,N_489);
xor U549 (N_549,N_497,N_456);
nor U550 (N_550,N_502,N_543);
xor U551 (N_551,N_522,N_506);
xor U552 (N_552,N_510,N_504);
and U553 (N_553,N_519,N_528);
nand U554 (N_554,N_541,N_545);
or U555 (N_555,N_534,N_513);
nor U556 (N_556,N_537,N_505);
and U557 (N_557,N_523,N_538);
xor U558 (N_558,N_503,N_531);
xnor U559 (N_559,N_540,N_517);
and U560 (N_560,N_500,N_526);
nor U561 (N_561,N_520,N_511);
or U562 (N_562,N_508,N_521);
and U563 (N_563,N_533,N_546);
nand U564 (N_564,N_524,N_544);
nor U565 (N_565,N_535,N_548);
and U566 (N_566,N_527,N_515);
nor U567 (N_567,N_532,N_530);
or U568 (N_568,N_539,N_525);
or U569 (N_569,N_549,N_536);
and U570 (N_570,N_516,N_547);
xor U571 (N_571,N_518,N_501);
and U572 (N_572,N_529,N_514);
nand U573 (N_573,N_509,N_507);
and U574 (N_574,N_542,N_512);
and U575 (N_575,N_526,N_512);
nand U576 (N_576,N_524,N_509);
and U577 (N_577,N_536,N_540);
xor U578 (N_578,N_505,N_519);
nand U579 (N_579,N_516,N_502);
and U580 (N_580,N_505,N_512);
xnor U581 (N_581,N_534,N_529);
nand U582 (N_582,N_548,N_522);
xor U583 (N_583,N_526,N_538);
and U584 (N_584,N_529,N_508);
nand U585 (N_585,N_530,N_505);
and U586 (N_586,N_539,N_511);
nor U587 (N_587,N_500,N_509);
xor U588 (N_588,N_517,N_509);
xnor U589 (N_589,N_504,N_518);
and U590 (N_590,N_530,N_501);
xor U591 (N_591,N_527,N_523);
nor U592 (N_592,N_521,N_534);
and U593 (N_593,N_523,N_528);
nor U594 (N_594,N_515,N_543);
xnor U595 (N_595,N_539,N_537);
xnor U596 (N_596,N_512,N_535);
nor U597 (N_597,N_537,N_517);
nand U598 (N_598,N_525,N_510);
xor U599 (N_599,N_535,N_528);
nor U600 (N_600,N_585,N_563);
nand U601 (N_601,N_582,N_587);
or U602 (N_602,N_573,N_588);
or U603 (N_603,N_555,N_579);
nand U604 (N_604,N_564,N_584);
nand U605 (N_605,N_591,N_586);
and U606 (N_606,N_596,N_556);
nor U607 (N_607,N_561,N_589);
nor U608 (N_608,N_595,N_558);
nor U609 (N_609,N_580,N_560);
nor U610 (N_610,N_553,N_552);
nor U611 (N_611,N_550,N_581);
and U612 (N_612,N_562,N_577);
nand U613 (N_613,N_565,N_578);
nor U614 (N_614,N_590,N_554);
xnor U615 (N_615,N_572,N_569);
nor U616 (N_616,N_566,N_571);
nor U617 (N_617,N_568,N_597);
nor U618 (N_618,N_598,N_574);
nor U619 (N_619,N_551,N_576);
and U620 (N_620,N_557,N_593);
xnor U621 (N_621,N_570,N_559);
and U622 (N_622,N_599,N_592);
and U623 (N_623,N_594,N_567);
nand U624 (N_624,N_583,N_575);
xor U625 (N_625,N_583,N_560);
nor U626 (N_626,N_581,N_565);
nor U627 (N_627,N_559,N_573);
or U628 (N_628,N_578,N_599);
and U629 (N_629,N_584,N_597);
xnor U630 (N_630,N_560,N_578);
xnor U631 (N_631,N_571,N_592);
and U632 (N_632,N_588,N_580);
nand U633 (N_633,N_597,N_574);
nor U634 (N_634,N_557,N_568);
xor U635 (N_635,N_566,N_597);
xor U636 (N_636,N_577,N_566);
nand U637 (N_637,N_572,N_577);
xnor U638 (N_638,N_585,N_555);
nand U639 (N_639,N_574,N_572);
and U640 (N_640,N_562,N_599);
xor U641 (N_641,N_593,N_555);
or U642 (N_642,N_573,N_574);
or U643 (N_643,N_589,N_554);
nand U644 (N_644,N_571,N_556);
or U645 (N_645,N_550,N_592);
or U646 (N_646,N_565,N_589);
xor U647 (N_647,N_595,N_594);
nand U648 (N_648,N_559,N_555);
and U649 (N_649,N_597,N_589);
or U650 (N_650,N_630,N_601);
nand U651 (N_651,N_619,N_616);
nor U652 (N_652,N_637,N_631);
xnor U653 (N_653,N_635,N_627);
xnor U654 (N_654,N_603,N_609);
or U655 (N_655,N_646,N_641);
nor U656 (N_656,N_639,N_602);
xnor U657 (N_657,N_615,N_605);
xnor U658 (N_658,N_618,N_617);
or U659 (N_659,N_612,N_640);
nor U660 (N_660,N_622,N_607);
and U661 (N_661,N_638,N_643);
nand U662 (N_662,N_620,N_606);
and U663 (N_663,N_633,N_621);
or U664 (N_664,N_613,N_608);
and U665 (N_665,N_614,N_642);
or U666 (N_666,N_623,N_629);
and U667 (N_667,N_632,N_600);
or U668 (N_668,N_611,N_649);
nand U669 (N_669,N_644,N_610);
and U670 (N_670,N_625,N_604);
xor U671 (N_671,N_645,N_647);
nor U672 (N_672,N_634,N_648);
or U673 (N_673,N_624,N_636);
or U674 (N_674,N_628,N_626);
nand U675 (N_675,N_621,N_630);
xor U676 (N_676,N_611,N_646);
xor U677 (N_677,N_610,N_619);
or U678 (N_678,N_624,N_616);
and U679 (N_679,N_646,N_631);
and U680 (N_680,N_638,N_642);
nand U681 (N_681,N_614,N_639);
or U682 (N_682,N_600,N_628);
xnor U683 (N_683,N_632,N_649);
xnor U684 (N_684,N_602,N_624);
nand U685 (N_685,N_610,N_641);
nor U686 (N_686,N_603,N_611);
nor U687 (N_687,N_637,N_605);
or U688 (N_688,N_636,N_640);
nand U689 (N_689,N_634,N_600);
nand U690 (N_690,N_605,N_626);
and U691 (N_691,N_601,N_602);
nand U692 (N_692,N_603,N_635);
and U693 (N_693,N_609,N_621);
xnor U694 (N_694,N_608,N_648);
and U695 (N_695,N_623,N_628);
xnor U696 (N_696,N_609,N_635);
xor U697 (N_697,N_630,N_634);
nor U698 (N_698,N_635,N_638);
or U699 (N_699,N_646,N_603);
or U700 (N_700,N_669,N_679);
and U701 (N_701,N_665,N_695);
nor U702 (N_702,N_650,N_682);
nor U703 (N_703,N_683,N_659);
nor U704 (N_704,N_686,N_653);
or U705 (N_705,N_671,N_664);
or U706 (N_706,N_661,N_680);
nand U707 (N_707,N_675,N_663);
or U708 (N_708,N_693,N_684);
and U709 (N_709,N_657,N_673);
or U710 (N_710,N_667,N_672);
nand U711 (N_711,N_689,N_688);
nand U712 (N_712,N_666,N_697);
nand U713 (N_713,N_692,N_658);
or U714 (N_714,N_696,N_685);
or U715 (N_715,N_670,N_681);
or U716 (N_716,N_652,N_687);
xnor U717 (N_717,N_698,N_651);
or U718 (N_718,N_656,N_676);
nand U719 (N_719,N_668,N_674);
and U720 (N_720,N_677,N_662);
nor U721 (N_721,N_699,N_690);
or U722 (N_722,N_654,N_678);
nand U723 (N_723,N_655,N_694);
nand U724 (N_724,N_660,N_691);
and U725 (N_725,N_674,N_666);
nor U726 (N_726,N_663,N_679);
or U727 (N_727,N_688,N_684);
xnor U728 (N_728,N_655,N_688);
nor U729 (N_729,N_670,N_656);
or U730 (N_730,N_674,N_695);
and U731 (N_731,N_671,N_694);
and U732 (N_732,N_693,N_692);
nand U733 (N_733,N_671,N_682);
nand U734 (N_734,N_659,N_670);
and U735 (N_735,N_674,N_673);
nand U736 (N_736,N_679,N_674);
nand U737 (N_737,N_650,N_689);
or U738 (N_738,N_656,N_652);
nand U739 (N_739,N_664,N_691);
or U740 (N_740,N_661,N_681);
or U741 (N_741,N_683,N_682);
xnor U742 (N_742,N_697,N_683);
xnor U743 (N_743,N_666,N_650);
nand U744 (N_744,N_686,N_656);
and U745 (N_745,N_655,N_690);
nand U746 (N_746,N_680,N_671);
or U747 (N_747,N_693,N_655);
and U748 (N_748,N_680,N_650);
or U749 (N_749,N_694,N_698);
nor U750 (N_750,N_708,N_740);
or U751 (N_751,N_736,N_706);
nand U752 (N_752,N_748,N_700);
xor U753 (N_753,N_723,N_743);
and U754 (N_754,N_709,N_734);
nand U755 (N_755,N_720,N_716);
nor U756 (N_756,N_738,N_733);
or U757 (N_757,N_712,N_725);
or U758 (N_758,N_721,N_702);
and U759 (N_759,N_704,N_727);
nand U760 (N_760,N_726,N_739);
xnor U761 (N_761,N_705,N_713);
nand U762 (N_762,N_724,N_735);
and U763 (N_763,N_707,N_729);
or U764 (N_764,N_742,N_737);
or U765 (N_765,N_745,N_722);
and U766 (N_766,N_728,N_703);
nand U767 (N_767,N_747,N_710);
or U768 (N_768,N_731,N_717);
nand U769 (N_769,N_732,N_701);
nor U770 (N_770,N_741,N_744);
or U771 (N_771,N_715,N_749);
or U772 (N_772,N_719,N_711);
nand U773 (N_773,N_730,N_714);
or U774 (N_774,N_746,N_718);
nor U775 (N_775,N_727,N_713);
and U776 (N_776,N_706,N_702);
xor U777 (N_777,N_712,N_704);
nor U778 (N_778,N_711,N_737);
nor U779 (N_779,N_729,N_735);
nor U780 (N_780,N_701,N_724);
xnor U781 (N_781,N_739,N_716);
or U782 (N_782,N_723,N_716);
and U783 (N_783,N_736,N_701);
and U784 (N_784,N_717,N_723);
nand U785 (N_785,N_734,N_738);
xnor U786 (N_786,N_703,N_704);
and U787 (N_787,N_730,N_711);
nand U788 (N_788,N_740,N_704);
xor U789 (N_789,N_730,N_700);
or U790 (N_790,N_738,N_707);
nand U791 (N_791,N_724,N_744);
or U792 (N_792,N_720,N_746);
or U793 (N_793,N_717,N_742);
and U794 (N_794,N_745,N_726);
nand U795 (N_795,N_716,N_728);
xnor U796 (N_796,N_744,N_702);
or U797 (N_797,N_745,N_730);
nand U798 (N_798,N_706,N_714);
or U799 (N_799,N_716,N_713);
nand U800 (N_800,N_770,N_764);
nor U801 (N_801,N_776,N_765);
or U802 (N_802,N_783,N_772);
or U803 (N_803,N_792,N_788);
and U804 (N_804,N_760,N_795);
and U805 (N_805,N_768,N_757);
nand U806 (N_806,N_754,N_791);
or U807 (N_807,N_785,N_777);
nor U808 (N_808,N_779,N_780);
or U809 (N_809,N_774,N_797);
or U810 (N_810,N_784,N_773);
nand U811 (N_811,N_793,N_787);
xor U812 (N_812,N_763,N_798);
nand U813 (N_813,N_781,N_761);
xnor U814 (N_814,N_769,N_758);
or U815 (N_815,N_778,N_755);
nand U816 (N_816,N_771,N_790);
nor U817 (N_817,N_750,N_759);
or U818 (N_818,N_753,N_756);
and U819 (N_819,N_762,N_799);
xor U820 (N_820,N_766,N_752);
and U821 (N_821,N_767,N_786);
xor U822 (N_822,N_775,N_796);
or U823 (N_823,N_782,N_794);
xor U824 (N_824,N_789,N_751);
and U825 (N_825,N_754,N_768);
xnor U826 (N_826,N_755,N_750);
or U827 (N_827,N_786,N_789);
xnor U828 (N_828,N_784,N_774);
xnor U829 (N_829,N_790,N_774);
and U830 (N_830,N_787,N_776);
nor U831 (N_831,N_798,N_754);
or U832 (N_832,N_790,N_788);
xnor U833 (N_833,N_786,N_791);
and U834 (N_834,N_780,N_750);
xor U835 (N_835,N_799,N_753);
nand U836 (N_836,N_754,N_789);
and U837 (N_837,N_770,N_778);
and U838 (N_838,N_773,N_791);
nor U839 (N_839,N_750,N_776);
nand U840 (N_840,N_763,N_753);
nand U841 (N_841,N_775,N_793);
or U842 (N_842,N_788,N_794);
nand U843 (N_843,N_751,N_785);
and U844 (N_844,N_778,N_783);
nand U845 (N_845,N_753,N_788);
or U846 (N_846,N_763,N_791);
or U847 (N_847,N_786,N_755);
nand U848 (N_848,N_766,N_782);
nor U849 (N_849,N_799,N_795);
nand U850 (N_850,N_834,N_804);
or U851 (N_851,N_822,N_821);
nor U852 (N_852,N_815,N_819);
nand U853 (N_853,N_835,N_842);
and U854 (N_854,N_838,N_848);
or U855 (N_855,N_812,N_826);
or U856 (N_856,N_846,N_832);
or U857 (N_857,N_823,N_829);
nand U858 (N_858,N_830,N_845);
nand U859 (N_859,N_816,N_800);
xor U860 (N_860,N_810,N_824);
or U861 (N_861,N_825,N_828);
nand U862 (N_862,N_849,N_837);
or U863 (N_863,N_806,N_843);
or U864 (N_864,N_801,N_820);
nor U865 (N_865,N_833,N_802);
nor U866 (N_866,N_803,N_827);
and U867 (N_867,N_809,N_805);
nand U868 (N_868,N_836,N_817);
nand U869 (N_869,N_831,N_844);
nor U870 (N_870,N_808,N_811);
xnor U871 (N_871,N_841,N_818);
nor U872 (N_872,N_814,N_847);
or U873 (N_873,N_813,N_839);
nand U874 (N_874,N_807,N_840);
or U875 (N_875,N_800,N_808);
nand U876 (N_876,N_825,N_843);
nand U877 (N_877,N_829,N_846);
xor U878 (N_878,N_849,N_841);
nand U879 (N_879,N_840,N_836);
or U880 (N_880,N_820,N_814);
xor U881 (N_881,N_822,N_802);
and U882 (N_882,N_802,N_814);
nor U883 (N_883,N_802,N_840);
nor U884 (N_884,N_840,N_834);
nor U885 (N_885,N_806,N_842);
or U886 (N_886,N_805,N_821);
nand U887 (N_887,N_803,N_839);
and U888 (N_888,N_814,N_828);
or U889 (N_889,N_831,N_849);
or U890 (N_890,N_845,N_809);
xor U891 (N_891,N_814,N_842);
nand U892 (N_892,N_804,N_827);
or U893 (N_893,N_828,N_819);
nand U894 (N_894,N_833,N_812);
and U895 (N_895,N_811,N_809);
xor U896 (N_896,N_849,N_804);
or U897 (N_897,N_841,N_822);
or U898 (N_898,N_840,N_829);
nand U899 (N_899,N_821,N_825);
nor U900 (N_900,N_867,N_894);
and U901 (N_901,N_896,N_874);
nand U902 (N_902,N_881,N_879);
nor U903 (N_903,N_890,N_859);
or U904 (N_904,N_891,N_878);
or U905 (N_905,N_863,N_858);
or U906 (N_906,N_862,N_856);
nor U907 (N_907,N_886,N_893);
and U908 (N_908,N_877,N_871);
or U909 (N_909,N_887,N_870);
or U910 (N_910,N_868,N_872);
nand U911 (N_911,N_885,N_857);
nand U912 (N_912,N_869,N_865);
nor U913 (N_913,N_873,N_875);
xor U914 (N_914,N_876,N_866);
xnor U915 (N_915,N_889,N_854);
xnor U916 (N_916,N_883,N_850);
nand U917 (N_917,N_884,N_851);
and U918 (N_918,N_882,N_899);
and U919 (N_919,N_861,N_852);
xnor U920 (N_920,N_898,N_892);
or U921 (N_921,N_888,N_897);
nor U922 (N_922,N_864,N_855);
and U923 (N_923,N_860,N_880);
and U924 (N_924,N_853,N_895);
and U925 (N_925,N_873,N_890);
nand U926 (N_926,N_850,N_860);
nand U927 (N_927,N_885,N_860);
or U928 (N_928,N_891,N_860);
xor U929 (N_929,N_878,N_862);
and U930 (N_930,N_853,N_857);
nor U931 (N_931,N_886,N_874);
xnor U932 (N_932,N_861,N_873);
and U933 (N_933,N_891,N_861);
and U934 (N_934,N_880,N_888);
and U935 (N_935,N_872,N_898);
xnor U936 (N_936,N_895,N_886);
or U937 (N_937,N_897,N_859);
nor U938 (N_938,N_890,N_853);
or U939 (N_939,N_861,N_856);
nand U940 (N_940,N_854,N_857);
or U941 (N_941,N_872,N_886);
nand U942 (N_942,N_877,N_880);
or U943 (N_943,N_885,N_855);
xnor U944 (N_944,N_859,N_855);
xnor U945 (N_945,N_862,N_877);
and U946 (N_946,N_854,N_895);
and U947 (N_947,N_893,N_855);
nand U948 (N_948,N_866,N_877);
or U949 (N_949,N_877,N_883);
nor U950 (N_950,N_919,N_943);
xnor U951 (N_951,N_904,N_935);
and U952 (N_952,N_921,N_933);
nor U953 (N_953,N_925,N_946);
nand U954 (N_954,N_907,N_909);
or U955 (N_955,N_932,N_949);
and U956 (N_956,N_927,N_939);
nor U957 (N_957,N_914,N_926);
xor U958 (N_958,N_929,N_901);
or U959 (N_959,N_902,N_918);
and U960 (N_960,N_913,N_947);
nor U961 (N_961,N_942,N_916);
or U962 (N_962,N_920,N_941);
xor U963 (N_963,N_928,N_917);
nand U964 (N_964,N_905,N_924);
or U965 (N_965,N_930,N_912);
nand U966 (N_966,N_910,N_934);
or U967 (N_967,N_945,N_923);
or U968 (N_968,N_944,N_940);
xor U969 (N_969,N_900,N_948);
or U970 (N_970,N_936,N_938);
nor U971 (N_971,N_937,N_903);
xnor U972 (N_972,N_915,N_908);
xor U973 (N_973,N_911,N_906);
nor U974 (N_974,N_931,N_922);
nand U975 (N_975,N_949,N_945);
and U976 (N_976,N_906,N_916);
and U977 (N_977,N_919,N_920);
nand U978 (N_978,N_917,N_913);
nor U979 (N_979,N_924,N_919);
xnor U980 (N_980,N_946,N_916);
nor U981 (N_981,N_936,N_933);
or U982 (N_982,N_921,N_929);
nand U983 (N_983,N_904,N_919);
nand U984 (N_984,N_924,N_901);
nand U985 (N_985,N_907,N_918);
or U986 (N_986,N_909,N_913);
and U987 (N_987,N_917,N_911);
nor U988 (N_988,N_932,N_925);
or U989 (N_989,N_922,N_917);
xor U990 (N_990,N_925,N_908);
xor U991 (N_991,N_914,N_933);
or U992 (N_992,N_947,N_941);
nor U993 (N_993,N_925,N_933);
nor U994 (N_994,N_916,N_937);
nor U995 (N_995,N_916,N_926);
nand U996 (N_996,N_935,N_927);
nand U997 (N_997,N_935,N_922);
nor U998 (N_998,N_901,N_928);
xnor U999 (N_999,N_946,N_933);
xor U1000 (N_1000,N_994,N_979);
xor U1001 (N_1001,N_980,N_951);
and U1002 (N_1002,N_989,N_965);
nand U1003 (N_1003,N_961,N_992);
xnor U1004 (N_1004,N_974,N_960);
nand U1005 (N_1005,N_978,N_964);
nor U1006 (N_1006,N_953,N_957);
nor U1007 (N_1007,N_950,N_976);
xor U1008 (N_1008,N_981,N_996);
nor U1009 (N_1009,N_970,N_998);
and U1010 (N_1010,N_956,N_983);
and U1011 (N_1011,N_969,N_954);
or U1012 (N_1012,N_966,N_968);
xnor U1013 (N_1013,N_959,N_999);
xor U1014 (N_1014,N_987,N_986);
and U1015 (N_1015,N_973,N_985);
or U1016 (N_1016,N_972,N_995);
and U1017 (N_1017,N_977,N_958);
and U1018 (N_1018,N_982,N_993);
nand U1019 (N_1019,N_952,N_984);
or U1020 (N_1020,N_971,N_991);
nand U1021 (N_1021,N_955,N_975);
xor U1022 (N_1022,N_988,N_962);
nor U1023 (N_1023,N_997,N_967);
or U1024 (N_1024,N_963,N_990);
nand U1025 (N_1025,N_971,N_989);
nand U1026 (N_1026,N_974,N_980);
nor U1027 (N_1027,N_952,N_994);
nand U1028 (N_1028,N_953,N_988);
nor U1029 (N_1029,N_975,N_954);
nor U1030 (N_1030,N_969,N_956);
or U1031 (N_1031,N_982,N_962);
nand U1032 (N_1032,N_988,N_974);
xor U1033 (N_1033,N_961,N_967);
or U1034 (N_1034,N_985,N_981);
nor U1035 (N_1035,N_995,N_959);
and U1036 (N_1036,N_996,N_995);
nand U1037 (N_1037,N_956,N_986);
nor U1038 (N_1038,N_962,N_991);
or U1039 (N_1039,N_976,N_987);
and U1040 (N_1040,N_979,N_983);
xnor U1041 (N_1041,N_951,N_967);
and U1042 (N_1042,N_962,N_972);
nand U1043 (N_1043,N_967,N_987);
xnor U1044 (N_1044,N_977,N_955);
nand U1045 (N_1045,N_953,N_975);
or U1046 (N_1046,N_972,N_983);
nand U1047 (N_1047,N_996,N_991);
or U1048 (N_1048,N_986,N_965);
or U1049 (N_1049,N_995,N_961);
or U1050 (N_1050,N_1031,N_1049);
nand U1051 (N_1051,N_1038,N_1021);
or U1052 (N_1052,N_1017,N_1012);
and U1053 (N_1053,N_1043,N_1029);
nand U1054 (N_1054,N_1048,N_1024);
and U1055 (N_1055,N_1045,N_1009);
or U1056 (N_1056,N_1016,N_1023);
and U1057 (N_1057,N_1025,N_1014);
and U1058 (N_1058,N_1015,N_1026);
and U1059 (N_1059,N_1046,N_1013);
and U1060 (N_1060,N_1039,N_1030);
nor U1061 (N_1061,N_1019,N_1010);
nand U1062 (N_1062,N_1003,N_1000);
and U1063 (N_1063,N_1005,N_1037);
xnor U1064 (N_1064,N_1040,N_1004);
xor U1065 (N_1065,N_1044,N_1008);
or U1066 (N_1066,N_1018,N_1034);
and U1067 (N_1067,N_1033,N_1006);
nor U1068 (N_1068,N_1027,N_1035);
nor U1069 (N_1069,N_1028,N_1032);
or U1070 (N_1070,N_1011,N_1007);
xnor U1071 (N_1071,N_1002,N_1001);
and U1072 (N_1072,N_1047,N_1036);
and U1073 (N_1073,N_1020,N_1042);
and U1074 (N_1074,N_1041,N_1022);
or U1075 (N_1075,N_1018,N_1021);
and U1076 (N_1076,N_1043,N_1035);
xnor U1077 (N_1077,N_1023,N_1036);
or U1078 (N_1078,N_1042,N_1014);
or U1079 (N_1079,N_1029,N_1006);
or U1080 (N_1080,N_1032,N_1045);
xor U1081 (N_1081,N_1047,N_1012);
and U1082 (N_1082,N_1046,N_1020);
nor U1083 (N_1083,N_1002,N_1045);
and U1084 (N_1084,N_1036,N_1020);
xor U1085 (N_1085,N_1031,N_1032);
nor U1086 (N_1086,N_1043,N_1012);
nor U1087 (N_1087,N_1023,N_1028);
nor U1088 (N_1088,N_1017,N_1013);
nor U1089 (N_1089,N_1038,N_1043);
nand U1090 (N_1090,N_1017,N_1041);
nor U1091 (N_1091,N_1001,N_1039);
nor U1092 (N_1092,N_1027,N_1020);
xor U1093 (N_1093,N_1037,N_1016);
and U1094 (N_1094,N_1040,N_1038);
xnor U1095 (N_1095,N_1012,N_1040);
and U1096 (N_1096,N_1009,N_1022);
nand U1097 (N_1097,N_1026,N_1024);
xor U1098 (N_1098,N_1009,N_1015);
or U1099 (N_1099,N_1025,N_1015);
and U1100 (N_1100,N_1078,N_1051);
and U1101 (N_1101,N_1082,N_1089);
or U1102 (N_1102,N_1098,N_1073);
and U1103 (N_1103,N_1099,N_1054);
nand U1104 (N_1104,N_1095,N_1093);
and U1105 (N_1105,N_1087,N_1074);
and U1106 (N_1106,N_1091,N_1080);
nand U1107 (N_1107,N_1063,N_1084);
or U1108 (N_1108,N_1053,N_1050);
xor U1109 (N_1109,N_1058,N_1097);
nor U1110 (N_1110,N_1061,N_1079);
or U1111 (N_1111,N_1075,N_1068);
nor U1112 (N_1112,N_1064,N_1055);
or U1113 (N_1113,N_1077,N_1062);
or U1114 (N_1114,N_1090,N_1052);
xor U1115 (N_1115,N_1094,N_1057);
nand U1116 (N_1116,N_1071,N_1067);
xnor U1117 (N_1117,N_1076,N_1066);
nand U1118 (N_1118,N_1092,N_1086);
nor U1119 (N_1119,N_1070,N_1081);
xnor U1120 (N_1120,N_1069,N_1059);
nand U1121 (N_1121,N_1096,N_1072);
or U1122 (N_1122,N_1056,N_1088);
and U1123 (N_1123,N_1060,N_1085);
nand U1124 (N_1124,N_1083,N_1065);
and U1125 (N_1125,N_1088,N_1050);
nor U1126 (N_1126,N_1093,N_1080);
nand U1127 (N_1127,N_1054,N_1067);
and U1128 (N_1128,N_1080,N_1068);
and U1129 (N_1129,N_1063,N_1068);
nand U1130 (N_1130,N_1096,N_1058);
nor U1131 (N_1131,N_1064,N_1054);
and U1132 (N_1132,N_1051,N_1062);
or U1133 (N_1133,N_1060,N_1083);
or U1134 (N_1134,N_1088,N_1079);
nand U1135 (N_1135,N_1088,N_1051);
and U1136 (N_1136,N_1098,N_1081);
or U1137 (N_1137,N_1070,N_1064);
or U1138 (N_1138,N_1068,N_1067);
nand U1139 (N_1139,N_1081,N_1083);
or U1140 (N_1140,N_1074,N_1099);
or U1141 (N_1141,N_1080,N_1077);
nand U1142 (N_1142,N_1070,N_1077);
nor U1143 (N_1143,N_1053,N_1063);
nor U1144 (N_1144,N_1061,N_1066);
xnor U1145 (N_1145,N_1053,N_1068);
nand U1146 (N_1146,N_1050,N_1097);
and U1147 (N_1147,N_1091,N_1056);
xor U1148 (N_1148,N_1056,N_1086);
and U1149 (N_1149,N_1055,N_1057);
and U1150 (N_1150,N_1143,N_1127);
and U1151 (N_1151,N_1114,N_1134);
xnor U1152 (N_1152,N_1109,N_1104);
xor U1153 (N_1153,N_1133,N_1106);
xnor U1154 (N_1154,N_1115,N_1112);
nor U1155 (N_1155,N_1118,N_1148);
and U1156 (N_1156,N_1113,N_1108);
xor U1157 (N_1157,N_1122,N_1100);
nand U1158 (N_1158,N_1132,N_1119);
or U1159 (N_1159,N_1110,N_1135);
and U1160 (N_1160,N_1138,N_1139);
or U1161 (N_1161,N_1149,N_1116);
xnor U1162 (N_1162,N_1120,N_1141);
and U1163 (N_1163,N_1105,N_1145);
or U1164 (N_1164,N_1102,N_1131);
nand U1165 (N_1165,N_1147,N_1128);
nand U1166 (N_1166,N_1103,N_1121);
and U1167 (N_1167,N_1142,N_1111);
and U1168 (N_1168,N_1107,N_1123);
and U1169 (N_1169,N_1144,N_1124);
and U1170 (N_1170,N_1117,N_1146);
xor U1171 (N_1171,N_1129,N_1136);
xor U1172 (N_1172,N_1126,N_1101);
nand U1173 (N_1173,N_1137,N_1125);
or U1174 (N_1174,N_1130,N_1140);
or U1175 (N_1175,N_1117,N_1147);
and U1176 (N_1176,N_1112,N_1129);
or U1177 (N_1177,N_1146,N_1109);
xnor U1178 (N_1178,N_1110,N_1149);
and U1179 (N_1179,N_1132,N_1139);
nor U1180 (N_1180,N_1141,N_1133);
nor U1181 (N_1181,N_1104,N_1135);
xor U1182 (N_1182,N_1140,N_1136);
nand U1183 (N_1183,N_1119,N_1127);
or U1184 (N_1184,N_1146,N_1105);
nor U1185 (N_1185,N_1108,N_1123);
nand U1186 (N_1186,N_1124,N_1109);
nor U1187 (N_1187,N_1107,N_1134);
or U1188 (N_1188,N_1125,N_1116);
xnor U1189 (N_1189,N_1111,N_1107);
and U1190 (N_1190,N_1127,N_1102);
xor U1191 (N_1191,N_1134,N_1129);
xnor U1192 (N_1192,N_1148,N_1116);
or U1193 (N_1193,N_1125,N_1147);
or U1194 (N_1194,N_1110,N_1128);
nor U1195 (N_1195,N_1148,N_1105);
nor U1196 (N_1196,N_1141,N_1108);
nand U1197 (N_1197,N_1130,N_1149);
nand U1198 (N_1198,N_1133,N_1111);
or U1199 (N_1199,N_1102,N_1144);
and U1200 (N_1200,N_1191,N_1194);
xor U1201 (N_1201,N_1190,N_1182);
nand U1202 (N_1202,N_1198,N_1179);
nor U1203 (N_1203,N_1199,N_1192);
xor U1204 (N_1204,N_1159,N_1173);
and U1205 (N_1205,N_1170,N_1165);
and U1206 (N_1206,N_1197,N_1186);
nor U1207 (N_1207,N_1189,N_1167);
or U1208 (N_1208,N_1187,N_1166);
nor U1209 (N_1209,N_1181,N_1193);
nor U1210 (N_1210,N_1188,N_1176);
and U1211 (N_1211,N_1178,N_1195);
nor U1212 (N_1212,N_1150,N_1151);
or U1213 (N_1213,N_1183,N_1162);
nor U1214 (N_1214,N_1175,N_1174);
and U1215 (N_1215,N_1184,N_1153);
and U1216 (N_1216,N_1157,N_1180);
nor U1217 (N_1217,N_1158,N_1156);
xnor U1218 (N_1218,N_1196,N_1154);
nor U1219 (N_1219,N_1160,N_1164);
and U1220 (N_1220,N_1168,N_1163);
or U1221 (N_1221,N_1155,N_1185);
and U1222 (N_1222,N_1169,N_1152);
or U1223 (N_1223,N_1172,N_1161);
and U1224 (N_1224,N_1171,N_1177);
or U1225 (N_1225,N_1172,N_1163);
nor U1226 (N_1226,N_1179,N_1158);
nor U1227 (N_1227,N_1185,N_1175);
nand U1228 (N_1228,N_1178,N_1156);
and U1229 (N_1229,N_1199,N_1185);
and U1230 (N_1230,N_1198,N_1180);
nand U1231 (N_1231,N_1160,N_1154);
nor U1232 (N_1232,N_1183,N_1172);
xor U1233 (N_1233,N_1156,N_1173);
and U1234 (N_1234,N_1153,N_1151);
nand U1235 (N_1235,N_1161,N_1169);
nand U1236 (N_1236,N_1180,N_1188);
xor U1237 (N_1237,N_1165,N_1168);
and U1238 (N_1238,N_1150,N_1182);
nor U1239 (N_1239,N_1189,N_1181);
and U1240 (N_1240,N_1172,N_1159);
nand U1241 (N_1241,N_1172,N_1197);
and U1242 (N_1242,N_1179,N_1182);
xnor U1243 (N_1243,N_1191,N_1171);
nor U1244 (N_1244,N_1168,N_1195);
nand U1245 (N_1245,N_1172,N_1162);
and U1246 (N_1246,N_1151,N_1159);
nor U1247 (N_1247,N_1193,N_1159);
or U1248 (N_1248,N_1177,N_1174);
and U1249 (N_1249,N_1157,N_1172);
nor U1250 (N_1250,N_1233,N_1224);
and U1251 (N_1251,N_1222,N_1229);
nand U1252 (N_1252,N_1209,N_1239);
and U1253 (N_1253,N_1236,N_1200);
nor U1254 (N_1254,N_1226,N_1230);
nor U1255 (N_1255,N_1214,N_1201);
xnor U1256 (N_1256,N_1207,N_1221);
xor U1257 (N_1257,N_1203,N_1242);
or U1258 (N_1258,N_1208,N_1235);
or U1259 (N_1259,N_1246,N_1237);
nor U1260 (N_1260,N_1205,N_1243);
xnor U1261 (N_1261,N_1210,N_1216);
and U1262 (N_1262,N_1213,N_1240);
nor U1263 (N_1263,N_1220,N_1244);
xor U1264 (N_1264,N_1232,N_1249);
nor U1265 (N_1265,N_1218,N_1248);
nor U1266 (N_1266,N_1211,N_1212);
nand U1267 (N_1267,N_1202,N_1217);
or U1268 (N_1268,N_1228,N_1245);
nand U1269 (N_1269,N_1219,N_1204);
and U1270 (N_1270,N_1238,N_1234);
or U1271 (N_1271,N_1215,N_1227);
or U1272 (N_1272,N_1206,N_1231);
nand U1273 (N_1273,N_1247,N_1225);
nor U1274 (N_1274,N_1241,N_1223);
nor U1275 (N_1275,N_1243,N_1241);
nor U1276 (N_1276,N_1230,N_1246);
and U1277 (N_1277,N_1242,N_1227);
and U1278 (N_1278,N_1246,N_1208);
nor U1279 (N_1279,N_1218,N_1209);
and U1280 (N_1280,N_1230,N_1224);
nand U1281 (N_1281,N_1225,N_1228);
and U1282 (N_1282,N_1218,N_1230);
nor U1283 (N_1283,N_1200,N_1238);
nand U1284 (N_1284,N_1205,N_1233);
or U1285 (N_1285,N_1207,N_1239);
nor U1286 (N_1286,N_1204,N_1228);
nor U1287 (N_1287,N_1248,N_1213);
nor U1288 (N_1288,N_1217,N_1241);
xor U1289 (N_1289,N_1233,N_1203);
and U1290 (N_1290,N_1209,N_1231);
nand U1291 (N_1291,N_1243,N_1235);
and U1292 (N_1292,N_1219,N_1234);
xor U1293 (N_1293,N_1221,N_1222);
nor U1294 (N_1294,N_1242,N_1216);
and U1295 (N_1295,N_1204,N_1225);
nand U1296 (N_1296,N_1206,N_1208);
or U1297 (N_1297,N_1209,N_1217);
xnor U1298 (N_1298,N_1243,N_1247);
nand U1299 (N_1299,N_1218,N_1201);
and U1300 (N_1300,N_1294,N_1269);
nor U1301 (N_1301,N_1265,N_1280);
and U1302 (N_1302,N_1263,N_1284);
and U1303 (N_1303,N_1253,N_1286);
nor U1304 (N_1304,N_1279,N_1293);
or U1305 (N_1305,N_1252,N_1272);
and U1306 (N_1306,N_1259,N_1268);
xnor U1307 (N_1307,N_1275,N_1281);
and U1308 (N_1308,N_1260,N_1256);
nand U1309 (N_1309,N_1297,N_1296);
xnor U1310 (N_1310,N_1274,N_1261);
or U1311 (N_1311,N_1288,N_1276);
and U1312 (N_1312,N_1251,N_1289);
nand U1313 (N_1313,N_1287,N_1254);
xnor U1314 (N_1314,N_1295,N_1267);
nand U1315 (N_1315,N_1278,N_1285);
xnor U1316 (N_1316,N_1257,N_1290);
and U1317 (N_1317,N_1292,N_1250);
and U1318 (N_1318,N_1273,N_1271);
or U1319 (N_1319,N_1299,N_1283);
xnor U1320 (N_1320,N_1282,N_1266);
and U1321 (N_1321,N_1262,N_1255);
nand U1322 (N_1322,N_1277,N_1264);
or U1323 (N_1323,N_1298,N_1270);
and U1324 (N_1324,N_1258,N_1291);
and U1325 (N_1325,N_1264,N_1286);
nor U1326 (N_1326,N_1296,N_1264);
nor U1327 (N_1327,N_1293,N_1287);
xor U1328 (N_1328,N_1285,N_1298);
xnor U1329 (N_1329,N_1268,N_1257);
nor U1330 (N_1330,N_1268,N_1273);
nand U1331 (N_1331,N_1250,N_1283);
nand U1332 (N_1332,N_1250,N_1260);
xnor U1333 (N_1333,N_1251,N_1271);
xor U1334 (N_1334,N_1295,N_1270);
nor U1335 (N_1335,N_1299,N_1272);
nor U1336 (N_1336,N_1262,N_1269);
nand U1337 (N_1337,N_1267,N_1251);
or U1338 (N_1338,N_1267,N_1273);
nand U1339 (N_1339,N_1291,N_1250);
nor U1340 (N_1340,N_1299,N_1250);
xnor U1341 (N_1341,N_1291,N_1266);
nor U1342 (N_1342,N_1282,N_1281);
or U1343 (N_1343,N_1268,N_1283);
or U1344 (N_1344,N_1279,N_1277);
nand U1345 (N_1345,N_1254,N_1285);
or U1346 (N_1346,N_1295,N_1256);
and U1347 (N_1347,N_1271,N_1283);
nand U1348 (N_1348,N_1289,N_1275);
xnor U1349 (N_1349,N_1294,N_1291);
and U1350 (N_1350,N_1334,N_1338);
nor U1351 (N_1351,N_1342,N_1318);
nand U1352 (N_1352,N_1308,N_1307);
and U1353 (N_1353,N_1317,N_1314);
and U1354 (N_1354,N_1333,N_1301);
and U1355 (N_1355,N_1348,N_1321);
and U1356 (N_1356,N_1336,N_1337);
nand U1357 (N_1357,N_1309,N_1347);
nand U1358 (N_1358,N_1329,N_1324);
nor U1359 (N_1359,N_1315,N_1320);
nor U1360 (N_1360,N_1322,N_1332);
or U1361 (N_1361,N_1304,N_1341);
nor U1362 (N_1362,N_1312,N_1326);
or U1363 (N_1363,N_1306,N_1319);
nor U1364 (N_1364,N_1331,N_1345);
nor U1365 (N_1365,N_1311,N_1330);
nand U1366 (N_1366,N_1313,N_1316);
and U1367 (N_1367,N_1310,N_1323);
xnor U1368 (N_1368,N_1349,N_1340);
nand U1369 (N_1369,N_1302,N_1325);
xor U1370 (N_1370,N_1300,N_1328);
nand U1371 (N_1371,N_1303,N_1327);
and U1372 (N_1372,N_1343,N_1344);
or U1373 (N_1373,N_1346,N_1335);
and U1374 (N_1374,N_1305,N_1339);
xnor U1375 (N_1375,N_1312,N_1338);
xor U1376 (N_1376,N_1330,N_1343);
xnor U1377 (N_1377,N_1311,N_1341);
nand U1378 (N_1378,N_1331,N_1303);
and U1379 (N_1379,N_1321,N_1333);
or U1380 (N_1380,N_1315,N_1304);
nor U1381 (N_1381,N_1339,N_1310);
nor U1382 (N_1382,N_1308,N_1329);
or U1383 (N_1383,N_1343,N_1341);
and U1384 (N_1384,N_1314,N_1308);
or U1385 (N_1385,N_1323,N_1346);
and U1386 (N_1386,N_1310,N_1306);
and U1387 (N_1387,N_1330,N_1320);
xnor U1388 (N_1388,N_1301,N_1328);
xor U1389 (N_1389,N_1309,N_1320);
nor U1390 (N_1390,N_1338,N_1326);
and U1391 (N_1391,N_1300,N_1324);
or U1392 (N_1392,N_1313,N_1303);
or U1393 (N_1393,N_1341,N_1336);
nand U1394 (N_1394,N_1336,N_1316);
nor U1395 (N_1395,N_1340,N_1347);
xnor U1396 (N_1396,N_1305,N_1338);
nor U1397 (N_1397,N_1323,N_1312);
and U1398 (N_1398,N_1312,N_1304);
nor U1399 (N_1399,N_1305,N_1308);
nor U1400 (N_1400,N_1385,N_1396);
nor U1401 (N_1401,N_1387,N_1393);
nor U1402 (N_1402,N_1356,N_1373);
nor U1403 (N_1403,N_1377,N_1350);
nand U1404 (N_1404,N_1355,N_1398);
or U1405 (N_1405,N_1380,N_1367);
xnor U1406 (N_1406,N_1384,N_1376);
nand U1407 (N_1407,N_1363,N_1353);
nor U1408 (N_1408,N_1352,N_1368);
and U1409 (N_1409,N_1383,N_1389);
or U1410 (N_1410,N_1388,N_1381);
nand U1411 (N_1411,N_1361,N_1360);
nand U1412 (N_1412,N_1359,N_1362);
or U1413 (N_1413,N_1397,N_1366);
xor U1414 (N_1414,N_1354,N_1369);
nor U1415 (N_1415,N_1364,N_1357);
or U1416 (N_1416,N_1372,N_1365);
nand U1417 (N_1417,N_1379,N_1394);
or U1418 (N_1418,N_1370,N_1358);
or U1419 (N_1419,N_1375,N_1392);
or U1420 (N_1420,N_1390,N_1399);
or U1421 (N_1421,N_1351,N_1382);
and U1422 (N_1422,N_1378,N_1395);
xor U1423 (N_1423,N_1386,N_1374);
or U1424 (N_1424,N_1371,N_1391);
and U1425 (N_1425,N_1374,N_1398);
xor U1426 (N_1426,N_1362,N_1371);
nand U1427 (N_1427,N_1392,N_1390);
or U1428 (N_1428,N_1387,N_1380);
xor U1429 (N_1429,N_1387,N_1361);
and U1430 (N_1430,N_1351,N_1388);
and U1431 (N_1431,N_1390,N_1386);
nand U1432 (N_1432,N_1388,N_1372);
nand U1433 (N_1433,N_1381,N_1373);
nand U1434 (N_1434,N_1393,N_1360);
and U1435 (N_1435,N_1370,N_1387);
or U1436 (N_1436,N_1385,N_1374);
xor U1437 (N_1437,N_1393,N_1374);
and U1438 (N_1438,N_1388,N_1359);
or U1439 (N_1439,N_1387,N_1365);
or U1440 (N_1440,N_1370,N_1359);
or U1441 (N_1441,N_1393,N_1383);
or U1442 (N_1442,N_1372,N_1389);
xnor U1443 (N_1443,N_1361,N_1351);
nand U1444 (N_1444,N_1353,N_1385);
xnor U1445 (N_1445,N_1374,N_1367);
xor U1446 (N_1446,N_1353,N_1362);
and U1447 (N_1447,N_1399,N_1369);
nor U1448 (N_1448,N_1364,N_1397);
nand U1449 (N_1449,N_1398,N_1393);
and U1450 (N_1450,N_1430,N_1408);
and U1451 (N_1451,N_1424,N_1401);
and U1452 (N_1452,N_1429,N_1441);
xnor U1453 (N_1453,N_1435,N_1420);
and U1454 (N_1454,N_1419,N_1445);
or U1455 (N_1455,N_1432,N_1442);
nand U1456 (N_1456,N_1436,N_1427);
nand U1457 (N_1457,N_1444,N_1413);
nor U1458 (N_1458,N_1404,N_1416);
nor U1459 (N_1459,N_1448,N_1434);
and U1460 (N_1460,N_1431,N_1449);
and U1461 (N_1461,N_1446,N_1423);
or U1462 (N_1462,N_1410,N_1426);
nand U1463 (N_1463,N_1433,N_1421);
and U1464 (N_1464,N_1447,N_1411);
nand U1465 (N_1465,N_1417,N_1443);
nor U1466 (N_1466,N_1437,N_1406);
nor U1467 (N_1467,N_1412,N_1414);
and U1468 (N_1468,N_1440,N_1418);
or U1469 (N_1469,N_1402,N_1405);
xor U1470 (N_1470,N_1438,N_1400);
nor U1471 (N_1471,N_1428,N_1439);
xnor U1472 (N_1472,N_1422,N_1415);
nor U1473 (N_1473,N_1425,N_1407);
or U1474 (N_1474,N_1403,N_1409);
and U1475 (N_1475,N_1435,N_1425);
xor U1476 (N_1476,N_1406,N_1402);
and U1477 (N_1477,N_1445,N_1447);
xor U1478 (N_1478,N_1401,N_1407);
nand U1479 (N_1479,N_1401,N_1413);
and U1480 (N_1480,N_1411,N_1446);
xnor U1481 (N_1481,N_1444,N_1443);
or U1482 (N_1482,N_1403,N_1439);
or U1483 (N_1483,N_1423,N_1445);
and U1484 (N_1484,N_1449,N_1426);
nand U1485 (N_1485,N_1412,N_1401);
xnor U1486 (N_1486,N_1447,N_1419);
and U1487 (N_1487,N_1443,N_1436);
and U1488 (N_1488,N_1426,N_1424);
nand U1489 (N_1489,N_1408,N_1427);
xnor U1490 (N_1490,N_1444,N_1449);
nor U1491 (N_1491,N_1449,N_1409);
xor U1492 (N_1492,N_1431,N_1430);
xor U1493 (N_1493,N_1430,N_1428);
xnor U1494 (N_1494,N_1405,N_1431);
nor U1495 (N_1495,N_1409,N_1429);
and U1496 (N_1496,N_1427,N_1438);
and U1497 (N_1497,N_1449,N_1402);
or U1498 (N_1498,N_1426,N_1401);
and U1499 (N_1499,N_1436,N_1441);
or U1500 (N_1500,N_1462,N_1459);
xnor U1501 (N_1501,N_1494,N_1452);
nand U1502 (N_1502,N_1461,N_1498);
nor U1503 (N_1503,N_1475,N_1484);
and U1504 (N_1504,N_1492,N_1483);
nand U1505 (N_1505,N_1476,N_1451);
or U1506 (N_1506,N_1474,N_1490);
nand U1507 (N_1507,N_1480,N_1472);
nor U1508 (N_1508,N_1481,N_1496);
xor U1509 (N_1509,N_1493,N_1465);
xor U1510 (N_1510,N_1454,N_1458);
nor U1511 (N_1511,N_1478,N_1467);
nand U1512 (N_1512,N_1466,N_1450);
nand U1513 (N_1513,N_1485,N_1463);
and U1514 (N_1514,N_1457,N_1479);
or U1515 (N_1515,N_1497,N_1489);
and U1516 (N_1516,N_1499,N_1491);
nor U1517 (N_1517,N_1482,N_1464);
nand U1518 (N_1518,N_1469,N_1487);
and U1519 (N_1519,N_1470,N_1488);
or U1520 (N_1520,N_1453,N_1473);
xor U1521 (N_1521,N_1460,N_1477);
nor U1522 (N_1522,N_1486,N_1456);
nor U1523 (N_1523,N_1471,N_1455);
and U1524 (N_1524,N_1495,N_1468);
nand U1525 (N_1525,N_1496,N_1478);
or U1526 (N_1526,N_1490,N_1452);
and U1527 (N_1527,N_1461,N_1489);
nor U1528 (N_1528,N_1484,N_1451);
xor U1529 (N_1529,N_1494,N_1481);
nor U1530 (N_1530,N_1475,N_1457);
nand U1531 (N_1531,N_1466,N_1498);
xor U1532 (N_1532,N_1451,N_1452);
xnor U1533 (N_1533,N_1496,N_1460);
nand U1534 (N_1534,N_1457,N_1468);
nor U1535 (N_1535,N_1461,N_1486);
nand U1536 (N_1536,N_1493,N_1480);
or U1537 (N_1537,N_1465,N_1490);
and U1538 (N_1538,N_1461,N_1458);
nand U1539 (N_1539,N_1460,N_1455);
or U1540 (N_1540,N_1480,N_1482);
nor U1541 (N_1541,N_1467,N_1486);
or U1542 (N_1542,N_1498,N_1467);
nor U1543 (N_1543,N_1490,N_1450);
nand U1544 (N_1544,N_1480,N_1497);
xor U1545 (N_1545,N_1456,N_1458);
nor U1546 (N_1546,N_1478,N_1464);
nor U1547 (N_1547,N_1472,N_1494);
or U1548 (N_1548,N_1499,N_1461);
and U1549 (N_1549,N_1490,N_1488);
and U1550 (N_1550,N_1535,N_1549);
or U1551 (N_1551,N_1500,N_1527);
xor U1552 (N_1552,N_1516,N_1544);
nand U1553 (N_1553,N_1501,N_1514);
xnor U1554 (N_1554,N_1507,N_1517);
and U1555 (N_1555,N_1543,N_1525);
nor U1556 (N_1556,N_1532,N_1529);
nand U1557 (N_1557,N_1531,N_1505);
and U1558 (N_1558,N_1546,N_1538);
xor U1559 (N_1559,N_1534,N_1536);
or U1560 (N_1560,N_1521,N_1530);
nor U1561 (N_1561,N_1524,N_1533);
and U1562 (N_1562,N_1541,N_1539);
or U1563 (N_1563,N_1545,N_1513);
or U1564 (N_1564,N_1512,N_1547);
nand U1565 (N_1565,N_1511,N_1540);
nand U1566 (N_1566,N_1502,N_1522);
nor U1567 (N_1567,N_1515,N_1537);
nor U1568 (N_1568,N_1518,N_1509);
nor U1569 (N_1569,N_1506,N_1548);
xor U1570 (N_1570,N_1508,N_1510);
and U1571 (N_1571,N_1520,N_1519);
nand U1572 (N_1572,N_1526,N_1528);
nand U1573 (N_1573,N_1504,N_1523);
or U1574 (N_1574,N_1542,N_1503);
nor U1575 (N_1575,N_1518,N_1519);
xor U1576 (N_1576,N_1503,N_1507);
xnor U1577 (N_1577,N_1513,N_1511);
or U1578 (N_1578,N_1514,N_1524);
nand U1579 (N_1579,N_1523,N_1503);
nor U1580 (N_1580,N_1538,N_1516);
or U1581 (N_1581,N_1531,N_1504);
xor U1582 (N_1582,N_1513,N_1517);
and U1583 (N_1583,N_1526,N_1523);
and U1584 (N_1584,N_1547,N_1534);
nor U1585 (N_1585,N_1531,N_1549);
nand U1586 (N_1586,N_1541,N_1516);
nand U1587 (N_1587,N_1532,N_1546);
xor U1588 (N_1588,N_1547,N_1543);
nand U1589 (N_1589,N_1534,N_1539);
nand U1590 (N_1590,N_1528,N_1514);
or U1591 (N_1591,N_1532,N_1541);
and U1592 (N_1592,N_1549,N_1502);
and U1593 (N_1593,N_1521,N_1531);
and U1594 (N_1594,N_1505,N_1513);
or U1595 (N_1595,N_1526,N_1545);
nor U1596 (N_1596,N_1532,N_1526);
nand U1597 (N_1597,N_1526,N_1505);
xnor U1598 (N_1598,N_1523,N_1500);
nand U1599 (N_1599,N_1536,N_1537);
and U1600 (N_1600,N_1570,N_1577);
or U1601 (N_1601,N_1593,N_1568);
nor U1602 (N_1602,N_1567,N_1563);
nand U1603 (N_1603,N_1589,N_1591);
xnor U1604 (N_1604,N_1588,N_1596);
or U1605 (N_1605,N_1587,N_1586);
nand U1606 (N_1606,N_1559,N_1564);
and U1607 (N_1607,N_1595,N_1553);
xor U1608 (N_1608,N_1572,N_1585);
or U1609 (N_1609,N_1566,N_1597);
or U1610 (N_1610,N_1554,N_1556);
xnor U1611 (N_1611,N_1574,N_1558);
nand U1612 (N_1612,N_1584,N_1550);
or U1613 (N_1613,N_1575,N_1561);
nand U1614 (N_1614,N_1590,N_1578);
or U1615 (N_1615,N_1580,N_1581);
and U1616 (N_1616,N_1598,N_1599);
nor U1617 (N_1617,N_1582,N_1579);
or U1618 (N_1618,N_1562,N_1583);
xor U1619 (N_1619,N_1551,N_1576);
xnor U1620 (N_1620,N_1557,N_1571);
nor U1621 (N_1621,N_1555,N_1552);
xor U1622 (N_1622,N_1594,N_1569);
nor U1623 (N_1623,N_1565,N_1592);
xor U1624 (N_1624,N_1560,N_1573);
nor U1625 (N_1625,N_1569,N_1579);
nand U1626 (N_1626,N_1584,N_1567);
nand U1627 (N_1627,N_1573,N_1584);
or U1628 (N_1628,N_1584,N_1568);
or U1629 (N_1629,N_1595,N_1562);
or U1630 (N_1630,N_1572,N_1555);
nor U1631 (N_1631,N_1574,N_1561);
nand U1632 (N_1632,N_1568,N_1560);
nor U1633 (N_1633,N_1552,N_1572);
xnor U1634 (N_1634,N_1558,N_1564);
nand U1635 (N_1635,N_1592,N_1590);
or U1636 (N_1636,N_1578,N_1569);
and U1637 (N_1637,N_1565,N_1554);
nor U1638 (N_1638,N_1552,N_1569);
and U1639 (N_1639,N_1563,N_1566);
or U1640 (N_1640,N_1583,N_1596);
nor U1641 (N_1641,N_1599,N_1571);
nor U1642 (N_1642,N_1587,N_1594);
nor U1643 (N_1643,N_1561,N_1583);
or U1644 (N_1644,N_1570,N_1550);
and U1645 (N_1645,N_1595,N_1560);
nor U1646 (N_1646,N_1581,N_1576);
or U1647 (N_1647,N_1579,N_1576);
xnor U1648 (N_1648,N_1568,N_1599);
nor U1649 (N_1649,N_1570,N_1597);
nor U1650 (N_1650,N_1619,N_1622);
nand U1651 (N_1651,N_1646,N_1623);
or U1652 (N_1652,N_1631,N_1603);
xnor U1653 (N_1653,N_1635,N_1638);
or U1654 (N_1654,N_1616,N_1620);
xnor U1655 (N_1655,N_1626,N_1610);
nand U1656 (N_1656,N_1628,N_1613);
or U1657 (N_1657,N_1641,N_1621);
and U1658 (N_1658,N_1637,N_1618);
nor U1659 (N_1659,N_1605,N_1649);
nand U1660 (N_1660,N_1608,N_1615);
nand U1661 (N_1661,N_1617,N_1612);
and U1662 (N_1662,N_1602,N_1609);
or U1663 (N_1663,N_1604,N_1624);
nand U1664 (N_1664,N_1634,N_1600);
and U1665 (N_1665,N_1644,N_1633);
nor U1666 (N_1666,N_1643,N_1648);
and U1667 (N_1667,N_1630,N_1629);
or U1668 (N_1668,N_1636,N_1625);
or U1669 (N_1669,N_1606,N_1645);
and U1670 (N_1670,N_1611,N_1632);
nand U1671 (N_1671,N_1627,N_1647);
nand U1672 (N_1672,N_1601,N_1640);
or U1673 (N_1673,N_1614,N_1639);
xnor U1674 (N_1674,N_1607,N_1642);
nand U1675 (N_1675,N_1628,N_1620);
and U1676 (N_1676,N_1621,N_1637);
nor U1677 (N_1677,N_1608,N_1646);
and U1678 (N_1678,N_1611,N_1634);
nand U1679 (N_1679,N_1637,N_1649);
and U1680 (N_1680,N_1624,N_1629);
or U1681 (N_1681,N_1626,N_1622);
or U1682 (N_1682,N_1621,N_1634);
or U1683 (N_1683,N_1645,N_1621);
xor U1684 (N_1684,N_1649,N_1622);
xnor U1685 (N_1685,N_1645,N_1641);
or U1686 (N_1686,N_1601,N_1638);
xor U1687 (N_1687,N_1638,N_1646);
and U1688 (N_1688,N_1600,N_1620);
or U1689 (N_1689,N_1627,N_1633);
nor U1690 (N_1690,N_1608,N_1604);
xnor U1691 (N_1691,N_1638,N_1600);
nor U1692 (N_1692,N_1635,N_1639);
xnor U1693 (N_1693,N_1648,N_1607);
nor U1694 (N_1694,N_1636,N_1646);
xor U1695 (N_1695,N_1608,N_1628);
xnor U1696 (N_1696,N_1623,N_1631);
nand U1697 (N_1697,N_1627,N_1611);
or U1698 (N_1698,N_1623,N_1635);
xnor U1699 (N_1699,N_1639,N_1642);
or U1700 (N_1700,N_1683,N_1685);
and U1701 (N_1701,N_1664,N_1672);
nand U1702 (N_1702,N_1688,N_1655);
and U1703 (N_1703,N_1671,N_1668);
nand U1704 (N_1704,N_1681,N_1670);
nor U1705 (N_1705,N_1656,N_1694);
or U1706 (N_1706,N_1689,N_1677);
nor U1707 (N_1707,N_1659,N_1690);
nand U1708 (N_1708,N_1658,N_1650);
or U1709 (N_1709,N_1682,N_1678);
and U1710 (N_1710,N_1691,N_1663);
and U1711 (N_1711,N_1680,N_1684);
or U1712 (N_1712,N_1676,N_1687);
and U1713 (N_1713,N_1657,N_1652);
or U1714 (N_1714,N_1665,N_1669);
xor U1715 (N_1715,N_1666,N_1661);
xor U1716 (N_1716,N_1686,N_1660);
xnor U1717 (N_1717,N_1692,N_1674);
nor U1718 (N_1718,N_1679,N_1654);
and U1719 (N_1719,N_1695,N_1696);
nor U1720 (N_1720,N_1667,N_1697);
or U1721 (N_1721,N_1675,N_1673);
or U1722 (N_1722,N_1662,N_1653);
and U1723 (N_1723,N_1693,N_1651);
nor U1724 (N_1724,N_1698,N_1699);
xor U1725 (N_1725,N_1683,N_1660);
nand U1726 (N_1726,N_1653,N_1682);
nor U1727 (N_1727,N_1689,N_1683);
nor U1728 (N_1728,N_1660,N_1666);
nand U1729 (N_1729,N_1650,N_1666);
nand U1730 (N_1730,N_1665,N_1678);
and U1731 (N_1731,N_1651,N_1689);
nor U1732 (N_1732,N_1659,N_1683);
and U1733 (N_1733,N_1659,N_1652);
nor U1734 (N_1734,N_1693,N_1684);
nand U1735 (N_1735,N_1663,N_1652);
and U1736 (N_1736,N_1666,N_1674);
xnor U1737 (N_1737,N_1677,N_1676);
xnor U1738 (N_1738,N_1694,N_1698);
and U1739 (N_1739,N_1653,N_1652);
nand U1740 (N_1740,N_1668,N_1699);
nand U1741 (N_1741,N_1678,N_1679);
nor U1742 (N_1742,N_1693,N_1664);
nor U1743 (N_1743,N_1657,N_1695);
or U1744 (N_1744,N_1687,N_1662);
or U1745 (N_1745,N_1657,N_1681);
nand U1746 (N_1746,N_1651,N_1697);
or U1747 (N_1747,N_1656,N_1661);
and U1748 (N_1748,N_1676,N_1679);
and U1749 (N_1749,N_1679,N_1664);
or U1750 (N_1750,N_1739,N_1701);
and U1751 (N_1751,N_1705,N_1706);
nor U1752 (N_1752,N_1719,N_1737);
and U1753 (N_1753,N_1703,N_1712);
nand U1754 (N_1754,N_1725,N_1732);
or U1755 (N_1755,N_1744,N_1715);
nor U1756 (N_1756,N_1711,N_1731);
and U1757 (N_1757,N_1704,N_1724);
xnor U1758 (N_1758,N_1738,N_1714);
and U1759 (N_1759,N_1718,N_1746);
nand U1760 (N_1760,N_1709,N_1710);
nand U1761 (N_1761,N_1702,N_1740);
or U1762 (N_1762,N_1708,N_1707);
nor U1763 (N_1763,N_1721,N_1747);
nor U1764 (N_1764,N_1736,N_1734);
and U1765 (N_1765,N_1727,N_1749);
xor U1766 (N_1766,N_1735,N_1720);
nor U1767 (N_1767,N_1726,N_1716);
or U1768 (N_1768,N_1722,N_1717);
nand U1769 (N_1769,N_1728,N_1748);
and U1770 (N_1770,N_1729,N_1745);
xnor U1771 (N_1771,N_1723,N_1730);
or U1772 (N_1772,N_1742,N_1741);
and U1773 (N_1773,N_1700,N_1713);
nor U1774 (N_1774,N_1733,N_1743);
xnor U1775 (N_1775,N_1701,N_1746);
and U1776 (N_1776,N_1747,N_1713);
xor U1777 (N_1777,N_1748,N_1739);
nand U1778 (N_1778,N_1733,N_1716);
nand U1779 (N_1779,N_1743,N_1724);
nor U1780 (N_1780,N_1705,N_1727);
nor U1781 (N_1781,N_1720,N_1704);
and U1782 (N_1782,N_1731,N_1701);
xnor U1783 (N_1783,N_1727,N_1731);
xnor U1784 (N_1784,N_1735,N_1701);
nor U1785 (N_1785,N_1744,N_1705);
and U1786 (N_1786,N_1721,N_1731);
and U1787 (N_1787,N_1717,N_1740);
or U1788 (N_1788,N_1739,N_1704);
xor U1789 (N_1789,N_1713,N_1738);
xor U1790 (N_1790,N_1748,N_1707);
xor U1791 (N_1791,N_1709,N_1706);
and U1792 (N_1792,N_1709,N_1745);
or U1793 (N_1793,N_1738,N_1716);
and U1794 (N_1794,N_1717,N_1742);
nand U1795 (N_1795,N_1722,N_1735);
or U1796 (N_1796,N_1737,N_1712);
or U1797 (N_1797,N_1710,N_1744);
nand U1798 (N_1798,N_1704,N_1721);
nand U1799 (N_1799,N_1735,N_1732);
nand U1800 (N_1800,N_1754,N_1783);
or U1801 (N_1801,N_1752,N_1785);
nand U1802 (N_1802,N_1789,N_1779);
and U1803 (N_1803,N_1778,N_1764);
nand U1804 (N_1804,N_1762,N_1784);
and U1805 (N_1805,N_1797,N_1794);
xor U1806 (N_1806,N_1773,N_1758);
nand U1807 (N_1807,N_1774,N_1786);
nor U1808 (N_1808,N_1775,N_1790);
and U1809 (N_1809,N_1799,N_1756);
or U1810 (N_1810,N_1770,N_1795);
xnor U1811 (N_1811,N_1780,N_1793);
nand U1812 (N_1812,N_1760,N_1755);
and U1813 (N_1813,N_1781,N_1759);
or U1814 (N_1814,N_1796,N_1798);
xor U1815 (N_1815,N_1766,N_1792);
or U1816 (N_1816,N_1751,N_1772);
nand U1817 (N_1817,N_1768,N_1765);
and U1818 (N_1818,N_1782,N_1791);
xor U1819 (N_1819,N_1769,N_1753);
nand U1820 (N_1820,N_1750,N_1777);
xor U1821 (N_1821,N_1763,N_1761);
or U1822 (N_1822,N_1787,N_1771);
nor U1823 (N_1823,N_1776,N_1767);
nand U1824 (N_1824,N_1788,N_1757);
and U1825 (N_1825,N_1769,N_1751);
nand U1826 (N_1826,N_1799,N_1795);
nor U1827 (N_1827,N_1787,N_1765);
or U1828 (N_1828,N_1799,N_1785);
nor U1829 (N_1829,N_1767,N_1785);
xor U1830 (N_1830,N_1792,N_1776);
nand U1831 (N_1831,N_1760,N_1751);
xnor U1832 (N_1832,N_1768,N_1791);
or U1833 (N_1833,N_1766,N_1760);
xor U1834 (N_1834,N_1763,N_1786);
and U1835 (N_1835,N_1793,N_1783);
nor U1836 (N_1836,N_1795,N_1758);
or U1837 (N_1837,N_1784,N_1795);
nor U1838 (N_1838,N_1798,N_1760);
xor U1839 (N_1839,N_1784,N_1780);
nand U1840 (N_1840,N_1754,N_1750);
nor U1841 (N_1841,N_1793,N_1787);
nor U1842 (N_1842,N_1789,N_1797);
xnor U1843 (N_1843,N_1764,N_1762);
xnor U1844 (N_1844,N_1763,N_1790);
nand U1845 (N_1845,N_1785,N_1780);
nand U1846 (N_1846,N_1750,N_1753);
and U1847 (N_1847,N_1793,N_1785);
nor U1848 (N_1848,N_1760,N_1783);
and U1849 (N_1849,N_1763,N_1785);
and U1850 (N_1850,N_1839,N_1824);
or U1851 (N_1851,N_1825,N_1829);
or U1852 (N_1852,N_1828,N_1817);
nand U1853 (N_1853,N_1811,N_1836);
xnor U1854 (N_1854,N_1831,N_1818);
or U1855 (N_1855,N_1822,N_1807);
xnor U1856 (N_1856,N_1840,N_1810);
nor U1857 (N_1857,N_1841,N_1845);
or U1858 (N_1858,N_1837,N_1830);
nand U1859 (N_1859,N_1842,N_1808);
nor U1860 (N_1860,N_1804,N_1844);
or U1861 (N_1861,N_1827,N_1816);
or U1862 (N_1862,N_1848,N_1832);
nand U1863 (N_1863,N_1820,N_1838);
and U1864 (N_1864,N_1802,N_1846);
xor U1865 (N_1865,N_1821,N_1805);
or U1866 (N_1866,N_1847,N_1823);
and U1867 (N_1867,N_1815,N_1835);
and U1868 (N_1868,N_1833,N_1849);
nor U1869 (N_1869,N_1812,N_1843);
xnor U1870 (N_1870,N_1801,N_1813);
xnor U1871 (N_1871,N_1806,N_1826);
and U1872 (N_1872,N_1809,N_1819);
xnor U1873 (N_1873,N_1803,N_1834);
and U1874 (N_1874,N_1800,N_1814);
or U1875 (N_1875,N_1816,N_1804);
nor U1876 (N_1876,N_1837,N_1847);
and U1877 (N_1877,N_1841,N_1837);
and U1878 (N_1878,N_1828,N_1802);
nand U1879 (N_1879,N_1835,N_1834);
and U1880 (N_1880,N_1818,N_1847);
xor U1881 (N_1881,N_1830,N_1849);
xnor U1882 (N_1882,N_1831,N_1812);
nor U1883 (N_1883,N_1800,N_1836);
nand U1884 (N_1884,N_1843,N_1841);
nand U1885 (N_1885,N_1847,N_1843);
nor U1886 (N_1886,N_1821,N_1820);
nand U1887 (N_1887,N_1845,N_1831);
nor U1888 (N_1888,N_1802,N_1824);
nand U1889 (N_1889,N_1848,N_1822);
and U1890 (N_1890,N_1821,N_1835);
and U1891 (N_1891,N_1813,N_1842);
nor U1892 (N_1892,N_1834,N_1825);
nor U1893 (N_1893,N_1837,N_1842);
nor U1894 (N_1894,N_1849,N_1822);
xor U1895 (N_1895,N_1826,N_1813);
and U1896 (N_1896,N_1823,N_1824);
and U1897 (N_1897,N_1823,N_1832);
nand U1898 (N_1898,N_1804,N_1807);
nor U1899 (N_1899,N_1842,N_1807);
and U1900 (N_1900,N_1852,N_1898);
nor U1901 (N_1901,N_1897,N_1860);
xnor U1902 (N_1902,N_1873,N_1883);
nor U1903 (N_1903,N_1892,N_1856);
nand U1904 (N_1904,N_1868,N_1896);
or U1905 (N_1905,N_1850,N_1869);
or U1906 (N_1906,N_1870,N_1880);
nand U1907 (N_1907,N_1889,N_1879);
nor U1908 (N_1908,N_1886,N_1872);
nand U1909 (N_1909,N_1853,N_1865);
nand U1910 (N_1910,N_1858,N_1863);
or U1911 (N_1911,N_1854,N_1871);
and U1912 (N_1912,N_1876,N_1882);
or U1913 (N_1913,N_1890,N_1893);
nor U1914 (N_1914,N_1877,N_1888);
xnor U1915 (N_1915,N_1864,N_1887);
nand U1916 (N_1916,N_1862,N_1881);
xor U1917 (N_1917,N_1899,N_1894);
xor U1918 (N_1918,N_1851,N_1857);
nor U1919 (N_1919,N_1895,N_1878);
or U1920 (N_1920,N_1874,N_1885);
and U1921 (N_1921,N_1866,N_1891);
xor U1922 (N_1922,N_1884,N_1875);
nand U1923 (N_1923,N_1861,N_1867);
or U1924 (N_1924,N_1859,N_1855);
nand U1925 (N_1925,N_1870,N_1877);
xor U1926 (N_1926,N_1856,N_1887);
or U1927 (N_1927,N_1878,N_1899);
nand U1928 (N_1928,N_1889,N_1887);
xnor U1929 (N_1929,N_1873,N_1889);
nand U1930 (N_1930,N_1856,N_1850);
xnor U1931 (N_1931,N_1851,N_1869);
nor U1932 (N_1932,N_1879,N_1852);
and U1933 (N_1933,N_1867,N_1886);
or U1934 (N_1934,N_1895,N_1860);
and U1935 (N_1935,N_1896,N_1893);
and U1936 (N_1936,N_1877,N_1892);
xor U1937 (N_1937,N_1874,N_1871);
xnor U1938 (N_1938,N_1873,N_1893);
xor U1939 (N_1939,N_1850,N_1876);
xor U1940 (N_1940,N_1896,N_1858);
nor U1941 (N_1941,N_1872,N_1853);
and U1942 (N_1942,N_1856,N_1854);
xnor U1943 (N_1943,N_1851,N_1882);
or U1944 (N_1944,N_1892,N_1894);
nand U1945 (N_1945,N_1881,N_1872);
and U1946 (N_1946,N_1886,N_1888);
nand U1947 (N_1947,N_1881,N_1880);
and U1948 (N_1948,N_1872,N_1883);
nor U1949 (N_1949,N_1899,N_1851);
nor U1950 (N_1950,N_1941,N_1917);
nand U1951 (N_1951,N_1948,N_1925);
xnor U1952 (N_1952,N_1936,N_1933);
nand U1953 (N_1953,N_1914,N_1928);
nand U1954 (N_1954,N_1920,N_1931);
nor U1955 (N_1955,N_1924,N_1921);
or U1956 (N_1956,N_1910,N_1942);
or U1957 (N_1957,N_1940,N_1923);
and U1958 (N_1958,N_1937,N_1944);
and U1959 (N_1959,N_1900,N_1911);
and U1960 (N_1960,N_1904,N_1945);
nand U1961 (N_1961,N_1932,N_1934);
xor U1962 (N_1962,N_1947,N_1922);
or U1963 (N_1963,N_1901,N_1915);
nor U1964 (N_1964,N_1902,N_1946);
nor U1965 (N_1965,N_1905,N_1919);
and U1966 (N_1966,N_1913,N_1908);
nor U1967 (N_1967,N_1949,N_1909);
xor U1968 (N_1968,N_1906,N_1912);
nand U1969 (N_1969,N_1939,N_1930);
nor U1970 (N_1970,N_1918,N_1935);
xor U1971 (N_1971,N_1927,N_1938);
or U1972 (N_1972,N_1916,N_1903);
nand U1973 (N_1973,N_1907,N_1943);
nand U1974 (N_1974,N_1929,N_1926);
and U1975 (N_1975,N_1912,N_1928);
or U1976 (N_1976,N_1944,N_1930);
nand U1977 (N_1977,N_1933,N_1904);
nor U1978 (N_1978,N_1944,N_1912);
nor U1979 (N_1979,N_1910,N_1927);
or U1980 (N_1980,N_1908,N_1944);
nor U1981 (N_1981,N_1942,N_1922);
nand U1982 (N_1982,N_1937,N_1941);
nor U1983 (N_1983,N_1948,N_1911);
and U1984 (N_1984,N_1932,N_1946);
nand U1985 (N_1985,N_1924,N_1915);
and U1986 (N_1986,N_1927,N_1944);
xor U1987 (N_1987,N_1930,N_1933);
nor U1988 (N_1988,N_1932,N_1928);
nor U1989 (N_1989,N_1908,N_1926);
nor U1990 (N_1990,N_1944,N_1906);
or U1991 (N_1991,N_1913,N_1909);
nand U1992 (N_1992,N_1933,N_1920);
xor U1993 (N_1993,N_1943,N_1927);
and U1994 (N_1994,N_1904,N_1905);
xnor U1995 (N_1995,N_1924,N_1907);
and U1996 (N_1996,N_1936,N_1929);
or U1997 (N_1997,N_1943,N_1933);
nand U1998 (N_1998,N_1943,N_1945);
nor U1999 (N_1999,N_1905,N_1933);
xnor U2000 (N_2000,N_1951,N_1953);
nor U2001 (N_2001,N_1955,N_1954);
xnor U2002 (N_2002,N_1996,N_1960);
nor U2003 (N_2003,N_1972,N_1976);
nand U2004 (N_2004,N_1962,N_1963);
or U2005 (N_2005,N_1979,N_1966);
xor U2006 (N_2006,N_1995,N_1974);
nand U2007 (N_2007,N_1970,N_1958);
xnor U2008 (N_2008,N_1977,N_1956);
nand U2009 (N_2009,N_1973,N_1990);
xor U2010 (N_2010,N_1998,N_1991);
or U2011 (N_2011,N_1984,N_1981);
xnor U2012 (N_2012,N_1952,N_1986);
nand U2013 (N_2013,N_1999,N_1978);
xor U2014 (N_2014,N_1968,N_1975);
nand U2015 (N_2015,N_1957,N_1994);
or U2016 (N_2016,N_1961,N_1971);
xor U2017 (N_2017,N_1969,N_1992);
nand U2018 (N_2018,N_1983,N_1950);
xor U2019 (N_2019,N_1988,N_1965);
xor U2020 (N_2020,N_1997,N_1980);
or U2021 (N_2021,N_1964,N_1982);
xor U2022 (N_2022,N_1989,N_1967);
nand U2023 (N_2023,N_1959,N_1993);
xnor U2024 (N_2024,N_1985,N_1987);
xnor U2025 (N_2025,N_1975,N_1952);
and U2026 (N_2026,N_1954,N_1958);
or U2027 (N_2027,N_1961,N_1953);
or U2028 (N_2028,N_1955,N_1998);
or U2029 (N_2029,N_1970,N_1955);
nor U2030 (N_2030,N_1999,N_1968);
and U2031 (N_2031,N_1985,N_1951);
nand U2032 (N_2032,N_1974,N_1960);
or U2033 (N_2033,N_1977,N_1985);
nor U2034 (N_2034,N_1973,N_1979);
nand U2035 (N_2035,N_1977,N_1955);
or U2036 (N_2036,N_1988,N_1967);
or U2037 (N_2037,N_1978,N_1984);
xor U2038 (N_2038,N_1968,N_1988);
and U2039 (N_2039,N_1970,N_1961);
or U2040 (N_2040,N_1983,N_1951);
or U2041 (N_2041,N_1974,N_1958);
or U2042 (N_2042,N_1954,N_1992);
and U2043 (N_2043,N_1981,N_1953);
nor U2044 (N_2044,N_1976,N_1950);
nor U2045 (N_2045,N_1969,N_1957);
and U2046 (N_2046,N_1983,N_1956);
nor U2047 (N_2047,N_1953,N_1992);
and U2048 (N_2048,N_1967,N_1968);
or U2049 (N_2049,N_1979,N_1994);
or U2050 (N_2050,N_2005,N_2019);
xor U2051 (N_2051,N_2021,N_2048);
or U2052 (N_2052,N_2013,N_2002);
xnor U2053 (N_2053,N_2025,N_2018);
nor U2054 (N_2054,N_2023,N_2036);
or U2055 (N_2055,N_2004,N_2009);
nand U2056 (N_2056,N_2047,N_2038);
nand U2057 (N_2057,N_2046,N_2044);
nand U2058 (N_2058,N_2039,N_2024);
nand U2059 (N_2059,N_2041,N_2034);
nand U2060 (N_2060,N_2017,N_2031);
or U2061 (N_2061,N_2012,N_2033);
nand U2062 (N_2062,N_2003,N_2008);
or U2063 (N_2063,N_2011,N_2026);
xnor U2064 (N_2064,N_2006,N_2049);
xnor U2065 (N_2065,N_2040,N_2010);
or U2066 (N_2066,N_2015,N_2042);
nor U2067 (N_2067,N_2016,N_2014);
or U2068 (N_2068,N_2001,N_2007);
and U2069 (N_2069,N_2020,N_2000);
or U2070 (N_2070,N_2030,N_2029);
or U2071 (N_2071,N_2043,N_2032);
nor U2072 (N_2072,N_2027,N_2037);
xor U2073 (N_2073,N_2035,N_2022);
nand U2074 (N_2074,N_2028,N_2045);
and U2075 (N_2075,N_2044,N_2000);
xnor U2076 (N_2076,N_2021,N_2025);
and U2077 (N_2077,N_2027,N_2022);
nand U2078 (N_2078,N_2018,N_2034);
nor U2079 (N_2079,N_2038,N_2018);
nand U2080 (N_2080,N_2012,N_2021);
nand U2081 (N_2081,N_2030,N_2043);
and U2082 (N_2082,N_2044,N_2048);
xnor U2083 (N_2083,N_2024,N_2001);
and U2084 (N_2084,N_2045,N_2011);
nor U2085 (N_2085,N_2032,N_2004);
and U2086 (N_2086,N_2029,N_2038);
or U2087 (N_2087,N_2010,N_2017);
and U2088 (N_2088,N_2013,N_2010);
nand U2089 (N_2089,N_2000,N_2012);
or U2090 (N_2090,N_2012,N_2045);
xnor U2091 (N_2091,N_2000,N_2030);
and U2092 (N_2092,N_2006,N_2034);
xnor U2093 (N_2093,N_2035,N_2037);
nand U2094 (N_2094,N_2007,N_2019);
xor U2095 (N_2095,N_2004,N_2048);
nand U2096 (N_2096,N_2030,N_2045);
nor U2097 (N_2097,N_2008,N_2016);
and U2098 (N_2098,N_2014,N_2046);
nand U2099 (N_2099,N_2044,N_2003);
nor U2100 (N_2100,N_2097,N_2080);
nand U2101 (N_2101,N_2089,N_2078);
xnor U2102 (N_2102,N_2059,N_2092);
and U2103 (N_2103,N_2067,N_2064);
nand U2104 (N_2104,N_2072,N_2096);
or U2105 (N_2105,N_2063,N_2090);
nor U2106 (N_2106,N_2056,N_2086);
or U2107 (N_2107,N_2075,N_2093);
and U2108 (N_2108,N_2091,N_2095);
nand U2109 (N_2109,N_2088,N_2060);
and U2110 (N_2110,N_2074,N_2083);
xor U2111 (N_2111,N_2058,N_2087);
xnor U2112 (N_2112,N_2077,N_2071);
nand U2113 (N_2113,N_2068,N_2079);
nand U2114 (N_2114,N_2062,N_2081);
xnor U2115 (N_2115,N_2050,N_2054);
or U2116 (N_2116,N_2098,N_2094);
and U2117 (N_2117,N_2057,N_2052);
nor U2118 (N_2118,N_2051,N_2055);
nor U2119 (N_2119,N_2073,N_2069);
xnor U2120 (N_2120,N_2070,N_2099);
xor U2121 (N_2121,N_2065,N_2082);
nand U2122 (N_2122,N_2061,N_2066);
nor U2123 (N_2123,N_2084,N_2076);
or U2124 (N_2124,N_2085,N_2053);
nand U2125 (N_2125,N_2064,N_2051);
and U2126 (N_2126,N_2056,N_2082);
nor U2127 (N_2127,N_2078,N_2097);
xnor U2128 (N_2128,N_2067,N_2054);
and U2129 (N_2129,N_2052,N_2078);
or U2130 (N_2130,N_2065,N_2076);
or U2131 (N_2131,N_2082,N_2052);
or U2132 (N_2132,N_2065,N_2094);
and U2133 (N_2133,N_2086,N_2076);
and U2134 (N_2134,N_2090,N_2092);
xor U2135 (N_2135,N_2052,N_2093);
xor U2136 (N_2136,N_2099,N_2058);
nand U2137 (N_2137,N_2077,N_2094);
nor U2138 (N_2138,N_2056,N_2091);
or U2139 (N_2139,N_2079,N_2098);
and U2140 (N_2140,N_2061,N_2076);
xor U2141 (N_2141,N_2068,N_2056);
nor U2142 (N_2142,N_2082,N_2075);
xor U2143 (N_2143,N_2087,N_2051);
and U2144 (N_2144,N_2071,N_2099);
nor U2145 (N_2145,N_2052,N_2056);
and U2146 (N_2146,N_2068,N_2095);
nor U2147 (N_2147,N_2073,N_2053);
or U2148 (N_2148,N_2080,N_2063);
xor U2149 (N_2149,N_2099,N_2066);
xor U2150 (N_2150,N_2128,N_2110);
and U2151 (N_2151,N_2109,N_2108);
xor U2152 (N_2152,N_2113,N_2147);
nor U2153 (N_2153,N_2136,N_2131);
xnor U2154 (N_2154,N_2135,N_2101);
or U2155 (N_2155,N_2143,N_2123);
or U2156 (N_2156,N_2132,N_2142);
nand U2157 (N_2157,N_2117,N_2116);
nor U2158 (N_2158,N_2124,N_2129);
nand U2159 (N_2159,N_2120,N_2140);
xnor U2160 (N_2160,N_2139,N_2146);
nand U2161 (N_2161,N_2114,N_2105);
and U2162 (N_2162,N_2112,N_2121);
nand U2163 (N_2163,N_2104,N_2134);
or U2164 (N_2164,N_2106,N_2148);
or U2165 (N_2165,N_2111,N_2119);
nor U2166 (N_2166,N_2122,N_2125);
nand U2167 (N_2167,N_2107,N_2138);
nand U2168 (N_2168,N_2126,N_2144);
xor U2169 (N_2169,N_2130,N_2118);
and U2170 (N_2170,N_2133,N_2102);
nand U2171 (N_2171,N_2103,N_2145);
xnor U2172 (N_2172,N_2137,N_2149);
nand U2173 (N_2173,N_2100,N_2115);
xor U2174 (N_2174,N_2141,N_2127);
or U2175 (N_2175,N_2124,N_2148);
and U2176 (N_2176,N_2124,N_2134);
or U2177 (N_2177,N_2123,N_2109);
or U2178 (N_2178,N_2113,N_2143);
xnor U2179 (N_2179,N_2100,N_2118);
xor U2180 (N_2180,N_2116,N_2128);
and U2181 (N_2181,N_2125,N_2146);
xnor U2182 (N_2182,N_2147,N_2105);
nor U2183 (N_2183,N_2123,N_2111);
and U2184 (N_2184,N_2129,N_2133);
xnor U2185 (N_2185,N_2149,N_2131);
nor U2186 (N_2186,N_2149,N_2102);
and U2187 (N_2187,N_2105,N_2123);
nand U2188 (N_2188,N_2106,N_2103);
nor U2189 (N_2189,N_2144,N_2101);
xnor U2190 (N_2190,N_2114,N_2148);
nor U2191 (N_2191,N_2147,N_2135);
and U2192 (N_2192,N_2126,N_2124);
xnor U2193 (N_2193,N_2111,N_2149);
and U2194 (N_2194,N_2132,N_2136);
or U2195 (N_2195,N_2107,N_2127);
xnor U2196 (N_2196,N_2128,N_2108);
nor U2197 (N_2197,N_2114,N_2132);
nor U2198 (N_2198,N_2109,N_2129);
or U2199 (N_2199,N_2123,N_2140);
nor U2200 (N_2200,N_2181,N_2161);
or U2201 (N_2201,N_2199,N_2186);
or U2202 (N_2202,N_2166,N_2183);
nor U2203 (N_2203,N_2179,N_2173);
nor U2204 (N_2204,N_2185,N_2187);
nand U2205 (N_2205,N_2157,N_2198);
nand U2206 (N_2206,N_2184,N_2158);
nor U2207 (N_2207,N_2195,N_2176);
nor U2208 (N_2208,N_2197,N_2156);
nor U2209 (N_2209,N_2193,N_2155);
xnor U2210 (N_2210,N_2154,N_2196);
xor U2211 (N_2211,N_2150,N_2170);
and U2212 (N_2212,N_2165,N_2153);
nand U2213 (N_2213,N_2163,N_2192);
or U2214 (N_2214,N_2152,N_2151);
nor U2215 (N_2215,N_2169,N_2167);
and U2216 (N_2216,N_2162,N_2190);
xor U2217 (N_2217,N_2189,N_2159);
and U2218 (N_2218,N_2177,N_2175);
nand U2219 (N_2219,N_2164,N_2168);
nand U2220 (N_2220,N_2194,N_2182);
and U2221 (N_2221,N_2178,N_2188);
nor U2222 (N_2222,N_2172,N_2160);
or U2223 (N_2223,N_2191,N_2180);
and U2224 (N_2224,N_2171,N_2174);
nand U2225 (N_2225,N_2185,N_2195);
nor U2226 (N_2226,N_2173,N_2193);
and U2227 (N_2227,N_2175,N_2181);
xnor U2228 (N_2228,N_2151,N_2164);
nand U2229 (N_2229,N_2198,N_2188);
nor U2230 (N_2230,N_2156,N_2180);
xnor U2231 (N_2231,N_2190,N_2178);
nor U2232 (N_2232,N_2193,N_2169);
and U2233 (N_2233,N_2177,N_2198);
or U2234 (N_2234,N_2180,N_2185);
xnor U2235 (N_2235,N_2198,N_2187);
and U2236 (N_2236,N_2167,N_2192);
nor U2237 (N_2237,N_2192,N_2181);
nor U2238 (N_2238,N_2174,N_2165);
nor U2239 (N_2239,N_2181,N_2168);
and U2240 (N_2240,N_2183,N_2161);
and U2241 (N_2241,N_2196,N_2185);
nor U2242 (N_2242,N_2178,N_2182);
and U2243 (N_2243,N_2194,N_2176);
and U2244 (N_2244,N_2167,N_2197);
nor U2245 (N_2245,N_2180,N_2187);
and U2246 (N_2246,N_2193,N_2150);
xnor U2247 (N_2247,N_2171,N_2188);
or U2248 (N_2248,N_2185,N_2150);
nor U2249 (N_2249,N_2169,N_2177);
xnor U2250 (N_2250,N_2236,N_2206);
nor U2251 (N_2251,N_2225,N_2229);
and U2252 (N_2252,N_2240,N_2241);
or U2253 (N_2253,N_2205,N_2239);
xnor U2254 (N_2254,N_2249,N_2234);
and U2255 (N_2255,N_2233,N_2211);
nand U2256 (N_2256,N_2235,N_2247);
and U2257 (N_2257,N_2203,N_2230);
nand U2258 (N_2258,N_2209,N_2231);
nor U2259 (N_2259,N_2227,N_2221);
xor U2260 (N_2260,N_2238,N_2207);
and U2261 (N_2261,N_2210,N_2242);
and U2262 (N_2262,N_2204,N_2246);
or U2263 (N_2263,N_2217,N_2226);
nor U2264 (N_2264,N_2215,N_2202);
nand U2265 (N_2265,N_2222,N_2218);
nand U2266 (N_2266,N_2224,N_2237);
xor U2267 (N_2267,N_2244,N_2220);
xor U2268 (N_2268,N_2232,N_2200);
nand U2269 (N_2269,N_2216,N_2223);
nand U2270 (N_2270,N_2212,N_2213);
and U2271 (N_2271,N_2214,N_2201);
or U2272 (N_2272,N_2243,N_2219);
nand U2273 (N_2273,N_2228,N_2248);
or U2274 (N_2274,N_2245,N_2208);
nor U2275 (N_2275,N_2203,N_2226);
xnor U2276 (N_2276,N_2215,N_2201);
and U2277 (N_2277,N_2230,N_2236);
and U2278 (N_2278,N_2225,N_2210);
nand U2279 (N_2279,N_2241,N_2200);
or U2280 (N_2280,N_2200,N_2218);
and U2281 (N_2281,N_2208,N_2227);
nor U2282 (N_2282,N_2225,N_2209);
or U2283 (N_2283,N_2244,N_2218);
or U2284 (N_2284,N_2204,N_2241);
or U2285 (N_2285,N_2203,N_2231);
xor U2286 (N_2286,N_2234,N_2200);
and U2287 (N_2287,N_2249,N_2210);
and U2288 (N_2288,N_2210,N_2232);
xnor U2289 (N_2289,N_2222,N_2206);
xor U2290 (N_2290,N_2220,N_2233);
and U2291 (N_2291,N_2203,N_2238);
nand U2292 (N_2292,N_2236,N_2227);
nor U2293 (N_2293,N_2220,N_2214);
xor U2294 (N_2294,N_2218,N_2214);
xnor U2295 (N_2295,N_2231,N_2224);
nor U2296 (N_2296,N_2200,N_2228);
nand U2297 (N_2297,N_2206,N_2245);
nand U2298 (N_2298,N_2218,N_2239);
or U2299 (N_2299,N_2238,N_2219);
xor U2300 (N_2300,N_2294,N_2284);
and U2301 (N_2301,N_2298,N_2292);
nand U2302 (N_2302,N_2285,N_2287);
or U2303 (N_2303,N_2279,N_2296);
xor U2304 (N_2304,N_2263,N_2266);
nand U2305 (N_2305,N_2261,N_2273);
nor U2306 (N_2306,N_2255,N_2270);
xor U2307 (N_2307,N_2299,N_2251);
or U2308 (N_2308,N_2276,N_2272);
and U2309 (N_2309,N_2280,N_2258);
or U2310 (N_2310,N_2271,N_2275);
nor U2311 (N_2311,N_2293,N_2253);
xor U2312 (N_2312,N_2281,N_2290);
or U2313 (N_2313,N_2297,N_2256);
or U2314 (N_2314,N_2250,N_2288);
nand U2315 (N_2315,N_2257,N_2262);
nand U2316 (N_2316,N_2274,N_2291);
or U2317 (N_2317,N_2260,N_2254);
and U2318 (N_2318,N_2265,N_2259);
nand U2319 (N_2319,N_2252,N_2268);
or U2320 (N_2320,N_2264,N_2282);
and U2321 (N_2321,N_2278,N_2267);
nor U2322 (N_2322,N_2283,N_2295);
nand U2323 (N_2323,N_2289,N_2277);
nand U2324 (N_2324,N_2286,N_2269);
and U2325 (N_2325,N_2275,N_2260);
and U2326 (N_2326,N_2276,N_2271);
nor U2327 (N_2327,N_2266,N_2283);
or U2328 (N_2328,N_2255,N_2289);
nor U2329 (N_2329,N_2262,N_2263);
xnor U2330 (N_2330,N_2274,N_2282);
nor U2331 (N_2331,N_2250,N_2299);
nor U2332 (N_2332,N_2268,N_2296);
nand U2333 (N_2333,N_2293,N_2288);
and U2334 (N_2334,N_2253,N_2267);
and U2335 (N_2335,N_2290,N_2271);
or U2336 (N_2336,N_2253,N_2269);
or U2337 (N_2337,N_2288,N_2252);
xnor U2338 (N_2338,N_2264,N_2293);
xor U2339 (N_2339,N_2284,N_2266);
and U2340 (N_2340,N_2273,N_2265);
and U2341 (N_2341,N_2251,N_2262);
or U2342 (N_2342,N_2264,N_2270);
xnor U2343 (N_2343,N_2273,N_2282);
nor U2344 (N_2344,N_2284,N_2283);
xor U2345 (N_2345,N_2284,N_2292);
or U2346 (N_2346,N_2274,N_2289);
nor U2347 (N_2347,N_2293,N_2285);
nand U2348 (N_2348,N_2299,N_2266);
nor U2349 (N_2349,N_2267,N_2287);
or U2350 (N_2350,N_2336,N_2318);
and U2351 (N_2351,N_2328,N_2330);
or U2352 (N_2352,N_2319,N_2332);
nand U2353 (N_2353,N_2302,N_2325);
xor U2354 (N_2354,N_2327,N_2317);
xor U2355 (N_2355,N_2315,N_2344);
xnor U2356 (N_2356,N_2304,N_2326);
and U2357 (N_2357,N_2335,N_2329);
xor U2358 (N_2358,N_2312,N_2337);
nor U2359 (N_2359,N_2320,N_2333);
nor U2360 (N_2360,N_2341,N_2306);
nand U2361 (N_2361,N_2347,N_2323);
xor U2362 (N_2362,N_2309,N_2331);
xnor U2363 (N_2363,N_2339,N_2343);
or U2364 (N_2364,N_2342,N_2349);
nand U2365 (N_2365,N_2316,N_2346);
or U2366 (N_2366,N_2322,N_2324);
nor U2367 (N_2367,N_2314,N_2321);
nor U2368 (N_2368,N_2305,N_2307);
nand U2369 (N_2369,N_2340,N_2311);
xnor U2370 (N_2370,N_2313,N_2338);
nand U2371 (N_2371,N_2310,N_2345);
xor U2372 (N_2372,N_2303,N_2300);
and U2373 (N_2373,N_2348,N_2301);
nand U2374 (N_2374,N_2308,N_2334);
or U2375 (N_2375,N_2317,N_2333);
or U2376 (N_2376,N_2329,N_2348);
and U2377 (N_2377,N_2349,N_2320);
xnor U2378 (N_2378,N_2349,N_2321);
xor U2379 (N_2379,N_2347,N_2336);
nor U2380 (N_2380,N_2343,N_2340);
nand U2381 (N_2381,N_2324,N_2331);
nand U2382 (N_2382,N_2319,N_2321);
nor U2383 (N_2383,N_2342,N_2313);
nand U2384 (N_2384,N_2318,N_2323);
nor U2385 (N_2385,N_2334,N_2303);
nand U2386 (N_2386,N_2317,N_2314);
nor U2387 (N_2387,N_2325,N_2315);
or U2388 (N_2388,N_2313,N_2330);
xor U2389 (N_2389,N_2342,N_2340);
and U2390 (N_2390,N_2322,N_2345);
nor U2391 (N_2391,N_2314,N_2337);
or U2392 (N_2392,N_2307,N_2314);
and U2393 (N_2393,N_2335,N_2327);
xor U2394 (N_2394,N_2308,N_2314);
nand U2395 (N_2395,N_2330,N_2336);
nand U2396 (N_2396,N_2349,N_2306);
nor U2397 (N_2397,N_2344,N_2310);
nor U2398 (N_2398,N_2320,N_2325);
xnor U2399 (N_2399,N_2306,N_2324);
nor U2400 (N_2400,N_2398,N_2374);
xnor U2401 (N_2401,N_2399,N_2364);
nand U2402 (N_2402,N_2389,N_2366);
xor U2403 (N_2403,N_2379,N_2353);
nand U2404 (N_2404,N_2357,N_2387);
nor U2405 (N_2405,N_2356,N_2397);
and U2406 (N_2406,N_2367,N_2361);
nand U2407 (N_2407,N_2362,N_2372);
and U2408 (N_2408,N_2376,N_2390);
xnor U2409 (N_2409,N_2385,N_2377);
nand U2410 (N_2410,N_2380,N_2368);
xnor U2411 (N_2411,N_2383,N_2378);
or U2412 (N_2412,N_2351,N_2392);
nor U2413 (N_2413,N_2354,N_2382);
or U2414 (N_2414,N_2375,N_2396);
xor U2415 (N_2415,N_2358,N_2371);
nand U2416 (N_2416,N_2388,N_2386);
or U2417 (N_2417,N_2350,N_2395);
and U2418 (N_2418,N_2391,N_2381);
or U2419 (N_2419,N_2369,N_2359);
xnor U2420 (N_2420,N_2373,N_2352);
nand U2421 (N_2421,N_2360,N_2394);
and U2422 (N_2422,N_2355,N_2370);
or U2423 (N_2423,N_2393,N_2365);
and U2424 (N_2424,N_2363,N_2384);
and U2425 (N_2425,N_2396,N_2360);
and U2426 (N_2426,N_2389,N_2380);
nand U2427 (N_2427,N_2372,N_2366);
nand U2428 (N_2428,N_2362,N_2350);
xor U2429 (N_2429,N_2375,N_2395);
xor U2430 (N_2430,N_2368,N_2363);
or U2431 (N_2431,N_2378,N_2384);
nor U2432 (N_2432,N_2388,N_2380);
and U2433 (N_2433,N_2361,N_2382);
and U2434 (N_2434,N_2398,N_2392);
nand U2435 (N_2435,N_2383,N_2362);
xnor U2436 (N_2436,N_2389,N_2354);
xor U2437 (N_2437,N_2353,N_2382);
xor U2438 (N_2438,N_2350,N_2392);
xnor U2439 (N_2439,N_2392,N_2354);
and U2440 (N_2440,N_2378,N_2370);
xor U2441 (N_2441,N_2356,N_2358);
xnor U2442 (N_2442,N_2362,N_2379);
and U2443 (N_2443,N_2352,N_2350);
xor U2444 (N_2444,N_2399,N_2385);
or U2445 (N_2445,N_2392,N_2363);
nor U2446 (N_2446,N_2361,N_2386);
or U2447 (N_2447,N_2359,N_2384);
nor U2448 (N_2448,N_2359,N_2385);
or U2449 (N_2449,N_2364,N_2354);
nor U2450 (N_2450,N_2447,N_2413);
nor U2451 (N_2451,N_2425,N_2407);
nand U2452 (N_2452,N_2434,N_2446);
xnor U2453 (N_2453,N_2412,N_2422);
and U2454 (N_2454,N_2420,N_2400);
xor U2455 (N_2455,N_2430,N_2445);
nand U2456 (N_2456,N_2411,N_2406);
and U2457 (N_2457,N_2416,N_2442);
and U2458 (N_2458,N_2432,N_2414);
nand U2459 (N_2459,N_2440,N_2418);
xnor U2460 (N_2460,N_2441,N_2424);
or U2461 (N_2461,N_2431,N_2437);
xnor U2462 (N_2462,N_2433,N_2405);
nand U2463 (N_2463,N_2449,N_2415);
and U2464 (N_2464,N_2438,N_2444);
and U2465 (N_2465,N_2436,N_2435);
xnor U2466 (N_2466,N_2404,N_2408);
nor U2467 (N_2467,N_2429,N_2419);
nor U2468 (N_2468,N_2403,N_2401);
and U2469 (N_2469,N_2402,N_2409);
and U2470 (N_2470,N_2410,N_2443);
nand U2471 (N_2471,N_2427,N_2439);
nand U2472 (N_2472,N_2426,N_2423);
nand U2473 (N_2473,N_2417,N_2428);
xor U2474 (N_2474,N_2421,N_2448);
xnor U2475 (N_2475,N_2443,N_2414);
and U2476 (N_2476,N_2424,N_2439);
and U2477 (N_2477,N_2415,N_2425);
and U2478 (N_2478,N_2439,N_2436);
and U2479 (N_2479,N_2413,N_2419);
nor U2480 (N_2480,N_2442,N_2407);
nor U2481 (N_2481,N_2439,N_2406);
xor U2482 (N_2482,N_2434,N_2408);
xor U2483 (N_2483,N_2422,N_2440);
or U2484 (N_2484,N_2422,N_2427);
xnor U2485 (N_2485,N_2445,N_2410);
nor U2486 (N_2486,N_2402,N_2446);
and U2487 (N_2487,N_2429,N_2436);
and U2488 (N_2488,N_2434,N_2417);
and U2489 (N_2489,N_2446,N_2407);
xor U2490 (N_2490,N_2425,N_2414);
xnor U2491 (N_2491,N_2437,N_2423);
or U2492 (N_2492,N_2434,N_2400);
or U2493 (N_2493,N_2413,N_2444);
and U2494 (N_2494,N_2428,N_2403);
nand U2495 (N_2495,N_2419,N_2409);
or U2496 (N_2496,N_2447,N_2429);
nand U2497 (N_2497,N_2402,N_2424);
or U2498 (N_2498,N_2419,N_2422);
nand U2499 (N_2499,N_2415,N_2421);
nor U2500 (N_2500,N_2464,N_2452);
xor U2501 (N_2501,N_2498,N_2454);
nor U2502 (N_2502,N_2470,N_2467);
nand U2503 (N_2503,N_2487,N_2473);
or U2504 (N_2504,N_2497,N_2475);
xor U2505 (N_2505,N_2469,N_2472);
nand U2506 (N_2506,N_2459,N_2485);
nand U2507 (N_2507,N_2474,N_2468);
nor U2508 (N_2508,N_2499,N_2457);
nor U2509 (N_2509,N_2471,N_2489);
xnor U2510 (N_2510,N_2491,N_2460);
nor U2511 (N_2511,N_2450,N_2483);
xnor U2512 (N_2512,N_2477,N_2453);
xnor U2513 (N_2513,N_2482,N_2461);
xor U2514 (N_2514,N_2481,N_2476);
nor U2515 (N_2515,N_2490,N_2458);
and U2516 (N_2516,N_2451,N_2456);
nor U2517 (N_2517,N_2496,N_2492);
xor U2518 (N_2518,N_2479,N_2486);
or U2519 (N_2519,N_2493,N_2455);
xor U2520 (N_2520,N_2465,N_2488);
xnor U2521 (N_2521,N_2462,N_2478);
or U2522 (N_2522,N_2494,N_2466);
xnor U2523 (N_2523,N_2484,N_2463);
xor U2524 (N_2524,N_2495,N_2480);
nor U2525 (N_2525,N_2496,N_2488);
nor U2526 (N_2526,N_2481,N_2472);
or U2527 (N_2527,N_2473,N_2498);
or U2528 (N_2528,N_2491,N_2463);
nand U2529 (N_2529,N_2481,N_2499);
nand U2530 (N_2530,N_2456,N_2476);
or U2531 (N_2531,N_2450,N_2484);
and U2532 (N_2532,N_2471,N_2452);
xnor U2533 (N_2533,N_2499,N_2453);
xnor U2534 (N_2534,N_2475,N_2489);
and U2535 (N_2535,N_2478,N_2488);
or U2536 (N_2536,N_2479,N_2459);
or U2537 (N_2537,N_2497,N_2450);
and U2538 (N_2538,N_2466,N_2454);
nand U2539 (N_2539,N_2493,N_2482);
and U2540 (N_2540,N_2461,N_2497);
nor U2541 (N_2541,N_2486,N_2469);
or U2542 (N_2542,N_2465,N_2497);
xnor U2543 (N_2543,N_2491,N_2458);
and U2544 (N_2544,N_2488,N_2457);
nor U2545 (N_2545,N_2492,N_2451);
nor U2546 (N_2546,N_2461,N_2493);
nor U2547 (N_2547,N_2455,N_2465);
nand U2548 (N_2548,N_2495,N_2488);
nand U2549 (N_2549,N_2472,N_2464);
and U2550 (N_2550,N_2534,N_2516);
or U2551 (N_2551,N_2530,N_2524);
and U2552 (N_2552,N_2541,N_2535);
nand U2553 (N_2553,N_2544,N_2543);
and U2554 (N_2554,N_2515,N_2528);
or U2555 (N_2555,N_2500,N_2521);
nor U2556 (N_2556,N_2548,N_2532);
nand U2557 (N_2557,N_2540,N_2504);
or U2558 (N_2558,N_2542,N_2526);
nor U2559 (N_2559,N_2546,N_2536);
or U2560 (N_2560,N_2501,N_2510);
and U2561 (N_2561,N_2511,N_2509);
xnor U2562 (N_2562,N_2529,N_2531);
and U2563 (N_2563,N_2503,N_2512);
and U2564 (N_2564,N_2549,N_2523);
nor U2565 (N_2565,N_2520,N_2513);
nor U2566 (N_2566,N_2517,N_2539);
nor U2567 (N_2567,N_2518,N_2538);
nor U2568 (N_2568,N_2506,N_2508);
and U2569 (N_2569,N_2547,N_2507);
nor U2570 (N_2570,N_2522,N_2533);
and U2571 (N_2571,N_2525,N_2527);
nor U2572 (N_2572,N_2537,N_2505);
and U2573 (N_2573,N_2514,N_2545);
xnor U2574 (N_2574,N_2502,N_2519);
nor U2575 (N_2575,N_2543,N_2535);
xor U2576 (N_2576,N_2511,N_2531);
nor U2577 (N_2577,N_2514,N_2531);
or U2578 (N_2578,N_2528,N_2533);
xnor U2579 (N_2579,N_2502,N_2524);
or U2580 (N_2580,N_2545,N_2511);
and U2581 (N_2581,N_2547,N_2549);
xnor U2582 (N_2582,N_2524,N_2515);
nor U2583 (N_2583,N_2507,N_2511);
or U2584 (N_2584,N_2533,N_2547);
nand U2585 (N_2585,N_2536,N_2541);
nor U2586 (N_2586,N_2539,N_2510);
nor U2587 (N_2587,N_2541,N_2510);
nor U2588 (N_2588,N_2547,N_2541);
and U2589 (N_2589,N_2525,N_2523);
and U2590 (N_2590,N_2509,N_2512);
or U2591 (N_2591,N_2545,N_2526);
or U2592 (N_2592,N_2531,N_2501);
or U2593 (N_2593,N_2504,N_2547);
or U2594 (N_2594,N_2515,N_2536);
nand U2595 (N_2595,N_2549,N_2504);
nand U2596 (N_2596,N_2544,N_2527);
or U2597 (N_2597,N_2544,N_2528);
or U2598 (N_2598,N_2513,N_2549);
nor U2599 (N_2599,N_2527,N_2517);
xnor U2600 (N_2600,N_2567,N_2559);
or U2601 (N_2601,N_2585,N_2595);
xor U2602 (N_2602,N_2577,N_2575);
xnor U2603 (N_2603,N_2554,N_2573);
xor U2604 (N_2604,N_2586,N_2553);
nor U2605 (N_2605,N_2561,N_2564);
or U2606 (N_2606,N_2588,N_2583);
nand U2607 (N_2607,N_2598,N_2580);
nand U2608 (N_2608,N_2557,N_2572);
and U2609 (N_2609,N_2599,N_2584);
xnor U2610 (N_2610,N_2594,N_2568);
xor U2611 (N_2611,N_2596,N_2562);
xor U2612 (N_2612,N_2551,N_2556);
xnor U2613 (N_2613,N_2571,N_2593);
nor U2614 (N_2614,N_2550,N_2578);
nor U2615 (N_2615,N_2597,N_2589);
xor U2616 (N_2616,N_2579,N_2574);
xnor U2617 (N_2617,N_2576,N_2563);
nor U2618 (N_2618,N_2570,N_2591);
or U2619 (N_2619,N_2569,N_2552);
xnor U2620 (N_2620,N_2560,N_2592);
or U2621 (N_2621,N_2566,N_2558);
xnor U2622 (N_2622,N_2582,N_2565);
nand U2623 (N_2623,N_2590,N_2587);
xnor U2624 (N_2624,N_2555,N_2581);
and U2625 (N_2625,N_2573,N_2587);
nand U2626 (N_2626,N_2564,N_2557);
or U2627 (N_2627,N_2585,N_2556);
xnor U2628 (N_2628,N_2590,N_2598);
nand U2629 (N_2629,N_2575,N_2594);
and U2630 (N_2630,N_2591,N_2556);
nand U2631 (N_2631,N_2599,N_2585);
nor U2632 (N_2632,N_2598,N_2577);
and U2633 (N_2633,N_2566,N_2594);
nor U2634 (N_2634,N_2588,N_2552);
nor U2635 (N_2635,N_2599,N_2595);
nor U2636 (N_2636,N_2587,N_2567);
nor U2637 (N_2637,N_2558,N_2595);
or U2638 (N_2638,N_2569,N_2572);
nor U2639 (N_2639,N_2584,N_2598);
nand U2640 (N_2640,N_2588,N_2595);
nand U2641 (N_2641,N_2592,N_2551);
nand U2642 (N_2642,N_2562,N_2553);
and U2643 (N_2643,N_2556,N_2589);
nand U2644 (N_2644,N_2557,N_2580);
nor U2645 (N_2645,N_2592,N_2583);
and U2646 (N_2646,N_2565,N_2563);
nand U2647 (N_2647,N_2587,N_2562);
nand U2648 (N_2648,N_2573,N_2574);
xnor U2649 (N_2649,N_2561,N_2560);
nor U2650 (N_2650,N_2641,N_2644);
nand U2651 (N_2651,N_2637,N_2649);
nand U2652 (N_2652,N_2601,N_2636);
nand U2653 (N_2653,N_2638,N_2602);
nor U2654 (N_2654,N_2600,N_2609);
and U2655 (N_2655,N_2645,N_2616);
and U2656 (N_2656,N_2608,N_2634);
xor U2657 (N_2657,N_2607,N_2631);
and U2658 (N_2658,N_2633,N_2627);
xnor U2659 (N_2659,N_2626,N_2619);
xnor U2660 (N_2660,N_2611,N_2606);
nor U2661 (N_2661,N_2603,N_2622);
xor U2662 (N_2662,N_2614,N_2646);
and U2663 (N_2663,N_2648,N_2618);
xnor U2664 (N_2664,N_2620,N_2604);
or U2665 (N_2665,N_2630,N_2615);
nand U2666 (N_2666,N_2612,N_2610);
or U2667 (N_2667,N_2635,N_2639);
nand U2668 (N_2668,N_2624,N_2621);
and U2669 (N_2669,N_2605,N_2632);
nor U2670 (N_2670,N_2628,N_2613);
or U2671 (N_2671,N_2629,N_2625);
or U2672 (N_2672,N_2617,N_2640);
xnor U2673 (N_2673,N_2643,N_2623);
and U2674 (N_2674,N_2642,N_2647);
or U2675 (N_2675,N_2624,N_2634);
nor U2676 (N_2676,N_2644,N_2610);
and U2677 (N_2677,N_2618,N_2640);
or U2678 (N_2678,N_2631,N_2600);
xor U2679 (N_2679,N_2613,N_2635);
and U2680 (N_2680,N_2647,N_2644);
xnor U2681 (N_2681,N_2613,N_2629);
and U2682 (N_2682,N_2642,N_2613);
nor U2683 (N_2683,N_2649,N_2602);
nand U2684 (N_2684,N_2642,N_2637);
xnor U2685 (N_2685,N_2618,N_2630);
nand U2686 (N_2686,N_2632,N_2614);
nand U2687 (N_2687,N_2611,N_2635);
and U2688 (N_2688,N_2631,N_2628);
or U2689 (N_2689,N_2609,N_2642);
and U2690 (N_2690,N_2645,N_2637);
and U2691 (N_2691,N_2608,N_2633);
nor U2692 (N_2692,N_2623,N_2628);
xor U2693 (N_2693,N_2633,N_2603);
xnor U2694 (N_2694,N_2631,N_2608);
and U2695 (N_2695,N_2626,N_2641);
nor U2696 (N_2696,N_2635,N_2619);
nor U2697 (N_2697,N_2630,N_2643);
or U2698 (N_2698,N_2623,N_2616);
xor U2699 (N_2699,N_2640,N_2648);
and U2700 (N_2700,N_2685,N_2659);
and U2701 (N_2701,N_2694,N_2653);
xor U2702 (N_2702,N_2660,N_2654);
and U2703 (N_2703,N_2667,N_2669);
nand U2704 (N_2704,N_2693,N_2672);
nor U2705 (N_2705,N_2697,N_2688);
and U2706 (N_2706,N_2695,N_2690);
nand U2707 (N_2707,N_2692,N_2668);
nor U2708 (N_2708,N_2691,N_2663);
and U2709 (N_2709,N_2658,N_2673);
nand U2710 (N_2710,N_2686,N_2679);
or U2711 (N_2711,N_2670,N_2656);
or U2712 (N_2712,N_2662,N_2696);
nand U2713 (N_2713,N_2681,N_2689);
xor U2714 (N_2714,N_2657,N_2665);
and U2715 (N_2715,N_2678,N_2683);
and U2716 (N_2716,N_2684,N_2664);
or U2717 (N_2717,N_2655,N_2676);
xnor U2718 (N_2718,N_2699,N_2677);
or U2719 (N_2719,N_2698,N_2674);
nor U2720 (N_2720,N_2650,N_2687);
and U2721 (N_2721,N_2671,N_2652);
or U2722 (N_2722,N_2661,N_2666);
nand U2723 (N_2723,N_2651,N_2675);
nand U2724 (N_2724,N_2680,N_2682);
and U2725 (N_2725,N_2650,N_2670);
nand U2726 (N_2726,N_2697,N_2686);
or U2727 (N_2727,N_2676,N_2658);
or U2728 (N_2728,N_2661,N_2683);
or U2729 (N_2729,N_2658,N_2651);
and U2730 (N_2730,N_2670,N_2669);
nor U2731 (N_2731,N_2695,N_2697);
xnor U2732 (N_2732,N_2686,N_2675);
and U2733 (N_2733,N_2685,N_2654);
nand U2734 (N_2734,N_2661,N_2660);
nand U2735 (N_2735,N_2676,N_2660);
nand U2736 (N_2736,N_2695,N_2658);
nor U2737 (N_2737,N_2667,N_2665);
or U2738 (N_2738,N_2659,N_2662);
nor U2739 (N_2739,N_2695,N_2687);
and U2740 (N_2740,N_2685,N_2696);
or U2741 (N_2741,N_2661,N_2689);
xor U2742 (N_2742,N_2684,N_2666);
or U2743 (N_2743,N_2671,N_2685);
or U2744 (N_2744,N_2687,N_2662);
xnor U2745 (N_2745,N_2698,N_2667);
or U2746 (N_2746,N_2654,N_2664);
and U2747 (N_2747,N_2674,N_2692);
and U2748 (N_2748,N_2668,N_2698);
and U2749 (N_2749,N_2653,N_2670);
and U2750 (N_2750,N_2705,N_2717);
nor U2751 (N_2751,N_2708,N_2741);
nor U2752 (N_2752,N_2719,N_2704);
xor U2753 (N_2753,N_2711,N_2718);
xnor U2754 (N_2754,N_2714,N_2710);
nor U2755 (N_2755,N_2736,N_2720);
or U2756 (N_2756,N_2727,N_2735);
and U2757 (N_2757,N_2746,N_2706);
and U2758 (N_2758,N_2728,N_2729);
or U2759 (N_2759,N_2738,N_2716);
and U2760 (N_2760,N_2749,N_2702);
nor U2761 (N_2761,N_2739,N_2703);
nor U2762 (N_2762,N_2747,N_2737);
nand U2763 (N_2763,N_2722,N_2743);
and U2764 (N_2764,N_2748,N_2732);
nor U2765 (N_2765,N_2745,N_2712);
nor U2766 (N_2766,N_2730,N_2726);
and U2767 (N_2767,N_2744,N_2724);
nor U2768 (N_2768,N_2715,N_2709);
xnor U2769 (N_2769,N_2734,N_2701);
or U2770 (N_2770,N_2733,N_2707);
nor U2771 (N_2771,N_2731,N_2725);
nand U2772 (N_2772,N_2700,N_2713);
nor U2773 (N_2773,N_2723,N_2742);
or U2774 (N_2774,N_2740,N_2721);
xnor U2775 (N_2775,N_2747,N_2725);
xor U2776 (N_2776,N_2717,N_2730);
or U2777 (N_2777,N_2724,N_2708);
and U2778 (N_2778,N_2747,N_2738);
or U2779 (N_2779,N_2711,N_2737);
nand U2780 (N_2780,N_2735,N_2709);
nor U2781 (N_2781,N_2704,N_2703);
nor U2782 (N_2782,N_2720,N_2734);
and U2783 (N_2783,N_2749,N_2747);
nand U2784 (N_2784,N_2746,N_2732);
nand U2785 (N_2785,N_2743,N_2714);
xnor U2786 (N_2786,N_2702,N_2716);
and U2787 (N_2787,N_2708,N_2726);
and U2788 (N_2788,N_2721,N_2724);
and U2789 (N_2789,N_2717,N_2728);
xor U2790 (N_2790,N_2736,N_2708);
and U2791 (N_2791,N_2730,N_2710);
nor U2792 (N_2792,N_2749,N_2743);
xnor U2793 (N_2793,N_2741,N_2738);
nor U2794 (N_2794,N_2735,N_2728);
nor U2795 (N_2795,N_2719,N_2737);
or U2796 (N_2796,N_2715,N_2739);
nor U2797 (N_2797,N_2748,N_2717);
and U2798 (N_2798,N_2738,N_2734);
nand U2799 (N_2799,N_2722,N_2735);
or U2800 (N_2800,N_2799,N_2753);
and U2801 (N_2801,N_2764,N_2758);
and U2802 (N_2802,N_2783,N_2777);
nor U2803 (N_2803,N_2778,N_2773);
nand U2804 (N_2804,N_2760,N_2772);
or U2805 (N_2805,N_2754,N_2796);
or U2806 (N_2806,N_2791,N_2756);
nand U2807 (N_2807,N_2781,N_2780);
xnor U2808 (N_2808,N_2788,N_2793);
nor U2809 (N_2809,N_2798,N_2759);
nor U2810 (N_2810,N_2782,N_2785);
and U2811 (N_2811,N_2792,N_2775);
nor U2812 (N_2812,N_2768,N_2789);
xor U2813 (N_2813,N_2784,N_2769);
xor U2814 (N_2814,N_2750,N_2795);
nand U2815 (N_2815,N_2757,N_2755);
or U2816 (N_2816,N_2761,N_2794);
nor U2817 (N_2817,N_2779,N_2774);
and U2818 (N_2818,N_2776,N_2762);
xor U2819 (N_2819,N_2790,N_2770);
nor U2820 (N_2820,N_2763,N_2765);
and U2821 (N_2821,N_2787,N_2766);
xor U2822 (N_2822,N_2752,N_2767);
nor U2823 (N_2823,N_2771,N_2786);
nand U2824 (N_2824,N_2797,N_2751);
nor U2825 (N_2825,N_2787,N_2798);
and U2826 (N_2826,N_2793,N_2767);
nor U2827 (N_2827,N_2758,N_2762);
or U2828 (N_2828,N_2787,N_2772);
nor U2829 (N_2829,N_2779,N_2780);
and U2830 (N_2830,N_2765,N_2783);
or U2831 (N_2831,N_2777,N_2790);
and U2832 (N_2832,N_2752,N_2797);
xor U2833 (N_2833,N_2776,N_2787);
nand U2834 (N_2834,N_2793,N_2773);
nor U2835 (N_2835,N_2774,N_2752);
xnor U2836 (N_2836,N_2796,N_2759);
nand U2837 (N_2837,N_2785,N_2761);
and U2838 (N_2838,N_2778,N_2783);
and U2839 (N_2839,N_2785,N_2750);
xor U2840 (N_2840,N_2790,N_2798);
nor U2841 (N_2841,N_2751,N_2788);
and U2842 (N_2842,N_2779,N_2761);
xnor U2843 (N_2843,N_2778,N_2780);
and U2844 (N_2844,N_2776,N_2778);
or U2845 (N_2845,N_2799,N_2779);
or U2846 (N_2846,N_2759,N_2791);
and U2847 (N_2847,N_2765,N_2761);
nand U2848 (N_2848,N_2755,N_2761);
or U2849 (N_2849,N_2751,N_2789);
or U2850 (N_2850,N_2825,N_2801);
nand U2851 (N_2851,N_2805,N_2830);
nor U2852 (N_2852,N_2810,N_2838);
and U2853 (N_2853,N_2816,N_2809);
nor U2854 (N_2854,N_2824,N_2821);
and U2855 (N_2855,N_2849,N_2840);
xor U2856 (N_2856,N_2826,N_2848);
and U2857 (N_2857,N_2820,N_2832);
nand U2858 (N_2858,N_2800,N_2845);
xnor U2859 (N_2859,N_2815,N_2807);
nor U2860 (N_2860,N_2836,N_2833);
xnor U2861 (N_2861,N_2827,N_2834);
nor U2862 (N_2862,N_2843,N_2839);
and U2863 (N_2863,N_2813,N_2837);
nor U2864 (N_2864,N_2812,N_2808);
or U2865 (N_2865,N_2802,N_2844);
xnor U2866 (N_2866,N_2829,N_2822);
nand U2867 (N_2867,N_2817,N_2841);
or U2868 (N_2868,N_2804,N_2811);
nand U2869 (N_2869,N_2831,N_2803);
or U2870 (N_2870,N_2835,N_2828);
or U2871 (N_2871,N_2806,N_2814);
nand U2872 (N_2872,N_2823,N_2846);
or U2873 (N_2873,N_2842,N_2818);
or U2874 (N_2874,N_2847,N_2819);
and U2875 (N_2875,N_2832,N_2837);
or U2876 (N_2876,N_2849,N_2838);
xor U2877 (N_2877,N_2827,N_2829);
nand U2878 (N_2878,N_2823,N_2842);
or U2879 (N_2879,N_2834,N_2844);
or U2880 (N_2880,N_2844,N_2832);
nand U2881 (N_2881,N_2808,N_2834);
and U2882 (N_2882,N_2834,N_2836);
xnor U2883 (N_2883,N_2816,N_2808);
xor U2884 (N_2884,N_2808,N_2825);
nand U2885 (N_2885,N_2833,N_2847);
or U2886 (N_2886,N_2833,N_2813);
nor U2887 (N_2887,N_2837,N_2831);
or U2888 (N_2888,N_2844,N_2823);
and U2889 (N_2889,N_2830,N_2847);
and U2890 (N_2890,N_2807,N_2837);
or U2891 (N_2891,N_2820,N_2826);
and U2892 (N_2892,N_2819,N_2835);
nand U2893 (N_2893,N_2807,N_2825);
xnor U2894 (N_2894,N_2804,N_2812);
xor U2895 (N_2895,N_2845,N_2825);
nand U2896 (N_2896,N_2810,N_2807);
and U2897 (N_2897,N_2817,N_2822);
xor U2898 (N_2898,N_2846,N_2812);
nand U2899 (N_2899,N_2844,N_2822);
or U2900 (N_2900,N_2857,N_2865);
and U2901 (N_2901,N_2852,N_2895);
and U2902 (N_2902,N_2871,N_2898);
nor U2903 (N_2903,N_2850,N_2873);
nand U2904 (N_2904,N_2867,N_2899);
nor U2905 (N_2905,N_2861,N_2879);
nor U2906 (N_2906,N_2863,N_2881);
nor U2907 (N_2907,N_2859,N_2856);
and U2908 (N_2908,N_2877,N_2892);
xor U2909 (N_2909,N_2894,N_2897);
nand U2910 (N_2910,N_2885,N_2882);
or U2911 (N_2911,N_2858,N_2880);
or U2912 (N_2912,N_2887,N_2872);
nand U2913 (N_2913,N_2874,N_2884);
nand U2914 (N_2914,N_2890,N_2883);
and U2915 (N_2915,N_2864,N_2891);
nor U2916 (N_2916,N_2868,N_2889);
xor U2917 (N_2917,N_2876,N_2878);
or U2918 (N_2918,N_2860,N_2855);
nand U2919 (N_2919,N_2862,N_2853);
and U2920 (N_2920,N_2888,N_2893);
nand U2921 (N_2921,N_2869,N_2896);
or U2922 (N_2922,N_2854,N_2875);
xor U2923 (N_2923,N_2870,N_2851);
nand U2924 (N_2924,N_2886,N_2866);
nor U2925 (N_2925,N_2887,N_2896);
nand U2926 (N_2926,N_2869,N_2854);
nor U2927 (N_2927,N_2851,N_2863);
xor U2928 (N_2928,N_2889,N_2881);
xor U2929 (N_2929,N_2864,N_2850);
or U2930 (N_2930,N_2898,N_2889);
and U2931 (N_2931,N_2869,N_2871);
xnor U2932 (N_2932,N_2871,N_2853);
or U2933 (N_2933,N_2868,N_2852);
nand U2934 (N_2934,N_2866,N_2889);
and U2935 (N_2935,N_2862,N_2863);
nand U2936 (N_2936,N_2868,N_2880);
nand U2937 (N_2937,N_2859,N_2854);
or U2938 (N_2938,N_2873,N_2871);
and U2939 (N_2939,N_2870,N_2886);
or U2940 (N_2940,N_2880,N_2859);
nor U2941 (N_2941,N_2892,N_2875);
nand U2942 (N_2942,N_2893,N_2857);
and U2943 (N_2943,N_2888,N_2880);
or U2944 (N_2944,N_2860,N_2875);
and U2945 (N_2945,N_2850,N_2863);
nor U2946 (N_2946,N_2873,N_2870);
or U2947 (N_2947,N_2866,N_2852);
xnor U2948 (N_2948,N_2887,N_2867);
nand U2949 (N_2949,N_2890,N_2895);
nor U2950 (N_2950,N_2926,N_2947);
nor U2951 (N_2951,N_2902,N_2928);
and U2952 (N_2952,N_2930,N_2906);
xor U2953 (N_2953,N_2921,N_2922);
nor U2954 (N_2954,N_2923,N_2944);
nor U2955 (N_2955,N_2912,N_2901);
or U2956 (N_2956,N_2911,N_2910);
nand U2957 (N_2957,N_2909,N_2933);
or U2958 (N_2958,N_2945,N_2939);
nor U2959 (N_2959,N_2946,N_2924);
or U2960 (N_2960,N_2934,N_2915);
nand U2961 (N_2961,N_2935,N_2929);
xor U2962 (N_2962,N_2938,N_2948);
xor U2963 (N_2963,N_2932,N_2907);
or U2964 (N_2964,N_2918,N_2900);
xor U2965 (N_2965,N_2905,N_2943);
nor U2966 (N_2966,N_2904,N_2940);
and U2967 (N_2967,N_2931,N_2949);
or U2968 (N_2968,N_2925,N_2916);
xnor U2969 (N_2969,N_2903,N_2936);
xnor U2970 (N_2970,N_2913,N_2942);
nand U2971 (N_2971,N_2914,N_2927);
nand U2972 (N_2972,N_2908,N_2917);
nand U2973 (N_2973,N_2919,N_2941);
and U2974 (N_2974,N_2937,N_2920);
xnor U2975 (N_2975,N_2937,N_2947);
or U2976 (N_2976,N_2945,N_2944);
nand U2977 (N_2977,N_2936,N_2914);
nor U2978 (N_2978,N_2907,N_2915);
nor U2979 (N_2979,N_2902,N_2935);
or U2980 (N_2980,N_2904,N_2942);
nor U2981 (N_2981,N_2937,N_2915);
nor U2982 (N_2982,N_2947,N_2908);
nor U2983 (N_2983,N_2941,N_2909);
and U2984 (N_2984,N_2929,N_2924);
or U2985 (N_2985,N_2930,N_2939);
and U2986 (N_2986,N_2939,N_2909);
nand U2987 (N_2987,N_2915,N_2927);
xnor U2988 (N_2988,N_2905,N_2908);
or U2989 (N_2989,N_2945,N_2946);
and U2990 (N_2990,N_2908,N_2926);
and U2991 (N_2991,N_2911,N_2907);
or U2992 (N_2992,N_2930,N_2931);
and U2993 (N_2993,N_2901,N_2940);
and U2994 (N_2994,N_2936,N_2935);
xor U2995 (N_2995,N_2915,N_2933);
and U2996 (N_2996,N_2944,N_2947);
nand U2997 (N_2997,N_2940,N_2918);
xnor U2998 (N_2998,N_2902,N_2919);
xnor U2999 (N_2999,N_2918,N_2919);
nor UO_0 (O_0,N_2973,N_2954);
nand UO_1 (O_1,N_2965,N_2967);
or UO_2 (O_2,N_2970,N_2950);
xnor UO_3 (O_3,N_2991,N_2996);
and UO_4 (O_4,N_2977,N_2953);
nand UO_5 (O_5,N_2980,N_2975);
nor UO_6 (O_6,N_2957,N_2987);
and UO_7 (O_7,N_2961,N_2968);
and UO_8 (O_8,N_2998,N_2969);
nand UO_9 (O_9,N_2972,N_2960);
and UO_10 (O_10,N_2955,N_2962);
nand UO_11 (O_11,N_2956,N_2958);
or UO_12 (O_12,N_2963,N_2990);
nor UO_13 (O_13,N_2993,N_2982);
or UO_14 (O_14,N_2994,N_2985);
nand UO_15 (O_15,N_2978,N_2959);
xor UO_16 (O_16,N_2997,N_2983);
or UO_17 (O_17,N_2966,N_2951);
nor UO_18 (O_18,N_2999,N_2979);
nand UO_19 (O_19,N_2971,N_2988);
and UO_20 (O_20,N_2992,N_2984);
or UO_21 (O_21,N_2986,N_2976);
nor UO_22 (O_22,N_2952,N_2964);
nand UO_23 (O_23,N_2981,N_2974);
nor UO_24 (O_24,N_2995,N_2989);
nand UO_25 (O_25,N_2996,N_2974);
nand UO_26 (O_26,N_2987,N_2966);
xor UO_27 (O_27,N_2977,N_2987);
nand UO_28 (O_28,N_2982,N_2954);
xor UO_29 (O_29,N_2957,N_2999);
nor UO_30 (O_30,N_2992,N_2988);
nor UO_31 (O_31,N_2993,N_2989);
or UO_32 (O_32,N_2986,N_2959);
xor UO_33 (O_33,N_2979,N_2965);
and UO_34 (O_34,N_2983,N_2971);
nor UO_35 (O_35,N_2967,N_2987);
nand UO_36 (O_36,N_2977,N_2997);
xor UO_37 (O_37,N_2999,N_2958);
nor UO_38 (O_38,N_2955,N_2997);
or UO_39 (O_39,N_2959,N_2970);
xor UO_40 (O_40,N_2980,N_2988);
or UO_41 (O_41,N_2958,N_2960);
or UO_42 (O_42,N_2950,N_2987);
xor UO_43 (O_43,N_2968,N_2977);
nor UO_44 (O_44,N_2994,N_2968);
or UO_45 (O_45,N_2955,N_2992);
or UO_46 (O_46,N_2997,N_2961);
nand UO_47 (O_47,N_2952,N_2985);
or UO_48 (O_48,N_2997,N_2950);
nor UO_49 (O_49,N_2969,N_2990);
or UO_50 (O_50,N_2989,N_2976);
xor UO_51 (O_51,N_2971,N_2982);
xnor UO_52 (O_52,N_2975,N_2997);
nand UO_53 (O_53,N_2992,N_2986);
nor UO_54 (O_54,N_2970,N_2979);
and UO_55 (O_55,N_2971,N_2978);
xnor UO_56 (O_56,N_2998,N_2954);
and UO_57 (O_57,N_2985,N_2960);
nand UO_58 (O_58,N_2993,N_2990);
xnor UO_59 (O_59,N_2998,N_2974);
nor UO_60 (O_60,N_2950,N_2985);
or UO_61 (O_61,N_2971,N_2990);
and UO_62 (O_62,N_2959,N_2963);
xnor UO_63 (O_63,N_2996,N_2988);
xor UO_64 (O_64,N_2960,N_2976);
nor UO_65 (O_65,N_2987,N_2959);
or UO_66 (O_66,N_2984,N_2969);
xnor UO_67 (O_67,N_2957,N_2965);
nor UO_68 (O_68,N_2965,N_2990);
or UO_69 (O_69,N_2988,N_2989);
or UO_70 (O_70,N_2952,N_2992);
or UO_71 (O_71,N_2989,N_2970);
nand UO_72 (O_72,N_2951,N_2978);
or UO_73 (O_73,N_2951,N_2954);
or UO_74 (O_74,N_2995,N_2955);
nand UO_75 (O_75,N_2974,N_2966);
nor UO_76 (O_76,N_2978,N_2985);
nor UO_77 (O_77,N_2999,N_2970);
xnor UO_78 (O_78,N_2983,N_2961);
xnor UO_79 (O_79,N_2988,N_2959);
xor UO_80 (O_80,N_2985,N_2996);
xnor UO_81 (O_81,N_2955,N_2950);
and UO_82 (O_82,N_2999,N_2974);
and UO_83 (O_83,N_2987,N_2999);
nor UO_84 (O_84,N_2955,N_2972);
nor UO_85 (O_85,N_2976,N_2953);
nand UO_86 (O_86,N_2989,N_2972);
and UO_87 (O_87,N_2994,N_2982);
and UO_88 (O_88,N_2976,N_2969);
nor UO_89 (O_89,N_2985,N_2968);
nand UO_90 (O_90,N_2969,N_2979);
and UO_91 (O_91,N_2953,N_2969);
nor UO_92 (O_92,N_2978,N_2980);
nand UO_93 (O_93,N_2951,N_2970);
xnor UO_94 (O_94,N_2962,N_2974);
or UO_95 (O_95,N_2999,N_2971);
nor UO_96 (O_96,N_2982,N_2957);
and UO_97 (O_97,N_2996,N_2978);
nand UO_98 (O_98,N_2964,N_2996);
nand UO_99 (O_99,N_2976,N_2988);
and UO_100 (O_100,N_2957,N_2953);
xor UO_101 (O_101,N_2956,N_2977);
and UO_102 (O_102,N_2953,N_2972);
and UO_103 (O_103,N_2954,N_2961);
or UO_104 (O_104,N_2958,N_2995);
or UO_105 (O_105,N_2964,N_2999);
or UO_106 (O_106,N_2956,N_2998);
and UO_107 (O_107,N_2969,N_2978);
or UO_108 (O_108,N_2999,N_2973);
and UO_109 (O_109,N_2971,N_2953);
nor UO_110 (O_110,N_2967,N_2956);
nor UO_111 (O_111,N_2991,N_2997);
nor UO_112 (O_112,N_2989,N_2966);
and UO_113 (O_113,N_2953,N_2970);
xnor UO_114 (O_114,N_2988,N_2968);
and UO_115 (O_115,N_2982,N_2966);
and UO_116 (O_116,N_2969,N_2973);
or UO_117 (O_117,N_2998,N_2960);
nor UO_118 (O_118,N_2973,N_2961);
xor UO_119 (O_119,N_2990,N_2956);
nor UO_120 (O_120,N_2974,N_2976);
or UO_121 (O_121,N_2982,N_2998);
nor UO_122 (O_122,N_2956,N_2999);
nor UO_123 (O_123,N_2969,N_2963);
nand UO_124 (O_124,N_2988,N_2958);
nor UO_125 (O_125,N_2984,N_2986);
nand UO_126 (O_126,N_2966,N_2984);
and UO_127 (O_127,N_2962,N_2990);
nand UO_128 (O_128,N_2985,N_2976);
or UO_129 (O_129,N_2999,N_2954);
xnor UO_130 (O_130,N_2978,N_2990);
nand UO_131 (O_131,N_2994,N_2977);
or UO_132 (O_132,N_2993,N_2997);
nor UO_133 (O_133,N_2957,N_2986);
nor UO_134 (O_134,N_2979,N_2956);
and UO_135 (O_135,N_2975,N_2968);
or UO_136 (O_136,N_2986,N_2956);
xor UO_137 (O_137,N_2980,N_2958);
or UO_138 (O_138,N_2976,N_2959);
nor UO_139 (O_139,N_2961,N_2956);
nand UO_140 (O_140,N_2955,N_2980);
or UO_141 (O_141,N_2951,N_2987);
xor UO_142 (O_142,N_2998,N_2951);
nor UO_143 (O_143,N_2986,N_2967);
or UO_144 (O_144,N_2951,N_2986);
xnor UO_145 (O_145,N_2950,N_2973);
nor UO_146 (O_146,N_2972,N_2984);
xnor UO_147 (O_147,N_2960,N_2964);
or UO_148 (O_148,N_2978,N_2963);
nand UO_149 (O_149,N_2970,N_2973);
or UO_150 (O_150,N_2951,N_2957);
nor UO_151 (O_151,N_2986,N_2982);
and UO_152 (O_152,N_2971,N_2979);
nor UO_153 (O_153,N_2958,N_2952);
or UO_154 (O_154,N_2950,N_2980);
nand UO_155 (O_155,N_2992,N_2981);
nand UO_156 (O_156,N_2989,N_2992);
or UO_157 (O_157,N_2992,N_2950);
or UO_158 (O_158,N_2994,N_2974);
nand UO_159 (O_159,N_2989,N_2999);
or UO_160 (O_160,N_2996,N_2973);
and UO_161 (O_161,N_2991,N_2994);
xor UO_162 (O_162,N_2993,N_2992);
nor UO_163 (O_163,N_2959,N_2980);
and UO_164 (O_164,N_2954,N_2994);
nor UO_165 (O_165,N_2962,N_2982);
or UO_166 (O_166,N_2962,N_2995);
xnor UO_167 (O_167,N_2971,N_2964);
and UO_168 (O_168,N_2983,N_2974);
xnor UO_169 (O_169,N_2988,N_2974);
nand UO_170 (O_170,N_2964,N_2951);
nand UO_171 (O_171,N_2959,N_2974);
xnor UO_172 (O_172,N_2957,N_2997);
nand UO_173 (O_173,N_2967,N_2950);
nand UO_174 (O_174,N_2964,N_2994);
and UO_175 (O_175,N_2986,N_2999);
nand UO_176 (O_176,N_2987,N_2983);
or UO_177 (O_177,N_2991,N_2988);
nand UO_178 (O_178,N_2958,N_2982);
nand UO_179 (O_179,N_2989,N_2968);
nor UO_180 (O_180,N_2978,N_2993);
xnor UO_181 (O_181,N_2994,N_2969);
xor UO_182 (O_182,N_2986,N_2965);
or UO_183 (O_183,N_2994,N_2959);
nand UO_184 (O_184,N_2972,N_2968);
nor UO_185 (O_185,N_2968,N_2979);
or UO_186 (O_186,N_2962,N_2986);
xor UO_187 (O_187,N_2962,N_2973);
xnor UO_188 (O_188,N_2967,N_2952);
nor UO_189 (O_189,N_2955,N_2957);
nor UO_190 (O_190,N_2960,N_2991);
nor UO_191 (O_191,N_2965,N_2972);
or UO_192 (O_192,N_2970,N_2958);
nand UO_193 (O_193,N_2975,N_2999);
or UO_194 (O_194,N_2957,N_2994);
and UO_195 (O_195,N_2957,N_2980);
and UO_196 (O_196,N_2986,N_2964);
and UO_197 (O_197,N_2950,N_2964);
and UO_198 (O_198,N_2967,N_2970);
nor UO_199 (O_199,N_2970,N_2990);
nand UO_200 (O_200,N_2953,N_2964);
or UO_201 (O_201,N_2956,N_2993);
and UO_202 (O_202,N_2989,N_2997);
or UO_203 (O_203,N_2953,N_2981);
nand UO_204 (O_204,N_2966,N_2978);
xor UO_205 (O_205,N_2969,N_2985);
nand UO_206 (O_206,N_2951,N_2994);
or UO_207 (O_207,N_2980,N_2971);
xor UO_208 (O_208,N_2992,N_2975);
nor UO_209 (O_209,N_2958,N_2964);
nor UO_210 (O_210,N_2972,N_2952);
nand UO_211 (O_211,N_2959,N_2955);
nor UO_212 (O_212,N_2968,N_2976);
nor UO_213 (O_213,N_2958,N_2953);
xor UO_214 (O_214,N_2979,N_2995);
and UO_215 (O_215,N_2977,N_2966);
xor UO_216 (O_216,N_2968,N_2973);
and UO_217 (O_217,N_2950,N_2966);
nand UO_218 (O_218,N_2973,N_2957);
and UO_219 (O_219,N_2982,N_2995);
nand UO_220 (O_220,N_2980,N_2969);
nor UO_221 (O_221,N_2977,N_2991);
nor UO_222 (O_222,N_2997,N_2992);
nand UO_223 (O_223,N_2977,N_2996);
or UO_224 (O_224,N_2981,N_2955);
nand UO_225 (O_225,N_2953,N_2994);
nand UO_226 (O_226,N_2973,N_2978);
nand UO_227 (O_227,N_2981,N_2977);
or UO_228 (O_228,N_2984,N_2973);
nor UO_229 (O_229,N_2996,N_2993);
or UO_230 (O_230,N_2958,N_2985);
nor UO_231 (O_231,N_2964,N_2966);
nor UO_232 (O_232,N_2998,N_2979);
xor UO_233 (O_233,N_2990,N_2961);
xnor UO_234 (O_234,N_2996,N_2959);
and UO_235 (O_235,N_2986,N_2972);
or UO_236 (O_236,N_2966,N_2988);
xor UO_237 (O_237,N_2968,N_2954);
xor UO_238 (O_238,N_2995,N_2952);
nand UO_239 (O_239,N_2982,N_2963);
xor UO_240 (O_240,N_2959,N_2989);
xnor UO_241 (O_241,N_2952,N_2998);
xnor UO_242 (O_242,N_2973,N_2952);
nor UO_243 (O_243,N_2962,N_2979);
nand UO_244 (O_244,N_2962,N_2969);
and UO_245 (O_245,N_2983,N_2964);
and UO_246 (O_246,N_2989,N_2962);
nand UO_247 (O_247,N_2976,N_2980);
nor UO_248 (O_248,N_2980,N_2960);
nand UO_249 (O_249,N_2951,N_2974);
nor UO_250 (O_250,N_2971,N_2975);
nor UO_251 (O_251,N_2954,N_2955);
and UO_252 (O_252,N_2998,N_2984);
or UO_253 (O_253,N_2956,N_2994);
nor UO_254 (O_254,N_2984,N_2990);
nor UO_255 (O_255,N_2963,N_2976);
nand UO_256 (O_256,N_2971,N_2991);
or UO_257 (O_257,N_2956,N_2983);
and UO_258 (O_258,N_2989,N_2985);
and UO_259 (O_259,N_2985,N_2986);
nor UO_260 (O_260,N_2978,N_2962);
nor UO_261 (O_261,N_2986,N_2968);
nor UO_262 (O_262,N_2964,N_2973);
nand UO_263 (O_263,N_2985,N_2987);
nor UO_264 (O_264,N_2993,N_2952);
and UO_265 (O_265,N_2963,N_2965);
or UO_266 (O_266,N_2950,N_2983);
xor UO_267 (O_267,N_2962,N_2988);
nand UO_268 (O_268,N_2995,N_2975);
nand UO_269 (O_269,N_2957,N_2989);
or UO_270 (O_270,N_2958,N_2990);
nand UO_271 (O_271,N_2958,N_2981);
xnor UO_272 (O_272,N_2960,N_2952);
or UO_273 (O_273,N_2967,N_2972);
nand UO_274 (O_274,N_2964,N_2997);
and UO_275 (O_275,N_2976,N_2965);
xor UO_276 (O_276,N_2996,N_2950);
xor UO_277 (O_277,N_2957,N_2981);
nand UO_278 (O_278,N_2978,N_2988);
nor UO_279 (O_279,N_2952,N_2962);
nor UO_280 (O_280,N_2977,N_2974);
xor UO_281 (O_281,N_2984,N_2955);
nor UO_282 (O_282,N_2956,N_2969);
nand UO_283 (O_283,N_2989,N_2984);
nor UO_284 (O_284,N_2991,N_2959);
and UO_285 (O_285,N_2995,N_2993);
nand UO_286 (O_286,N_2998,N_2970);
and UO_287 (O_287,N_2977,N_2999);
nor UO_288 (O_288,N_2956,N_2991);
and UO_289 (O_289,N_2985,N_2982);
or UO_290 (O_290,N_2991,N_2974);
nand UO_291 (O_291,N_2951,N_2965);
or UO_292 (O_292,N_2987,N_2963);
xnor UO_293 (O_293,N_2965,N_2966);
nand UO_294 (O_294,N_2985,N_2981);
xnor UO_295 (O_295,N_2983,N_2984);
and UO_296 (O_296,N_2995,N_2972);
or UO_297 (O_297,N_2984,N_2991);
xor UO_298 (O_298,N_2968,N_2987);
nand UO_299 (O_299,N_2979,N_2975);
xor UO_300 (O_300,N_2981,N_2967);
nand UO_301 (O_301,N_2988,N_2981);
nor UO_302 (O_302,N_2969,N_2970);
xor UO_303 (O_303,N_2972,N_2962);
nor UO_304 (O_304,N_2969,N_2972);
xor UO_305 (O_305,N_2979,N_2984);
nand UO_306 (O_306,N_2968,N_2983);
xor UO_307 (O_307,N_2978,N_2970);
or UO_308 (O_308,N_2964,N_2988);
xnor UO_309 (O_309,N_2983,N_2986);
nor UO_310 (O_310,N_2982,N_2970);
and UO_311 (O_311,N_2969,N_2983);
xor UO_312 (O_312,N_2968,N_2971);
xor UO_313 (O_313,N_2990,N_2985);
nand UO_314 (O_314,N_2972,N_2998);
xnor UO_315 (O_315,N_2978,N_2967);
and UO_316 (O_316,N_2952,N_2971);
xnor UO_317 (O_317,N_2966,N_2961);
or UO_318 (O_318,N_2956,N_2981);
nor UO_319 (O_319,N_2961,N_2960);
and UO_320 (O_320,N_2991,N_2975);
nor UO_321 (O_321,N_2970,N_2988);
nand UO_322 (O_322,N_2966,N_2990);
and UO_323 (O_323,N_2974,N_2971);
nand UO_324 (O_324,N_2969,N_2965);
and UO_325 (O_325,N_2951,N_2980);
or UO_326 (O_326,N_2953,N_2962);
nor UO_327 (O_327,N_2978,N_2999);
or UO_328 (O_328,N_2988,N_2984);
xor UO_329 (O_329,N_2960,N_2988);
nor UO_330 (O_330,N_2971,N_2977);
nand UO_331 (O_331,N_2985,N_2963);
nand UO_332 (O_332,N_2998,N_2983);
xor UO_333 (O_333,N_2960,N_2951);
nor UO_334 (O_334,N_2992,N_2980);
nor UO_335 (O_335,N_2958,N_2954);
nand UO_336 (O_336,N_2994,N_2986);
or UO_337 (O_337,N_2959,N_2992);
and UO_338 (O_338,N_2981,N_2966);
xor UO_339 (O_339,N_2954,N_2977);
nand UO_340 (O_340,N_2981,N_2987);
or UO_341 (O_341,N_2953,N_2961);
xnor UO_342 (O_342,N_2996,N_2982);
and UO_343 (O_343,N_2974,N_2980);
xnor UO_344 (O_344,N_2983,N_2965);
nand UO_345 (O_345,N_2995,N_2998);
nand UO_346 (O_346,N_2962,N_2958);
xnor UO_347 (O_347,N_2970,N_2976);
xor UO_348 (O_348,N_2972,N_2988);
nand UO_349 (O_349,N_2984,N_2980);
xor UO_350 (O_350,N_2982,N_2952);
nor UO_351 (O_351,N_2984,N_2964);
nor UO_352 (O_352,N_2974,N_2967);
nand UO_353 (O_353,N_2993,N_2967);
nor UO_354 (O_354,N_2958,N_2978);
nand UO_355 (O_355,N_2993,N_2999);
nand UO_356 (O_356,N_2986,N_2990);
nand UO_357 (O_357,N_2981,N_2963);
nor UO_358 (O_358,N_2981,N_2982);
and UO_359 (O_359,N_2982,N_2961);
nand UO_360 (O_360,N_2955,N_2961);
nor UO_361 (O_361,N_2973,N_2959);
and UO_362 (O_362,N_2955,N_2956);
nand UO_363 (O_363,N_2953,N_2973);
nor UO_364 (O_364,N_2995,N_2960);
or UO_365 (O_365,N_2985,N_2973);
nor UO_366 (O_366,N_2975,N_2974);
and UO_367 (O_367,N_2978,N_2984);
xor UO_368 (O_368,N_2961,N_2986);
nor UO_369 (O_369,N_2988,N_2969);
xnor UO_370 (O_370,N_2954,N_2988);
or UO_371 (O_371,N_2954,N_2953);
nand UO_372 (O_372,N_2977,N_2982);
and UO_373 (O_373,N_2992,N_2960);
or UO_374 (O_374,N_2990,N_2982);
xnor UO_375 (O_375,N_2969,N_2989);
xnor UO_376 (O_376,N_2998,N_2971);
nor UO_377 (O_377,N_2992,N_2966);
nand UO_378 (O_378,N_2991,N_2979);
or UO_379 (O_379,N_2954,N_2978);
nor UO_380 (O_380,N_2963,N_2977);
nand UO_381 (O_381,N_2955,N_2983);
and UO_382 (O_382,N_2952,N_2996);
nor UO_383 (O_383,N_2980,N_2991);
nand UO_384 (O_384,N_2969,N_2954);
nand UO_385 (O_385,N_2972,N_2974);
nor UO_386 (O_386,N_2970,N_2981);
xor UO_387 (O_387,N_2975,N_2967);
or UO_388 (O_388,N_2960,N_2953);
or UO_389 (O_389,N_2995,N_2973);
and UO_390 (O_390,N_2977,N_2984);
and UO_391 (O_391,N_2983,N_2966);
and UO_392 (O_392,N_2968,N_2970);
nand UO_393 (O_393,N_2983,N_2960);
nand UO_394 (O_394,N_2993,N_2971);
nor UO_395 (O_395,N_2978,N_2998);
or UO_396 (O_396,N_2991,N_2955);
or UO_397 (O_397,N_2974,N_2953);
nor UO_398 (O_398,N_2990,N_2991);
nor UO_399 (O_399,N_2954,N_2971);
nand UO_400 (O_400,N_2954,N_2995);
nand UO_401 (O_401,N_2956,N_2957);
or UO_402 (O_402,N_2969,N_2982);
or UO_403 (O_403,N_2978,N_2955);
and UO_404 (O_404,N_2954,N_2962);
nor UO_405 (O_405,N_2961,N_2952);
or UO_406 (O_406,N_2990,N_2950);
xnor UO_407 (O_407,N_2990,N_2968);
and UO_408 (O_408,N_2981,N_2964);
and UO_409 (O_409,N_2996,N_2971);
nand UO_410 (O_410,N_2979,N_2963);
and UO_411 (O_411,N_2954,N_2979);
or UO_412 (O_412,N_2957,N_2976);
nor UO_413 (O_413,N_2963,N_2951);
and UO_414 (O_414,N_2988,N_2983);
nand UO_415 (O_415,N_2956,N_2964);
nand UO_416 (O_416,N_2988,N_2961);
nor UO_417 (O_417,N_2979,N_2994);
and UO_418 (O_418,N_2999,N_2951);
or UO_419 (O_419,N_2961,N_2958);
nor UO_420 (O_420,N_2975,N_2963);
nand UO_421 (O_421,N_2985,N_2997);
xnor UO_422 (O_422,N_2978,N_2950);
or UO_423 (O_423,N_2961,N_2972);
nand UO_424 (O_424,N_2957,N_2984);
nand UO_425 (O_425,N_2955,N_2966);
nor UO_426 (O_426,N_2990,N_2960);
and UO_427 (O_427,N_2983,N_2972);
nand UO_428 (O_428,N_2955,N_2982);
nor UO_429 (O_429,N_2951,N_2979);
or UO_430 (O_430,N_2960,N_2984);
nor UO_431 (O_431,N_2961,N_2978);
or UO_432 (O_432,N_2961,N_2964);
nor UO_433 (O_433,N_2976,N_2955);
nor UO_434 (O_434,N_2998,N_2975);
nor UO_435 (O_435,N_2999,N_2963);
nand UO_436 (O_436,N_2998,N_2988);
or UO_437 (O_437,N_2967,N_2959);
nor UO_438 (O_438,N_2969,N_2966);
xnor UO_439 (O_439,N_2982,N_2984);
nor UO_440 (O_440,N_2998,N_2980);
xor UO_441 (O_441,N_2971,N_2965);
or UO_442 (O_442,N_2975,N_2976);
xnor UO_443 (O_443,N_2977,N_2955);
nand UO_444 (O_444,N_2957,N_2993);
and UO_445 (O_445,N_2981,N_2976);
xnor UO_446 (O_446,N_2950,N_2994);
nand UO_447 (O_447,N_2983,N_2973);
xor UO_448 (O_448,N_2957,N_2968);
nand UO_449 (O_449,N_2990,N_2989);
and UO_450 (O_450,N_2975,N_2986);
nor UO_451 (O_451,N_2975,N_2984);
and UO_452 (O_452,N_2982,N_2980);
nor UO_453 (O_453,N_2986,N_2973);
xor UO_454 (O_454,N_2996,N_2968);
and UO_455 (O_455,N_2975,N_2977);
nand UO_456 (O_456,N_2965,N_2954);
xnor UO_457 (O_457,N_2989,N_2977);
nor UO_458 (O_458,N_2990,N_2987);
nor UO_459 (O_459,N_2954,N_2957);
xnor UO_460 (O_460,N_2969,N_2981);
and UO_461 (O_461,N_2964,N_2990);
and UO_462 (O_462,N_2970,N_2955);
xnor UO_463 (O_463,N_2957,N_2995);
and UO_464 (O_464,N_2967,N_2966);
xor UO_465 (O_465,N_2980,N_2985);
or UO_466 (O_466,N_2958,N_2997);
xnor UO_467 (O_467,N_2991,N_2961);
and UO_468 (O_468,N_2967,N_2958);
or UO_469 (O_469,N_2983,N_2953);
and UO_470 (O_470,N_2968,N_2955);
or UO_471 (O_471,N_2982,N_2960);
or UO_472 (O_472,N_2974,N_2985);
or UO_473 (O_473,N_2962,N_2981);
nand UO_474 (O_474,N_2970,N_2964);
nor UO_475 (O_475,N_2978,N_2987);
nand UO_476 (O_476,N_2990,N_2967);
and UO_477 (O_477,N_2958,N_2977);
and UO_478 (O_478,N_2965,N_2991);
xor UO_479 (O_479,N_2971,N_2981);
and UO_480 (O_480,N_2959,N_2962);
and UO_481 (O_481,N_2987,N_2996);
nor UO_482 (O_482,N_2954,N_2991);
and UO_483 (O_483,N_2959,N_2964);
and UO_484 (O_484,N_2965,N_2999);
and UO_485 (O_485,N_2979,N_2967);
nor UO_486 (O_486,N_2953,N_2959);
nand UO_487 (O_487,N_2991,N_2992);
nor UO_488 (O_488,N_2952,N_2999);
and UO_489 (O_489,N_2953,N_2984);
or UO_490 (O_490,N_2959,N_2954);
or UO_491 (O_491,N_2978,N_2991);
or UO_492 (O_492,N_2984,N_2981);
or UO_493 (O_493,N_2961,N_2998);
or UO_494 (O_494,N_2994,N_2967);
nand UO_495 (O_495,N_2950,N_2971);
xnor UO_496 (O_496,N_2954,N_2972);
xnor UO_497 (O_497,N_2975,N_2978);
nor UO_498 (O_498,N_2957,N_2967);
or UO_499 (O_499,N_2955,N_2974);
endmodule