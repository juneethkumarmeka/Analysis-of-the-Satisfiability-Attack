module basic_1500_15000_2000_5_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_18,In_1400);
and U1 (N_1,In_1252,In_1160);
or U2 (N_2,In_1446,In_986);
nand U3 (N_3,In_219,In_879);
xor U4 (N_4,In_1310,In_677);
xnor U5 (N_5,In_822,In_443);
and U6 (N_6,In_440,In_70);
or U7 (N_7,In_305,In_373);
nand U8 (N_8,In_1012,In_1347);
nor U9 (N_9,In_390,In_3);
or U10 (N_10,In_1179,In_728);
or U11 (N_11,In_1052,In_617);
nand U12 (N_12,In_169,In_422);
or U13 (N_13,In_1321,In_332);
nand U14 (N_14,In_831,In_635);
and U15 (N_15,In_551,In_1144);
nand U16 (N_16,In_476,In_323);
nor U17 (N_17,In_1061,In_752);
or U18 (N_18,In_241,In_381);
nor U19 (N_19,In_172,In_526);
or U20 (N_20,In_60,In_1381);
xor U21 (N_21,In_1011,In_571);
or U22 (N_22,In_200,In_1067);
and U23 (N_23,In_1247,In_912);
nand U24 (N_24,In_162,In_100);
and U25 (N_25,In_818,In_410);
nand U26 (N_26,In_953,In_7);
and U27 (N_27,In_956,In_507);
nor U28 (N_28,In_700,In_606);
and U29 (N_29,In_924,In_345);
nor U30 (N_30,In_302,In_969);
nand U31 (N_31,In_512,In_846);
and U32 (N_32,In_59,In_1178);
nand U33 (N_33,In_599,In_480);
nand U34 (N_34,In_73,In_431);
nand U35 (N_35,In_152,In_828);
or U36 (N_36,In_459,In_922);
nand U37 (N_37,In_511,In_616);
nand U38 (N_38,In_984,In_790);
and U39 (N_39,In_1435,In_519);
and U40 (N_40,In_21,In_52);
xnor U41 (N_41,In_38,In_191);
xor U42 (N_42,In_954,In_259);
nor U43 (N_43,In_117,In_399);
or U44 (N_44,In_707,In_646);
or U45 (N_45,In_868,In_449);
nor U46 (N_46,In_216,In_1239);
xor U47 (N_47,In_1173,In_1390);
or U48 (N_48,In_209,In_656);
nand U49 (N_49,In_29,In_1250);
or U50 (N_50,In_958,In_861);
and U51 (N_51,In_1357,In_1209);
or U52 (N_52,In_553,In_1298);
or U53 (N_53,In_126,In_1208);
nand U54 (N_54,In_321,In_691);
nand U55 (N_55,In_246,In_1242);
and U56 (N_56,In_139,In_327);
and U57 (N_57,In_939,In_962);
and U58 (N_58,In_185,In_638);
or U59 (N_59,In_583,In_252);
nor U60 (N_60,In_562,In_849);
or U61 (N_61,In_411,In_826);
and U62 (N_62,In_1385,In_625);
and U63 (N_63,In_769,In_1387);
nor U64 (N_64,In_362,In_1037);
xnor U65 (N_65,In_1189,In_400);
and U66 (N_66,In_539,In_417);
and U67 (N_67,In_749,In_781);
xor U68 (N_68,In_28,In_518);
or U69 (N_69,In_785,In_1266);
nand U70 (N_70,In_1030,In_223);
or U71 (N_71,In_166,In_1223);
nor U72 (N_72,In_670,In_1312);
nor U73 (N_73,In_723,In_63);
nor U74 (N_74,In_387,In_397);
or U75 (N_75,In_739,In_1262);
nand U76 (N_76,In_19,In_217);
nor U77 (N_77,In_1380,In_1422);
nand U78 (N_78,In_1459,In_1001);
and U79 (N_79,In_1318,In_347);
xnor U80 (N_80,In_573,In_832);
or U81 (N_81,In_661,In_914);
nor U82 (N_82,In_1485,In_726);
nor U83 (N_83,In_446,In_1075);
nand U84 (N_84,In_1218,In_243);
or U85 (N_85,In_1194,In_477);
and U86 (N_86,In_27,In_86);
nand U87 (N_87,In_655,In_565);
or U88 (N_88,In_313,In_1103);
nand U89 (N_89,In_1113,In_307);
nand U90 (N_90,In_469,In_970);
nor U91 (N_91,In_1366,In_467);
nand U92 (N_92,In_1344,In_42);
and U93 (N_93,In_508,In_1311);
nand U94 (N_94,In_1039,In_667);
and U95 (N_95,In_479,In_394);
nand U96 (N_96,In_1276,In_1292);
or U97 (N_97,In_917,In_325);
or U98 (N_98,In_1222,In_577);
and U99 (N_99,In_567,In_342);
nor U100 (N_100,In_1376,In_466);
or U101 (N_101,In_45,In_890);
and U102 (N_102,In_344,In_1049);
xor U103 (N_103,In_1120,In_475);
nand U104 (N_104,In_665,In_392);
or U105 (N_105,In_231,In_1035);
nand U106 (N_106,In_955,In_1442);
xor U107 (N_107,In_483,In_1154);
xnor U108 (N_108,In_201,In_1460);
and U109 (N_109,In_1201,In_555);
or U110 (N_110,In_1115,In_93);
nand U111 (N_111,In_836,In_759);
nand U112 (N_112,In_488,In_94);
nor U113 (N_113,In_77,In_1207);
nor U114 (N_114,In_393,In_340);
nand U115 (N_115,In_552,In_160);
or U116 (N_116,In_1349,In_1101);
nor U117 (N_117,In_1232,In_840);
or U118 (N_118,In_894,In_1394);
and U119 (N_119,In_647,In_258);
and U120 (N_120,In_242,In_963);
xnor U121 (N_121,In_951,In_751);
nor U122 (N_122,In_1413,In_238);
nand U123 (N_123,In_529,In_330);
and U124 (N_124,In_983,In_87);
nand U125 (N_125,In_343,In_1068);
nor U126 (N_126,In_1082,In_1213);
nand U127 (N_127,In_870,In_1433);
xnor U128 (N_128,In_904,In_1352);
nor U129 (N_129,In_1185,In_947);
nor U130 (N_130,In_99,In_1341);
and U131 (N_131,In_319,In_782);
and U132 (N_132,In_391,In_192);
nor U133 (N_133,In_1140,In_370);
or U134 (N_134,In_515,In_379);
nand U135 (N_135,In_196,In_1305);
and U136 (N_136,In_1184,In_1405);
or U137 (N_137,In_893,In_816);
nor U138 (N_138,In_992,In_31);
or U139 (N_139,In_468,In_1116);
nand U140 (N_140,In_128,In_1267);
or U141 (N_141,In_273,In_652);
or U142 (N_142,In_709,In_744);
and U143 (N_143,In_1156,In_1466);
or U144 (N_144,In_694,In_909);
and U145 (N_145,In_1461,In_1203);
or U146 (N_146,In_1444,In_1322);
or U147 (N_147,In_388,In_1475);
nand U148 (N_148,In_470,In_1470);
and U149 (N_149,In_1097,In_355);
nor U150 (N_150,In_680,In_1000);
nor U151 (N_151,In_239,In_1026);
xor U152 (N_152,In_1043,In_1240);
or U153 (N_153,In_442,In_973);
nor U154 (N_154,In_1355,In_280);
or U155 (N_155,In_1482,In_1086);
or U156 (N_156,In_1147,In_805);
xor U157 (N_157,In_47,In_741);
and U158 (N_158,In_386,In_1439);
and U159 (N_159,In_1278,In_1332);
and U160 (N_160,In_1010,In_352);
nand U161 (N_161,In_804,In_815);
and U162 (N_162,In_1118,In_717);
and U163 (N_163,In_1462,In_131);
nand U164 (N_164,In_1083,In_761);
or U165 (N_165,In_919,In_1195);
nor U166 (N_166,In_229,In_704);
or U167 (N_167,In_841,In_11);
nor U168 (N_168,In_982,In_213);
nand U169 (N_169,In_452,In_506);
nor U170 (N_170,In_257,In_1112);
or U171 (N_171,In_620,In_1265);
nand U172 (N_172,In_734,In_1196);
and U173 (N_173,In_1469,In_499);
nand U174 (N_174,In_996,In_684);
nand U175 (N_175,In_722,In_1443);
or U176 (N_176,In_718,In_1338);
or U177 (N_177,In_548,In_309);
or U178 (N_178,In_136,In_92);
and U179 (N_179,In_474,In_800);
and U180 (N_180,In_502,In_899);
or U181 (N_181,In_1393,In_773);
or U182 (N_182,In_170,In_1333);
nand U183 (N_183,In_1361,In_1453);
or U184 (N_184,In_275,In_409);
and U185 (N_185,In_224,In_1397);
and U186 (N_186,In_811,In_630);
nand U187 (N_187,In_1428,In_845);
xor U188 (N_188,In_750,In_654);
and U189 (N_189,In_64,In_703);
nor U190 (N_190,In_141,In_101);
or U191 (N_191,In_51,In_1170);
nand U192 (N_192,In_1077,In_13);
xor U193 (N_193,In_426,In_1127);
or U194 (N_194,In_1345,In_582);
and U195 (N_195,In_82,In_1161);
and U196 (N_196,In_966,In_1020);
or U197 (N_197,In_663,In_1259);
nor U198 (N_198,In_335,In_850);
nand U199 (N_199,In_1215,In_780);
xnor U200 (N_200,In_1430,In_1457);
nand U201 (N_201,In_487,In_928);
and U202 (N_202,In_1414,In_568);
or U203 (N_203,In_1448,In_642);
nor U204 (N_204,In_820,In_1210);
nand U205 (N_205,In_43,In_1018);
nand U206 (N_206,In_481,In_1078);
or U207 (N_207,In_455,In_603);
xnor U208 (N_208,In_883,In_33);
nand U209 (N_209,In_184,In_1374);
xnor U210 (N_210,In_1014,In_294);
or U211 (N_211,In_1495,In_1135);
and U212 (N_212,In_851,In_287);
or U213 (N_213,In_376,In_1166);
nor U214 (N_214,In_1382,In_1139);
or U215 (N_215,In_424,In_834);
nor U216 (N_216,In_181,In_318);
nand U217 (N_217,In_1155,In_934);
nand U218 (N_218,In_807,In_255);
or U219 (N_219,In_103,In_407);
or U220 (N_220,In_610,In_317);
nor U221 (N_221,In_639,In_199);
nand U222 (N_222,In_1050,In_176);
nor U223 (N_223,In_6,In_1377);
nor U224 (N_224,In_687,In_268);
nor U225 (N_225,In_501,In_1488);
nor U226 (N_226,In_1283,In_1133);
nand U227 (N_227,In_801,In_1163);
and U228 (N_228,In_971,In_1085);
or U229 (N_229,In_173,In_460);
and U230 (N_230,In_1299,In_1406);
xnor U231 (N_231,In_607,In_916);
nand U232 (N_232,In_668,In_1481);
nand U233 (N_233,In_897,In_648);
or U234 (N_234,In_1251,In_1188);
nand U235 (N_235,In_1301,In_1192);
and U236 (N_236,In_799,In_1108);
nor U237 (N_237,In_398,In_1330);
nand U238 (N_238,In_1263,In_1130);
and U239 (N_239,In_67,In_299);
nand U240 (N_240,In_1107,In_587);
nand U241 (N_241,In_806,In_1193);
nor U242 (N_242,In_492,In_858);
nor U243 (N_243,In_39,In_368);
nand U244 (N_244,In_1304,In_533);
and U245 (N_245,In_1069,In_1412);
and U246 (N_246,In_119,In_1307);
and U247 (N_247,In_1114,In_353);
or U248 (N_248,In_1104,In_1256);
nor U249 (N_249,In_1105,In_133);
nand U250 (N_250,In_68,In_366);
nand U251 (N_251,In_719,In_920);
nand U252 (N_252,In_632,In_197);
nor U253 (N_253,In_685,In_776);
xnor U254 (N_254,In_835,In_1151);
nand U255 (N_255,In_1497,In_696);
nand U256 (N_256,In_159,In_143);
nand U257 (N_257,In_608,In_447);
nand U258 (N_258,In_1248,In_1226);
or U259 (N_259,In_1099,In_389);
nor U260 (N_260,In_585,In_532);
and U261 (N_261,In_1423,In_227);
xnor U262 (N_262,In_17,In_1031);
or U263 (N_263,In_521,In_580);
and U264 (N_264,In_1190,In_406);
and U265 (N_265,In_416,In_165);
xor U266 (N_266,In_618,In_471);
nor U267 (N_267,In_102,In_1230);
nor U268 (N_268,In_936,In_732);
nor U269 (N_269,In_847,In_121);
and U270 (N_270,In_1490,In_848);
nor U271 (N_271,In_303,In_896);
nand U272 (N_272,In_793,In_743);
xnor U273 (N_273,In_784,In_277);
nor U274 (N_274,In_183,In_786);
or U275 (N_275,In_724,In_348);
or U276 (N_276,In_930,In_423);
nor U277 (N_277,In_1290,In_1062);
nor U278 (N_278,In_1360,In_1125);
or U279 (N_279,In_1295,In_421);
or U280 (N_280,In_425,In_1093);
or U281 (N_281,In_864,In_214);
xnor U282 (N_282,In_1362,In_637);
nand U283 (N_283,In_276,In_1306);
xnor U284 (N_284,In_337,In_931);
nor U285 (N_285,In_15,In_1261);
nor U286 (N_286,In_803,In_365);
nand U287 (N_287,In_178,In_633);
nand U288 (N_288,In_1021,In_53);
nor U289 (N_289,In_1288,In_1053);
nand U290 (N_290,In_0,In_251);
or U291 (N_291,In_46,In_377);
nand U292 (N_292,In_856,In_730);
xor U293 (N_293,In_641,In_977);
nor U294 (N_294,In_225,In_1006);
xor U295 (N_295,In_116,In_1445);
nand U296 (N_296,In_911,In_900);
nor U297 (N_297,In_232,In_413);
nor U298 (N_298,In_731,In_1205);
or U299 (N_299,In_1415,In_293);
or U300 (N_300,In_360,In_774);
nand U301 (N_301,In_282,In_1016);
and U302 (N_302,In_320,In_753);
nand U303 (N_303,In_435,In_634);
or U304 (N_304,In_1253,In_693);
and U305 (N_305,In_324,In_952);
nand U306 (N_306,In_1257,In_586);
or U307 (N_307,In_1491,In_1432);
and U308 (N_308,In_81,In_540);
nand U309 (N_309,In_813,In_26);
or U310 (N_310,In_742,In_714);
nand U311 (N_311,In_371,In_706);
nor U312 (N_312,In_829,In_1024);
or U313 (N_313,In_572,In_1369);
nand U314 (N_314,In_1143,In_333);
or U315 (N_315,In_619,In_1065);
xor U316 (N_316,In_1157,In_910);
or U317 (N_317,In_1227,In_1073);
nor U318 (N_318,In_609,In_578);
and U319 (N_319,In_270,In_927);
nand U320 (N_320,In_817,In_1167);
nand U321 (N_321,In_796,In_1424);
nor U322 (N_322,In_2,In_1383);
nand U323 (N_323,In_69,In_892);
xnor U324 (N_324,In_589,In_943);
nor U325 (N_325,In_1449,In_867);
nor U326 (N_326,In_1089,In_702);
nand U327 (N_327,In_510,In_929);
nand U328 (N_328,In_1176,In_998);
nor U329 (N_329,In_686,In_1291);
nor U330 (N_330,In_795,In_576);
nor U331 (N_331,In_1142,In_626);
and U332 (N_332,In_146,In_1229);
nand U333 (N_333,In_535,In_1111);
nor U334 (N_334,In_358,In_498);
nor U335 (N_335,In_1088,In_188);
xor U336 (N_336,In_1174,In_274);
and U337 (N_337,In_80,In_1465);
xor U338 (N_338,In_1055,In_1109);
or U339 (N_339,In_808,In_193);
nand U340 (N_340,In_810,In_249);
or U341 (N_341,In_177,In_266);
or U342 (N_342,In_1463,In_402);
nand U343 (N_343,In_210,In_175);
xnor U344 (N_344,In_1302,In_14);
and U345 (N_345,In_190,In_240);
nand U346 (N_346,In_374,In_737);
or U347 (N_347,In_1081,In_701);
nand U348 (N_348,In_109,In_1447);
nand U349 (N_349,In_1441,In_1395);
or U350 (N_350,In_575,In_1241);
and U351 (N_351,In_1181,In_860);
xnor U352 (N_352,In_437,In_78);
or U353 (N_353,In_1489,In_244);
nor U354 (N_354,In_1379,In_297);
and U355 (N_355,In_945,In_142);
nor U356 (N_356,In_1426,In_558);
nor U357 (N_357,In_1429,In_604);
and U358 (N_358,In_418,In_689);
and U359 (N_359,In_260,In_182);
nor U360 (N_360,In_300,In_334);
and U361 (N_361,In_1198,In_311);
nand U362 (N_362,In_401,In_1007);
xor U363 (N_363,In_125,In_1060);
nor U364 (N_364,In_1402,In_1388);
and U365 (N_365,In_872,In_821);
nor U366 (N_366,In_88,In_1389);
or U367 (N_367,In_1420,In_179);
and U368 (N_368,In_1280,In_1315);
xnor U369 (N_369,In_279,In_819);
and U370 (N_370,In_948,In_1177);
or U371 (N_371,In_1294,In_1408);
nand U372 (N_372,In_1323,In_155);
or U373 (N_373,In_91,In_461);
nor U374 (N_374,In_1100,In_1047);
or U375 (N_375,In_130,In_150);
or U376 (N_376,In_1375,In_740);
nor U377 (N_377,In_1172,In_1246);
and U378 (N_378,In_509,In_738);
and U379 (N_379,In_908,In_1492);
nor U380 (N_380,In_600,In_1214);
and U381 (N_381,In_531,In_935);
nand U382 (N_382,In_754,In_1152);
or U383 (N_383,In_1498,In_494);
nor U384 (N_384,In_1045,In_1244);
and U385 (N_385,In_913,In_1199);
and U386 (N_386,In_859,In_420);
nand U387 (N_387,In_843,In_195);
and U388 (N_388,In_71,In_35);
nor U389 (N_389,In_888,In_322);
and U390 (N_390,In_112,In_676);
and U391 (N_391,In_104,In_151);
and U392 (N_392,In_1245,In_651);
and U393 (N_393,In_154,In_415);
and U394 (N_394,In_653,In_37);
nand U395 (N_395,In_797,In_308);
and U396 (N_396,In_118,In_84);
nand U397 (N_397,In_329,In_1386);
and U398 (N_398,In_108,In_264);
nand U399 (N_399,In_180,In_1028);
and U400 (N_400,In_156,In_538);
or U401 (N_401,In_1437,In_1450);
nand U402 (N_402,In_853,In_1141);
nand U403 (N_403,In_1277,In_697);
xor U404 (N_404,In_1496,In_1219);
or U405 (N_405,In_234,In_906);
or U406 (N_406,In_9,In_588);
and U407 (N_407,In_877,In_158);
and U408 (N_408,In_987,In_1233);
and U409 (N_409,In_32,In_884);
and U410 (N_410,In_48,In_298);
nand U411 (N_411,In_1326,In_783);
nand U412 (N_412,In_202,In_1478);
nand U413 (N_413,In_1058,In_439);
xnor U414 (N_414,In_1027,In_341);
nand U415 (N_415,In_1396,In_1421);
nor U416 (N_416,In_1087,In_645);
and U417 (N_417,In_525,In_901);
nor U418 (N_418,In_369,In_865);
or U419 (N_419,In_764,In_1074);
and U420 (N_420,In_1317,In_825);
nand U421 (N_421,In_1419,In_1216);
xnor U422 (N_422,In_57,In_683);
and U423 (N_423,In_1162,In_1427);
or U424 (N_424,In_50,In_1336);
nand U425 (N_425,In_596,In_1407);
and U426 (N_426,In_157,In_316);
nand U427 (N_427,In_451,In_1458);
nand U428 (N_428,In_1409,In_198);
or U429 (N_429,In_1499,In_950);
nor U430 (N_430,In_594,In_729);
nor U431 (N_431,In_4,In_679);
or U432 (N_432,In_756,In_1098);
nor U433 (N_433,In_1095,In_623);
nand U434 (N_434,In_824,In_1042);
or U435 (N_435,In_1009,In_543);
or U436 (N_436,In_946,In_611);
nand U437 (N_437,In_1002,In_1325);
xnor U438 (N_438,In_854,In_263);
or U439 (N_439,In_412,In_1080);
xnor U440 (N_440,In_1313,In_852);
xor U441 (N_441,In_777,In_1316);
nand U442 (N_442,In_755,In_563);
nor U443 (N_443,In_285,In_1057);
xnor U444 (N_444,In_968,In_331);
or U445 (N_445,In_1234,In_1476);
nand U446 (N_446,In_380,In_484);
and U447 (N_447,In_602,In_289);
or U448 (N_448,In_561,In_83);
nor U449 (N_449,In_438,In_363);
and U450 (N_450,In_505,In_716);
nor U451 (N_451,In_886,In_122);
nor U452 (N_452,In_1070,In_1356);
nor U453 (N_453,In_627,In_113);
and U454 (N_454,In_105,In_855);
or U455 (N_455,In_1134,In_145);
and U456 (N_456,In_1328,In_1486);
and U457 (N_457,In_964,In_495);
nand U458 (N_458,In_1410,In_1372);
and U459 (N_459,In_1048,In_721);
and U460 (N_460,In_493,In_1046);
nor U461 (N_461,In_725,In_995);
xnor U462 (N_462,In_235,In_74);
nor U463 (N_463,In_1110,In_763);
xnor U464 (N_464,In_34,In_304);
and U465 (N_465,In_591,In_905);
nor U466 (N_466,In_336,In_889);
or U467 (N_467,In_699,In_328);
and U468 (N_468,In_557,In_823);
nand U469 (N_469,In_658,In_1044);
and U470 (N_470,In_1271,In_1335);
nor U471 (N_471,In_514,In_473);
nor U472 (N_472,In_1417,In_339);
nand U473 (N_473,In_253,In_1017);
or U474 (N_474,In_288,In_1260);
or U475 (N_475,In_1436,In_839);
nor U476 (N_476,In_1090,In_915);
or U477 (N_477,In_727,In_350);
nor U478 (N_478,In_713,In_115);
and U479 (N_479,In_712,In_351);
nor U480 (N_480,In_1249,In_593);
nor U481 (N_481,In_1091,In_622);
nor U482 (N_482,In_798,In_189);
nor U483 (N_483,In_144,In_463);
nand U484 (N_484,In_1025,In_650);
nand U485 (N_485,In_207,In_1308);
nor U486 (N_486,In_1149,In_942);
and U487 (N_487,In_1084,In_569);
nand U488 (N_488,In_75,In_838);
and U489 (N_489,In_628,In_1473);
or U490 (N_490,In_444,In_644);
xnor U491 (N_491,In_1454,In_748);
nand U492 (N_492,In_54,In_215);
or U493 (N_493,In_1314,In_1059);
and U494 (N_494,In_978,In_462);
nor U495 (N_495,In_385,In_1353);
or U496 (N_496,In_1106,In_513);
and U497 (N_497,In_736,In_430);
nor U498 (N_498,In_1368,In_527);
nor U499 (N_499,In_296,In_186);
nor U500 (N_500,In_486,In_1224);
or U501 (N_501,In_1153,In_698);
nor U502 (N_502,In_1286,In_1279);
or U503 (N_503,In_1183,In_873);
nor U504 (N_504,In_812,In_1164);
and U505 (N_505,In_1411,In_419);
and U506 (N_506,In_564,In_862);
or U507 (N_507,In_124,In_349);
nand U508 (N_508,In_613,In_20);
xor U509 (N_509,In_408,In_944);
nand U510 (N_510,In_990,In_882);
or U511 (N_511,In_671,In_1434);
and U512 (N_512,In_1339,In_708);
nor U513 (N_513,In_1029,In_1348);
and U514 (N_514,In_290,In_649);
nand U515 (N_515,In_378,In_876);
nand U516 (N_516,In_866,In_250);
nand U517 (N_517,In_1094,In_1236);
and U518 (N_518,In_516,In_211);
and U519 (N_519,In_695,In_937);
xor U520 (N_520,In_1136,In_546);
or U521 (N_521,In_1275,In_269);
and U522 (N_522,In_584,In_1398);
nand U523 (N_523,In_1220,In_167);
or U524 (N_524,In_1054,In_1354);
and U525 (N_525,In_1200,In_659);
nor U526 (N_526,In_1455,In_833);
or U527 (N_527,In_536,In_590);
nor U528 (N_528,In_541,In_1479);
xnor U529 (N_529,In_448,In_520);
xnor U530 (N_530,In_1342,In_1324);
nand U531 (N_531,In_779,In_1350);
and U532 (N_532,In_770,In_135);
nand U533 (N_533,In_1180,In_504);
or U534 (N_534,In_95,In_1358);
nor U535 (N_535,In_1119,In_1063);
nand U536 (N_536,In_1272,In_36);
or U537 (N_537,In_291,In_262);
and U538 (N_538,In_985,In_674);
or U539 (N_539,In_842,In_1129);
nor U540 (N_540,In_961,In_1487);
nor U541 (N_541,In_989,In_1367);
nand U542 (N_542,In_972,In_1126);
nand U543 (N_543,In_496,In_140);
and U544 (N_544,In_1329,In_517);
nor U545 (N_545,In_168,In_148);
and U546 (N_546,In_1484,In_107);
and U547 (N_547,In_147,In_1269);
nor U548 (N_548,In_1401,In_1072);
xnor U549 (N_549,In_560,In_1165);
and U550 (N_550,In_857,In_1480);
nor U551 (N_551,In_710,In_1483);
and U552 (N_552,In_891,In_433);
nand U553 (N_553,In_236,In_1289);
nand U554 (N_554,In_615,In_132);
and U555 (N_555,In_967,In_534);
or U556 (N_556,In_1132,In_161);
or U557 (N_557,In_90,In_346);
or U558 (N_558,In_1363,In_705);
and U559 (N_559,In_903,In_1243);
nand U560 (N_560,In_310,In_844);
nor U561 (N_561,In_434,In_720);
nor U562 (N_562,In_1211,In_1254);
and U563 (N_563,In_994,In_907);
nand U564 (N_564,In_745,In_1171);
nor U565 (N_565,In_138,In_601);
and U566 (N_566,In_1471,In_1346);
and U567 (N_567,In_869,In_222);
and U568 (N_568,In_1221,In_690);
and U569 (N_569,In_1191,In_1327);
nand U570 (N_570,In_1255,In_85);
nor U571 (N_571,In_267,In_163);
and U572 (N_572,In_233,In_675);
and U573 (N_573,In_292,In_621);
or U574 (N_574,In_1258,In_1225);
or U575 (N_575,In_237,In_871);
nor U576 (N_576,In_523,In_212);
nor U577 (N_577,In_528,In_164);
or U578 (N_578,In_688,In_566);
nand U579 (N_579,In_1399,In_1452);
and U580 (N_580,In_56,In_1);
nor U581 (N_581,In_809,In_522);
nor U582 (N_582,In_55,In_491);
nand U583 (N_583,In_1138,In_10);
nor U584 (N_584,In_450,In_1300);
xor U585 (N_585,In_356,In_208);
or U586 (N_586,In_12,In_1015);
xnor U587 (N_587,In_441,In_457);
nor U588 (N_588,In_1343,In_1197);
nor U589 (N_589,In_993,In_367);
nor U590 (N_590,In_1022,In_1071);
nand U591 (N_591,In_1123,In_794);
and U592 (N_592,In_428,In_789);
and U593 (N_593,In_62,In_624);
and U594 (N_594,In_134,In_1212);
nor U595 (N_595,In_542,In_89);
and U596 (N_596,In_106,In_432);
and U597 (N_597,In_997,In_454);
nor U598 (N_598,In_326,In_581);
or U599 (N_599,In_8,In_361);
nor U600 (N_600,In_220,In_1494);
and U601 (N_601,In_925,In_1217);
xnor U602 (N_602,In_66,In_1187);
nand U603 (N_603,In_550,In_1403);
nor U604 (N_604,In_762,In_1128);
nand U605 (N_605,In_1370,In_315);
or U606 (N_606,In_758,In_666);
nand U607 (N_607,In_429,In_1092);
or U608 (N_608,In_1040,In_747);
and U609 (N_609,In_1145,In_1231);
and U610 (N_610,In_306,In_1285);
or U611 (N_611,In_791,In_248);
nor U612 (N_612,In_382,In_384);
or U613 (N_613,In_271,In_187);
nor U614 (N_614,In_364,In_1122);
nand U615 (N_615,In_123,In_1204);
and U616 (N_616,In_874,In_383);
or U617 (N_617,In_61,In_940);
nand U618 (N_618,In_711,In_281);
xnor U619 (N_619,In_957,In_1438);
and U620 (N_620,In_1264,In_312);
xnor U621 (N_621,In_1303,In_1340);
or U622 (N_622,In_1051,In_228);
or U623 (N_623,In_544,In_549);
nor U624 (N_624,In_1202,In_44);
xnor U625 (N_625,In_746,In_283);
and U626 (N_626,In_359,In_733);
or U627 (N_627,In_489,In_1175);
xnor U628 (N_628,In_1418,In_926);
nor U629 (N_629,In_129,In_1472);
nor U630 (N_630,In_837,In_204);
or U631 (N_631,In_1391,In_1284);
or U632 (N_632,In_111,In_49);
and U633 (N_633,In_1359,In_120);
or U634 (N_634,In_265,In_1431);
nand U635 (N_635,In_629,In_556);
nand U636 (N_636,In_1159,In_1331);
nand U637 (N_637,In_640,In_975);
xnor U638 (N_638,In_482,In_41);
and U639 (N_639,In_1451,In_1066);
nand U640 (N_640,In_301,In_830);
or U641 (N_641,In_547,In_1038);
and U642 (N_642,In_40,In_918);
or U643 (N_643,In_203,In_1079);
and U644 (N_644,In_1287,In_1493);
nand U645 (N_645,In_863,In_921);
or U646 (N_646,In_295,In_881);
xor U647 (N_647,In_631,In_110);
xor U648 (N_648,In_194,In_692);
nor U649 (N_649,In_660,In_885);
and U650 (N_650,In_938,In_974);
nor U651 (N_651,In_715,In_765);
or U652 (N_652,In_375,In_114);
and U653 (N_653,In_1003,In_999);
nand U654 (N_654,In_30,In_261);
nand U655 (N_655,In_1425,In_403);
nor U656 (N_656,In_24,In_1169);
nor U657 (N_657,In_1293,In_22);
and U658 (N_658,In_254,In_286);
nand U659 (N_659,In_991,In_127);
and U660 (N_660,In_1309,In_153);
nand U661 (N_661,In_1228,In_875);
nand U662 (N_662,In_595,In_965);
and U663 (N_663,In_636,In_988);
nand U664 (N_664,In_664,In_775);
nand U665 (N_665,In_338,In_554);
nand U666 (N_666,In_767,In_579);
nor U667 (N_667,In_1131,In_1270);
nand U668 (N_668,In_23,In_643);
and U669 (N_669,In_902,In_1036);
nand U670 (N_670,In_574,In_768);
nor U671 (N_671,In_1158,In_778);
or U672 (N_672,In_478,In_669);
or U673 (N_673,In_980,In_171);
and U674 (N_674,In_1182,In_396);
and U675 (N_675,In_456,In_1206);
nand U676 (N_676,In_221,In_445);
nor U677 (N_677,In_682,In_976);
nand U678 (N_678,In_1416,In_949);
nor U679 (N_679,In_612,In_827);
nor U680 (N_680,In_58,In_1351);
or U681 (N_681,In_772,In_1296);
nor U682 (N_682,In_500,In_1013);
nor U683 (N_683,In_530,In_464);
nor U684 (N_684,In_771,In_1373);
xor U685 (N_685,In_149,In_757);
nor U686 (N_686,In_284,In_1032);
and U687 (N_687,In_404,In_497);
and U688 (N_688,In_1237,In_357);
and U689 (N_689,In_206,In_933);
nand U690 (N_690,In_1281,In_1004);
and U691 (N_691,In_979,In_657);
nand U692 (N_692,In_941,In_614);
and U693 (N_693,In_1467,In_545);
nand U694 (N_694,In_1121,In_354);
nand U695 (N_695,In_272,In_960);
or U696 (N_696,In_959,In_1364);
nand U697 (N_697,In_72,In_1137);
or U698 (N_698,In_25,In_1477);
nand U699 (N_699,In_559,In_880);
nor U700 (N_700,In_1273,In_205);
nand U701 (N_701,In_1034,In_247);
nand U702 (N_702,In_458,In_1392);
nand U703 (N_703,In_1238,In_898);
nor U704 (N_704,In_1186,In_1235);
nor U705 (N_705,In_1056,In_1384);
or U706 (N_706,In_1023,In_485);
nor U707 (N_707,In_5,In_218);
and U708 (N_708,In_1365,In_878);
and U709 (N_709,In_681,In_673);
or U710 (N_710,In_372,In_1041);
nor U711 (N_711,In_1168,In_1378);
or U712 (N_712,In_490,In_453);
nor U713 (N_713,In_1096,In_570);
or U714 (N_714,In_1297,In_1456);
nand U715 (N_715,In_662,In_1076);
nand U716 (N_716,In_735,In_1117);
xnor U717 (N_717,In_245,In_766);
and U718 (N_718,In_598,In_1064);
nor U719 (N_719,In_923,In_932);
or U720 (N_720,In_1019,In_792);
xor U721 (N_721,In_1033,In_1146);
or U722 (N_722,In_314,In_1468);
nor U723 (N_723,In_788,In_678);
and U724 (N_724,In_592,In_76);
nor U725 (N_725,In_98,In_524);
nand U726 (N_726,In_16,In_802);
and U727 (N_727,In_760,In_405);
or U728 (N_728,In_472,In_465);
or U729 (N_729,In_605,In_137);
and U730 (N_730,In_1268,In_278);
nor U731 (N_731,In_814,In_981);
and U732 (N_732,In_256,In_65);
and U733 (N_733,In_503,In_1474);
or U734 (N_734,In_1150,In_1320);
nor U735 (N_735,In_1371,In_414);
and U736 (N_736,In_427,In_895);
nand U737 (N_737,In_1319,In_174);
nand U738 (N_738,In_1404,In_537);
nand U739 (N_739,In_1124,In_230);
or U740 (N_740,In_395,In_1005);
nand U741 (N_741,In_1440,In_1008);
and U742 (N_742,In_1334,In_597);
nand U743 (N_743,In_97,In_1337);
or U744 (N_744,In_226,In_787);
or U745 (N_745,In_1464,In_1148);
nor U746 (N_746,In_672,In_79);
xnor U747 (N_747,In_96,In_1282);
xnor U748 (N_748,In_436,In_887);
nor U749 (N_749,In_1274,In_1102);
or U750 (N_750,In_506,In_576);
and U751 (N_751,In_1335,In_851);
or U752 (N_752,In_427,In_617);
or U753 (N_753,In_114,In_941);
nand U754 (N_754,In_1069,In_848);
or U755 (N_755,In_271,In_243);
or U756 (N_756,In_445,In_460);
or U757 (N_757,In_688,In_1451);
and U758 (N_758,In_928,In_836);
and U759 (N_759,In_1288,In_1138);
or U760 (N_760,In_114,In_276);
and U761 (N_761,In_743,In_990);
or U762 (N_762,In_882,In_323);
and U763 (N_763,In_25,In_514);
xor U764 (N_764,In_1110,In_276);
nand U765 (N_765,In_1483,In_1309);
nor U766 (N_766,In_21,In_1285);
nor U767 (N_767,In_94,In_1092);
xnor U768 (N_768,In_1332,In_1060);
or U769 (N_769,In_327,In_23);
nor U770 (N_770,In_916,In_593);
and U771 (N_771,In_580,In_1169);
nand U772 (N_772,In_1266,In_225);
or U773 (N_773,In_456,In_335);
xnor U774 (N_774,In_1042,In_16);
and U775 (N_775,In_1027,In_133);
or U776 (N_776,In_617,In_1196);
or U777 (N_777,In_898,In_115);
or U778 (N_778,In_577,In_287);
nor U779 (N_779,In_923,In_567);
and U780 (N_780,In_16,In_1091);
and U781 (N_781,In_105,In_1270);
nor U782 (N_782,In_445,In_1063);
xnor U783 (N_783,In_406,In_229);
and U784 (N_784,In_50,In_250);
xor U785 (N_785,In_1055,In_575);
nand U786 (N_786,In_1018,In_1118);
nand U787 (N_787,In_959,In_373);
and U788 (N_788,In_936,In_492);
and U789 (N_789,In_680,In_1313);
xor U790 (N_790,In_946,In_1257);
and U791 (N_791,In_1167,In_1092);
nand U792 (N_792,In_1005,In_782);
nand U793 (N_793,In_512,In_174);
xor U794 (N_794,In_1325,In_1226);
or U795 (N_795,In_1113,In_1398);
nand U796 (N_796,In_1313,In_922);
and U797 (N_797,In_332,In_1266);
or U798 (N_798,In_431,In_708);
and U799 (N_799,In_887,In_180);
nand U800 (N_800,In_309,In_839);
nand U801 (N_801,In_156,In_967);
nand U802 (N_802,In_658,In_605);
nor U803 (N_803,In_1387,In_465);
nand U804 (N_804,In_1329,In_576);
xor U805 (N_805,In_580,In_638);
and U806 (N_806,In_148,In_1185);
nand U807 (N_807,In_538,In_735);
and U808 (N_808,In_613,In_931);
nor U809 (N_809,In_650,In_1092);
or U810 (N_810,In_155,In_818);
nand U811 (N_811,In_1486,In_761);
and U812 (N_812,In_874,In_1326);
and U813 (N_813,In_399,In_1107);
nand U814 (N_814,In_1138,In_692);
or U815 (N_815,In_873,In_1402);
nand U816 (N_816,In_1132,In_991);
xnor U817 (N_817,In_568,In_1221);
nor U818 (N_818,In_64,In_1215);
nor U819 (N_819,In_986,In_1077);
and U820 (N_820,In_559,In_30);
and U821 (N_821,In_289,In_1167);
or U822 (N_822,In_1465,In_297);
nand U823 (N_823,In_1364,In_1160);
or U824 (N_824,In_1305,In_855);
nor U825 (N_825,In_1316,In_656);
and U826 (N_826,In_1165,In_697);
and U827 (N_827,In_563,In_1448);
nor U828 (N_828,In_1200,In_589);
and U829 (N_829,In_244,In_841);
nand U830 (N_830,In_636,In_340);
nand U831 (N_831,In_1449,In_1433);
and U832 (N_832,In_545,In_754);
or U833 (N_833,In_910,In_1213);
nand U834 (N_834,In_563,In_1379);
and U835 (N_835,In_1378,In_407);
and U836 (N_836,In_1195,In_319);
and U837 (N_837,In_31,In_926);
nand U838 (N_838,In_38,In_680);
xor U839 (N_839,In_203,In_783);
or U840 (N_840,In_45,In_1394);
and U841 (N_841,In_1375,In_1287);
nand U842 (N_842,In_1154,In_1097);
and U843 (N_843,In_535,In_146);
nand U844 (N_844,In_299,In_839);
nand U845 (N_845,In_911,In_1058);
or U846 (N_846,In_1311,In_318);
and U847 (N_847,In_879,In_352);
nand U848 (N_848,In_703,In_832);
or U849 (N_849,In_1027,In_935);
nor U850 (N_850,In_1278,In_694);
nand U851 (N_851,In_586,In_617);
and U852 (N_852,In_756,In_619);
and U853 (N_853,In_613,In_1314);
nor U854 (N_854,In_618,In_714);
nand U855 (N_855,In_790,In_230);
xnor U856 (N_856,In_556,In_634);
nand U857 (N_857,In_1230,In_82);
nand U858 (N_858,In_1038,In_1121);
or U859 (N_859,In_808,In_251);
nand U860 (N_860,In_718,In_1261);
and U861 (N_861,In_1044,In_298);
and U862 (N_862,In_828,In_958);
and U863 (N_863,In_1484,In_961);
or U864 (N_864,In_140,In_395);
xnor U865 (N_865,In_276,In_226);
or U866 (N_866,In_597,In_1322);
or U867 (N_867,In_914,In_345);
or U868 (N_868,In_1181,In_63);
nor U869 (N_869,In_444,In_100);
xor U870 (N_870,In_118,In_1340);
nand U871 (N_871,In_1026,In_783);
nor U872 (N_872,In_454,In_422);
nand U873 (N_873,In_797,In_68);
nand U874 (N_874,In_1283,In_181);
xor U875 (N_875,In_561,In_248);
nand U876 (N_876,In_1222,In_1114);
xnor U877 (N_877,In_1161,In_576);
nand U878 (N_878,In_949,In_1224);
or U879 (N_879,In_1061,In_743);
nand U880 (N_880,In_291,In_1415);
or U881 (N_881,In_233,In_1353);
nand U882 (N_882,In_906,In_731);
nand U883 (N_883,In_945,In_175);
or U884 (N_884,In_573,In_1102);
xor U885 (N_885,In_850,In_268);
or U886 (N_886,In_1180,In_1342);
or U887 (N_887,In_1471,In_1031);
or U888 (N_888,In_1244,In_592);
or U889 (N_889,In_1184,In_1333);
and U890 (N_890,In_614,In_38);
nor U891 (N_891,In_269,In_916);
nand U892 (N_892,In_878,In_6);
and U893 (N_893,In_895,In_960);
nor U894 (N_894,In_1201,In_936);
nor U895 (N_895,In_11,In_1014);
and U896 (N_896,In_604,In_1341);
xor U897 (N_897,In_833,In_1347);
and U898 (N_898,In_1474,In_848);
nor U899 (N_899,In_307,In_111);
nor U900 (N_900,In_624,In_189);
nor U901 (N_901,In_735,In_751);
nand U902 (N_902,In_1087,In_523);
nand U903 (N_903,In_1256,In_955);
nand U904 (N_904,In_123,In_1112);
and U905 (N_905,In_137,In_382);
and U906 (N_906,In_139,In_1286);
and U907 (N_907,In_1318,In_1277);
nor U908 (N_908,In_128,In_277);
nor U909 (N_909,In_677,In_164);
xnor U910 (N_910,In_1274,In_1366);
and U911 (N_911,In_942,In_579);
or U912 (N_912,In_1333,In_423);
nor U913 (N_913,In_1283,In_1048);
nand U914 (N_914,In_1472,In_110);
and U915 (N_915,In_1446,In_163);
and U916 (N_916,In_164,In_425);
or U917 (N_917,In_451,In_779);
nand U918 (N_918,In_1426,In_936);
xnor U919 (N_919,In_685,In_348);
nand U920 (N_920,In_509,In_697);
nand U921 (N_921,In_776,In_1149);
nand U922 (N_922,In_1163,In_1027);
nand U923 (N_923,In_1497,In_140);
and U924 (N_924,In_269,In_784);
or U925 (N_925,In_1394,In_1071);
and U926 (N_926,In_163,In_1031);
nor U927 (N_927,In_1176,In_1414);
and U928 (N_928,In_1393,In_1142);
and U929 (N_929,In_1147,In_625);
or U930 (N_930,In_1139,In_256);
nor U931 (N_931,In_618,In_727);
nand U932 (N_932,In_25,In_159);
nor U933 (N_933,In_260,In_1390);
nor U934 (N_934,In_122,In_815);
xnor U935 (N_935,In_794,In_930);
nand U936 (N_936,In_158,In_1150);
nor U937 (N_937,In_140,In_1060);
nand U938 (N_938,In_357,In_1282);
or U939 (N_939,In_232,In_62);
nor U940 (N_940,In_386,In_547);
or U941 (N_941,In_404,In_1226);
or U942 (N_942,In_1328,In_1464);
nor U943 (N_943,In_1489,In_82);
xor U944 (N_944,In_1264,In_1027);
nor U945 (N_945,In_889,In_193);
or U946 (N_946,In_1077,In_329);
nor U947 (N_947,In_1317,In_891);
or U948 (N_948,In_833,In_204);
and U949 (N_949,In_386,In_530);
nor U950 (N_950,In_1103,In_117);
nand U951 (N_951,In_1008,In_149);
or U952 (N_952,In_947,In_224);
nand U953 (N_953,In_485,In_223);
nor U954 (N_954,In_1285,In_1000);
nor U955 (N_955,In_1283,In_473);
or U956 (N_956,In_1154,In_1359);
nand U957 (N_957,In_694,In_319);
or U958 (N_958,In_941,In_1016);
and U959 (N_959,In_692,In_1120);
or U960 (N_960,In_417,In_1431);
or U961 (N_961,In_1260,In_1471);
xor U962 (N_962,In_307,In_599);
nor U963 (N_963,In_635,In_1296);
or U964 (N_964,In_1006,In_1171);
and U965 (N_965,In_1103,In_1122);
and U966 (N_966,In_900,In_1402);
or U967 (N_967,In_1179,In_1082);
and U968 (N_968,In_1480,In_816);
nand U969 (N_969,In_449,In_983);
or U970 (N_970,In_1237,In_248);
nor U971 (N_971,In_577,In_532);
or U972 (N_972,In_1445,In_391);
nand U973 (N_973,In_1278,In_835);
or U974 (N_974,In_630,In_1450);
nand U975 (N_975,In_128,In_126);
nand U976 (N_976,In_1436,In_986);
nand U977 (N_977,In_797,In_449);
nand U978 (N_978,In_1113,In_100);
nor U979 (N_979,In_504,In_334);
and U980 (N_980,In_1094,In_411);
xor U981 (N_981,In_366,In_430);
or U982 (N_982,In_342,In_624);
or U983 (N_983,In_1306,In_332);
xnor U984 (N_984,In_1380,In_1264);
nand U985 (N_985,In_491,In_598);
nand U986 (N_986,In_1088,In_151);
nor U987 (N_987,In_87,In_101);
nand U988 (N_988,In_939,In_1217);
nand U989 (N_989,In_1134,In_1200);
or U990 (N_990,In_943,In_1313);
xor U991 (N_991,In_1149,In_1057);
and U992 (N_992,In_1222,In_617);
and U993 (N_993,In_397,In_181);
nand U994 (N_994,In_376,In_1410);
nor U995 (N_995,In_1250,In_1327);
nand U996 (N_996,In_1176,In_949);
nand U997 (N_997,In_511,In_631);
or U998 (N_998,In_614,In_450);
nand U999 (N_999,In_116,In_1185);
nand U1000 (N_1000,In_1438,In_869);
or U1001 (N_1001,In_323,In_705);
or U1002 (N_1002,In_625,In_648);
nand U1003 (N_1003,In_1197,In_122);
nor U1004 (N_1004,In_474,In_538);
nand U1005 (N_1005,In_1355,In_409);
nor U1006 (N_1006,In_214,In_156);
and U1007 (N_1007,In_862,In_264);
or U1008 (N_1008,In_1157,In_1400);
or U1009 (N_1009,In_599,In_1165);
and U1010 (N_1010,In_801,In_945);
and U1011 (N_1011,In_1011,In_379);
nor U1012 (N_1012,In_338,In_250);
nor U1013 (N_1013,In_1434,In_539);
nand U1014 (N_1014,In_641,In_20);
nor U1015 (N_1015,In_230,In_842);
nand U1016 (N_1016,In_1117,In_82);
or U1017 (N_1017,In_487,In_210);
nor U1018 (N_1018,In_539,In_95);
nor U1019 (N_1019,In_357,In_1236);
xnor U1020 (N_1020,In_442,In_386);
and U1021 (N_1021,In_1276,In_581);
or U1022 (N_1022,In_191,In_682);
or U1023 (N_1023,In_40,In_561);
and U1024 (N_1024,In_269,In_199);
nor U1025 (N_1025,In_165,In_753);
nor U1026 (N_1026,In_1462,In_462);
or U1027 (N_1027,In_84,In_953);
nand U1028 (N_1028,In_824,In_1270);
nand U1029 (N_1029,In_1030,In_969);
nand U1030 (N_1030,In_813,In_603);
nor U1031 (N_1031,In_163,In_1285);
nand U1032 (N_1032,In_733,In_102);
or U1033 (N_1033,In_862,In_1305);
nor U1034 (N_1034,In_1429,In_91);
and U1035 (N_1035,In_148,In_998);
nand U1036 (N_1036,In_956,In_1376);
and U1037 (N_1037,In_240,In_711);
nor U1038 (N_1038,In_1070,In_458);
and U1039 (N_1039,In_957,In_479);
and U1040 (N_1040,In_415,In_610);
or U1041 (N_1041,In_390,In_1498);
nand U1042 (N_1042,In_1184,In_251);
or U1043 (N_1043,In_961,In_1126);
nand U1044 (N_1044,In_1276,In_616);
nor U1045 (N_1045,In_236,In_371);
nand U1046 (N_1046,In_1132,In_273);
xnor U1047 (N_1047,In_385,In_1);
nor U1048 (N_1048,In_1324,In_960);
or U1049 (N_1049,In_1210,In_269);
and U1050 (N_1050,In_762,In_60);
or U1051 (N_1051,In_199,In_448);
and U1052 (N_1052,In_102,In_340);
or U1053 (N_1053,In_1304,In_472);
nor U1054 (N_1054,In_1443,In_918);
and U1055 (N_1055,In_1060,In_178);
or U1056 (N_1056,In_654,In_1309);
or U1057 (N_1057,In_1175,In_354);
and U1058 (N_1058,In_455,In_947);
nand U1059 (N_1059,In_1489,In_238);
nand U1060 (N_1060,In_812,In_471);
nor U1061 (N_1061,In_1316,In_451);
nand U1062 (N_1062,In_313,In_1262);
nor U1063 (N_1063,In_1381,In_341);
nand U1064 (N_1064,In_444,In_342);
and U1065 (N_1065,In_311,In_332);
or U1066 (N_1066,In_58,In_470);
nor U1067 (N_1067,In_601,In_1123);
or U1068 (N_1068,In_449,In_712);
or U1069 (N_1069,In_1265,In_1231);
nor U1070 (N_1070,In_919,In_1422);
xnor U1071 (N_1071,In_985,In_521);
nand U1072 (N_1072,In_1403,In_959);
nand U1073 (N_1073,In_466,In_790);
xnor U1074 (N_1074,In_121,In_1248);
nand U1075 (N_1075,In_486,In_414);
xor U1076 (N_1076,In_1230,In_405);
or U1077 (N_1077,In_1169,In_821);
xnor U1078 (N_1078,In_802,In_78);
and U1079 (N_1079,In_1290,In_783);
and U1080 (N_1080,In_413,In_576);
nor U1081 (N_1081,In_151,In_509);
or U1082 (N_1082,In_1278,In_160);
or U1083 (N_1083,In_137,In_1317);
nor U1084 (N_1084,In_1200,In_1067);
nor U1085 (N_1085,In_1335,In_1466);
and U1086 (N_1086,In_924,In_1366);
nor U1087 (N_1087,In_1146,In_234);
or U1088 (N_1088,In_240,In_1350);
and U1089 (N_1089,In_433,In_764);
nor U1090 (N_1090,In_1099,In_608);
nor U1091 (N_1091,In_1164,In_14);
and U1092 (N_1092,In_1168,In_397);
nor U1093 (N_1093,In_273,In_658);
nor U1094 (N_1094,In_1404,In_312);
and U1095 (N_1095,In_204,In_112);
or U1096 (N_1096,In_646,In_378);
nor U1097 (N_1097,In_405,In_957);
or U1098 (N_1098,In_32,In_356);
or U1099 (N_1099,In_18,In_26);
or U1100 (N_1100,In_1364,In_1412);
nor U1101 (N_1101,In_16,In_1458);
nand U1102 (N_1102,In_444,In_329);
nand U1103 (N_1103,In_1452,In_328);
and U1104 (N_1104,In_1180,In_960);
nor U1105 (N_1105,In_973,In_26);
nor U1106 (N_1106,In_136,In_85);
or U1107 (N_1107,In_611,In_1348);
nor U1108 (N_1108,In_933,In_804);
and U1109 (N_1109,In_299,In_495);
nor U1110 (N_1110,In_355,In_1278);
and U1111 (N_1111,In_969,In_1314);
nand U1112 (N_1112,In_218,In_247);
and U1113 (N_1113,In_1190,In_1445);
nand U1114 (N_1114,In_473,In_943);
nand U1115 (N_1115,In_394,In_798);
nand U1116 (N_1116,In_193,In_602);
and U1117 (N_1117,In_566,In_403);
or U1118 (N_1118,In_1004,In_1186);
or U1119 (N_1119,In_774,In_464);
or U1120 (N_1120,In_1149,In_398);
nor U1121 (N_1121,In_803,In_336);
nand U1122 (N_1122,In_764,In_823);
or U1123 (N_1123,In_278,In_1467);
and U1124 (N_1124,In_1298,In_864);
or U1125 (N_1125,In_226,In_1330);
and U1126 (N_1126,In_1248,In_333);
or U1127 (N_1127,In_121,In_284);
nand U1128 (N_1128,In_737,In_1231);
or U1129 (N_1129,In_634,In_1158);
or U1130 (N_1130,In_552,In_489);
and U1131 (N_1131,In_161,In_1280);
xnor U1132 (N_1132,In_901,In_1084);
nand U1133 (N_1133,In_866,In_1449);
nand U1134 (N_1134,In_490,In_1347);
or U1135 (N_1135,In_654,In_577);
and U1136 (N_1136,In_1255,In_1286);
nand U1137 (N_1137,In_517,In_785);
nor U1138 (N_1138,In_378,In_302);
and U1139 (N_1139,In_1168,In_998);
nor U1140 (N_1140,In_434,In_1267);
xnor U1141 (N_1141,In_148,In_1458);
or U1142 (N_1142,In_307,In_364);
and U1143 (N_1143,In_550,In_1074);
and U1144 (N_1144,In_1378,In_520);
or U1145 (N_1145,In_1462,In_1233);
nor U1146 (N_1146,In_521,In_540);
nor U1147 (N_1147,In_495,In_1112);
nand U1148 (N_1148,In_653,In_563);
nor U1149 (N_1149,In_1341,In_1428);
and U1150 (N_1150,In_473,In_1350);
and U1151 (N_1151,In_1144,In_989);
nor U1152 (N_1152,In_993,In_133);
nor U1153 (N_1153,In_741,In_1409);
or U1154 (N_1154,In_125,In_456);
nand U1155 (N_1155,In_1165,In_778);
and U1156 (N_1156,In_227,In_739);
or U1157 (N_1157,In_662,In_1017);
nand U1158 (N_1158,In_76,In_1431);
and U1159 (N_1159,In_76,In_1019);
or U1160 (N_1160,In_925,In_633);
and U1161 (N_1161,In_1390,In_1463);
xnor U1162 (N_1162,In_1181,In_1068);
nor U1163 (N_1163,In_1344,In_761);
and U1164 (N_1164,In_1173,In_588);
nor U1165 (N_1165,In_1494,In_436);
and U1166 (N_1166,In_1202,In_120);
and U1167 (N_1167,In_648,In_1108);
and U1168 (N_1168,In_1275,In_1044);
and U1169 (N_1169,In_1426,In_1499);
xnor U1170 (N_1170,In_1318,In_1360);
nor U1171 (N_1171,In_530,In_595);
or U1172 (N_1172,In_1217,In_84);
nand U1173 (N_1173,In_1101,In_1157);
and U1174 (N_1174,In_897,In_827);
nand U1175 (N_1175,In_320,In_1225);
nor U1176 (N_1176,In_222,In_200);
or U1177 (N_1177,In_1326,In_1361);
xor U1178 (N_1178,In_1345,In_82);
nand U1179 (N_1179,In_196,In_1209);
nor U1180 (N_1180,In_877,In_1419);
or U1181 (N_1181,In_1312,In_1332);
nand U1182 (N_1182,In_494,In_1163);
or U1183 (N_1183,In_511,In_472);
or U1184 (N_1184,In_837,In_1153);
nand U1185 (N_1185,In_1129,In_1113);
xnor U1186 (N_1186,In_312,In_1020);
xor U1187 (N_1187,In_1211,In_321);
or U1188 (N_1188,In_738,In_595);
nand U1189 (N_1189,In_363,In_263);
nor U1190 (N_1190,In_1048,In_908);
nor U1191 (N_1191,In_824,In_776);
and U1192 (N_1192,In_126,In_508);
and U1193 (N_1193,In_212,In_1015);
or U1194 (N_1194,In_1461,In_368);
nand U1195 (N_1195,In_704,In_1054);
and U1196 (N_1196,In_163,In_1039);
nand U1197 (N_1197,In_1091,In_1282);
xnor U1198 (N_1198,In_1143,In_792);
and U1199 (N_1199,In_848,In_138);
and U1200 (N_1200,In_1495,In_1410);
or U1201 (N_1201,In_102,In_1458);
nor U1202 (N_1202,In_588,In_346);
xor U1203 (N_1203,In_312,In_319);
nor U1204 (N_1204,In_1064,In_548);
nor U1205 (N_1205,In_19,In_924);
nor U1206 (N_1206,In_1185,In_473);
or U1207 (N_1207,In_1011,In_1493);
and U1208 (N_1208,In_938,In_878);
nand U1209 (N_1209,In_228,In_339);
and U1210 (N_1210,In_724,In_600);
and U1211 (N_1211,In_1159,In_12);
and U1212 (N_1212,In_1008,In_1477);
nand U1213 (N_1213,In_1365,In_341);
nor U1214 (N_1214,In_386,In_19);
and U1215 (N_1215,In_1211,In_1369);
and U1216 (N_1216,In_766,In_697);
nand U1217 (N_1217,In_1250,In_431);
xor U1218 (N_1218,In_129,In_107);
nor U1219 (N_1219,In_209,In_324);
and U1220 (N_1220,In_828,In_242);
and U1221 (N_1221,In_263,In_62);
nor U1222 (N_1222,In_1198,In_1199);
and U1223 (N_1223,In_1191,In_1383);
or U1224 (N_1224,In_1365,In_106);
nor U1225 (N_1225,In_736,In_1413);
or U1226 (N_1226,In_1073,In_1365);
nand U1227 (N_1227,In_287,In_818);
nor U1228 (N_1228,In_289,In_1276);
and U1229 (N_1229,In_634,In_612);
or U1230 (N_1230,In_660,In_1220);
nor U1231 (N_1231,In_1097,In_1292);
or U1232 (N_1232,In_341,In_1447);
xor U1233 (N_1233,In_1063,In_55);
nand U1234 (N_1234,In_1089,In_1346);
and U1235 (N_1235,In_1054,In_423);
or U1236 (N_1236,In_166,In_1046);
and U1237 (N_1237,In_354,In_739);
or U1238 (N_1238,In_1390,In_1349);
nor U1239 (N_1239,In_1389,In_856);
nand U1240 (N_1240,In_667,In_1191);
or U1241 (N_1241,In_903,In_1332);
nand U1242 (N_1242,In_1376,In_1378);
and U1243 (N_1243,In_1171,In_456);
nor U1244 (N_1244,In_1022,In_635);
and U1245 (N_1245,In_850,In_171);
nand U1246 (N_1246,In_1016,In_1242);
and U1247 (N_1247,In_1403,In_1368);
or U1248 (N_1248,In_758,In_1219);
nor U1249 (N_1249,In_409,In_320);
or U1250 (N_1250,In_317,In_629);
or U1251 (N_1251,In_888,In_193);
nor U1252 (N_1252,In_807,In_427);
nand U1253 (N_1253,In_481,In_238);
nor U1254 (N_1254,In_1127,In_186);
and U1255 (N_1255,In_146,In_687);
nor U1256 (N_1256,In_87,In_1401);
or U1257 (N_1257,In_1146,In_765);
and U1258 (N_1258,In_506,In_81);
nand U1259 (N_1259,In_108,In_1224);
and U1260 (N_1260,In_115,In_858);
or U1261 (N_1261,In_319,In_1413);
nand U1262 (N_1262,In_559,In_1451);
nor U1263 (N_1263,In_711,In_620);
or U1264 (N_1264,In_1097,In_705);
and U1265 (N_1265,In_815,In_238);
nor U1266 (N_1266,In_152,In_661);
nor U1267 (N_1267,In_951,In_132);
and U1268 (N_1268,In_688,In_45);
nor U1269 (N_1269,In_311,In_418);
or U1270 (N_1270,In_1104,In_1397);
nor U1271 (N_1271,In_1230,In_472);
nand U1272 (N_1272,In_1214,In_1108);
or U1273 (N_1273,In_1421,In_1262);
and U1274 (N_1274,In_387,In_1423);
or U1275 (N_1275,In_985,In_667);
xor U1276 (N_1276,In_373,In_461);
and U1277 (N_1277,In_1386,In_577);
and U1278 (N_1278,In_805,In_494);
nor U1279 (N_1279,In_1025,In_865);
and U1280 (N_1280,In_278,In_158);
xnor U1281 (N_1281,In_401,In_1194);
nor U1282 (N_1282,In_302,In_718);
nor U1283 (N_1283,In_1013,In_381);
nand U1284 (N_1284,In_1103,In_659);
or U1285 (N_1285,In_872,In_473);
nor U1286 (N_1286,In_1474,In_729);
and U1287 (N_1287,In_271,In_442);
and U1288 (N_1288,In_119,In_287);
or U1289 (N_1289,In_198,In_696);
or U1290 (N_1290,In_587,In_1458);
xnor U1291 (N_1291,In_687,In_1242);
and U1292 (N_1292,In_1115,In_1057);
or U1293 (N_1293,In_324,In_474);
nor U1294 (N_1294,In_998,In_85);
nand U1295 (N_1295,In_1227,In_725);
nor U1296 (N_1296,In_405,In_919);
nor U1297 (N_1297,In_142,In_38);
or U1298 (N_1298,In_540,In_152);
xor U1299 (N_1299,In_653,In_364);
nor U1300 (N_1300,In_1146,In_1172);
nor U1301 (N_1301,In_1334,In_34);
and U1302 (N_1302,In_123,In_1088);
nand U1303 (N_1303,In_1415,In_1160);
or U1304 (N_1304,In_1100,In_1024);
nor U1305 (N_1305,In_855,In_1260);
or U1306 (N_1306,In_997,In_1366);
nand U1307 (N_1307,In_915,In_1496);
or U1308 (N_1308,In_568,In_165);
nand U1309 (N_1309,In_301,In_605);
xnor U1310 (N_1310,In_47,In_1265);
or U1311 (N_1311,In_1123,In_508);
and U1312 (N_1312,In_816,In_111);
nor U1313 (N_1313,In_327,In_292);
xor U1314 (N_1314,In_596,In_250);
nor U1315 (N_1315,In_746,In_335);
or U1316 (N_1316,In_1475,In_471);
or U1317 (N_1317,In_867,In_1111);
nand U1318 (N_1318,In_608,In_563);
or U1319 (N_1319,In_812,In_1037);
or U1320 (N_1320,In_554,In_634);
and U1321 (N_1321,In_72,In_441);
nand U1322 (N_1322,In_1297,In_1442);
nand U1323 (N_1323,In_25,In_1065);
or U1324 (N_1324,In_438,In_1499);
and U1325 (N_1325,In_1447,In_993);
or U1326 (N_1326,In_1476,In_616);
and U1327 (N_1327,In_264,In_891);
nor U1328 (N_1328,In_878,In_1218);
and U1329 (N_1329,In_1122,In_1258);
and U1330 (N_1330,In_404,In_804);
nor U1331 (N_1331,In_933,In_993);
nor U1332 (N_1332,In_1373,In_690);
and U1333 (N_1333,In_1161,In_230);
nand U1334 (N_1334,In_885,In_1236);
or U1335 (N_1335,In_1355,In_234);
nand U1336 (N_1336,In_1330,In_237);
or U1337 (N_1337,In_1252,In_1166);
nor U1338 (N_1338,In_177,In_233);
and U1339 (N_1339,In_57,In_578);
nand U1340 (N_1340,In_1389,In_1117);
nand U1341 (N_1341,In_376,In_367);
or U1342 (N_1342,In_843,In_744);
or U1343 (N_1343,In_107,In_627);
or U1344 (N_1344,In_375,In_729);
and U1345 (N_1345,In_668,In_1375);
and U1346 (N_1346,In_1367,In_278);
nor U1347 (N_1347,In_1377,In_1012);
and U1348 (N_1348,In_1269,In_1464);
or U1349 (N_1349,In_111,In_712);
and U1350 (N_1350,In_168,In_618);
and U1351 (N_1351,In_679,In_1045);
and U1352 (N_1352,In_73,In_1176);
nor U1353 (N_1353,In_530,In_1437);
nor U1354 (N_1354,In_1183,In_1118);
xnor U1355 (N_1355,In_1359,In_556);
nor U1356 (N_1356,In_487,In_973);
xnor U1357 (N_1357,In_643,In_1345);
and U1358 (N_1358,In_360,In_1411);
xor U1359 (N_1359,In_686,In_407);
or U1360 (N_1360,In_101,In_544);
nor U1361 (N_1361,In_436,In_1136);
xnor U1362 (N_1362,In_48,In_967);
nand U1363 (N_1363,In_538,In_243);
nand U1364 (N_1364,In_56,In_55);
or U1365 (N_1365,In_203,In_256);
nor U1366 (N_1366,In_1075,In_1108);
nor U1367 (N_1367,In_1395,In_1445);
and U1368 (N_1368,In_1066,In_141);
nand U1369 (N_1369,In_504,In_1432);
and U1370 (N_1370,In_367,In_382);
xnor U1371 (N_1371,In_1367,In_342);
and U1372 (N_1372,In_784,In_432);
and U1373 (N_1373,In_1257,In_967);
and U1374 (N_1374,In_1084,In_1293);
or U1375 (N_1375,In_261,In_385);
and U1376 (N_1376,In_1464,In_990);
nor U1377 (N_1377,In_81,In_1484);
nand U1378 (N_1378,In_1312,In_1226);
xnor U1379 (N_1379,In_302,In_200);
and U1380 (N_1380,In_1210,In_275);
nand U1381 (N_1381,In_10,In_249);
and U1382 (N_1382,In_614,In_330);
nand U1383 (N_1383,In_1496,In_854);
nand U1384 (N_1384,In_493,In_212);
nand U1385 (N_1385,In_647,In_1322);
xnor U1386 (N_1386,In_124,In_16);
xor U1387 (N_1387,In_195,In_340);
and U1388 (N_1388,In_844,In_1457);
nand U1389 (N_1389,In_743,In_27);
nor U1390 (N_1390,In_1457,In_284);
xor U1391 (N_1391,In_1266,In_717);
nor U1392 (N_1392,In_776,In_1122);
or U1393 (N_1393,In_1180,In_749);
xnor U1394 (N_1394,In_32,In_1039);
and U1395 (N_1395,In_547,In_862);
and U1396 (N_1396,In_432,In_1236);
xor U1397 (N_1397,In_1291,In_257);
nor U1398 (N_1398,In_988,In_362);
nand U1399 (N_1399,In_628,In_528);
nand U1400 (N_1400,In_112,In_383);
and U1401 (N_1401,In_459,In_899);
and U1402 (N_1402,In_417,In_807);
and U1403 (N_1403,In_1182,In_130);
nand U1404 (N_1404,In_733,In_625);
nor U1405 (N_1405,In_863,In_284);
or U1406 (N_1406,In_1479,In_978);
and U1407 (N_1407,In_59,In_1064);
nand U1408 (N_1408,In_449,In_755);
nand U1409 (N_1409,In_1283,In_493);
xor U1410 (N_1410,In_1251,In_1090);
and U1411 (N_1411,In_25,In_1403);
nor U1412 (N_1412,In_1012,In_198);
and U1413 (N_1413,In_667,In_1051);
nand U1414 (N_1414,In_109,In_868);
and U1415 (N_1415,In_478,In_1443);
nand U1416 (N_1416,In_793,In_988);
and U1417 (N_1417,In_893,In_651);
xnor U1418 (N_1418,In_1071,In_535);
nand U1419 (N_1419,In_267,In_662);
and U1420 (N_1420,In_1030,In_98);
nand U1421 (N_1421,In_347,In_1390);
xnor U1422 (N_1422,In_17,In_196);
or U1423 (N_1423,In_543,In_1037);
or U1424 (N_1424,In_1025,In_1496);
and U1425 (N_1425,In_133,In_1200);
nand U1426 (N_1426,In_1095,In_906);
or U1427 (N_1427,In_569,In_543);
nor U1428 (N_1428,In_1080,In_190);
or U1429 (N_1429,In_742,In_474);
or U1430 (N_1430,In_768,In_108);
or U1431 (N_1431,In_581,In_458);
and U1432 (N_1432,In_1113,In_1316);
nor U1433 (N_1433,In_1369,In_558);
xnor U1434 (N_1434,In_937,In_1358);
nand U1435 (N_1435,In_1126,In_777);
or U1436 (N_1436,In_199,In_538);
nor U1437 (N_1437,In_1327,In_419);
nor U1438 (N_1438,In_1338,In_664);
or U1439 (N_1439,In_982,In_1451);
nor U1440 (N_1440,In_553,In_875);
and U1441 (N_1441,In_601,In_972);
or U1442 (N_1442,In_914,In_596);
nor U1443 (N_1443,In_10,In_788);
or U1444 (N_1444,In_1311,In_688);
and U1445 (N_1445,In_699,In_1054);
nand U1446 (N_1446,In_786,In_175);
and U1447 (N_1447,In_1098,In_900);
or U1448 (N_1448,In_715,In_883);
nand U1449 (N_1449,In_1298,In_12);
or U1450 (N_1450,In_1088,In_1368);
xor U1451 (N_1451,In_1191,In_550);
nor U1452 (N_1452,In_497,In_1309);
or U1453 (N_1453,In_415,In_564);
and U1454 (N_1454,In_1110,In_835);
xor U1455 (N_1455,In_913,In_297);
and U1456 (N_1456,In_479,In_236);
or U1457 (N_1457,In_326,In_1139);
nor U1458 (N_1458,In_1309,In_491);
nand U1459 (N_1459,In_1373,In_563);
and U1460 (N_1460,In_908,In_1483);
or U1461 (N_1461,In_327,In_1307);
or U1462 (N_1462,In_227,In_807);
nor U1463 (N_1463,In_1039,In_576);
and U1464 (N_1464,In_1227,In_397);
nor U1465 (N_1465,In_176,In_1033);
nand U1466 (N_1466,In_322,In_711);
xor U1467 (N_1467,In_686,In_452);
nor U1468 (N_1468,In_576,In_900);
or U1469 (N_1469,In_1180,In_492);
xor U1470 (N_1470,In_315,In_1022);
and U1471 (N_1471,In_1273,In_64);
or U1472 (N_1472,In_694,In_499);
nor U1473 (N_1473,In_574,In_837);
and U1474 (N_1474,In_817,In_1407);
or U1475 (N_1475,In_694,In_816);
or U1476 (N_1476,In_1218,In_1313);
xor U1477 (N_1477,In_286,In_235);
and U1478 (N_1478,In_1210,In_581);
nor U1479 (N_1479,In_467,In_1256);
or U1480 (N_1480,In_730,In_102);
and U1481 (N_1481,In_757,In_1227);
and U1482 (N_1482,In_237,In_1339);
xnor U1483 (N_1483,In_110,In_577);
nand U1484 (N_1484,In_301,In_1377);
or U1485 (N_1485,In_325,In_403);
and U1486 (N_1486,In_681,In_205);
nor U1487 (N_1487,In_1215,In_109);
nor U1488 (N_1488,In_1047,In_648);
nor U1489 (N_1489,In_82,In_90);
nand U1490 (N_1490,In_648,In_734);
nand U1491 (N_1491,In_1027,In_1258);
or U1492 (N_1492,In_303,In_1380);
nor U1493 (N_1493,In_605,In_1137);
or U1494 (N_1494,In_931,In_898);
and U1495 (N_1495,In_1066,In_11);
and U1496 (N_1496,In_570,In_747);
xnor U1497 (N_1497,In_323,In_816);
and U1498 (N_1498,In_1329,In_317);
nor U1499 (N_1499,In_1343,In_450);
nor U1500 (N_1500,In_801,In_694);
and U1501 (N_1501,In_1099,In_144);
nand U1502 (N_1502,In_1050,In_1235);
or U1503 (N_1503,In_850,In_1093);
and U1504 (N_1504,In_1312,In_554);
xor U1505 (N_1505,In_518,In_980);
nand U1506 (N_1506,In_272,In_290);
xnor U1507 (N_1507,In_686,In_1464);
or U1508 (N_1508,In_323,In_606);
nand U1509 (N_1509,In_237,In_193);
and U1510 (N_1510,In_580,In_968);
or U1511 (N_1511,In_831,In_46);
and U1512 (N_1512,In_1240,In_817);
or U1513 (N_1513,In_1331,In_72);
nand U1514 (N_1514,In_1380,In_1452);
nand U1515 (N_1515,In_172,In_51);
xnor U1516 (N_1516,In_336,In_1372);
or U1517 (N_1517,In_1429,In_1448);
nor U1518 (N_1518,In_1344,In_1377);
xor U1519 (N_1519,In_1038,In_800);
nand U1520 (N_1520,In_207,In_1375);
or U1521 (N_1521,In_734,In_1389);
or U1522 (N_1522,In_475,In_827);
or U1523 (N_1523,In_211,In_361);
or U1524 (N_1524,In_1181,In_102);
and U1525 (N_1525,In_1044,In_842);
nor U1526 (N_1526,In_354,In_1488);
nor U1527 (N_1527,In_605,In_1175);
and U1528 (N_1528,In_516,In_1172);
or U1529 (N_1529,In_6,In_1196);
nand U1530 (N_1530,In_629,In_135);
and U1531 (N_1531,In_194,In_1487);
and U1532 (N_1532,In_513,In_324);
nand U1533 (N_1533,In_94,In_0);
and U1534 (N_1534,In_1305,In_368);
or U1535 (N_1535,In_17,In_876);
nand U1536 (N_1536,In_207,In_1287);
and U1537 (N_1537,In_622,In_1228);
nor U1538 (N_1538,In_1269,In_1463);
and U1539 (N_1539,In_215,In_160);
and U1540 (N_1540,In_1276,In_920);
or U1541 (N_1541,In_650,In_983);
xnor U1542 (N_1542,In_1075,In_244);
and U1543 (N_1543,In_757,In_841);
nand U1544 (N_1544,In_980,In_850);
nor U1545 (N_1545,In_360,In_1159);
nor U1546 (N_1546,In_1133,In_316);
nand U1547 (N_1547,In_381,In_1135);
nand U1548 (N_1548,In_1180,In_855);
nor U1549 (N_1549,In_198,In_574);
nand U1550 (N_1550,In_442,In_155);
or U1551 (N_1551,In_809,In_68);
or U1552 (N_1552,In_978,In_28);
or U1553 (N_1553,In_80,In_42);
nor U1554 (N_1554,In_277,In_582);
nand U1555 (N_1555,In_880,In_1265);
and U1556 (N_1556,In_439,In_296);
nand U1557 (N_1557,In_334,In_415);
nor U1558 (N_1558,In_535,In_949);
or U1559 (N_1559,In_1257,In_463);
nor U1560 (N_1560,In_270,In_1122);
or U1561 (N_1561,In_1291,In_571);
or U1562 (N_1562,In_405,In_981);
or U1563 (N_1563,In_337,In_444);
nand U1564 (N_1564,In_426,In_83);
nor U1565 (N_1565,In_1188,In_797);
nand U1566 (N_1566,In_941,In_197);
or U1567 (N_1567,In_610,In_335);
and U1568 (N_1568,In_681,In_1034);
and U1569 (N_1569,In_428,In_516);
nand U1570 (N_1570,In_156,In_972);
nor U1571 (N_1571,In_973,In_48);
nand U1572 (N_1572,In_522,In_392);
nor U1573 (N_1573,In_1423,In_1169);
and U1574 (N_1574,In_784,In_707);
nand U1575 (N_1575,In_830,In_558);
or U1576 (N_1576,In_302,In_1434);
nand U1577 (N_1577,In_1285,In_98);
nand U1578 (N_1578,In_1362,In_1135);
nand U1579 (N_1579,In_83,In_1242);
nand U1580 (N_1580,In_577,In_935);
or U1581 (N_1581,In_725,In_1010);
nand U1582 (N_1582,In_1111,In_478);
or U1583 (N_1583,In_509,In_726);
or U1584 (N_1584,In_701,In_139);
and U1585 (N_1585,In_825,In_627);
and U1586 (N_1586,In_1067,In_1116);
and U1587 (N_1587,In_178,In_543);
xor U1588 (N_1588,In_808,In_1075);
nor U1589 (N_1589,In_863,In_463);
and U1590 (N_1590,In_1350,In_967);
nor U1591 (N_1591,In_43,In_1397);
xnor U1592 (N_1592,In_360,In_486);
or U1593 (N_1593,In_584,In_162);
or U1594 (N_1594,In_324,In_1102);
and U1595 (N_1595,In_159,In_1403);
or U1596 (N_1596,In_1137,In_414);
nor U1597 (N_1597,In_622,In_258);
nor U1598 (N_1598,In_524,In_772);
or U1599 (N_1599,In_991,In_1416);
nand U1600 (N_1600,In_988,In_617);
and U1601 (N_1601,In_782,In_260);
and U1602 (N_1602,In_1239,In_353);
or U1603 (N_1603,In_418,In_343);
nand U1604 (N_1604,In_128,In_583);
or U1605 (N_1605,In_1114,In_477);
nor U1606 (N_1606,In_948,In_1184);
nor U1607 (N_1607,In_1199,In_60);
and U1608 (N_1608,In_1359,In_439);
or U1609 (N_1609,In_994,In_416);
nor U1610 (N_1610,In_611,In_1095);
nand U1611 (N_1611,In_385,In_93);
nor U1612 (N_1612,In_1023,In_1356);
or U1613 (N_1613,In_90,In_648);
and U1614 (N_1614,In_206,In_420);
nand U1615 (N_1615,In_1309,In_956);
and U1616 (N_1616,In_153,In_1228);
and U1617 (N_1617,In_683,In_1499);
nor U1618 (N_1618,In_331,In_312);
nor U1619 (N_1619,In_1059,In_1377);
or U1620 (N_1620,In_40,In_1219);
and U1621 (N_1621,In_1092,In_389);
nor U1622 (N_1622,In_1438,In_134);
xor U1623 (N_1623,In_1201,In_1121);
nand U1624 (N_1624,In_1363,In_80);
nand U1625 (N_1625,In_849,In_687);
or U1626 (N_1626,In_845,In_1342);
or U1627 (N_1627,In_713,In_229);
nor U1628 (N_1628,In_935,In_372);
or U1629 (N_1629,In_532,In_683);
or U1630 (N_1630,In_348,In_1246);
and U1631 (N_1631,In_854,In_400);
or U1632 (N_1632,In_408,In_967);
or U1633 (N_1633,In_973,In_1435);
xor U1634 (N_1634,In_781,In_260);
nor U1635 (N_1635,In_179,In_859);
nand U1636 (N_1636,In_195,In_471);
nor U1637 (N_1637,In_573,In_683);
and U1638 (N_1638,In_176,In_1219);
and U1639 (N_1639,In_498,In_530);
nor U1640 (N_1640,In_882,In_218);
or U1641 (N_1641,In_220,In_1095);
nand U1642 (N_1642,In_256,In_40);
nor U1643 (N_1643,In_1049,In_784);
or U1644 (N_1644,In_863,In_375);
nor U1645 (N_1645,In_104,In_1103);
nand U1646 (N_1646,In_1147,In_750);
nand U1647 (N_1647,In_907,In_852);
nand U1648 (N_1648,In_671,In_166);
nor U1649 (N_1649,In_1169,In_648);
nand U1650 (N_1650,In_45,In_1099);
and U1651 (N_1651,In_1492,In_691);
nand U1652 (N_1652,In_569,In_310);
or U1653 (N_1653,In_715,In_710);
nor U1654 (N_1654,In_1241,In_1002);
and U1655 (N_1655,In_990,In_125);
nor U1656 (N_1656,In_373,In_389);
nor U1657 (N_1657,In_128,In_961);
or U1658 (N_1658,In_1028,In_105);
nand U1659 (N_1659,In_812,In_1070);
and U1660 (N_1660,In_1259,In_401);
xnor U1661 (N_1661,In_1225,In_1244);
xnor U1662 (N_1662,In_939,In_1155);
nand U1663 (N_1663,In_1044,In_787);
nand U1664 (N_1664,In_374,In_732);
nor U1665 (N_1665,In_212,In_1393);
nor U1666 (N_1666,In_1331,In_660);
and U1667 (N_1667,In_728,In_775);
and U1668 (N_1668,In_711,In_591);
or U1669 (N_1669,In_5,In_1023);
xor U1670 (N_1670,In_466,In_794);
or U1671 (N_1671,In_1276,In_49);
nand U1672 (N_1672,In_1189,In_134);
nand U1673 (N_1673,In_1000,In_1421);
nor U1674 (N_1674,In_1201,In_240);
and U1675 (N_1675,In_122,In_684);
or U1676 (N_1676,In_74,In_929);
and U1677 (N_1677,In_628,In_317);
or U1678 (N_1678,In_972,In_481);
nor U1679 (N_1679,In_795,In_396);
and U1680 (N_1680,In_1185,In_862);
and U1681 (N_1681,In_1452,In_1248);
nand U1682 (N_1682,In_275,In_786);
nor U1683 (N_1683,In_1286,In_690);
nand U1684 (N_1684,In_169,In_698);
nand U1685 (N_1685,In_1000,In_853);
nor U1686 (N_1686,In_1185,In_370);
nand U1687 (N_1687,In_159,In_732);
xnor U1688 (N_1688,In_125,In_1402);
or U1689 (N_1689,In_1377,In_1252);
and U1690 (N_1690,In_678,In_1489);
nand U1691 (N_1691,In_1047,In_417);
nor U1692 (N_1692,In_1169,In_431);
nand U1693 (N_1693,In_477,In_185);
nor U1694 (N_1694,In_1384,In_374);
or U1695 (N_1695,In_1069,In_888);
nor U1696 (N_1696,In_925,In_587);
nand U1697 (N_1697,In_1031,In_750);
nand U1698 (N_1698,In_824,In_379);
and U1699 (N_1699,In_406,In_1484);
nand U1700 (N_1700,In_1390,In_1150);
nand U1701 (N_1701,In_315,In_1077);
nor U1702 (N_1702,In_162,In_717);
nand U1703 (N_1703,In_1004,In_646);
nand U1704 (N_1704,In_135,In_831);
or U1705 (N_1705,In_816,In_603);
nand U1706 (N_1706,In_763,In_1269);
or U1707 (N_1707,In_521,In_185);
nand U1708 (N_1708,In_924,In_1018);
nor U1709 (N_1709,In_487,In_1149);
or U1710 (N_1710,In_1275,In_936);
xnor U1711 (N_1711,In_403,In_451);
nand U1712 (N_1712,In_1434,In_591);
and U1713 (N_1713,In_517,In_410);
xnor U1714 (N_1714,In_746,In_1463);
and U1715 (N_1715,In_578,In_849);
xnor U1716 (N_1716,In_1385,In_146);
nand U1717 (N_1717,In_1288,In_584);
nor U1718 (N_1718,In_867,In_405);
nand U1719 (N_1719,In_48,In_960);
nor U1720 (N_1720,In_52,In_65);
nor U1721 (N_1721,In_450,In_53);
and U1722 (N_1722,In_387,In_499);
nand U1723 (N_1723,In_151,In_1314);
and U1724 (N_1724,In_991,In_976);
or U1725 (N_1725,In_965,In_158);
nor U1726 (N_1726,In_1014,In_419);
or U1727 (N_1727,In_213,In_1400);
nor U1728 (N_1728,In_527,In_1124);
and U1729 (N_1729,In_39,In_1278);
nor U1730 (N_1730,In_12,In_149);
nor U1731 (N_1731,In_792,In_693);
and U1732 (N_1732,In_974,In_94);
nor U1733 (N_1733,In_1428,In_541);
and U1734 (N_1734,In_528,In_533);
and U1735 (N_1735,In_601,In_215);
or U1736 (N_1736,In_1021,In_348);
nand U1737 (N_1737,In_917,In_646);
nand U1738 (N_1738,In_901,In_296);
and U1739 (N_1739,In_785,In_1364);
nand U1740 (N_1740,In_180,In_44);
nand U1741 (N_1741,In_1239,In_194);
nor U1742 (N_1742,In_693,In_1356);
or U1743 (N_1743,In_1433,In_292);
nand U1744 (N_1744,In_486,In_834);
and U1745 (N_1745,In_928,In_701);
and U1746 (N_1746,In_1134,In_1358);
nor U1747 (N_1747,In_122,In_1243);
xor U1748 (N_1748,In_834,In_1393);
and U1749 (N_1749,In_360,In_518);
nand U1750 (N_1750,In_1489,In_729);
nor U1751 (N_1751,In_389,In_438);
nor U1752 (N_1752,In_1067,In_683);
xnor U1753 (N_1753,In_638,In_1250);
nor U1754 (N_1754,In_1256,In_663);
or U1755 (N_1755,In_161,In_1348);
or U1756 (N_1756,In_875,In_846);
nor U1757 (N_1757,In_564,In_947);
nor U1758 (N_1758,In_314,In_41);
nand U1759 (N_1759,In_43,In_1334);
xor U1760 (N_1760,In_1325,In_1180);
and U1761 (N_1761,In_550,In_392);
xor U1762 (N_1762,In_771,In_225);
xor U1763 (N_1763,In_708,In_123);
and U1764 (N_1764,In_798,In_230);
xor U1765 (N_1765,In_689,In_165);
or U1766 (N_1766,In_865,In_230);
nor U1767 (N_1767,In_1209,In_1086);
and U1768 (N_1768,In_1415,In_495);
nand U1769 (N_1769,In_684,In_364);
xor U1770 (N_1770,In_1158,In_530);
nor U1771 (N_1771,In_1446,In_988);
nand U1772 (N_1772,In_567,In_1192);
nand U1773 (N_1773,In_784,In_1405);
nand U1774 (N_1774,In_1221,In_412);
and U1775 (N_1775,In_44,In_297);
and U1776 (N_1776,In_1061,In_722);
nand U1777 (N_1777,In_1332,In_1334);
and U1778 (N_1778,In_1139,In_500);
nor U1779 (N_1779,In_850,In_605);
nand U1780 (N_1780,In_1385,In_291);
nand U1781 (N_1781,In_852,In_319);
or U1782 (N_1782,In_286,In_894);
and U1783 (N_1783,In_913,In_1323);
or U1784 (N_1784,In_748,In_859);
or U1785 (N_1785,In_1393,In_1047);
and U1786 (N_1786,In_322,In_1407);
nor U1787 (N_1787,In_1316,In_1060);
and U1788 (N_1788,In_868,In_1086);
nor U1789 (N_1789,In_1316,In_622);
and U1790 (N_1790,In_783,In_1167);
nand U1791 (N_1791,In_1126,In_1103);
nand U1792 (N_1792,In_209,In_986);
nor U1793 (N_1793,In_541,In_400);
and U1794 (N_1794,In_837,In_1451);
nand U1795 (N_1795,In_7,In_1231);
nor U1796 (N_1796,In_698,In_1284);
and U1797 (N_1797,In_1087,In_1098);
nand U1798 (N_1798,In_326,In_1286);
nor U1799 (N_1799,In_1188,In_300);
or U1800 (N_1800,In_1487,In_772);
xor U1801 (N_1801,In_290,In_792);
nand U1802 (N_1802,In_1060,In_1322);
and U1803 (N_1803,In_1344,In_1363);
nand U1804 (N_1804,In_313,In_1454);
or U1805 (N_1805,In_342,In_110);
and U1806 (N_1806,In_138,In_1196);
and U1807 (N_1807,In_45,In_27);
and U1808 (N_1808,In_702,In_1054);
and U1809 (N_1809,In_819,In_1301);
nand U1810 (N_1810,In_220,In_934);
and U1811 (N_1811,In_608,In_269);
nand U1812 (N_1812,In_869,In_485);
and U1813 (N_1813,In_1239,In_1023);
nand U1814 (N_1814,In_1421,In_666);
and U1815 (N_1815,In_1087,In_555);
or U1816 (N_1816,In_1355,In_1379);
and U1817 (N_1817,In_308,In_270);
xor U1818 (N_1818,In_1448,In_649);
xor U1819 (N_1819,In_1244,In_1341);
nand U1820 (N_1820,In_499,In_1173);
nand U1821 (N_1821,In_1430,In_173);
and U1822 (N_1822,In_1197,In_941);
nand U1823 (N_1823,In_1179,In_498);
and U1824 (N_1824,In_1075,In_1154);
and U1825 (N_1825,In_434,In_921);
or U1826 (N_1826,In_261,In_1215);
nor U1827 (N_1827,In_770,In_430);
nand U1828 (N_1828,In_1023,In_926);
and U1829 (N_1829,In_521,In_638);
or U1830 (N_1830,In_575,In_408);
and U1831 (N_1831,In_302,In_132);
nand U1832 (N_1832,In_228,In_584);
and U1833 (N_1833,In_644,In_1122);
or U1834 (N_1834,In_366,In_567);
and U1835 (N_1835,In_946,In_1418);
or U1836 (N_1836,In_1124,In_1397);
nor U1837 (N_1837,In_1270,In_256);
nand U1838 (N_1838,In_181,In_753);
or U1839 (N_1839,In_434,In_890);
nor U1840 (N_1840,In_541,In_7);
and U1841 (N_1841,In_218,In_521);
nor U1842 (N_1842,In_1177,In_447);
nor U1843 (N_1843,In_409,In_211);
or U1844 (N_1844,In_590,In_850);
nor U1845 (N_1845,In_983,In_894);
nand U1846 (N_1846,In_1386,In_945);
nor U1847 (N_1847,In_329,In_535);
xor U1848 (N_1848,In_278,In_75);
nand U1849 (N_1849,In_445,In_425);
and U1850 (N_1850,In_366,In_1069);
or U1851 (N_1851,In_773,In_1178);
nand U1852 (N_1852,In_617,In_1447);
or U1853 (N_1853,In_1490,In_1208);
and U1854 (N_1854,In_1350,In_1313);
nand U1855 (N_1855,In_269,In_65);
nor U1856 (N_1856,In_460,In_315);
nor U1857 (N_1857,In_1229,In_1165);
or U1858 (N_1858,In_14,In_884);
nand U1859 (N_1859,In_1368,In_185);
and U1860 (N_1860,In_975,In_121);
or U1861 (N_1861,In_1130,In_124);
and U1862 (N_1862,In_956,In_40);
and U1863 (N_1863,In_1354,In_1035);
xnor U1864 (N_1864,In_386,In_575);
and U1865 (N_1865,In_754,In_1105);
nor U1866 (N_1866,In_278,In_324);
nand U1867 (N_1867,In_429,In_669);
nor U1868 (N_1868,In_332,In_1109);
nand U1869 (N_1869,In_1300,In_1296);
xnor U1870 (N_1870,In_728,In_571);
nand U1871 (N_1871,In_1493,In_1476);
nand U1872 (N_1872,In_742,In_879);
nand U1873 (N_1873,In_167,In_1453);
nor U1874 (N_1874,In_194,In_471);
and U1875 (N_1875,In_821,In_414);
nor U1876 (N_1876,In_1437,In_606);
or U1877 (N_1877,In_750,In_1427);
or U1878 (N_1878,In_75,In_560);
or U1879 (N_1879,In_139,In_230);
xor U1880 (N_1880,In_1146,In_125);
nor U1881 (N_1881,In_1062,In_1381);
nor U1882 (N_1882,In_994,In_122);
and U1883 (N_1883,In_186,In_522);
or U1884 (N_1884,In_1219,In_163);
nand U1885 (N_1885,In_333,In_473);
nand U1886 (N_1886,In_506,In_785);
nor U1887 (N_1887,In_879,In_1397);
nor U1888 (N_1888,In_96,In_1034);
nand U1889 (N_1889,In_1220,In_543);
and U1890 (N_1890,In_1474,In_1296);
nor U1891 (N_1891,In_834,In_741);
and U1892 (N_1892,In_824,In_53);
or U1893 (N_1893,In_474,In_822);
nor U1894 (N_1894,In_1010,In_732);
nor U1895 (N_1895,In_1406,In_796);
xor U1896 (N_1896,In_360,In_1264);
xor U1897 (N_1897,In_1260,In_37);
and U1898 (N_1898,In_345,In_121);
and U1899 (N_1899,In_833,In_1293);
xnor U1900 (N_1900,In_767,In_413);
nor U1901 (N_1901,In_1371,In_1076);
nand U1902 (N_1902,In_1230,In_1212);
or U1903 (N_1903,In_686,In_331);
and U1904 (N_1904,In_1463,In_138);
and U1905 (N_1905,In_585,In_636);
nand U1906 (N_1906,In_766,In_194);
or U1907 (N_1907,In_1237,In_817);
or U1908 (N_1908,In_821,In_36);
nor U1909 (N_1909,In_1393,In_703);
nand U1910 (N_1910,In_738,In_1272);
and U1911 (N_1911,In_663,In_518);
nand U1912 (N_1912,In_266,In_953);
and U1913 (N_1913,In_1292,In_1231);
or U1914 (N_1914,In_228,In_70);
nand U1915 (N_1915,In_1103,In_776);
nand U1916 (N_1916,In_1206,In_280);
nand U1917 (N_1917,In_1002,In_309);
and U1918 (N_1918,In_721,In_912);
or U1919 (N_1919,In_1467,In_636);
nand U1920 (N_1920,In_408,In_9);
or U1921 (N_1921,In_353,In_329);
or U1922 (N_1922,In_985,In_1499);
nor U1923 (N_1923,In_915,In_526);
and U1924 (N_1924,In_434,In_1400);
nor U1925 (N_1925,In_671,In_1268);
nand U1926 (N_1926,In_286,In_675);
and U1927 (N_1927,In_479,In_653);
or U1928 (N_1928,In_1321,In_917);
nor U1929 (N_1929,In_1045,In_348);
and U1930 (N_1930,In_544,In_1128);
or U1931 (N_1931,In_42,In_267);
nor U1932 (N_1932,In_1214,In_1473);
or U1933 (N_1933,In_249,In_86);
and U1934 (N_1934,In_1495,In_258);
nor U1935 (N_1935,In_370,In_919);
xnor U1936 (N_1936,In_1188,In_212);
nand U1937 (N_1937,In_257,In_1396);
xnor U1938 (N_1938,In_101,In_1037);
nor U1939 (N_1939,In_1273,In_1130);
and U1940 (N_1940,In_92,In_1229);
xnor U1941 (N_1941,In_1123,In_1234);
and U1942 (N_1942,In_1309,In_113);
nor U1943 (N_1943,In_529,In_284);
nor U1944 (N_1944,In_616,In_916);
xor U1945 (N_1945,In_875,In_974);
xnor U1946 (N_1946,In_22,In_1054);
nor U1947 (N_1947,In_1346,In_1358);
and U1948 (N_1948,In_1052,In_229);
nand U1949 (N_1949,In_1234,In_332);
nor U1950 (N_1950,In_775,In_806);
and U1951 (N_1951,In_1228,In_1207);
and U1952 (N_1952,In_839,In_56);
nand U1953 (N_1953,In_1300,In_1169);
nor U1954 (N_1954,In_181,In_1393);
xor U1955 (N_1955,In_939,In_375);
nand U1956 (N_1956,In_66,In_574);
nor U1957 (N_1957,In_86,In_1002);
nand U1958 (N_1958,In_142,In_1002);
nand U1959 (N_1959,In_126,In_957);
nand U1960 (N_1960,In_1032,In_277);
nand U1961 (N_1961,In_917,In_1332);
nor U1962 (N_1962,In_708,In_1417);
and U1963 (N_1963,In_1218,In_1495);
or U1964 (N_1964,In_1215,In_149);
nor U1965 (N_1965,In_444,In_610);
or U1966 (N_1966,In_1228,In_451);
or U1967 (N_1967,In_267,In_470);
and U1968 (N_1968,In_985,In_1151);
xor U1969 (N_1969,In_855,In_699);
nand U1970 (N_1970,In_200,In_1263);
or U1971 (N_1971,In_1418,In_249);
or U1972 (N_1972,In_1158,In_284);
nand U1973 (N_1973,In_1313,In_538);
and U1974 (N_1974,In_1237,In_1174);
nand U1975 (N_1975,In_337,In_1456);
nor U1976 (N_1976,In_436,In_1042);
or U1977 (N_1977,In_746,In_564);
xor U1978 (N_1978,In_1129,In_314);
and U1979 (N_1979,In_445,In_1206);
nor U1980 (N_1980,In_380,In_167);
nand U1981 (N_1981,In_199,In_66);
nor U1982 (N_1982,In_605,In_383);
nor U1983 (N_1983,In_956,In_341);
and U1984 (N_1984,In_1437,In_153);
and U1985 (N_1985,In_1259,In_1246);
nor U1986 (N_1986,In_253,In_1372);
nor U1987 (N_1987,In_82,In_162);
and U1988 (N_1988,In_839,In_1465);
or U1989 (N_1989,In_105,In_479);
xnor U1990 (N_1990,In_1445,In_1034);
nand U1991 (N_1991,In_471,In_619);
or U1992 (N_1992,In_649,In_1096);
nand U1993 (N_1993,In_388,In_619);
nor U1994 (N_1994,In_72,In_606);
nand U1995 (N_1995,In_111,In_1435);
or U1996 (N_1996,In_804,In_578);
or U1997 (N_1997,In_1374,In_1219);
or U1998 (N_1998,In_342,In_1218);
and U1999 (N_1999,In_400,In_546);
nand U2000 (N_2000,In_55,In_0);
nand U2001 (N_2001,In_777,In_1192);
xnor U2002 (N_2002,In_519,In_1418);
nand U2003 (N_2003,In_852,In_517);
or U2004 (N_2004,In_722,In_1354);
xor U2005 (N_2005,In_1046,In_224);
and U2006 (N_2006,In_1495,In_1099);
or U2007 (N_2007,In_235,In_463);
nand U2008 (N_2008,In_1312,In_1466);
or U2009 (N_2009,In_882,In_1158);
or U2010 (N_2010,In_1487,In_999);
and U2011 (N_2011,In_1047,In_740);
nand U2012 (N_2012,In_1206,In_792);
nor U2013 (N_2013,In_522,In_1029);
nand U2014 (N_2014,In_219,In_1040);
and U2015 (N_2015,In_1255,In_292);
xor U2016 (N_2016,In_1196,In_713);
or U2017 (N_2017,In_248,In_286);
nand U2018 (N_2018,In_575,In_1315);
and U2019 (N_2019,In_710,In_1273);
and U2020 (N_2020,In_706,In_1148);
and U2021 (N_2021,In_975,In_291);
xor U2022 (N_2022,In_707,In_887);
xnor U2023 (N_2023,In_892,In_1045);
nor U2024 (N_2024,In_684,In_1404);
nor U2025 (N_2025,In_942,In_64);
nor U2026 (N_2026,In_209,In_165);
xnor U2027 (N_2027,In_1298,In_958);
or U2028 (N_2028,In_750,In_687);
nor U2029 (N_2029,In_1344,In_765);
nor U2030 (N_2030,In_1477,In_144);
or U2031 (N_2031,In_1001,In_773);
nand U2032 (N_2032,In_1214,In_315);
nand U2033 (N_2033,In_210,In_225);
or U2034 (N_2034,In_1002,In_705);
or U2035 (N_2035,In_626,In_1375);
nor U2036 (N_2036,In_802,In_695);
and U2037 (N_2037,In_520,In_1056);
or U2038 (N_2038,In_1047,In_660);
xor U2039 (N_2039,In_848,In_54);
nor U2040 (N_2040,In_1025,In_1260);
nand U2041 (N_2041,In_1188,In_808);
or U2042 (N_2042,In_519,In_1170);
or U2043 (N_2043,In_274,In_850);
xnor U2044 (N_2044,In_970,In_875);
nor U2045 (N_2045,In_631,In_1041);
and U2046 (N_2046,In_369,In_1443);
or U2047 (N_2047,In_1264,In_1206);
nand U2048 (N_2048,In_1012,In_383);
xnor U2049 (N_2049,In_1482,In_637);
or U2050 (N_2050,In_474,In_981);
xor U2051 (N_2051,In_929,In_535);
or U2052 (N_2052,In_1159,In_1008);
and U2053 (N_2053,In_1395,In_643);
or U2054 (N_2054,In_1280,In_1136);
or U2055 (N_2055,In_1075,In_215);
or U2056 (N_2056,In_337,In_692);
xnor U2057 (N_2057,In_935,In_218);
nand U2058 (N_2058,In_411,In_196);
or U2059 (N_2059,In_1360,In_198);
or U2060 (N_2060,In_1110,In_346);
or U2061 (N_2061,In_1054,In_168);
or U2062 (N_2062,In_1363,In_1109);
nor U2063 (N_2063,In_856,In_293);
nor U2064 (N_2064,In_1051,In_370);
xnor U2065 (N_2065,In_363,In_65);
nor U2066 (N_2066,In_469,In_1153);
or U2067 (N_2067,In_134,In_626);
or U2068 (N_2068,In_1172,In_15);
xor U2069 (N_2069,In_1334,In_1315);
nand U2070 (N_2070,In_147,In_924);
nand U2071 (N_2071,In_1245,In_271);
or U2072 (N_2072,In_994,In_838);
or U2073 (N_2073,In_766,In_1444);
or U2074 (N_2074,In_1047,In_343);
and U2075 (N_2075,In_165,In_1090);
and U2076 (N_2076,In_223,In_1232);
xnor U2077 (N_2077,In_146,In_428);
and U2078 (N_2078,In_774,In_518);
nor U2079 (N_2079,In_203,In_94);
and U2080 (N_2080,In_154,In_130);
nor U2081 (N_2081,In_594,In_901);
nand U2082 (N_2082,In_885,In_545);
nand U2083 (N_2083,In_915,In_897);
and U2084 (N_2084,In_878,In_1042);
or U2085 (N_2085,In_1226,In_725);
or U2086 (N_2086,In_645,In_872);
and U2087 (N_2087,In_1406,In_168);
nand U2088 (N_2088,In_904,In_1400);
nor U2089 (N_2089,In_572,In_705);
and U2090 (N_2090,In_767,In_402);
nor U2091 (N_2091,In_985,In_340);
and U2092 (N_2092,In_809,In_676);
and U2093 (N_2093,In_384,In_1234);
and U2094 (N_2094,In_1457,In_1253);
nand U2095 (N_2095,In_612,In_949);
and U2096 (N_2096,In_993,In_598);
nor U2097 (N_2097,In_480,In_1120);
nand U2098 (N_2098,In_155,In_1150);
or U2099 (N_2099,In_299,In_810);
xor U2100 (N_2100,In_898,In_434);
and U2101 (N_2101,In_184,In_227);
and U2102 (N_2102,In_249,In_1479);
and U2103 (N_2103,In_100,In_29);
or U2104 (N_2104,In_178,In_149);
or U2105 (N_2105,In_425,In_821);
nand U2106 (N_2106,In_251,In_1452);
or U2107 (N_2107,In_1019,In_92);
or U2108 (N_2108,In_1228,In_549);
xor U2109 (N_2109,In_1208,In_1169);
nand U2110 (N_2110,In_388,In_342);
and U2111 (N_2111,In_811,In_858);
xnor U2112 (N_2112,In_926,In_1077);
nand U2113 (N_2113,In_963,In_163);
nor U2114 (N_2114,In_1395,In_1160);
xor U2115 (N_2115,In_12,In_1106);
nand U2116 (N_2116,In_601,In_304);
nor U2117 (N_2117,In_258,In_721);
and U2118 (N_2118,In_288,In_608);
nand U2119 (N_2119,In_353,In_1414);
nand U2120 (N_2120,In_1373,In_1232);
nor U2121 (N_2121,In_718,In_1312);
xnor U2122 (N_2122,In_1332,In_75);
nor U2123 (N_2123,In_1219,In_918);
and U2124 (N_2124,In_1118,In_229);
nand U2125 (N_2125,In_807,In_599);
nand U2126 (N_2126,In_876,In_481);
or U2127 (N_2127,In_380,In_1309);
nor U2128 (N_2128,In_596,In_1242);
or U2129 (N_2129,In_334,In_62);
nand U2130 (N_2130,In_965,In_1407);
nor U2131 (N_2131,In_749,In_1007);
and U2132 (N_2132,In_60,In_873);
and U2133 (N_2133,In_1366,In_754);
and U2134 (N_2134,In_963,In_1201);
nor U2135 (N_2135,In_696,In_506);
xnor U2136 (N_2136,In_819,In_950);
or U2137 (N_2137,In_856,In_381);
nand U2138 (N_2138,In_409,In_1308);
xnor U2139 (N_2139,In_443,In_841);
or U2140 (N_2140,In_241,In_1169);
nor U2141 (N_2141,In_100,In_208);
and U2142 (N_2142,In_606,In_1408);
or U2143 (N_2143,In_4,In_1207);
or U2144 (N_2144,In_864,In_1103);
nand U2145 (N_2145,In_34,In_1299);
or U2146 (N_2146,In_824,In_440);
and U2147 (N_2147,In_1143,In_391);
nor U2148 (N_2148,In_1179,In_1021);
and U2149 (N_2149,In_158,In_835);
nor U2150 (N_2150,In_1136,In_1462);
or U2151 (N_2151,In_206,In_725);
nand U2152 (N_2152,In_113,In_44);
and U2153 (N_2153,In_808,In_373);
and U2154 (N_2154,In_1310,In_406);
or U2155 (N_2155,In_407,In_1031);
nand U2156 (N_2156,In_886,In_774);
nand U2157 (N_2157,In_1414,In_1270);
or U2158 (N_2158,In_994,In_1263);
nor U2159 (N_2159,In_579,In_207);
xnor U2160 (N_2160,In_674,In_601);
or U2161 (N_2161,In_1136,In_67);
or U2162 (N_2162,In_1360,In_1210);
xor U2163 (N_2163,In_272,In_1159);
and U2164 (N_2164,In_1169,In_388);
and U2165 (N_2165,In_1191,In_1258);
or U2166 (N_2166,In_321,In_326);
and U2167 (N_2167,In_796,In_451);
nor U2168 (N_2168,In_1161,In_202);
nor U2169 (N_2169,In_1043,In_449);
or U2170 (N_2170,In_178,In_1068);
and U2171 (N_2171,In_872,In_30);
or U2172 (N_2172,In_1182,In_902);
nor U2173 (N_2173,In_1499,In_7);
and U2174 (N_2174,In_384,In_1270);
xor U2175 (N_2175,In_160,In_1445);
nand U2176 (N_2176,In_1086,In_26);
nor U2177 (N_2177,In_1070,In_766);
or U2178 (N_2178,In_150,In_143);
and U2179 (N_2179,In_817,In_502);
and U2180 (N_2180,In_1029,In_1406);
and U2181 (N_2181,In_1337,In_594);
nand U2182 (N_2182,In_785,In_990);
nand U2183 (N_2183,In_1431,In_36);
or U2184 (N_2184,In_940,In_874);
or U2185 (N_2185,In_1271,In_888);
and U2186 (N_2186,In_93,In_7);
xnor U2187 (N_2187,In_980,In_280);
and U2188 (N_2188,In_1184,In_736);
or U2189 (N_2189,In_84,In_379);
nand U2190 (N_2190,In_1292,In_589);
and U2191 (N_2191,In_339,In_1120);
nand U2192 (N_2192,In_935,In_714);
or U2193 (N_2193,In_895,In_628);
or U2194 (N_2194,In_131,In_507);
and U2195 (N_2195,In_550,In_1485);
and U2196 (N_2196,In_25,In_417);
nand U2197 (N_2197,In_867,In_155);
nor U2198 (N_2198,In_1432,In_923);
and U2199 (N_2199,In_1107,In_1179);
or U2200 (N_2200,In_1195,In_1270);
nand U2201 (N_2201,In_418,In_437);
or U2202 (N_2202,In_916,In_892);
and U2203 (N_2203,In_712,In_680);
nand U2204 (N_2204,In_873,In_837);
nor U2205 (N_2205,In_1430,In_1213);
nor U2206 (N_2206,In_1092,In_43);
and U2207 (N_2207,In_1368,In_1303);
nand U2208 (N_2208,In_217,In_0);
and U2209 (N_2209,In_516,In_1497);
nand U2210 (N_2210,In_1189,In_899);
nand U2211 (N_2211,In_30,In_1123);
nor U2212 (N_2212,In_210,In_299);
nor U2213 (N_2213,In_1020,In_646);
nor U2214 (N_2214,In_278,In_1069);
or U2215 (N_2215,In_1379,In_979);
nand U2216 (N_2216,In_1003,In_1368);
nor U2217 (N_2217,In_1183,In_999);
or U2218 (N_2218,In_518,In_12);
nor U2219 (N_2219,In_412,In_12);
xor U2220 (N_2220,In_1204,In_1029);
nor U2221 (N_2221,In_881,In_591);
nand U2222 (N_2222,In_1297,In_367);
or U2223 (N_2223,In_1015,In_437);
and U2224 (N_2224,In_1260,In_731);
or U2225 (N_2225,In_153,In_44);
xnor U2226 (N_2226,In_719,In_891);
nor U2227 (N_2227,In_834,In_538);
or U2228 (N_2228,In_345,In_1096);
nor U2229 (N_2229,In_1279,In_236);
nand U2230 (N_2230,In_1469,In_524);
nand U2231 (N_2231,In_229,In_258);
nor U2232 (N_2232,In_1207,In_970);
nor U2233 (N_2233,In_826,In_382);
nor U2234 (N_2234,In_1288,In_61);
xnor U2235 (N_2235,In_1232,In_1417);
nor U2236 (N_2236,In_341,In_1384);
or U2237 (N_2237,In_234,In_427);
nor U2238 (N_2238,In_364,In_1413);
nor U2239 (N_2239,In_1438,In_1460);
or U2240 (N_2240,In_739,In_882);
and U2241 (N_2241,In_196,In_88);
or U2242 (N_2242,In_26,In_1127);
xnor U2243 (N_2243,In_804,In_341);
nand U2244 (N_2244,In_1286,In_1408);
nand U2245 (N_2245,In_652,In_129);
nand U2246 (N_2246,In_1468,In_349);
nor U2247 (N_2247,In_1220,In_1135);
or U2248 (N_2248,In_354,In_868);
and U2249 (N_2249,In_156,In_445);
xor U2250 (N_2250,In_321,In_674);
and U2251 (N_2251,In_1099,In_1386);
xnor U2252 (N_2252,In_1334,In_270);
or U2253 (N_2253,In_715,In_176);
xnor U2254 (N_2254,In_1082,In_346);
nor U2255 (N_2255,In_1495,In_1009);
xnor U2256 (N_2256,In_1032,In_1086);
nor U2257 (N_2257,In_1351,In_1107);
or U2258 (N_2258,In_426,In_1144);
nor U2259 (N_2259,In_169,In_325);
nand U2260 (N_2260,In_1370,In_623);
nand U2261 (N_2261,In_806,In_516);
or U2262 (N_2262,In_861,In_718);
nor U2263 (N_2263,In_744,In_643);
and U2264 (N_2264,In_1411,In_1126);
or U2265 (N_2265,In_1450,In_561);
and U2266 (N_2266,In_917,In_1374);
nand U2267 (N_2267,In_1312,In_1327);
nand U2268 (N_2268,In_496,In_438);
nand U2269 (N_2269,In_1244,In_1127);
and U2270 (N_2270,In_1472,In_319);
nand U2271 (N_2271,In_1221,In_89);
nor U2272 (N_2272,In_40,In_529);
xnor U2273 (N_2273,In_535,In_784);
or U2274 (N_2274,In_75,In_280);
nor U2275 (N_2275,In_613,In_1075);
xor U2276 (N_2276,In_1013,In_979);
or U2277 (N_2277,In_1447,In_540);
nor U2278 (N_2278,In_568,In_199);
nand U2279 (N_2279,In_1245,In_437);
xnor U2280 (N_2280,In_517,In_940);
nand U2281 (N_2281,In_794,In_573);
nand U2282 (N_2282,In_116,In_719);
and U2283 (N_2283,In_994,In_454);
nor U2284 (N_2284,In_1266,In_95);
xor U2285 (N_2285,In_879,In_1259);
nand U2286 (N_2286,In_296,In_44);
and U2287 (N_2287,In_993,In_891);
nor U2288 (N_2288,In_515,In_889);
or U2289 (N_2289,In_1329,In_121);
or U2290 (N_2290,In_77,In_1406);
or U2291 (N_2291,In_22,In_1349);
or U2292 (N_2292,In_1485,In_265);
and U2293 (N_2293,In_7,In_688);
or U2294 (N_2294,In_984,In_537);
and U2295 (N_2295,In_481,In_356);
nor U2296 (N_2296,In_26,In_286);
and U2297 (N_2297,In_769,In_841);
and U2298 (N_2298,In_404,In_417);
nor U2299 (N_2299,In_1408,In_35);
nand U2300 (N_2300,In_1070,In_1463);
nand U2301 (N_2301,In_946,In_1073);
nor U2302 (N_2302,In_440,In_97);
nor U2303 (N_2303,In_5,In_1467);
or U2304 (N_2304,In_542,In_92);
nor U2305 (N_2305,In_486,In_211);
nor U2306 (N_2306,In_188,In_299);
nor U2307 (N_2307,In_532,In_1243);
or U2308 (N_2308,In_182,In_270);
and U2309 (N_2309,In_437,In_696);
and U2310 (N_2310,In_1178,In_347);
nor U2311 (N_2311,In_1463,In_1029);
and U2312 (N_2312,In_208,In_459);
nand U2313 (N_2313,In_813,In_325);
or U2314 (N_2314,In_1262,In_199);
or U2315 (N_2315,In_1204,In_1107);
nor U2316 (N_2316,In_1281,In_1044);
nor U2317 (N_2317,In_468,In_1302);
or U2318 (N_2318,In_454,In_999);
xor U2319 (N_2319,In_295,In_632);
and U2320 (N_2320,In_692,In_165);
and U2321 (N_2321,In_923,In_56);
xnor U2322 (N_2322,In_872,In_996);
xnor U2323 (N_2323,In_1291,In_1164);
or U2324 (N_2324,In_316,In_905);
or U2325 (N_2325,In_560,In_200);
xnor U2326 (N_2326,In_394,In_978);
and U2327 (N_2327,In_1079,In_1227);
xnor U2328 (N_2328,In_145,In_760);
and U2329 (N_2329,In_1010,In_592);
nor U2330 (N_2330,In_1408,In_1431);
nor U2331 (N_2331,In_611,In_1241);
nand U2332 (N_2332,In_806,In_360);
and U2333 (N_2333,In_1089,In_506);
nor U2334 (N_2334,In_1016,In_648);
and U2335 (N_2335,In_965,In_1232);
nand U2336 (N_2336,In_1353,In_1242);
and U2337 (N_2337,In_336,In_155);
nor U2338 (N_2338,In_1266,In_491);
xnor U2339 (N_2339,In_1248,In_284);
nor U2340 (N_2340,In_408,In_537);
and U2341 (N_2341,In_381,In_714);
and U2342 (N_2342,In_832,In_470);
nor U2343 (N_2343,In_327,In_264);
nand U2344 (N_2344,In_162,In_146);
or U2345 (N_2345,In_727,In_273);
or U2346 (N_2346,In_343,In_959);
nor U2347 (N_2347,In_678,In_202);
and U2348 (N_2348,In_1468,In_637);
xor U2349 (N_2349,In_112,In_465);
and U2350 (N_2350,In_260,In_1475);
nand U2351 (N_2351,In_8,In_1262);
and U2352 (N_2352,In_486,In_1089);
and U2353 (N_2353,In_630,In_524);
or U2354 (N_2354,In_370,In_608);
or U2355 (N_2355,In_715,In_495);
and U2356 (N_2356,In_1308,In_255);
or U2357 (N_2357,In_721,In_990);
nand U2358 (N_2358,In_1071,In_1082);
or U2359 (N_2359,In_557,In_370);
or U2360 (N_2360,In_717,In_1220);
nor U2361 (N_2361,In_417,In_97);
or U2362 (N_2362,In_857,In_1289);
nand U2363 (N_2363,In_87,In_1055);
xor U2364 (N_2364,In_815,In_932);
nand U2365 (N_2365,In_1078,In_876);
and U2366 (N_2366,In_1314,In_475);
or U2367 (N_2367,In_704,In_733);
or U2368 (N_2368,In_483,In_521);
or U2369 (N_2369,In_565,In_66);
nand U2370 (N_2370,In_1051,In_895);
and U2371 (N_2371,In_1457,In_499);
nand U2372 (N_2372,In_293,In_1490);
nor U2373 (N_2373,In_815,In_537);
or U2374 (N_2374,In_1061,In_663);
and U2375 (N_2375,In_942,In_258);
nor U2376 (N_2376,In_209,In_252);
or U2377 (N_2377,In_1048,In_1108);
xor U2378 (N_2378,In_697,In_1316);
nand U2379 (N_2379,In_195,In_1097);
nor U2380 (N_2380,In_754,In_1206);
or U2381 (N_2381,In_85,In_345);
nand U2382 (N_2382,In_431,In_1329);
and U2383 (N_2383,In_379,In_1352);
nand U2384 (N_2384,In_901,In_395);
and U2385 (N_2385,In_1225,In_1222);
xor U2386 (N_2386,In_40,In_921);
nand U2387 (N_2387,In_1060,In_1478);
or U2388 (N_2388,In_1372,In_88);
nor U2389 (N_2389,In_513,In_1089);
nand U2390 (N_2390,In_1337,In_37);
nand U2391 (N_2391,In_892,In_1024);
nand U2392 (N_2392,In_1272,In_114);
and U2393 (N_2393,In_821,In_1249);
nor U2394 (N_2394,In_1078,In_303);
xnor U2395 (N_2395,In_909,In_674);
nor U2396 (N_2396,In_1165,In_949);
nand U2397 (N_2397,In_702,In_251);
xnor U2398 (N_2398,In_1104,In_756);
nand U2399 (N_2399,In_453,In_945);
nor U2400 (N_2400,In_915,In_1201);
nand U2401 (N_2401,In_824,In_467);
xnor U2402 (N_2402,In_554,In_1248);
nor U2403 (N_2403,In_1411,In_222);
xnor U2404 (N_2404,In_1022,In_963);
nor U2405 (N_2405,In_87,In_784);
or U2406 (N_2406,In_1301,In_610);
or U2407 (N_2407,In_1170,In_472);
nand U2408 (N_2408,In_1416,In_120);
nor U2409 (N_2409,In_128,In_600);
nor U2410 (N_2410,In_159,In_731);
nand U2411 (N_2411,In_757,In_738);
nand U2412 (N_2412,In_43,In_541);
or U2413 (N_2413,In_1186,In_1);
and U2414 (N_2414,In_1357,In_1322);
and U2415 (N_2415,In_1128,In_1044);
nand U2416 (N_2416,In_1162,In_1298);
and U2417 (N_2417,In_101,In_592);
or U2418 (N_2418,In_753,In_269);
nor U2419 (N_2419,In_832,In_775);
xnor U2420 (N_2420,In_492,In_804);
or U2421 (N_2421,In_93,In_226);
nand U2422 (N_2422,In_405,In_230);
nand U2423 (N_2423,In_149,In_604);
and U2424 (N_2424,In_1098,In_663);
nand U2425 (N_2425,In_466,In_1102);
nor U2426 (N_2426,In_1381,In_1080);
nor U2427 (N_2427,In_27,In_727);
nor U2428 (N_2428,In_1272,In_901);
or U2429 (N_2429,In_1057,In_1401);
nand U2430 (N_2430,In_460,In_1234);
xor U2431 (N_2431,In_811,In_269);
nor U2432 (N_2432,In_1213,In_1186);
nand U2433 (N_2433,In_938,In_521);
nor U2434 (N_2434,In_729,In_1049);
or U2435 (N_2435,In_1148,In_1420);
xor U2436 (N_2436,In_579,In_1297);
xor U2437 (N_2437,In_1155,In_309);
or U2438 (N_2438,In_303,In_827);
or U2439 (N_2439,In_614,In_587);
nor U2440 (N_2440,In_497,In_281);
nand U2441 (N_2441,In_1328,In_970);
xnor U2442 (N_2442,In_905,In_327);
nor U2443 (N_2443,In_977,In_1122);
nand U2444 (N_2444,In_430,In_900);
or U2445 (N_2445,In_840,In_1477);
and U2446 (N_2446,In_715,In_747);
and U2447 (N_2447,In_1421,In_216);
and U2448 (N_2448,In_787,In_857);
and U2449 (N_2449,In_436,In_920);
nand U2450 (N_2450,In_419,In_1063);
or U2451 (N_2451,In_836,In_1060);
nor U2452 (N_2452,In_464,In_894);
nor U2453 (N_2453,In_902,In_1076);
or U2454 (N_2454,In_364,In_406);
or U2455 (N_2455,In_314,In_1481);
nor U2456 (N_2456,In_513,In_1432);
nand U2457 (N_2457,In_696,In_229);
and U2458 (N_2458,In_1194,In_709);
nor U2459 (N_2459,In_1267,In_806);
nand U2460 (N_2460,In_307,In_1259);
or U2461 (N_2461,In_1395,In_916);
xnor U2462 (N_2462,In_783,In_1387);
nand U2463 (N_2463,In_1032,In_1416);
nor U2464 (N_2464,In_499,In_1369);
xor U2465 (N_2465,In_726,In_236);
xnor U2466 (N_2466,In_838,In_738);
nor U2467 (N_2467,In_990,In_1231);
and U2468 (N_2468,In_1207,In_492);
nand U2469 (N_2469,In_153,In_1165);
and U2470 (N_2470,In_683,In_739);
nor U2471 (N_2471,In_383,In_1279);
and U2472 (N_2472,In_234,In_1088);
or U2473 (N_2473,In_171,In_40);
or U2474 (N_2474,In_121,In_880);
xnor U2475 (N_2475,In_534,In_422);
nand U2476 (N_2476,In_512,In_1100);
or U2477 (N_2477,In_878,In_1400);
and U2478 (N_2478,In_1494,In_856);
nand U2479 (N_2479,In_215,In_1114);
nand U2480 (N_2480,In_1007,In_417);
nand U2481 (N_2481,In_265,In_96);
nand U2482 (N_2482,In_697,In_1033);
nor U2483 (N_2483,In_202,In_767);
or U2484 (N_2484,In_36,In_201);
or U2485 (N_2485,In_1205,In_376);
or U2486 (N_2486,In_272,In_1453);
or U2487 (N_2487,In_279,In_1205);
and U2488 (N_2488,In_973,In_1233);
nor U2489 (N_2489,In_96,In_1080);
nand U2490 (N_2490,In_264,In_529);
nand U2491 (N_2491,In_912,In_185);
and U2492 (N_2492,In_937,In_216);
and U2493 (N_2493,In_1028,In_529);
nor U2494 (N_2494,In_69,In_1443);
nand U2495 (N_2495,In_591,In_1463);
or U2496 (N_2496,In_776,In_1001);
or U2497 (N_2497,In_214,In_335);
xor U2498 (N_2498,In_1458,In_604);
and U2499 (N_2499,In_1094,In_365);
xnor U2500 (N_2500,In_1404,In_2);
or U2501 (N_2501,In_813,In_17);
nor U2502 (N_2502,In_1435,In_1402);
nand U2503 (N_2503,In_583,In_560);
or U2504 (N_2504,In_370,In_316);
nor U2505 (N_2505,In_926,In_185);
and U2506 (N_2506,In_1187,In_267);
nand U2507 (N_2507,In_1005,In_949);
and U2508 (N_2508,In_438,In_366);
nand U2509 (N_2509,In_477,In_1300);
nand U2510 (N_2510,In_116,In_836);
xor U2511 (N_2511,In_757,In_748);
or U2512 (N_2512,In_508,In_914);
nor U2513 (N_2513,In_1015,In_920);
nand U2514 (N_2514,In_1272,In_1201);
or U2515 (N_2515,In_608,In_1247);
or U2516 (N_2516,In_1322,In_925);
xor U2517 (N_2517,In_863,In_888);
nand U2518 (N_2518,In_422,In_363);
or U2519 (N_2519,In_523,In_127);
xor U2520 (N_2520,In_492,In_863);
nand U2521 (N_2521,In_401,In_759);
nor U2522 (N_2522,In_1040,In_1128);
nand U2523 (N_2523,In_949,In_183);
nor U2524 (N_2524,In_1045,In_131);
or U2525 (N_2525,In_1480,In_756);
nor U2526 (N_2526,In_1171,In_1191);
xor U2527 (N_2527,In_929,In_58);
xor U2528 (N_2528,In_615,In_1049);
and U2529 (N_2529,In_850,In_640);
and U2530 (N_2530,In_257,In_376);
nand U2531 (N_2531,In_579,In_294);
nor U2532 (N_2532,In_1385,In_840);
xor U2533 (N_2533,In_380,In_1273);
nand U2534 (N_2534,In_348,In_1253);
nor U2535 (N_2535,In_921,In_778);
nand U2536 (N_2536,In_1259,In_545);
nand U2537 (N_2537,In_826,In_999);
xnor U2538 (N_2538,In_692,In_820);
nor U2539 (N_2539,In_109,In_1452);
nor U2540 (N_2540,In_622,In_723);
or U2541 (N_2541,In_1461,In_1428);
nand U2542 (N_2542,In_195,In_66);
nand U2543 (N_2543,In_774,In_1206);
nand U2544 (N_2544,In_168,In_140);
nor U2545 (N_2545,In_665,In_420);
or U2546 (N_2546,In_295,In_698);
and U2547 (N_2547,In_946,In_1359);
nand U2548 (N_2548,In_1423,In_1478);
or U2549 (N_2549,In_1248,In_1339);
and U2550 (N_2550,In_194,In_1133);
and U2551 (N_2551,In_315,In_422);
nor U2552 (N_2552,In_1365,In_204);
and U2553 (N_2553,In_1087,In_669);
or U2554 (N_2554,In_1384,In_1409);
nand U2555 (N_2555,In_379,In_444);
nand U2556 (N_2556,In_1320,In_2);
or U2557 (N_2557,In_1085,In_160);
or U2558 (N_2558,In_652,In_550);
and U2559 (N_2559,In_261,In_421);
nand U2560 (N_2560,In_584,In_851);
and U2561 (N_2561,In_62,In_1252);
nand U2562 (N_2562,In_1490,In_511);
or U2563 (N_2563,In_942,In_393);
nand U2564 (N_2564,In_292,In_462);
nand U2565 (N_2565,In_1362,In_1065);
or U2566 (N_2566,In_683,In_104);
nor U2567 (N_2567,In_1239,In_1224);
nand U2568 (N_2568,In_1494,In_979);
and U2569 (N_2569,In_712,In_699);
or U2570 (N_2570,In_1262,In_684);
nand U2571 (N_2571,In_163,In_110);
nand U2572 (N_2572,In_709,In_806);
nor U2573 (N_2573,In_1485,In_888);
or U2574 (N_2574,In_1487,In_1329);
nor U2575 (N_2575,In_1213,In_629);
nor U2576 (N_2576,In_33,In_248);
nand U2577 (N_2577,In_344,In_1408);
or U2578 (N_2578,In_1366,In_1333);
and U2579 (N_2579,In_1438,In_335);
and U2580 (N_2580,In_766,In_358);
nand U2581 (N_2581,In_492,In_514);
and U2582 (N_2582,In_936,In_63);
xnor U2583 (N_2583,In_345,In_1175);
nor U2584 (N_2584,In_1204,In_448);
nand U2585 (N_2585,In_195,In_776);
and U2586 (N_2586,In_37,In_1185);
or U2587 (N_2587,In_642,In_432);
or U2588 (N_2588,In_907,In_985);
nor U2589 (N_2589,In_670,In_963);
nand U2590 (N_2590,In_1188,In_6);
and U2591 (N_2591,In_923,In_557);
nor U2592 (N_2592,In_1325,In_859);
and U2593 (N_2593,In_9,In_1443);
or U2594 (N_2594,In_245,In_50);
nor U2595 (N_2595,In_1093,In_844);
and U2596 (N_2596,In_721,In_428);
nor U2597 (N_2597,In_392,In_1068);
nand U2598 (N_2598,In_1398,In_480);
nor U2599 (N_2599,In_1003,In_854);
or U2600 (N_2600,In_573,In_526);
and U2601 (N_2601,In_753,In_1009);
nor U2602 (N_2602,In_1498,In_1223);
or U2603 (N_2603,In_1460,In_7);
xnor U2604 (N_2604,In_715,In_718);
nor U2605 (N_2605,In_937,In_596);
and U2606 (N_2606,In_280,In_1095);
xnor U2607 (N_2607,In_1371,In_249);
nor U2608 (N_2608,In_1345,In_1169);
nor U2609 (N_2609,In_547,In_299);
nand U2610 (N_2610,In_1426,In_303);
and U2611 (N_2611,In_770,In_1249);
nand U2612 (N_2612,In_1412,In_5);
nor U2613 (N_2613,In_720,In_1082);
and U2614 (N_2614,In_980,In_942);
xor U2615 (N_2615,In_331,In_1000);
or U2616 (N_2616,In_961,In_183);
nand U2617 (N_2617,In_255,In_550);
and U2618 (N_2618,In_1051,In_360);
and U2619 (N_2619,In_1008,In_604);
xnor U2620 (N_2620,In_273,In_219);
or U2621 (N_2621,In_276,In_1403);
or U2622 (N_2622,In_103,In_150);
xnor U2623 (N_2623,In_1168,In_213);
xnor U2624 (N_2624,In_493,In_726);
or U2625 (N_2625,In_20,In_1438);
nor U2626 (N_2626,In_1137,In_1261);
xnor U2627 (N_2627,In_1096,In_1023);
and U2628 (N_2628,In_380,In_973);
nor U2629 (N_2629,In_1431,In_419);
and U2630 (N_2630,In_1018,In_10);
and U2631 (N_2631,In_858,In_1387);
and U2632 (N_2632,In_1168,In_483);
nand U2633 (N_2633,In_718,In_789);
or U2634 (N_2634,In_1188,In_182);
nor U2635 (N_2635,In_127,In_1230);
nor U2636 (N_2636,In_868,In_339);
nand U2637 (N_2637,In_1125,In_1280);
nand U2638 (N_2638,In_439,In_523);
nand U2639 (N_2639,In_881,In_1436);
and U2640 (N_2640,In_1233,In_512);
nand U2641 (N_2641,In_798,In_1267);
nor U2642 (N_2642,In_261,In_1036);
xnor U2643 (N_2643,In_178,In_349);
nand U2644 (N_2644,In_1158,In_349);
nand U2645 (N_2645,In_20,In_416);
and U2646 (N_2646,In_220,In_1050);
nor U2647 (N_2647,In_1045,In_149);
nand U2648 (N_2648,In_971,In_629);
and U2649 (N_2649,In_1459,In_713);
nor U2650 (N_2650,In_66,In_1494);
xnor U2651 (N_2651,In_293,In_1482);
or U2652 (N_2652,In_1397,In_729);
nand U2653 (N_2653,In_1279,In_1282);
nor U2654 (N_2654,In_1196,In_1496);
nor U2655 (N_2655,In_1044,In_234);
nand U2656 (N_2656,In_1117,In_356);
nor U2657 (N_2657,In_731,In_951);
nor U2658 (N_2658,In_792,In_104);
or U2659 (N_2659,In_1153,In_946);
xnor U2660 (N_2660,In_545,In_1348);
nand U2661 (N_2661,In_13,In_361);
or U2662 (N_2662,In_120,In_1029);
or U2663 (N_2663,In_1108,In_466);
nor U2664 (N_2664,In_1383,In_514);
and U2665 (N_2665,In_479,In_1127);
nand U2666 (N_2666,In_1005,In_622);
nand U2667 (N_2667,In_1099,In_797);
nor U2668 (N_2668,In_1384,In_420);
and U2669 (N_2669,In_235,In_308);
xnor U2670 (N_2670,In_990,In_330);
and U2671 (N_2671,In_901,In_1490);
or U2672 (N_2672,In_466,In_1349);
xor U2673 (N_2673,In_407,In_504);
nor U2674 (N_2674,In_514,In_711);
or U2675 (N_2675,In_1257,In_513);
nand U2676 (N_2676,In_435,In_1063);
nor U2677 (N_2677,In_537,In_1008);
nor U2678 (N_2678,In_1286,In_314);
nor U2679 (N_2679,In_503,In_105);
or U2680 (N_2680,In_197,In_1143);
or U2681 (N_2681,In_526,In_515);
nor U2682 (N_2682,In_1343,In_4);
nor U2683 (N_2683,In_555,In_667);
nor U2684 (N_2684,In_1159,In_468);
and U2685 (N_2685,In_1264,In_900);
or U2686 (N_2686,In_49,In_716);
and U2687 (N_2687,In_859,In_891);
or U2688 (N_2688,In_706,In_430);
nor U2689 (N_2689,In_1174,In_302);
nor U2690 (N_2690,In_1078,In_528);
nand U2691 (N_2691,In_848,In_559);
xor U2692 (N_2692,In_121,In_1339);
nand U2693 (N_2693,In_111,In_330);
nor U2694 (N_2694,In_89,In_818);
xor U2695 (N_2695,In_908,In_1324);
nor U2696 (N_2696,In_1102,In_65);
or U2697 (N_2697,In_752,In_1408);
or U2698 (N_2698,In_456,In_1254);
nand U2699 (N_2699,In_842,In_1336);
nor U2700 (N_2700,In_624,In_248);
and U2701 (N_2701,In_46,In_55);
or U2702 (N_2702,In_1033,In_675);
nor U2703 (N_2703,In_61,In_804);
nor U2704 (N_2704,In_1167,In_350);
and U2705 (N_2705,In_164,In_83);
nand U2706 (N_2706,In_713,In_164);
or U2707 (N_2707,In_435,In_459);
nand U2708 (N_2708,In_1049,In_387);
nand U2709 (N_2709,In_11,In_958);
nand U2710 (N_2710,In_767,In_1391);
and U2711 (N_2711,In_15,In_608);
or U2712 (N_2712,In_1182,In_1114);
and U2713 (N_2713,In_750,In_709);
and U2714 (N_2714,In_1431,In_67);
and U2715 (N_2715,In_666,In_407);
nand U2716 (N_2716,In_931,In_1246);
nand U2717 (N_2717,In_296,In_1482);
nor U2718 (N_2718,In_6,In_314);
nor U2719 (N_2719,In_233,In_1206);
or U2720 (N_2720,In_1379,In_150);
or U2721 (N_2721,In_857,In_264);
and U2722 (N_2722,In_1481,In_1004);
xnor U2723 (N_2723,In_930,In_1343);
nand U2724 (N_2724,In_1096,In_1158);
nand U2725 (N_2725,In_789,In_279);
nor U2726 (N_2726,In_119,In_1393);
xor U2727 (N_2727,In_740,In_808);
or U2728 (N_2728,In_525,In_1371);
or U2729 (N_2729,In_441,In_1483);
or U2730 (N_2730,In_337,In_1363);
nor U2731 (N_2731,In_629,In_499);
or U2732 (N_2732,In_1236,In_838);
nand U2733 (N_2733,In_1111,In_258);
nand U2734 (N_2734,In_23,In_1088);
nand U2735 (N_2735,In_48,In_1317);
or U2736 (N_2736,In_84,In_96);
nand U2737 (N_2737,In_1309,In_1363);
or U2738 (N_2738,In_127,In_110);
nand U2739 (N_2739,In_45,In_1149);
and U2740 (N_2740,In_244,In_305);
or U2741 (N_2741,In_440,In_390);
or U2742 (N_2742,In_952,In_418);
or U2743 (N_2743,In_611,In_1087);
nor U2744 (N_2744,In_47,In_631);
and U2745 (N_2745,In_852,In_324);
and U2746 (N_2746,In_994,In_342);
nor U2747 (N_2747,In_763,In_861);
nor U2748 (N_2748,In_1277,In_163);
xnor U2749 (N_2749,In_385,In_1281);
nand U2750 (N_2750,In_394,In_210);
and U2751 (N_2751,In_1188,In_1434);
nor U2752 (N_2752,In_1321,In_816);
and U2753 (N_2753,In_968,In_571);
and U2754 (N_2754,In_512,In_1179);
nand U2755 (N_2755,In_1245,In_667);
nor U2756 (N_2756,In_946,In_528);
and U2757 (N_2757,In_948,In_193);
or U2758 (N_2758,In_708,In_1301);
or U2759 (N_2759,In_1402,In_1328);
nand U2760 (N_2760,In_1275,In_317);
and U2761 (N_2761,In_963,In_745);
or U2762 (N_2762,In_1399,In_841);
nand U2763 (N_2763,In_413,In_1239);
nor U2764 (N_2764,In_199,In_16);
or U2765 (N_2765,In_1444,In_1334);
nor U2766 (N_2766,In_724,In_27);
or U2767 (N_2767,In_921,In_590);
nor U2768 (N_2768,In_1454,In_856);
and U2769 (N_2769,In_1426,In_749);
or U2770 (N_2770,In_285,In_983);
or U2771 (N_2771,In_1097,In_95);
and U2772 (N_2772,In_589,In_190);
nor U2773 (N_2773,In_193,In_46);
and U2774 (N_2774,In_89,In_1434);
nand U2775 (N_2775,In_1395,In_1226);
nor U2776 (N_2776,In_186,In_907);
nand U2777 (N_2777,In_409,In_1061);
nor U2778 (N_2778,In_281,In_1341);
nor U2779 (N_2779,In_148,In_941);
nor U2780 (N_2780,In_435,In_1396);
nor U2781 (N_2781,In_1316,In_493);
and U2782 (N_2782,In_1449,In_811);
xor U2783 (N_2783,In_580,In_103);
or U2784 (N_2784,In_399,In_1180);
nand U2785 (N_2785,In_649,In_206);
nand U2786 (N_2786,In_405,In_684);
nand U2787 (N_2787,In_8,In_201);
or U2788 (N_2788,In_1177,In_254);
nor U2789 (N_2789,In_53,In_1192);
xor U2790 (N_2790,In_1352,In_253);
xor U2791 (N_2791,In_729,In_148);
nand U2792 (N_2792,In_6,In_548);
nand U2793 (N_2793,In_1156,In_1277);
xnor U2794 (N_2794,In_778,In_356);
nand U2795 (N_2795,In_321,In_908);
or U2796 (N_2796,In_888,In_814);
and U2797 (N_2797,In_550,In_1097);
or U2798 (N_2798,In_868,In_916);
nand U2799 (N_2799,In_564,In_832);
or U2800 (N_2800,In_660,In_661);
or U2801 (N_2801,In_128,In_174);
xor U2802 (N_2802,In_195,In_1391);
and U2803 (N_2803,In_1195,In_717);
or U2804 (N_2804,In_228,In_737);
and U2805 (N_2805,In_20,In_859);
nor U2806 (N_2806,In_131,In_774);
nand U2807 (N_2807,In_717,In_1369);
or U2808 (N_2808,In_537,In_1119);
nand U2809 (N_2809,In_1396,In_1030);
or U2810 (N_2810,In_1254,In_766);
or U2811 (N_2811,In_1237,In_1274);
or U2812 (N_2812,In_660,In_614);
or U2813 (N_2813,In_273,In_791);
nor U2814 (N_2814,In_909,In_734);
nand U2815 (N_2815,In_1235,In_1123);
xor U2816 (N_2816,In_1154,In_1402);
nor U2817 (N_2817,In_173,In_601);
and U2818 (N_2818,In_141,In_752);
nand U2819 (N_2819,In_536,In_235);
and U2820 (N_2820,In_771,In_1020);
nor U2821 (N_2821,In_1476,In_579);
nand U2822 (N_2822,In_223,In_670);
nand U2823 (N_2823,In_1144,In_687);
or U2824 (N_2824,In_149,In_1146);
xor U2825 (N_2825,In_478,In_894);
nand U2826 (N_2826,In_178,In_603);
and U2827 (N_2827,In_1271,In_1026);
or U2828 (N_2828,In_55,In_356);
or U2829 (N_2829,In_351,In_693);
nand U2830 (N_2830,In_436,In_338);
and U2831 (N_2831,In_765,In_120);
and U2832 (N_2832,In_672,In_502);
or U2833 (N_2833,In_1215,In_744);
nand U2834 (N_2834,In_1294,In_643);
or U2835 (N_2835,In_953,In_687);
and U2836 (N_2836,In_818,In_1206);
nand U2837 (N_2837,In_247,In_750);
nor U2838 (N_2838,In_849,In_1294);
nand U2839 (N_2839,In_1422,In_967);
and U2840 (N_2840,In_168,In_1109);
nor U2841 (N_2841,In_242,In_157);
nor U2842 (N_2842,In_42,In_634);
xnor U2843 (N_2843,In_1249,In_155);
or U2844 (N_2844,In_324,In_1080);
nor U2845 (N_2845,In_205,In_88);
and U2846 (N_2846,In_359,In_846);
nor U2847 (N_2847,In_611,In_261);
nor U2848 (N_2848,In_762,In_1124);
and U2849 (N_2849,In_868,In_1260);
xnor U2850 (N_2850,In_1307,In_1114);
xor U2851 (N_2851,In_134,In_218);
nand U2852 (N_2852,In_1406,In_533);
or U2853 (N_2853,In_388,In_1038);
nor U2854 (N_2854,In_871,In_670);
nand U2855 (N_2855,In_1389,In_942);
nor U2856 (N_2856,In_48,In_851);
or U2857 (N_2857,In_951,In_72);
and U2858 (N_2858,In_1249,In_227);
and U2859 (N_2859,In_20,In_1180);
nand U2860 (N_2860,In_957,In_398);
or U2861 (N_2861,In_1097,In_387);
and U2862 (N_2862,In_1099,In_586);
and U2863 (N_2863,In_916,In_182);
and U2864 (N_2864,In_502,In_1229);
nor U2865 (N_2865,In_865,In_55);
nor U2866 (N_2866,In_373,In_1099);
or U2867 (N_2867,In_718,In_298);
nand U2868 (N_2868,In_84,In_210);
nand U2869 (N_2869,In_1405,In_1245);
and U2870 (N_2870,In_936,In_1309);
and U2871 (N_2871,In_956,In_1076);
nand U2872 (N_2872,In_523,In_1033);
nand U2873 (N_2873,In_1293,In_500);
or U2874 (N_2874,In_1116,In_452);
xor U2875 (N_2875,In_1174,In_546);
nor U2876 (N_2876,In_274,In_303);
xnor U2877 (N_2877,In_382,In_613);
or U2878 (N_2878,In_1384,In_511);
and U2879 (N_2879,In_399,In_791);
and U2880 (N_2880,In_6,In_769);
or U2881 (N_2881,In_1051,In_1353);
or U2882 (N_2882,In_1057,In_1177);
nor U2883 (N_2883,In_889,In_639);
or U2884 (N_2884,In_1088,In_1394);
nor U2885 (N_2885,In_1450,In_787);
nand U2886 (N_2886,In_1234,In_424);
or U2887 (N_2887,In_106,In_25);
nor U2888 (N_2888,In_457,In_195);
or U2889 (N_2889,In_547,In_1323);
nor U2890 (N_2890,In_999,In_203);
and U2891 (N_2891,In_70,In_964);
nor U2892 (N_2892,In_902,In_426);
nor U2893 (N_2893,In_707,In_199);
nor U2894 (N_2894,In_724,In_1443);
or U2895 (N_2895,In_486,In_520);
or U2896 (N_2896,In_954,In_1298);
and U2897 (N_2897,In_1312,In_1211);
xnor U2898 (N_2898,In_278,In_869);
xnor U2899 (N_2899,In_1482,In_1006);
or U2900 (N_2900,In_301,In_1361);
nand U2901 (N_2901,In_549,In_1441);
nor U2902 (N_2902,In_749,In_70);
and U2903 (N_2903,In_1315,In_852);
or U2904 (N_2904,In_495,In_1311);
or U2905 (N_2905,In_44,In_1430);
nor U2906 (N_2906,In_439,In_1083);
nand U2907 (N_2907,In_1276,In_1151);
and U2908 (N_2908,In_700,In_812);
nor U2909 (N_2909,In_124,In_1267);
nand U2910 (N_2910,In_1497,In_237);
and U2911 (N_2911,In_1205,In_1123);
nand U2912 (N_2912,In_884,In_990);
or U2913 (N_2913,In_315,In_411);
and U2914 (N_2914,In_435,In_691);
or U2915 (N_2915,In_721,In_1454);
nor U2916 (N_2916,In_890,In_455);
nand U2917 (N_2917,In_1195,In_745);
or U2918 (N_2918,In_1006,In_483);
nand U2919 (N_2919,In_1240,In_854);
nand U2920 (N_2920,In_1158,In_211);
nand U2921 (N_2921,In_150,In_958);
nand U2922 (N_2922,In_914,In_185);
nor U2923 (N_2923,In_522,In_409);
nor U2924 (N_2924,In_86,In_726);
nand U2925 (N_2925,In_556,In_570);
and U2926 (N_2926,In_278,In_1040);
xor U2927 (N_2927,In_1270,In_889);
and U2928 (N_2928,In_952,In_320);
and U2929 (N_2929,In_496,In_1465);
nor U2930 (N_2930,In_228,In_726);
nor U2931 (N_2931,In_1135,In_1210);
nor U2932 (N_2932,In_891,In_927);
and U2933 (N_2933,In_37,In_482);
nand U2934 (N_2934,In_352,In_1113);
or U2935 (N_2935,In_1412,In_1325);
nor U2936 (N_2936,In_473,In_110);
or U2937 (N_2937,In_260,In_475);
nand U2938 (N_2938,In_275,In_857);
nor U2939 (N_2939,In_1081,In_696);
nor U2940 (N_2940,In_431,In_821);
and U2941 (N_2941,In_506,In_342);
and U2942 (N_2942,In_773,In_1445);
nor U2943 (N_2943,In_228,In_81);
nor U2944 (N_2944,In_615,In_1308);
nand U2945 (N_2945,In_1104,In_267);
xor U2946 (N_2946,In_257,In_358);
nor U2947 (N_2947,In_1166,In_944);
nand U2948 (N_2948,In_869,In_715);
nor U2949 (N_2949,In_821,In_1374);
and U2950 (N_2950,In_629,In_552);
nor U2951 (N_2951,In_84,In_1376);
and U2952 (N_2952,In_1177,In_1051);
nor U2953 (N_2953,In_621,In_119);
xor U2954 (N_2954,In_116,In_813);
and U2955 (N_2955,In_1156,In_1170);
and U2956 (N_2956,In_635,In_335);
nand U2957 (N_2957,In_1404,In_438);
nor U2958 (N_2958,In_1141,In_898);
or U2959 (N_2959,In_373,In_1170);
and U2960 (N_2960,In_769,In_106);
nand U2961 (N_2961,In_330,In_1015);
nor U2962 (N_2962,In_1432,In_993);
nand U2963 (N_2963,In_1208,In_1407);
or U2964 (N_2964,In_284,In_155);
xnor U2965 (N_2965,In_148,In_488);
nor U2966 (N_2966,In_740,In_1410);
or U2967 (N_2967,In_318,In_1039);
or U2968 (N_2968,In_395,In_426);
or U2969 (N_2969,In_1320,In_1431);
or U2970 (N_2970,In_1126,In_1188);
and U2971 (N_2971,In_1013,In_98);
or U2972 (N_2972,In_391,In_856);
nand U2973 (N_2973,In_1204,In_716);
nor U2974 (N_2974,In_1089,In_377);
or U2975 (N_2975,In_758,In_699);
or U2976 (N_2976,In_789,In_189);
nor U2977 (N_2977,In_404,In_1120);
or U2978 (N_2978,In_600,In_588);
nand U2979 (N_2979,In_1063,In_1377);
nor U2980 (N_2980,In_1225,In_485);
and U2981 (N_2981,In_371,In_574);
xor U2982 (N_2982,In_146,In_1339);
xnor U2983 (N_2983,In_762,In_1037);
and U2984 (N_2984,In_689,In_668);
nand U2985 (N_2985,In_976,In_854);
or U2986 (N_2986,In_325,In_1050);
nor U2987 (N_2987,In_371,In_1168);
xnor U2988 (N_2988,In_735,In_842);
nand U2989 (N_2989,In_167,In_482);
and U2990 (N_2990,In_43,In_118);
xnor U2991 (N_2991,In_680,In_1068);
nor U2992 (N_2992,In_110,In_1483);
and U2993 (N_2993,In_945,In_1132);
or U2994 (N_2994,In_615,In_1080);
and U2995 (N_2995,In_49,In_525);
nand U2996 (N_2996,In_962,In_1087);
nand U2997 (N_2997,In_642,In_616);
xnor U2998 (N_2998,In_1394,In_821);
and U2999 (N_2999,In_5,In_677);
xnor U3000 (N_3000,N_525,N_2201);
nor U3001 (N_3001,N_1911,N_697);
nand U3002 (N_3002,N_2322,N_107);
and U3003 (N_3003,N_1220,N_433);
nand U3004 (N_3004,N_2332,N_2946);
nand U3005 (N_3005,N_298,N_1265);
nand U3006 (N_3006,N_1039,N_2816);
nand U3007 (N_3007,N_2141,N_1653);
or U3008 (N_3008,N_1584,N_1199);
and U3009 (N_3009,N_2503,N_402);
nand U3010 (N_3010,N_1908,N_2040);
and U3011 (N_3011,N_508,N_1967);
nand U3012 (N_3012,N_350,N_2694);
nand U3013 (N_3013,N_2840,N_2776);
or U3014 (N_3014,N_757,N_1375);
and U3015 (N_3015,N_2680,N_2249);
nor U3016 (N_3016,N_2510,N_1001);
nand U3017 (N_3017,N_2357,N_1172);
and U3018 (N_3018,N_84,N_554);
and U3019 (N_3019,N_2127,N_1512);
and U3020 (N_3020,N_1500,N_1705);
nor U3021 (N_3021,N_1390,N_2793);
xnor U3022 (N_3022,N_516,N_2049);
and U3023 (N_3023,N_2482,N_2651);
and U3024 (N_3024,N_122,N_224);
and U3025 (N_3025,N_2595,N_1515);
nand U3026 (N_3026,N_507,N_2956);
xor U3027 (N_3027,N_1591,N_1429);
nand U3028 (N_3028,N_174,N_502);
and U3029 (N_3029,N_247,N_943);
and U3030 (N_3030,N_2571,N_1754);
nand U3031 (N_3031,N_1863,N_2874);
or U3032 (N_3032,N_932,N_1791);
nand U3033 (N_3033,N_2847,N_1054);
nand U3034 (N_3034,N_2205,N_2262);
xnor U3035 (N_3035,N_801,N_1113);
nand U3036 (N_3036,N_1816,N_130);
and U3037 (N_3037,N_2621,N_1782);
nand U3038 (N_3038,N_2354,N_810);
or U3039 (N_3039,N_1813,N_445);
and U3040 (N_3040,N_2137,N_116);
and U3041 (N_3041,N_483,N_2033);
and U3042 (N_3042,N_2182,N_1477);
xnor U3043 (N_3043,N_1872,N_836);
nand U3044 (N_3044,N_578,N_2740);
nor U3045 (N_3045,N_1451,N_2626);
or U3046 (N_3046,N_1472,N_1431);
nand U3047 (N_3047,N_2094,N_2412);
nor U3048 (N_3048,N_990,N_944);
nor U3049 (N_3049,N_1481,N_2544);
and U3050 (N_3050,N_2574,N_1651);
xor U3051 (N_3051,N_2446,N_1005);
or U3052 (N_3052,N_1049,N_119);
and U3053 (N_3053,N_2071,N_1819);
nand U3054 (N_3054,N_2032,N_1264);
or U3055 (N_3055,N_1938,N_1405);
or U3056 (N_3056,N_2752,N_667);
or U3057 (N_3057,N_1915,N_475);
nor U3058 (N_3058,N_115,N_2742);
nor U3059 (N_3059,N_2778,N_329);
or U3060 (N_3060,N_925,N_745);
nor U3061 (N_3061,N_55,N_538);
nor U3062 (N_3062,N_933,N_887);
nor U3063 (N_3063,N_539,N_735);
and U3064 (N_3064,N_2416,N_297);
xnor U3065 (N_3065,N_480,N_684);
nand U3066 (N_3066,N_2961,N_2817);
and U3067 (N_3067,N_1457,N_573);
nand U3068 (N_3068,N_821,N_1288);
or U3069 (N_3069,N_2132,N_491);
and U3070 (N_3070,N_2393,N_63);
nand U3071 (N_3071,N_1870,N_518);
nand U3072 (N_3072,N_2161,N_861);
nor U3073 (N_3073,N_909,N_2430);
xor U3074 (N_3074,N_1180,N_775);
and U3075 (N_3075,N_929,N_1256);
or U3076 (N_3076,N_565,N_2226);
or U3077 (N_3077,N_2538,N_1888);
nor U3078 (N_3078,N_30,N_551);
nand U3079 (N_3079,N_172,N_1469);
nor U3080 (N_3080,N_1459,N_1885);
or U3081 (N_3081,N_64,N_2310);
or U3082 (N_3082,N_2466,N_1369);
or U3083 (N_3083,N_737,N_526);
nand U3084 (N_3084,N_1035,N_1984);
or U3085 (N_3085,N_1499,N_1421);
or U3086 (N_3086,N_278,N_210);
and U3087 (N_3087,N_1731,N_779);
and U3088 (N_3088,N_1023,N_16);
and U3089 (N_3089,N_979,N_1823);
nor U3090 (N_3090,N_147,N_270);
nor U3091 (N_3091,N_1510,N_2986);
nand U3092 (N_3092,N_1461,N_1218);
nand U3093 (N_3093,N_1917,N_666);
and U3094 (N_3094,N_957,N_2819);
and U3095 (N_3095,N_1935,N_830);
nand U3096 (N_3096,N_2667,N_2689);
nand U3097 (N_3097,N_1024,N_837);
nor U3098 (N_3098,N_1126,N_2663);
and U3099 (N_3099,N_2285,N_2916);
nand U3100 (N_3100,N_785,N_2359);
nor U3101 (N_3101,N_2758,N_780);
xor U3102 (N_3102,N_82,N_1835);
or U3103 (N_3103,N_953,N_2634);
xnor U3104 (N_3104,N_1290,N_56);
and U3105 (N_3105,N_2494,N_1815);
or U3106 (N_3106,N_2060,N_1799);
nor U3107 (N_3107,N_2418,N_2832);
nand U3108 (N_3108,N_704,N_62);
or U3109 (N_3109,N_2526,N_257);
or U3110 (N_3110,N_1620,N_308);
nand U3111 (N_3111,N_342,N_593);
nor U3112 (N_3112,N_1454,N_1777);
nor U3113 (N_3113,N_2435,N_1190);
xnor U3114 (N_3114,N_2933,N_739);
or U3115 (N_3115,N_1261,N_146);
nor U3116 (N_3116,N_668,N_1797);
and U3117 (N_3117,N_2330,N_1743);
and U3118 (N_3118,N_1853,N_1843);
nand U3119 (N_3119,N_412,N_1950);
or U3120 (N_3120,N_2400,N_2247);
nand U3121 (N_3121,N_42,N_2575);
and U3122 (N_3122,N_101,N_2318);
and U3123 (N_3123,N_1167,N_2893);
nand U3124 (N_3124,N_838,N_898);
and U3125 (N_3125,N_288,N_1013);
and U3126 (N_3126,N_817,N_2973);
or U3127 (N_3127,N_723,N_1123);
nand U3128 (N_3128,N_1478,N_1166);
nor U3129 (N_3129,N_2671,N_2925);
nand U3130 (N_3130,N_339,N_818);
nand U3131 (N_3131,N_1897,N_2851);
and U3132 (N_3132,N_309,N_422);
and U3133 (N_3133,N_2200,N_27);
nor U3134 (N_3134,N_499,N_613);
nor U3135 (N_3135,N_1525,N_141);
xor U3136 (N_3136,N_908,N_897);
nor U3137 (N_3137,N_2438,N_131);
or U3138 (N_3138,N_450,N_819);
or U3139 (N_3139,N_2347,N_1131);
nor U3140 (N_3140,N_425,N_1466);
and U3141 (N_3141,N_1845,N_826);
and U3142 (N_3142,N_2422,N_1331);
or U3143 (N_3143,N_1277,N_2950);
nor U3144 (N_3144,N_2399,N_2809);
and U3145 (N_3145,N_1505,N_2241);
nor U3146 (N_3146,N_2949,N_2609);
nor U3147 (N_3147,N_2209,N_547);
nor U3148 (N_3148,N_2484,N_157);
or U3149 (N_3149,N_1953,N_2186);
nor U3150 (N_3150,N_2815,N_2214);
and U3151 (N_3151,N_768,N_520);
and U3152 (N_3152,N_1271,N_594);
and U3153 (N_3153,N_7,N_1255);
and U3154 (N_3154,N_2632,N_687);
nor U3155 (N_3155,N_2193,N_1934);
and U3156 (N_3156,N_2918,N_2644);
and U3157 (N_3157,N_604,N_992);
and U3158 (N_3158,N_2829,N_514);
and U3159 (N_3159,N_1895,N_1055);
nor U3160 (N_3160,N_243,N_2795);
or U3161 (N_3161,N_2647,N_1502);
and U3162 (N_3162,N_345,N_2695);
nor U3163 (N_3163,N_1086,N_1089);
and U3164 (N_3164,N_653,N_2566);
nand U3165 (N_3165,N_2867,N_344);
or U3166 (N_3166,N_1877,N_476);
and U3167 (N_3167,N_1043,N_2062);
or U3168 (N_3168,N_2869,N_474);
or U3169 (N_3169,N_1419,N_2042);
nand U3170 (N_3170,N_1983,N_1031);
or U3171 (N_3171,N_1338,N_1606);
nor U3172 (N_3172,N_874,N_572);
and U3173 (N_3173,N_2501,N_189);
and U3174 (N_3174,N_2424,N_2581);
nand U3175 (N_3175,N_1626,N_948);
nor U3176 (N_3176,N_2089,N_788);
nor U3177 (N_3177,N_198,N_2230);
or U3178 (N_3178,N_2618,N_2822);
nor U3179 (N_3179,N_2155,N_873);
and U3180 (N_3180,N_466,N_41);
or U3181 (N_3181,N_936,N_2602);
nor U3182 (N_3182,N_1156,N_451);
or U3183 (N_3183,N_2272,N_1016);
or U3184 (N_3184,N_2520,N_1268);
and U3185 (N_3185,N_1458,N_1471);
nor U3186 (N_3186,N_2459,N_1857);
and U3187 (N_3187,N_418,N_2716);
nand U3188 (N_3188,N_2440,N_1137);
or U3189 (N_3189,N_428,N_2004);
xor U3190 (N_3190,N_877,N_472);
nand U3191 (N_3191,N_2135,N_982);
and U3192 (N_3192,N_1337,N_1786);
nand U3193 (N_3193,N_652,N_2326);
and U3194 (N_3194,N_915,N_232);
nand U3195 (N_3195,N_678,N_235);
and U3196 (N_3196,N_1493,N_803);
nand U3197 (N_3197,N_1990,N_439);
nand U3198 (N_3198,N_1922,N_732);
nor U3199 (N_3199,N_204,N_1600);
nand U3200 (N_3200,N_1683,N_2468);
nand U3201 (N_3201,N_252,N_1794);
and U3202 (N_3202,N_2288,N_1107);
nor U3203 (N_3203,N_1298,N_2368);
xor U3204 (N_3204,N_2331,N_1412);
and U3205 (N_3205,N_1132,N_2294);
nand U3206 (N_3206,N_1989,N_2080);
nor U3207 (N_3207,N_2997,N_1355);
nor U3208 (N_3208,N_1809,N_1102);
nor U3209 (N_3209,N_1859,N_748);
and U3210 (N_3210,N_1291,N_512);
or U3211 (N_3211,N_2382,N_2843);
and U3212 (N_3212,N_2989,N_2050);
or U3213 (N_3213,N_1785,N_799);
or U3214 (N_3214,N_1974,N_1424);
nand U3215 (N_3215,N_105,N_2369);
or U3216 (N_3216,N_1221,N_1836);
nor U3217 (N_3217,N_2572,N_470);
nand U3218 (N_3218,N_1657,N_1962);
xor U3219 (N_3219,N_2649,N_113);
and U3220 (N_3220,N_1345,N_1691);
nand U3221 (N_3221,N_31,N_1322);
nand U3222 (N_3222,N_2396,N_556);
and U3223 (N_3223,N_1452,N_1904);
nor U3224 (N_3224,N_506,N_2124);
and U3225 (N_3225,N_2990,N_614);
nor U3226 (N_3226,N_1028,N_383);
and U3227 (N_3227,N_2523,N_2407);
nand U3228 (N_3228,N_487,N_711);
nor U3229 (N_3229,N_588,N_1728);
or U3230 (N_3230,N_2748,N_1844);
nand U3231 (N_3231,N_872,N_2115);
xnor U3232 (N_3232,N_1425,N_2111);
or U3233 (N_3233,N_44,N_277);
or U3234 (N_3234,N_820,N_380);
or U3235 (N_3235,N_2473,N_746);
nor U3236 (N_3236,N_2275,N_1491);
or U3237 (N_3237,N_2022,N_1002);
xnor U3238 (N_3238,N_1427,N_2163);
nor U3239 (N_3239,N_665,N_1432);
nor U3240 (N_3240,N_1931,N_1656);
nor U3241 (N_3241,N_592,N_1630);
and U3242 (N_3242,N_2063,N_579);
nor U3243 (N_3243,N_435,N_2592);
nand U3244 (N_3244,N_164,N_2336);
nand U3245 (N_3245,N_1542,N_1968);
or U3246 (N_3246,N_2659,N_2530);
nor U3247 (N_3247,N_2653,N_231);
or U3248 (N_3248,N_1940,N_1475);
or U3249 (N_3249,N_314,N_2219);
nand U3250 (N_3250,N_2968,N_844);
nand U3251 (N_3251,N_1926,N_1352);
or U3252 (N_3252,N_1531,N_2577);
and U3253 (N_3253,N_2614,N_2560);
or U3254 (N_3254,N_619,N_2029);
or U3255 (N_3255,N_1581,N_1849);
nor U3256 (N_3256,N_1108,N_1313);
or U3257 (N_3257,N_2547,N_1894);
nor U3258 (N_3258,N_1441,N_906);
nor U3259 (N_3259,N_1018,N_2008);
or U3260 (N_3260,N_712,N_1411);
or U3261 (N_3261,N_279,N_1456);
nor U3262 (N_3262,N_2669,N_2744);
and U3263 (N_3263,N_1530,N_557);
or U3264 (N_3264,N_2512,N_813);
or U3265 (N_3265,N_2162,N_1186);
or U3266 (N_3266,N_1391,N_201);
nor U3267 (N_3267,N_13,N_59);
xor U3268 (N_3268,N_1566,N_609);
or U3269 (N_3269,N_706,N_312);
nand U3270 (N_3270,N_276,N_2091);
and U3271 (N_3271,N_1747,N_1360);
nand U3272 (N_3272,N_1476,N_617);
xor U3273 (N_3273,N_913,N_217);
and U3274 (N_3274,N_1628,N_726);
nand U3275 (N_3275,N_1947,N_2725);
or U3276 (N_3276,N_2180,N_2909);
and U3277 (N_3277,N_2726,N_354);
or U3278 (N_3278,N_376,N_1029);
nand U3279 (N_3279,N_1992,N_134);
nand U3280 (N_3280,N_756,N_750);
and U3281 (N_3281,N_1160,N_1625);
nor U3282 (N_3282,N_2700,N_169);
or U3283 (N_3283,N_2979,N_2567);
xor U3284 (N_3284,N_1960,N_2048);
or U3285 (N_3285,N_644,N_1608);
nor U3286 (N_3286,N_2849,N_1539);
or U3287 (N_3287,N_2858,N_950);
nor U3288 (N_3288,N_2442,N_2969);
nor U3289 (N_3289,N_390,N_1346);
and U3290 (N_3290,N_494,N_2761);
nand U3291 (N_3291,N_1563,N_103);
nand U3292 (N_3292,N_632,N_2100);
and U3293 (N_3293,N_2388,N_50);
nor U3294 (N_3294,N_2786,N_178);
or U3295 (N_3295,N_1891,N_151);
and U3296 (N_3296,N_88,N_2469);
and U3297 (N_3297,N_1184,N_1715);
and U3298 (N_3298,N_362,N_2421);
or U3299 (N_3299,N_533,N_1116);
nand U3300 (N_3300,N_2084,N_1623);
or U3301 (N_3301,N_1202,N_2806);
nor U3302 (N_3302,N_1096,N_2590);
and U3303 (N_3303,N_2065,N_2184);
nor U3304 (N_3304,N_548,N_2178);
and U3305 (N_3305,N_2707,N_2114);
or U3306 (N_3306,N_424,N_771);
and U3307 (N_3307,N_1003,N_66);
nand U3308 (N_3308,N_2565,N_701);
nor U3309 (N_3309,N_1052,N_2537);
nand U3310 (N_3310,N_1504,N_1253);
or U3311 (N_3311,N_688,N_2967);
or U3312 (N_3312,N_2489,N_870);
and U3313 (N_3313,N_927,N_2225);
or U3314 (N_3314,N_1660,N_1701);
nor U3315 (N_3315,N_1364,N_355);
nand U3316 (N_3316,N_500,N_1604);
nor U3317 (N_3317,N_1730,N_2656);
nand U3318 (N_3318,N_1293,N_1388);
and U3319 (N_3319,N_2931,N_2677);
nand U3320 (N_3320,N_2894,N_148);
nor U3321 (N_3321,N_370,N_484);
and U3322 (N_3322,N_1286,N_1263);
nand U3323 (N_3323,N_2823,N_2055);
and U3324 (N_3324,N_521,N_485);
and U3325 (N_3325,N_1729,N_479);
and U3326 (N_3326,N_2,N_2585);
nand U3327 (N_3327,N_1215,N_2044);
nor U3328 (N_3328,N_2386,N_2349);
and U3329 (N_3329,N_248,N_2682);
xor U3330 (N_3330,N_1841,N_1529);
nand U3331 (N_3331,N_2499,N_1341);
nand U3332 (N_3332,N_2522,N_938);
and U3333 (N_3333,N_843,N_316);
nand U3334 (N_3334,N_2911,N_2654);
or U3335 (N_3335,N_332,N_1666);
xnor U3336 (N_3336,N_1042,N_156);
nor U3337 (N_3337,N_2687,N_498);
and U3338 (N_3338,N_659,N_1828);
nand U3339 (N_3339,N_132,N_2298);
nor U3340 (N_3340,N_2692,N_997);
and U3341 (N_3341,N_1485,N_2899);
or U3342 (N_3342,N_2491,N_33);
or U3343 (N_3343,N_274,N_2658);
and U3344 (N_3344,N_1925,N_2160);
nand U3345 (N_3345,N_2710,N_2437);
nand U3346 (N_3346,N_335,N_2953);
or U3347 (N_3347,N_1796,N_1074);
and U3348 (N_3348,N_2199,N_2945);
or U3349 (N_3349,N_19,N_2263);
and U3350 (N_3350,N_582,N_850);
or U3351 (N_3351,N_2993,N_1898);
xor U3352 (N_3352,N_2943,N_1060);
or U3353 (N_3353,N_2756,N_1362);
or U3354 (N_3354,N_411,N_97);
nor U3355 (N_3355,N_2037,N_456);
or U3356 (N_3356,N_2980,N_1348);
and U3357 (N_3357,N_1101,N_2923);
xor U3358 (N_3358,N_437,N_2739);
xor U3359 (N_3359,N_2777,N_2690);
or U3360 (N_3360,N_2377,N_2248);
and U3361 (N_3361,N_2939,N_1304);
nor U3362 (N_3362,N_2176,N_1862);
and U3363 (N_3363,N_1704,N_1387);
or U3364 (N_3364,N_1463,N_696);
nor U3365 (N_3365,N_1899,N_919);
nand U3366 (N_3366,N_391,N_2836);
and U3367 (N_3367,N_1244,N_399);
nor U3368 (N_3368,N_1150,N_2106);
and U3369 (N_3369,N_2373,N_692);
nor U3370 (N_3370,N_1098,N_777);
or U3371 (N_3371,N_1027,N_1311);
and U3372 (N_3372,N_37,N_2625);
and U3373 (N_3373,N_2211,N_1869);
or U3374 (N_3374,N_5,N_2947);
or U3375 (N_3375,N_845,N_2720);
and U3376 (N_3376,N_1945,N_2951);
nand U3377 (N_3377,N_2165,N_715);
nor U3378 (N_3378,N_2741,N_2808);
or U3379 (N_3379,N_2676,N_2315);
and U3380 (N_3380,N_1490,N_1384);
xor U3381 (N_3381,N_2427,N_2884);
nor U3382 (N_3382,N_2928,N_1295);
nor U3383 (N_3383,N_1713,N_2805);
or U3384 (N_3384,N_333,N_705);
xor U3385 (N_3385,N_2492,N_1336);
and U3386 (N_3386,N_461,N_952);
and U3387 (N_3387,N_612,N_51);
and U3388 (N_3388,N_623,N_1408);
and U3389 (N_3389,N_1112,N_544);
or U3390 (N_3390,N_607,N_2245);
or U3391 (N_3391,N_2172,N_2696);
nor U3392 (N_3392,N_1639,N_420);
nand U3393 (N_3393,N_1981,N_2559);
and U3394 (N_3394,N_2835,N_2151);
xor U3395 (N_3395,N_860,N_1738);
and U3396 (N_3396,N_1280,N_94);
or U3397 (N_3397,N_2324,N_1946);
nand U3398 (N_3398,N_2637,N_1978);
or U3399 (N_3399,N_1414,N_438);
nand U3400 (N_3400,N_834,N_2167);
nand U3401 (N_3401,N_1114,N_382);
or U3402 (N_3402,N_1309,N_2088);
and U3403 (N_3403,N_1335,N_1072);
xnor U3404 (N_3404,N_2238,N_1225);
nand U3405 (N_3405,N_2675,N_357);
xor U3406 (N_3406,N_2477,N_2803);
nand U3407 (N_3407,N_2086,N_328);
and U3408 (N_3408,N_313,N_1171);
and U3409 (N_3409,N_2766,N_492);
nor U3410 (N_3410,N_1178,N_2028);
nand U3411 (N_3411,N_1846,N_244);
or U3412 (N_3412,N_2098,N_1874);
nand U3413 (N_3413,N_2255,N_1544);
nand U3414 (N_3414,N_1327,N_326);
nor U3415 (N_3415,N_1679,N_2759);
or U3416 (N_3416,N_2092,N_440);
or U3417 (N_3417,N_2150,N_2066);
nor U3418 (N_3418,N_1567,N_2011);
or U3419 (N_3419,N_1987,N_310);
and U3420 (N_3420,N_2453,N_1507);
and U3421 (N_3421,N_912,N_2772);
or U3422 (N_3422,N_2838,N_2578);
nor U3423 (N_3423,N_2233,N_1995);
or U3424 (N_3424,N_2171,N_2307);
xor U3425 (N_3425,N_2356,N_2306);
nor U3426 (N_3426,N_1927,N_1251);
nor U3427 (N_3427,N_441,N_1808);
nor U3428 (N_3428,N_1189,N_585);
nand U3429 (N_3429,N_1370,N_2814);
and U3430 (N_3430,N_1564,N_2058);
or U3431 (N_3431,N_1445,N_1855);
or U3432 (N_3432,N_2215,N_1323);
or U3433 (N_3433,N_2846,N_1206);
nand U3434 (N_3434,N_2765,N_1622);
or U3435 (N_3435,N_208,N_2449);
nor U3436 (N_3436,N_2735,N_1587);
and U3437 (N_3437,N_258,N_1737);
or U3438 (N_3438,N_1867,N_1208);
or U3439 (N_3439,N_11,N_1589);
or U3440 (N_3440,N_852,N_1550);
and U3441 (N_3441,N_2964,N_1964);
or U3442 (N_3442,N_2379,N_2591);
nand U3443 (N_3443,N_1140,N_1183);
xnor U3444 (N_3444,N_1484,N_1736);
or U3445 (N_3445,N_904,N_597);
and U3446 (N_3446,N_2782,N_2246);
nand U3447 (N_3447,N_1068,N_1514);
nor U3448 (N_3448,N_626,N_136);
nor U3449 (N_3449,N_738,N_117);
nand U3450 (N_3450,N_2952,N_975);
nand U3451 (N_3451,N_1822,N_513);
nor U3452 (N_3452,N_656,N_1325);
and U3453 (N_3453,N_459,N_846);
xor U3454 (N_3454,N_793,N_1278);
nor U3455 (N_3455,N_2932,N_1793);
and U3456 (N_3456,N_1924,N_1257);
nor U3457 (N_3457,N_2987,N_1125);
nand U3458 (N_3458,N_1032,N_1821);
or U3459 (N_3459,N_956,N_1385);
or U3460 (N_3460,N_2763,N_985);
xnor U3461 (N_3461,N_48,N_2441);
or U3462 (N_3462,N_2563,N_2069);
or U3463 (N_3463,N_1267,N_2075);
nand U3464 (N_3464,N_21,N_1501);
or U3465 (N_3465,N_336,N_2717);
nand U3466 (N_3466,N_1076,N_2460);
nor U3467 (N_3467,N_2960,N_108);
xor U3468 (N_3468,N_2363,N_758);
nand U3469 (N_3469,N_2733,N_662);
or U3470 (N_3470,N_976,N_1465);
or U3471 (N_3471,N_2768,N_2751);
and U3472 (N_3472,N_2606,N_2804);
nand U3473 (N_3473,N_416,N_2556);
and U3474 (N_3474,N_1426,N_892);
or U3475 (N_3475,N_220,N_1443);
nor U3476 (N_3476,N_522,N_849);
nand U3477 (N_3477,N_1307,N_75);
and U3478 (N_3478,N_2206,N_960);
and U3479 (N_3479,N_546,N_2589);
nor U3480 (N_3480,N_67,N_1590);
nor U3481 (N_3481,N_1741,N_1854);
and U3482 (N_3482,N_2593,N_1858);
and U3483 (N_3483,N_57,N_1109);
or U3484 (N_3484,N_303,N_2660);
nor U3485 (N_3485,N_1966,N_2096);
or U3486 (N_3486,N_1674,N_401);
or U3487 (N_3487,N_713,N_2021);
and U3488 (N_3488,N_1332,N_2301);
nor U3489 (N_3489,N_528,N_888);
nand U3490 (N_3490,N_2810,N_1528);
xor U3491 (N_3491,N_504,N_866);
and U3492 (N_3492,N_176,N_797);
nand U3493 (N_3493,N_924,N_1672);
or U3494 (N_3494,N_1410,N_882);
nor U3495 (N_3495,N_1795,N_414);
or U3496 (N_3496,N_2149,N_2177);
or U3497 (N_3497,N_1040,N_2885);
and U3498 (N_3498,N_807,N_2630);
and U3499 (N_3499,N_2865,N_2333);
nor U3500 (N_3500,N_47,N_2857);
xnor U3501 (N_3501,N_847,N_740);
xor U3502 (N_3502,N_2540,N_690);
nor U3503 (N_3503,N_2546,N_381);
nand U3504 (N_3504,N_1866,N_1138);
xnor U3505 (N_3505,N_2221,N_1876);
nand U3506 (N_3506,N_962,N_629);
and U3507 (N_3507,N_4,N_1297);
or U3508 (N_3508,N_417,N_2103);
and U3509 (N_3509,N_2254,N_2024);
and U3510 (N_3510,N_1686,N_2862);
or U3511 (N_3511,N_1861,N_1474);
or U3512 (N_3512,N_2072,N_226);
or U3513 (N_3513,N_165,N_2600);
xor U3514 (N_3514,N_2619,N_2746);
or U3515 (N_3515,N_1779,N_2788);
nor U3516 (N_3516,N_123,N_2616);
nand U3517 (N_3517,N_1618,N_1269);
or U3518 (N_3518,N_2320,N_24);
or U3519 (N_3519,N_1727,N_1605);
nand U3520 (N_3520,N_856,N_222);
or U3521 (N_3521,N_2374,N_1554);
nand U3522 (N_3522,N_100,N_2723);
or U3523 (N_3523,N_2411,N_763);
nand U3524 (N_3524,N_1204,N_2929);
nor U3525 (N_3525,N_2216,N_2038);
or U3526 (N_3526,N_398,N_1763);
xnor U3527 (N_3527,N_1046,N_2352);
nand U3528 (N_3528,N_1033,N_1243);
and U3529 (N_3529,N_851,N_2470);
nor U3530 (N_3530,N_240,N_2371);
and U3531 (N_3531,N_2991,N_266);
or U3532 (N_3532,N_163,N_1996);
and U3533 (N_3533,N_970,N_549);
nand U3534 (N_3534,N_1889,N_1670);
and U3535 (N_3535,N_1752,N_343);
nand U3536 (N_3536,N_2429,N_2534);
and U3537 (N_3537,N_651,N_1732);
nor U3538 (N_3538,N_1181,N_1585);
xnor U3539 (N_3539,N_2433,N_2325);
or U3540 (N_3540,N_2615,N_2781);
nor U3541 (N_3541,N_1025,N_2047);
or U3542 (N_3542,N_1582,N_273);
or U3543 (N_3543,N_90,N_2224);
nand U3544 (N_3544,N_1609,N_940);
or U3545 (N_3545,N_1668,N_25);
nor U3546 (N_3546,N_1308,N_159);
and U3547 (N_3547,N_2490,N_2525);
nor U3548 (N_3548,N_2164,N_2513);
and U3549 (N_3549,N_1942,N_670);
nand U3550 (N_3550,N_559,N_640);
or U3551 (N_3551,N_1214,N_1367);
and U3552 (N_3552,N_893,N_937);
nand U3553 (N_3553,N_294,N_1494);
or U3554 (N_3554,N_2025,N_1326);
and U3555 (N_3555,N_2866,N_2749);
nand U3556 (N_3556,N_1229,N_1928);
or U3557 (N_3557,N_229,N_1759);
or U3558 (N_3558,N_718,N_36);
xor U3559 (N_3559,N_1073,N_1266);
or U3560 (N_3560,N_2476,N_2841);
nand U3561 (N_3561,N_388,N_2212);
nand U3562 (N_3562,N_1416,N_1179);
nand U3563 (N_3563,N_2284,N_1742);
nand U3564 (N_3564,N_1239,N_2539);
nor U3565 (N_3565,N_964,N_537);
nor U3566 (N_3566,N_2498,N_2934);
nor U3567 (N_3567,N_15,N_1919);
and U3568 (N_3568,N_465,N_2295);
nor U3569 (N_3569,N_1780,N_1580);
nand U3570 (N_3570,N_1547,N_349);
and U3571 (N_3571,N_430,N_1087);
or U3572 (N_3572,N_322,N_809);
or U3573 (N_3573,N_1555,N_591);
nand U3574 (N_3574,N_1690,N_1506);
xnor U3575 (N_3575,N_595,N_2718);
xnor U3576 (N_3576,N_52,N_1805);
xor U3577 (N_3577,N_1062,N_2236);
or U3578 (N_3578,N_1932,N_2531);
and U3579 (N_3579,N_2773,N_1051);
and U3580 (N_3580,N_1305,N_463);
or U3581 (N_3581,N_262,N_1719);
nand U3582 (N_3582,N_816,N_2235);
xor U3583 (N_3583,N_228,N_543);
xor U3584 (N_3584,N_2147,N_2023);
nor U3585 (N_3585,N_452,N_389);
or U3586 (N_3586,N_875,N_2890);
and U3587 (N_3587,N_2289,N_2903);
nand U3588 (N_3588,N_1083,N_947);
or U3589 (N_3589,N_647,N_324);
or U3590 (N_3590,N_734,N_2445);
xnor U3591 (N_3591,N_2688,N_20);
or U3592 (N_3592,N_2678,N_1744);
nor U3593 (N_3593,N_783,N_550);
or U3594 (N_3594,N_280,N_1467);
and U3595 (N_3595,N_1053,N_1274);
and U3596 (N_3596,N_170,N_2978);
nand U3597 (N_3597,N_410,N_1115);
and U3598 (N_3598,N_2902,N_2603);
nand U3599 (N_3599,N_2737,N_722);
xnor U3600 (N_3600,N_2919,N_1397);
nor U3601 (N_3601,N_621,N_1464);
nor U3602 (N_3602,N_1883,N_1147);
or U3603 (N_3603,N_1110,N_1201);
nand U3604 (N_3604,N_1586,N_1971);
or U3605 (N_3605,N_2850,N_2981);
xor U3606 (N_3606,N_842,N_752);
nand U3607 (N_3607,N_1723,N_1698);
and U3608 (N_3608,N_1203,N_618);
nor U3609 (N_3609,N_1703,N_1428);
nand U3610 (N_3610,N_2936,N_731);
nand U3611 (N_3611,N_2533,N_2018);
or U3612 (N_3612,N_2260,N_152);
and U3613 (N_3613,N_2256,N_987);
nor U3614 (N_3614,N_1347,N_1120);
nor U3615 (N_3615,N_2300,N_1839);
and U3616 (N_3616,N_1603,N_1285);
nor U3617 (N_3617,N_2784,N_1058);
nor U3618 (N_3618,N_1879,N_584);
nand U3619 (N_3619,N_1447,N_1975);
and U3620 (N_3620,N_239,N_1673);
nand U3621 (N_3621,N_2913,N_2714);
or U3622 (N_3622,N_679,N_2633);
nand U3623 (N_3623,N_2118,N_832);
and U3624 (N_3624,N_2561,N_1568);
nor U3625 (N_3625,N_1216,N_2014);
xnor U3626 (N_3626,N_8,N_2830);
and U3627 (N_3627,N_996,N_2905);
nand U3628 (N_3628,N_1881,N_1219);
nor U3629 (N_3629,N_2940,N_2397);
and U3630 (N_3630,N_1556,N_635);
or U3631 (N_3631,N_900,N_129);
nand U3632 (N_3632,N_2994,N_300);
nor U3633 (N_3633,N_473,N_2787);
or U3634 (N_3634,N_736,N_2095);
nand U3635 (N_3635,N_1430,N_869);
nand U3636 (N_3636,N_1064,N_268);
or U3637 (N_3637,N_369,N_1914);
nor U3638 (N_3638,N_2504,N_2194);
or U3639 (N_3639,N_1814,N_202);
nor U3640 (N_3640,N_2521,N_415);
or U3641 (N_3641,N_1551,N_2582);
nand U3642 (N_3642,N_986,N_356);
and U3643 (N_3643,N_1511,N_918);
and U3644 (N_3644,N_978,N_2408);
or U3645 (N_3645,N_1050,N_1185);
nand U3646 (N_3646,N_1470,N_808);
nand U3647 (N_3647,N_787,N_2110);
and U3648 (N_3648,N_1404,N_2821);
or U3649 (N_3649,N_2785,N_2444);
and U3650 (N_3650,N_287,N_1575);
nor U3651 (N_3651,N_2030,N_1198);
nor U3652 (N_3652,N_2853,N_2061);
and U3653 (N_3653,N_917,N_2188);
or U3654 (N_3654,N_187,N_397);
nand U3655 (N_3655,N_1342,N_495);
nor U3656 (N_3656,N_1148,N_1127);
or U3657 (N_3657,N_2478,N_2910);
or U3658 (N_3658,N_2031,N_1733);
nand U3659 (N_3659,N_1571,N_454);
or U3660 (N_3660,N_137,N_2767);
nor U3661 (N_3661,N_2887,N_2281);
or U3662 (N_3662,N_2010,N_1757);
nor U3663 (N_3663,N_1383,N_1007);
and U3664 (N_3664,N_386,N_2204);
nor U3665 (N_3665,N_951,N_221);
nor U3666 (N_3666,N_432,N_998);
and U3667 (N_3667,N_1205,N_1906);
or U3668 (N_3668,N_1248,N_2922);
and U3669 (N_3669,N_2056,N_2057);
xnor U3670 (N_3670,N_227,N_773);
nand U3671 (N_3671,N_2898,N_74);
nand U3672 (N_3672,N_1661,N_1143);
and U3673 (N_3673,N_1306,N_2493);
or U3674 (N_3674,N_2738,N_1488);
or U3675 (N_3675,N_2629,N_606);
nand U3676 (N_3676,N_643,N_1078);
nor U3677 (N_3677,N_1769,N_1276);
or U3678 (N_3678,N_1831,N_2988);
or U3679 (N_3679,N_2834,N_1489);
nand U3680 (N_3680,N_1636,N_519);
or U3681 (N_3681,N_695,N_1070);
nand U3682 (N_3682,N_2000,N_2129);
and U3683 (N_3683,N_1923,N_1047);
nand U3684 (N_3684,N_804,N_1617);
nand U3685 (N_3685,N_2303,N_2750);
or U3686 (N_3686,N_1324,N_2068);
nor U3687 (N_3687,N_2328,N_2611);
nor U3688 (N_3688,N_1258,N_86);
or U3689 (N_3689,N_2941,N_884);
nor U3690 (N_3690,N_1233,N_1252);
nand U3691 (N_3691,N_1873,N_194);
xor U3692 (N_3692,N_2456,N_192);
or U3693 (N_3693,N_2975,N_963);
and U3694 (N_3694,N_1030,N_1545);
and U3695 (N_3695,N_2406,N_2562);
and U3696 (N_3696,N_1155,N_744);
nand U3697 (N_3697,N_291,N_1356);
and U3698 (N_3698,N_286,N_2554);
or U3699 (N_3699,N_1784,N_1483);
nor U3700 (N_3700,N_2101,N_1021);
nand U3701 (N_3701,N_419,N_1537);
and U3702 (N_3702,N_2580,N_802);
and U3703 (N_3703,N_2192,N_2342);
nand U3704 (N_3704,N_633,N_2278);
or U3705 (N_3705,N_2244,N_1788);
nor U3706 (N_3706,N_2855,N_2610);
nand U3707 (N_3707,N_223,N_1170);
and U3708 (N_3708,N_2265,N_587);
nand U3709 (N_3709,N_2142,N_589);
xnor U3710 (N_3710,N_1842,N_879);
xnor U3711 (N_3711,N_2190,N_1260);
nor U3712 (N_3712,N_1826,N_2121);
nor U3713 (N_3713,N_2705,N_2143);
and U3714 (N_3714,N_765,N_1209);
and U3715 (N_3715,N_246,N_1245);
or U3716 (N_3716,N_2640,N_2535);
xor U3717 (N_3717,N_1817,N_73);
xor U3718 (N_3718,N_2730,N_827);
and U3719 (N_3719,N_1213,N_2511);
nand U3720 (N_3720,N_2848,N_1720);
nand U3721 (N_3721,N_2348,N_2824);
nand U3722 (N_3722,N_958,N_988);
nand U3723 (N_3723,N_158,N_2579);
nand U3724 (N_3724,N_1634,N_1085);
nor U3725 (N_3725,N_1583,N_1632);
and U3726 (N_3726,N_1599,N_120);
or U3727 (N_3727,N_2413,N_1077);
nand U3728 (N_3728,N_1242,N_1572);
or U3729 (N_3729,N_2461,N_2297);
nand U3730 (N_3730,N_1921,N_1569);
nand U3731 (N_3731,N_2641,N_1624);
and U3732 (N_3732,N_1868,N_786);
and U3733 (N_3733,N_1136,N_181);
nor U3734 (N_3734,N_798,N_1746);
or U3735 (N_3735,N_1294,N_449);
or U3736 (N_3736,N_12,N_2553);
or U3737 (N_3737,N_1864,N_1798);
nor U3738 (N_3738,N_1303,N_1241);
nand U3739 (N_3739,N_2087,N_1118);
or U3740 (N_3740,N_207,N_586);
or U3741 (N_3741,N_1880,N_571);
nand U3742 (N_3742,N_654,N_2704);
and U3743 (N_3743,N_2157,N_2475);
nor U3744 (N_3744,N_175,N_1357);
nand U3745 (N_3745,N_72,N_1659);
and U3746 (N_3746,N_469,N_676);
or U3747 (N_3747,N_2870,N_2509);
nor U3748 (N_3748,N_1772,N_236);
nand U3749 (N_3749,N_570,N_2207);
nand U3750 (N_3750,N_1075,N_1273);
and U3751 (N_3751,N_1161,N_1549);
nor U3752 (N_3752,N_505,N_702);
nand U3753 (N_3753,N_250,N_2208);
nor U3754 (N_3754,N_1958,N_886);
and U3755 (N_3755,N_2666,N_177);
or U3756 (N_3756,N_2912,N_2131);
nor U3757 (N_3757,N_2027,N_878);
and U3758 (N_3758,N_1224,N_1415);
nand U3759 (N_3759,N_1223,N_1177);
nand U3760 (N_3760,N_1909,N_1850);
nor U3761 (N_3761,N_2410,N_1037);
nand U3762 (N_3762,N_1768,N_576);
xnor U3763 (N_3763,N_1407,N_1396);
or U3764 (N_3764,N_144,N_980);
nor U3765 (N_3765,N_2405,N_35);
and U3766 (N_3766,N_359,N_2181);
xor U3767 (N_3767,N_2126,N_2812);
xor U3768 (N_3768,N_206,N_1588);
nor U3769 (N_3769,N_2875,N_1401);
nor U3770 (N_3770,N_2555,N_2077);
and U3771 (N_3771,N_263,N_1665);
or U3772 (N_3772,N_2134,N_1576);
or U3773 (N_3773,N_447,N_1259);
nand U3774 (N_3774,N_1988,N_230);
nor U3775 (N_3775,N_1593,N_2826);
and U3776 (N_3776,N_261,N_2001);
and U3777 (N_3777,N_608,N_199);
xnor U3778 (N_3778,N_800,N_1044);
and U3779 (N_3779,N_899,N_2251);
nand U3780 (N_3780,N_658,N_1806);
or U3781 (N_3781,N_741,N_211);
and U3782 (N_3782,N_1339,N_1);
and U3783 (N_3783,N_1755,N_602);
and U3784 (N_3784,N_1562,N_2351);
and U3785 (N_3785,N_2528,N_969);
and U3786 (N_3786,N_2770,N_2218);
xnor U3787 (N_3787,N_531,N_290);
or U3788 (N_3788,N_1372,N_2296);
and U3789 (N_3789,N_2112,N_1020);
nor U3790 (N_3790,N_2223,N_161);
nand U3791 (N_3791,N_1022,N_2334);
nand U3792 (N_3792,N_2573,N_625);
nand U3793 (N_3793,N_2557,N_693);
or U3794 (N_3794,N_2668,N_1106);
nand U3795 (N_3795,N_1226,N_2291);
and U3796 (N_3796,N_868,N_876);
nor U3797 (N_3797,N_1236,N_1192);
or U3798 (N_3798,N_489,N_880);
or U3799 (N_3799,N_1492,N_1283);
or U3800 (N_3800,N_599,N_1423);
or U3801 (N_3801,N_155,N_254);
or U3802 (N_3802,N_806,N_1133);
nand U3803 (N_3803,N_2078,N_2724);
and U3804 (N_3804,N_45,N_2409);
or U3805 (N_3805,N_1538,N_2628);
nor U3806 (N_3806,N_2802,N_2856);
and U3807 (N_3807,N_149,N_2719);
and U3808 (N_3808,N_2257,N_1418);
nor U3809 (N_3809,N_1103,N_1460);
or U3810 (N_3810,N_2496,N_2465);
nor U3811 (N_3811,N_353,N_1145);
nor U3812 (N_3812,N_1232,N_2425);
and U3813 (N_3813,N_1319,N_1976);
and U3814 (N_3814,N_360,N_2684);
or U3815 (N_3815,N_2158,N_663);
nor U3816 (N_3816,N_3,N_2385);
nand U3817 (N_3817,N_2882,N_1056);
xor U3818 (N_3818,N_510,N_2003);
and U3819 (N_3819,N_1655,N_2026);
nor U3820 (N_3820,N_128,N_1212);
or U3821 (N_3821,N_2107,N_2426);
and U3822 (N_3822,N_2116,N_385);
and U3823 (N_3823,N_1641,N_2587);
nand U3824 (N_3824,N_1227,N_515);
nand U3825 (N_3825,N_1152,N_373);
nand U3826 (N_3826,N_49,N_2760);
xnor U3827 (N_3827,N_1980,N_43);
xnor U3828 (N_3828,N_458,N_1559);
or U3829 (N_3829,N_1902,N_2395);
or U3830 (N_3830,N_1393,N_596);
nor U3831 (N_3831,N_703,N_271);
or U3832 (N_3832,N_2273,N_318);
or U3833 (N_3833,N_2139,N_2650);
or U3834 (N_3834,N_2959,N_2012);
and U3835 (N_3835,N_444,N_2588);
nor U3836 (N_3836,N_1144,N_1520);
and U3837 (N_3837,N_1262,N_1353);
and U3838 (N_3838,N_2358,N_384);
or U3839 (N_3839,N_2102,N_2319);
or U3840 (N_3840,N_755,N_209);
and U3841 (N_3841,N_2471,N_1678);
nand U3842 (N_3842,N_815,N_1986);
nand U3843 (N_3843,N_503,N_581);
and U3844 (N_3844,N_1081,N_1767);
nor U3845 (N_3845,N_1896,N_848);
xnor U3846 (N_3846,N_529,N_1724);
and U3847 (N_3847,N_1057,N_2861);
nor U3848 (N_3848,N_2217,N_193);
or U3849 (N_3849,N_1321,N_1395);
nand U3850 (N_3850,N_541,N_54);
and U3851 (N_3851,N_724,N_2655);
and U3852 (N_3852,N_2683,N_1941);
xor U3853 (N_3853,N_1972,N_972);
nor U3854 (N_3854,N_1579,N_896);
nand U3855 (N_3855,N_770,N_1139);
xor U3856 (N_3856,N_1893,N_902);
xor U3857 (N_3857,N_1508,N_2712);
or U3858 (N_3858,N_138,N_2376);
xor U3859 (N_3859,N_1616,N_1693);
xor U3860 (N_3860,N_674,N_2779);
nand U3861 (N_3861,N_2799,N_1129);
and U3862 (N_3862,N_1099,N_781);
nand U3863 (N_3863,N_1820,N_2963);
xnor U3864 (N_3864,N_1371,N_1437);
xnor U3865 (N_3865,N_14,N_2860);
nor U3866 (N_3866,N_197,N_1642);
and U3867 (N_3867,N_2569,N_761);
nor U3868 (N_3868,N_1237,N_2790);
and U3869 (N_3869,N_2506,N_1540);
nand U3870 (N_3870,N_1800,N_2937);
nand U3871 (N_3871,N_2213,N_1270);
xor U3872 (N_3872,N_2627,N_1749);
and U3873 (N_3873,N_367,N_1829);
nor U3874 (N_3874,N_1333,N_1453);
xnor U3875 (N_3875,N_1851,N_81);
and U3876 (N_3876,N_302,N_946);
or U3877 (N_3877,N_611,N_2189);
nor U3878 (N_3878,N_1756,N_96);
or U3879 (N_3879,N_1598,N_173);
nor U3880 (N_3880,N_1210,N_1350);
or U3881 (N_3881,N_524,N_791);
nand U3882 (N_3882,N_2148,N_1887);
nand U3883 (N_3883,N_1541,N_824);
and U3884 (N_3884,N_311,N_76);
nand U3885 (N_3885,N_1830,N_446);
nor U3886 (N_3886,N_1789,N_1045);
xnor U3887 (N_3887,N_2039,N_2881);
xnor U3888 (N_3888,N_2896,N_363);
nor U3889 (N_3889,N_624,N_2043);
and U3890 (N_3890,N_1649,N_2594);
and U3891 (N_3891,N_1761,N_2839);
xor U3892 (N_3892,N_2232,N_1930);
and U3893 (N_3893,N_1631,N_2747);
nand U3894 (N_3894,N_497,N_1182);
nand U3895 (N_3895,N_1197,N_2117);
and U3896 (N_3896,N_1310,N_1300);
nor U3897 (N_3897,N_2403,N_760);
or U3898 (N_3898,N_2791,N_1597);
nand U3899 (N_3899,N_403,N_920);
nor U3900 (N_3900,N_2495,N_2125);
nor U3901 (N_3901,N_1231,N_1543);
nor U3902 (N_3902,N_2317,N_2541);
or U3903 (N_3903,N_2920,N_1495);
or U3904 (N_3904,N_1771,N_478);
or U3905 (N_3905,N_396,N_493);
or U3906 (N_3906,N_1066,N_2900);
and U3907 (N_3907,N_1695,N_1517);
or U3908 (N_3908,N_708,N_2305);
xor U3909 (N_3909,N_2620,N_1006);
or U3910 (N_3910,N_1105,N_139);
nor U3911 (N_3911,N_1963,N_1694);
xnor U3912 (N_3912,N_1944,N_545);
or U3913 (N_3913,N_330,N_1847);
and U3914 (N_3914,N_93,N_145);
xnor U3915 (N_3915,N_664,N_1281);
nand U3916 (N_3916,N_2570,N_1234);
and U3917 (N_3917,N_337,N_2105);
nor U3918 (N_3918,N_1943,N_2813);
nand U3919 (N_3919,N_2321,N_404);
nor U3920 (N_3920,N_561,N_162);
or U3921 (N_3921,N_590,N_99);
nand U3922 (N_3922,N_393,N_2601);
and U3923 (N_3923,N_2327,N_1711);
nand U3924 (N_3924,N_320,N_2360);
nand U3925 (N_3925,N_392,N_2505);
nor U3926 (N_3926,N_2992,N_9);
nand U3927 (N_3927,N_2145,N_1692);
or U3928 (N_3928,N_2998,N_188);
nor U3929 (N_3929,N_1832,N_1366);
or U3930 (N_3930,N_2984,N_575);
xor U3931 (N_3931,N_2392,N_184);
and U3932 (N_3932,N_1142,N_253);
or U3933 (N_3933,N_365,N_1833);
nand U3934 (N_3934,N_2662,N_2895);
nor U3935 (N_3935,N_1340,N_218);
or U3936 (N_3936,N_930,N_778);
or U3937 (N_3937,N_1977,N_1982);
nand U3938 (N_3938,N_1296,N_34);
nand U3939 (N_3939,N_238,N_22);
or U3940 (N_3940,N_1707,N_601);
or U3941 (N_3941,N_429,N_1065);
nor U3942 (N_3942,N_889,N_364);
xor U3943 (N_3943,N_2119,N_1328);
and U3944 (N_3944,N_2097,N_2271);
or U3945 (N_3945,N_1765,N_2970);
or U3946 (N_3946,N_1314,N_1522);
xor U3947 (N_3947,N_1937,N_338);
and U3948 (N_3948,N_1361,N_792);
xnor U3949 (N_3949,N_457,N_2380);
nor U3950 (N_3950,N_812,N_1527);
and U3951 (N_3951,N_1557,N_2367);
or U3952 (N_3952,N_2108,N_126);
xnor U3953 (N_3953,N_615,N_1739);
nor U3954 (N_3954,N_1676,N_2133);
nand U3955 (N_3955,N_2703,N_776);
nand U3956 (N_3956,N_822,N_1552);
nor U3957 (N_3957,N_1222,N_981);
nand U3958 (N_3958,N_883,N_1573);
and U3959 (N_3959,N_733,N_2227);
nand U3960 (N_3960,N_179,N_2195);
nor U3961 (N_3961,N_839,N_2277);
and U3962 (N_3962,N_2697,N_124);
or U3963 (N_3963,N_2381,N_413);
or U3964 (N_3964,N_1792,N_2954);
or U3965 (N_3965,N_1991,N_219);
or U3966 (N_3966,N_1810,N_1196);
nand U3967 (N_3967,N_180,N_1647);
nor U3968 (N_3968,N_2921,N_2329);
nand U3969 (N_3969,N_1011,N_2169);
nor U3970 (N_3970,N_1351,N_1207);
nor U3971 (N_3971,N_1449,N_1838);
or U3972 (N_3972,N_104,N_1230);
and U3973 (N_3973,N_2082,N_2372);
or U3974 (N_3974,N_1498,N_2283);
xor U3975 (N_3975,N_1521,N_2877);
xnor U3976 (N_3976,N_259,N_482);
or U3977 (N_3977,N_2203,N_2977);
or U3978 (N_3978,N_2123,N_2982);
and U3979 (N_3979,N_577,N_167);
nand U3980 (N_3980,N_2889,N_2335);
xor U3981 (N_3981,N_1164,N_2389);
nand U3982 (N_3982,N_1700,N_2996);
nand U3983 (N_3983,N_2079,N_1709);
and U3984 (N_3984,N_1000,N_1654);
nand U3985 (N_3985,N_1292,N_1019);
xor U3986 (N_3986,N_1999,N_999);
xor U3987 (N_3987,N_863,N_1985);
nor U3988 (N_3988,N_1677,N_2480);
nor U3989 (N_3989,N_2183,N_1718);
and U3990 (N_3990,N_346,N_2146);
nor U3991 (N_3991,N_2443,N_366);
or U3992 (N_3992,N_1959,N_828);
or U3993 (N_3993,N_1168,N_954);
nor U3994 (N_3994,N_1955,N_304);
or U3995 (N_3995,N_1135,N_407);
xor U3996 (N_3996,N_347,N_754);
or U3997 (N_3997,N_1740,N_1905);
nand U3998 (N_3998,N_1750,N_923);
nor U3999 (N_3999,N_1299,N_749);
xor U4000 (N_4000,N_191,N_694);
nand U4001 (N_4001,N_2780,N_1710);
nor U4002 (N_4002,N_881,N_295);
nand U4003 (N_4003,N_677,N_2170);
or U4004 (N_4004,N_443,N_1778);
and U4005 (N_4005,N_1358,N_2099);
xor U4006 (N_4006,N_2551,N_2883);
or U4007 (N_4007,N_2323,N_967);
nand U4008 (N_4008,N_2999,N_2144);
nor U4009 (N_4009,N_2398,N_150);
nand U4010 (N_4010,N_968,N_1059);
nand U4011 (N_4011,N_1302,N_566);
and U4012 (N_4012,N_2309,N_2801);
xnor U4013 (N_4013,N_657,N_1920);
nor U4014 (N_4014,N_1157,N_305);
nand U4015 (N_4015,N_455,N_2607);
nand U4016 (N_4016,N_1134,N_2552);
and U4017 (N_4017,N_991,N_1667);
nor U4018 (N_4018,N_1650,N_558);
xnor U4019 (N_4019,N_995,N_1807);
nor U4020 (N_4020,N_0,N_564);
xnor U4021 (N_4021,N_2753,N_1712);
or U4022 (N_4022,N_325,N_1381);
nor U4023 (N_4023,N_683,N_2820);
and U4024 (N_4024,N_1442,N_971);
or U4025 (N_4025,N_2995,N_2545);
or U4026 (N_4026,N_2891,N_321);
nand U4027 (N_4027,N_477,N_642);
nand U4028 (N_4028,N_2486,N_2173);
and U4029 (N_4029,N_2239,N_922);
or U4030 (N_4030,N_784,N_2652);
xor U4031 (N_4031,N_1706,N_2414);
nand U4032 (N_4032,N_2210,N_2016);
and U4033 (N_4033,N_1316,N_1368);
or U4034 (N_4034,N_1061,N_2269);
or U4035 (N_4035,N_1516,N_17);
and U4036 (N_4036,N_864,N_2090);
nor U4037 (N_4037,N_984,N_111);
nor U4038 (N_4038,N_1910,N_377);
or U4039 (N_4039,N_2153,N_1901);
xnor U4040 (N_4040,N_460,N_112);
nand U4041 (N_4041,N_2279,N_2231);
nor U4042 (N_4042,N_2596,N_1574);
nor U4043 (N_4043,N_481,N_1722);
and U4044 (N_4044,N_2673,N_1970);
nand U4045 (N_4045,N_2643,N_2798);
nor U4046 (N_4046,N_2985,N_1448);
or U4047 (N_4047,N_1014,N_2341);
nand U4048 (N_4048,N_2657,N_1373);
nand U4049 (N_4049,N_2314,N_620);
nand U4050 (N_4050,N_2054,N_2002);
nor U4051 (N_4051,N_301,N_2892);
nor U4052 (N_4052,N_1592,N_368);
or U4053 (N_4053,N_65,N_2745);
and U4054 (N_4054,N_2196,N_1803);
nand U4055 (N_4055,N_2485,N_2093);
xor U4056 (N_4056,N_840,N_2965);
nor U4057 (N_4057,N_2104,N_1612);
or U4058 (N_4058,N_661,N_2337);
nor U4059 (N_4059,N_1824,N_1455);
and U4060 (N_4060,N_2454,N_1533);
nand U4061 (N_4061,N_1629,N_2428);
or U4062 (N_4062,N_2052,N_1675);
nand U4063 (N_4063,N_2159,N_1249);
or U4064 (N_4064,N_1645,N_1633);
nor U4065 (N_4065,N_80,N_939);
and U4066 (N_4066,N_841,N_833);
nor U4067 (N_4067,N_2664,N_1041);
or U4068 (N_4068,N_2051,N_1088);
and U4069 (N_4069,N_352,N_645);
nand U4070 (N_4070,N_636,N_907);
nand U4071 (N_4071,N_1903,N_372);
nor U4072 (N_4072,N_2311,N_378);
nand U4073 (N_4073,N_2962,N_598);
or U4074 (N_4074,N_2420,N_98);
nand U4075 (N_4075,N_1526,N_1957);
nand U4076 (N_4076,N_2914,N_1536);
nor U4077 (N_4077,N_110,N_671);
nor U4078 (N_4078,N_2757,N_2293);
or U4079 (N_4079,N_1907,N_421);
and U4080 (N_4080,N_1162,N_2417);
and U4081 (N_4081,N_700,N_102);
and U4082 (N_4082,N_672,N_1638);
nor U4083 (N_4083,N_1403,N_1151);
nand U4084 (N_4084,N_1848,N_265);
nor U4085 (N_4085,N_160,N_1601);
or U4086 (N_4086,N_941,N_2355);
and U4087 (N_4087,N_2722,N_2743);
and U4088 (N_4088,N_2136,N_2185);
xor U4089 (N_4089,N_2796,N_2604);
xor U4090 (N_4090,N_935,N_905);
nor U4091 (N_4091,N_1334,N_2524);
and U4092 (N_4092,N_1827,N_2344);
nand U4093 (N_4093,N_709,N_1195);
nand U4094 (N_4094,N_1121,N_379);
nor U4095 (N_4095,N_2672,N_1697);
xnor U4096 (N_4096,N_315,N_1865);
and U4097 (N_4097,N_1735,N_721);
or U4098 (N_4098,N_1091,N_2457);
nand U4099 (N_4099,N_2481,N_1398);
nand U4100 (N_4100,N_1900,N_154);
and U4101 (N_4101,N_264,N_1696);
and U4102 (N_4102,N_1015,N_517);
nand U4103 (N_4103,N_540,N_2729);
and U4104 (N_4104,N_2191,N_707);
nand U4105 (N_4105,N_38,N_1409);
and U4106 (N_4106,N_2709,N_1714);
xor U4107 (N_4107,N_955,N_1320);
nor U4108 (N_4108,N_1936,N_1892);
nor U4109 (N_4109,N_1104,N_1169);
nand U4110 (N_4110,N_583,N_2548);
and U4111 (N_4111,N_1496,N_2081);
and U4112 (N_4112,N_993,N_560);
or U4113 (N_4113,N_1615,N_1801);
and U4114 (N_4114,N_2007,N_2362);
or U4115 (N_4115,N_2507,N_2699);
nor U4116 (N_4116,N_249,N_1389);
nor U4117 (N_4117,N_2873,N_1402);
or U4118 (N_4118,N_2701,N_2762);
or U4119 (N_4119,N_1450,N_2175);
or U4120 (N_4120,N_53,N_2904);
or U4121 (N_4121,N_2234,N_448);
nand U4122 (N_4122,N_1652,N_974);
nor U4123 (N_4123,N_1417,N_361);
nand U4124 (N_4124,N_1317,N_2179);
or U4125 (N_4125,N_1648,N_648);
or U4126 (N_4126,N_753,N_2833);
xor U4127 (N_4127,N_921,N_2338);
or U4128 (N_4128,N_1916,N_1509);
and U4129 (N_4129,N_2292,N_959);
nor U4130 (N_4130,N_1565,N_1595);
nor U4131 (N_4131,N_1535,N_2927);
or U4132 (N_4132,N_1688,N_23);
and U4133 (N_4133,N_2586,N_1446);
or U4134 (N_4134,N_299,N_2035);
and U4135 (N_4135,N_1486,N_1191);
or U4136 (N_4136,N_2648,N_2187);
or U4137 (N_4137,N_1376,N_2728);
nor U4138 (N_4138,N_789,N_2955);
nor U4139 (N_4139,N_1282,N_1558);
nor U4140 (N_4140,N_727,N_1093);
and U4141 (N_4141,N_2019,N_2597);
or U4142 (N_4142,N_772,N_1094);
or U4143 (N_4143,N_168,N_2844);
xor U4144 (N_4144,N_743,N_1699);
nand U4145 (N_4145,N_2783,N_1238);
nor U4146 (N_4146,N_2827,N_341);
nor U4147 (N_4147,N_977,N_1762);
and U4148 (N_4148,N_427,N_486);
xnor U4149 (N_4149,N_1764,N_2755);
nor U4150 (N_4150,N_2034,N_109);
nor U4151 (N_4151,N_1523,N_1122);
nand U4152 (N_4152,N_686,N_1951);
and U4153 (N_4153,N_1344,N_140);
nor U4154 (N_4154,N_532,N_408);
xnor U4155 (N_4155,N_282,N_1751);
nor U4156 (N_4156,N_2229,N_2431);
or U4157 (N_4157,N_916,N_1130);
nand U4158 (N_4158,N_1067,N_1154);
or U4159 (N_4159,N_1664,N_1969);
xor U4160 (N_4160,N_2842,N_961);
nand U4161 (N_4161,N_603,N_1561);
nor U4162 (N_4162,N_1774,N_825);
nor U4163 (N_4163,N_319,N_1682);
nor U4164 (N_4164,N_1240,N_2972);
nor U4165 (N_4165,N_296,N_1753);
or U4166 (N_4166,N_2711,N_2713);
and U4167 (N_4167,N_2365,N_2450);
xnor U4168 (N_4168,N_32,N_2930);
nand U4169 (N_4169,N_1413,N_2876);
and U4170 (N_4170,N_2901,N_1596);
nor U4171 (N_4171,N_256,N_855);
and U4172 (N_4172,N_867,N_10);
or U4173 (N_4173,N_1287,N_1518);
nand U4174 (N_4174,N_1783,N_1790);
and U4175 (N_4175,N_2415,N_2543);
nand U4176 (N_4176,N_1149,N_18);
xor U4177 (N_4177,N_153,N_1359);
xnor U4178 (N_4178,N_405,N_717);
or U4179 (N_4179,N_2584,N_747);
or U4180 (N_4180,N_2886,N_1163);
and U4181 (N_4181,N_2064,N_1702);
xnor U4182 (N_4182,N_1017,N_1100);
or U4183 (N_4183,N_351,N_2983);
and U4184 (N_4184,N_69,N_2474);
nor U4185 (N_4185,N_2613,N_1433);
or U4186 (N_4186,N_1912,N_28);
and U4187 (N_4187,N_2464,N_814);
nand U4188 (N_4188,N_2774,N_340);
and U4189 (N_4189,N_2661,N_1128);
and U4190 (N_4190,N_859,N_135);
nor U4191 (N_4191,N_689,N_1482);
nand U4192 (N_4192,N_1284,N_895);
or U4193 (N_4193,N_2390,N_1374);
or U4194 (N_4194,N_306,N_1856);
or U4195 (N_4195,N_1117,N_200);
and U4196 (N_4196,N_2732,N_2837);
and U4197 (N_4197,N_655,N_1330);
nand U4198 (N_4198,N_1708,N_1194);
nor U4199 (N_4199,N_2370,N_216);
or U4200 (N_4200,N_2154,N_2974);
or U4201 (N_4201,N_1619,N_2353);
and U4202 (N_4202,N_1519,N_1009);
nand U4203 (N_4203,N_2863,N_2452);
nand U4204 (N_4204,N_805,N_829);
or U4205 (N_4205,N_1658,N_2908);
nor U4206 (N_4206,N_1246,N_2448);
and U4207 (N_4207,N_196,N_2635);
nand U4208 (N_4208,N_2483,N_431);
xor U4209 (N_4209,N_1663,N_2623);
or U4210 (N_4210,N_2966,N_317);
nor U4211 (N_4211,N_1614,N_1200);
or U4212 (N_4212,N_555,N_78);
nand U4213 (N_4213,N_2375,N_2859);
and U4214 (N_4214,N_1513,N_1272);
nand U4215 (N_4215,N_83,N_1949);
and U4216 (N_4216,N_1534,N_2488);
nor U4217 (N_4217,N_1973,N_1008);
nor U4218 (N_4218,N_374,N_142);
or U4219 (N_4219,N_1097,N_1392);
nand U4220 (N_4220,N_2879,N_2702);
nor U4221 (N_4221,N_2514,N_2053);
nor U4222 (N_4222,N_2915,N_2394);
and U4223 (N_4223,N_2558,N_616);
or U4224 (N_4224,N_699,N_1175);
nor U4225 (N_4225,N_1468,N_1837);
and U4226 (N_4226,N_2447,N_1479);
nand U4227 (N_4227,N_2423,N_1546);
or U4228 (N_4228,N_2598,N_1420);
xor U4229 (N_4229,N_2515,N_2685);
nand U4230 (N_4230,N_2576,N_910);
nor U4231 (N_4231,N_501,N_2532);
nand U4232 (N_4232,N_600,N_2828);
xnor U4233 (N_4233,N_2605,N_1716);
or U4234 (N_4234,N_1153,N_911);
nand U4235 (N_4235,N_1725,N_488);
and U4236 (N_4236,N_1480,N_1146);
or U4237 (N_4237,N_2267,N_835);
or U4238 (N_4238,N_719,N_213);
or U4239 (N_4239,N_2202,N_2721);
and U4240 (N_4240,N_2878,N_794);
nor U4241 (N_4241,N_534,N_2674);
and U4242 (N_4242,N_1217,N_552);
xor U4243 (N_4243,N_2073,N_903);
nor U4244 (N_4244,N_1254,N_536);
and U4245 (N_4245,N_2706,N_641);
and U4246 (N_4246,N_1802,N_530);
and U4247 (N_4247,N_1082,N_2854);
nand U4248 (N_4248,N_436,N_1607);
nor U4249 (N_4249,N_1315,N_2599);
and U4250 (N_4250,N_1174,N_1825);
nand U4251 (N_4251,N_39,N_2339);
or U4252 (N_4252,N_1954,N_1685);
and U4253 (N_4253,N_2764,N_2487);
nand U4254 (N_4254,N_1621,N_2006);
or U4255 (N_4255,N_255,N_638);
and U4256 (N_4256,N_966,N_1637);
nand U4257 (N_4257,N_2222,N_2617);
or U4258 (N_4258,N_2612,N_395);
nor U4259 (N_4259,N_2736,N_118);
or U4260 (N_4260,N_1929,N_680);
xor U4261 (N_4261,N_490,N_2451);
or U4262 (N_4262,N_1884,N_622);
and U4263 (N_4263,N_720,N_2518);
nor U4264 (N_4264,N_1804,N_133);
nor U4265 (N_4265,N_26,N_2304);
or U4266 (N_4266,N_272,N_865);
nand U4267 (N_4267,N_1886,N_237);
and U4268 (N_4268,N_1635,N_1524);
nor U4269 (N_4269,N_462,N_2316);
xnor U4270 (N_4270,N_2845,N_2638);
or U4271 (N_4271,N_1188,N_1090);
and U4272 (N_4272,N_2009,N_1379);
xnor U4273 (N_4273,N_2734,N_1627);
xor U4274 (N_4274,N_831,N_891);
nand U4275 (N_4275,N_471,N_1279);
and U4276 (N_4276,N_2872,N_1497);
nand U4277 (N_4277,N_1875,N_2387);
or U4278 (N_4278,N_190,N_2715);
nor U4279 (N_4279,N_2350,N_1435);
xor U4280 (N_4280,N_1594,N_375);
nand U4281 (N_4281,N_2698,N_468);
and U4282 (N_4282,N_2020,N_2120);
nor U4283 (N_4283,N_60,N_269);
nand U4284 (N_4284,N_496,N_2313);
nand U4285 (N_4285,N_2497,N_650);
nor U4286 (N_4286,N_1578,N_2013);
and U4287 (N_4287,N_2463,N_1503);
and U4288 (N_4288,N_2691,N_1644);
nand U4289 (N_4289,N_1878,N_2608);
and U4290 (N_4290,N_2926,N_2168);
and U4291 (N_4291,N_1165,N_234);
nand U4292 (N_4292,N_2264,N_774);
and U4293 (N_4293,N_1689,N_853);
nand U4294 (N_4294,N_1979,N_1250);
nand U4295 (N_4295,N_1462,N_669);
nand U4296 (N_4296,N_225,N_914);
or U4297 (N_4297,N_2220,N_2130);
or U4298 (N_4298,N_1553,N_1438);
nand U4299 (N_4299,N_2152,N_553);
nand U4300 (N_4300,N_2243,N_759);
nand U4301 (N_4301,N_1187,N_1770);
nor U4302 (N_4302,N_762,N_2280);
and U4303 (N_4303,N_1948,N_795);
xor U4304 (N_4304,N_289,N_2516);
and U4305 (N_4305,N_989,N_728);
xnor U4306 (N_4306,N_426,N_1956);
and U4307 (N_4307,N_1961,N_1444);
or U4308 (N_4308,N_2258,N_467);
xor U4309 (N_4309,N_673,N_1646);
xor U4310 (N_4310,N_215,N_2059);
or U4311 (N_4311,N_2138,N_2266);
nor U4312 (N_4312,N_2083,N_790);
nor U4313 (N_4313,N_2686,N_2825);
nor U4314 (N_4314,N_631,N_371);
and U4315 (N_4315,N_2174,N_2868);
nand U4316 (N_4316,N_394,N_1748);
nor U4317 (N_4317,N_2361,N_2871);
nor U4318 (N_4318,N_1812,N_885);
or U4319 (N_4319,N_2378,N_284);
nand U4320 (N_4320,N_2383,N_241);
nor U4321 (N_4321,N_681,N_1548);
and U4322 (N_4322,N_767,N_2268);
nand U4323 (N_4323,N_730,N_1610);
or U4324 (N_4324,N_1193,N_1684);
xor U4325 (N_4325,N_29,N_567);
and U4326 (N_4326,N_1235,N_195);
or U4327 (N_4327,N_2402,N_1671);
nand U4328 (N_4328,N_1734,N_358);
xor U4329 (N_4329,N_143,N_949);
or U4330 (N_4330,N_327,N_983);
nor U4331 (N_4331,N_2679,N_2888);
nor U4332 (N_4332,N_1834,N_1173);
xnor U4333 (N_4333,N_2419,N_2287);
nand U4334 (N_4334,N_166,N_2754);
and U4335 (N_4335,N_2642,N_334);
nand U4336 (N_4336,N_2957,N_2665);
nor U4337 (N_4337,N_2794,N_1775);
nand U4338 (N_4338,N_58,N_1010);
and U4339 (N_4339,N_61,N_2113);
xor U4340 (N_4340,N_1998,N_2924);
nor U4341 (N_4341,N_2166,N_203);
xnor U4342 (N_4342,N_890,N_68);
nand U4343 (N_4343,N_2976,N_580);
nor U4344 (N_4344,N_823,N_1939);
xor U4345 (N_4345,N_1643,N_934);
nor U4346 (N_4346,N_639,N_1092);
or U4347 (N_4347,N_1434,N_1965);
and U4348 (N_4348,N_1758,N_1997);
nand U4349 (N_4349,N_2631,N_2681);
xor U4350 (N_4350,N_1602,N_2343);
and U4351 (N_4351,N_894,N_857);
and U4352 (N_4352,N_2636,N_562);
nor U4353 (N_4353,N_260,N_453);
nand U4354 (N_4354,N_1890,N_1852);
nand U4355 (N_4355,N_742,N_2364);
and U4356 (N_4356,N_183,N_91);
xnor U4357 (N_4357,N_2775,N_423);
nor U4358 (N_4358,N_2404,N_928);
or U4359 (N_4359,N_307,N_214);
nor U4360 (N_4360,N_2237,N_637);
or U4361 (N_4361,N_1726,N_542);
and U4362 (N_4362,N_2645,N_574);
nand U4363 (N_4363,N_2340,N_2076);
or U4364 (N_4364,N_1487,N_46);
or U4365 (N_4365,N_2302,N_464);
nand U4366 (N_4366,N_2693,N_2384);
and U4367 (N_4367,N_710,N_2252);
nor U4368 (N_4368,N_1386,N_71);
or U4369 (N_4369,N_527,N_1577);
and U4370 (N_4370,N_114,N_1918);
and U4371 (N_4371,N_901,N_2017);
and U4372 (N_4372,N_2731,N_523);
xnor U4373 (N_4373,N_2458,N_660);
and U4374 (N_4374,N_2308,N_2529);
nand U4375 (N_4375,N_1312,N_2938);
or U4376 (N_4376,N_2439,N_186);
nor U4377 (N_4377,N_610,N_1613);
or U4378 (N_4378,N_1993,N_2198);
or U4379 (N_4379,N_926,N_1004);
nand U4380 (N_4380,N_2550,N_2831);
nand U4381 (N_4381,N_2942,N_275);
and U4382 (N_4382,N_1611,N_1080);
or U4383 (N_4383,N_942,N_92);
and U4384 (N_4384,N_858,N_1781);
and U4385 (N_4385,N_682,N_2128);
xnor U4386 (N_4386,N_2519,N_2299);
and U4387 (N_4387,N_2036,N_994);
nor U4388 (N_4388,N_1399,N_2261);
nand U4389 (N_4389,N_563,N_2789);
nor U4390 (N_4390,N_675,N_764);
nor U4391 (N_4391,N_1840,N_267);
and U4392 (N_4392,N_442,N_945);
xnor U4393 (N_4393,N_1721,N_2800);
or U4394 (N_4394,N_568,N_2276);
nand U4395 (N_4395,N_2622,N_1681);
and U4396 (N_4396,N_605,N_2771);
xor U4397 (N_4397,N_1380,N_811);
and U4398 (N_4398,N_283,N_2240);
nand U4399 (N_4399,N_2290,N_1176);
or U4400 (N_4400,N_125,N_1394);
and U4401 (N_4401,N_2436,N_106);
or U4402 (N_4402,N_1913,N_2253);
or U4403 (N_4403,N_127,N_281);
or U4404 (N_4404,N_1211,N_2517);
nand U4405 (N_4405,N_1119,N_1071);
or U4406 (N_4406,N_2479,N_2907);
and U4407 (N_4407,N_1012,N_348);
nand U4408 (N_4408,N_698,N_1141);
nand U4409 (N_4409,N_1329,N_2864);
or U4410 (N_4410,N_40,N_766);
nor U4411 (N_4411,N_649,N_2568);
nor U4412 (N_4412,N_2472,N_2624);
or U4413 (N_4413,N_2259,N_628);
nor U4414 (N_4414,N_2250,N_2639);
xor U4415 (N_4415,N_95,N_1994);
or U4416 (N_4416,N_182,N_1034);
or U4417 (N_4417,N_2462,N_716);
and U4418 (N_4418,N_725,N_511);
or U4419 (N_4419,N_871,N_87);
or U4420 (N_4420,N_1773,N_2797);
xnor U4421 (N_4421,N_1158,N_714);
nor U4422 (N_4422,N_2811,N_2041);
and U4423 (N_4423,N_2852,N_1378);
nand U4424 (N_4424,N_1063,N_2046);
and U4425 (N_4425,N_245,N_2727);
nor U4426 (N_4426,N_627,N_2432);
nor U4427 (N_4427,N_1440,N_1640);
nand U4428 (N_4428,N_1301,N_1289);
nor U4429 (N_4429,N_171,N_1473);
nand U4430 (N_4430,N_2508,N_2897);
nand U4431 (N_4431,N_1084,N_205);
nand U4432 (N_4432,N_434,N_233);
or U4433 (N_4433,N_2536,N_751);
nand U4434 (N_4434,N_2286,N_2906);
nor U4435 (N_4435,N_2346,N_2807);
nand U4436 (N_4436,N_1745,N_1687);
nor U4437 (N_4437,N_2045,N_729);
and U4438 (N_4438,N_691,N_409);
nor U4439 (N_4439,N_185,N_1069);
nor U4440 (N_4440,N_931,N_1669);
nand U4441 (N_4441,N_1882,N_1662);
or U4442 (N_4442,N_1382,N_85);
nand U4443 (N_4443,N_2564,N_2401);
nor U4444 (N_4444,N_1532,N_1026);
nand U4445 (N_4445,N_2282,N_569);
or U4446 (N_4446,N_1787,N_1247);
nor U4447 (N_4447,N_400,N_212);
nor U4448 (N_4448,N_1570,N_1871);
nor U4449 (N_4449,N_2958,N_769);
or U4450 (N_4450,N_2228,N_2074);
xor U4451 (N_4451,N_1048,N_2274);
and U4452 (N_4452,N_973,N_1349);
and U4453 (N_4453,N_77,N_6);
or U4454 (N_4454,N_2197,N_285);
or U4455 (N_4455,N_646,N_1228);
and U4456 (N_4456,N_2366,N_2917);
nor U4457 (N_4457,N_2542,N_1159);
nand U4458 (N_4458,N_1038,N_2391);
and U4459 (N_4459,N_2502,N_2769);
nand U4460 (N_4460,N_685,N_634);
nand U4461 (N_4461,N_1377,N_965);
or U4462 (N_4462,N_854,N_1363);
nor U4463 (N_4463,N_535,N_1406);
or U4464 (N_4464,N_1343,N_292);
or U4465 (N_4465,N_2242,N_331);
nand U4466 (N_4466,N_1776,N_387);
and U4467 (N_4467,N_293,N_2085);
nand U4468 (N_4468,N_1760,N_1933);
nor U4469 (N_4469,N_2109,N_1365);
nand U4470 (N_4470,N_796,N_1818);
xnor U4471 (N_4471,N_2944,N_2270);
and U4472 (N_4472,N_251,N_70);
or U4473 (N_4473,N_782,N_1318);
nor U4474 (N_4474,N_1354,N_2005);
and U4475 (N_4475,N_323,N_1079);
and U4476 (N_4476,N_2583,N_2156);
or U4477 (N_4477,N_2880,N_1811);
nor U4478 (N_4478,N_2015,N_1680);
xnor U4479 (N_4479,N_1124,N_1560);
nand U4480 (N_4480,N_1766,N_1400);
nand U4481 (N_4481,N_242,N_509);
or U4482 (N_4482,N_2070,N_89);
and U4483 (N_4483,N_2971,N_406);
or U4484 (N_4484,N_79,N_2948);
or U4485 (N_4485,N_2935,N_2708);
nor U4486 (N_4486,N_2345,N_1095);
or U4487 (N_4487,N_1952,N_862);
and U4488 (N_4488,N_1036,N_630);
and U4489 (N_4489,N_1436,N_1111);
nand U4490 (N_4490,N_2122,N_2067);
nor U4491 (N_4491,N_2455,N_1422);
nand U4492 (N_4492,N_2500,N_2140);
nand U4493 (N_4493,N_2434,N_2670);
or U4494 (N_4494,N_2549,N_1860);
or U4495 (N_4495,N_2527,N_1717);
nor U4496 (N_4496,N_2818,N_2792);
or U4497 (N_4497,N_121,N_2312);
nand U4498 (N_4498,N_2646,N_1275);
nor U4499 (N_4499,N_2467,N_1439);
nor U4500 (N_4500,N_1953,N_1253);
nand U4501 (N_4501,N_1419,N_2808);
nand U4502 (N_4502,N_1090,N_2378);
or U4503 (N_4503,N_92,N_2014);
and U4504 (N_4504,N_334,N_176);
or U4505 (N_4505,N_2279,N_1143);
or U4506 (N_4506,N_323,N_304);
xnor U4507 (N_4507,N_2156,N_1382);
nor U4508 (N_4508,N_2534,N_1695);
and U4509 (N_4509,N_485,N_2986);
nor U4510 (N_4510,N_164,N_2500);
xnor U4511 (N_4511,N_999,N_1133);
nand U4512 (N_4512,N_115,N_2271);
nor U4513 (N_4513,N_1935,N_2803);
or U4514 (N_4514,N_257,N_2562);
and U4515 (N_4515,N_330,N_2640);
nor U4516 (N_4516,N_977,N_874);
nand U4517 (N_4517,N_917,N_1498);
and U4518 (N_4518,N_949,N_1347);
xnor U4519 (N_4519,N_238,N_2828);
and U4520 (N_4520,N_99,N_2461);
nor U4521 (N_4521,N_1977,N_1468);
and U4522 (N_4522,N_2379,N_1754);
nor U4523 (N_4523,N_1745,N_589);
nor U4524 (N_4524,N_2125,N_2801);
nand U4525 (N_4525,N_181,N_2844);
xor U4526 (N_4526,N_1295,N_773);
or U4527 (N_4527,N_1901,N_838);
and U4528 (N_4528,N_465,N_1697);
xnor U4529 (N_4529,N_2465,N_2396);
and U4530 (N_4530,N_585,N_1169);
nand U4531 (N_4531,N_393,N_2806);
nor U4532 (N_4532,N_529,N_354);
or U4533 (N_4533,N_588,N_1310);
nand U4534 (N_4534,N_2544,N_405);
nand U4535 (N_4535,N_125,N_2078);
nor U4536 (N_4536,N_2153,N_1741);
and U4537 (N_4537,N_1507,N_1549);
nor U4538 (N_4538,N_156,N_2252);
or U4539 (N_4539,N_1666,N_144);
and U4540 (N_4540,N_794,N_1042);
nand U4541 (N_4541,N_2011,N_2645);
or U4542 (N_4542,N_453,N_1307);
or U4543 (N_4543,N_2551,N_1677);
and U4544 (N_4544,N_2595,N_2031);
nand U4545 (N_4545,N_1356,N_1848);
and U4546 (N_4546,N_2028,N_732);
nor U4547 (N_4547,N_1612,N_1173);
xor U4548 (N_4548,N_944,N_461);
or U4549 (N_4549,N_558,N_2997);
nor U4550 (N_4550,N_1164,N_869);
or U4551 (N_4551,N_162,N_1552);
nor U4552 (N_4552,N_437,N_128);
nor U4553 (N_4553,N_1182,N_605);
nor U4554 (N_4554,N_1838,N_2067);
nor U4555 (N_4555,N_193,N_1637);
xnor U4556 (N_4556,N_1474,N_2715);
nand U4557 (N_4557,N_912,N_1606);
nand U4558 (N_4558,N_2712,N_1093);
and U4559 (N_4559,N_2142,N_1005);
nand U4560 (N_4560,N_2509,N_2614);
nand U4561 (N_4561,N_1036,N_2211);
xor U4562 (N_4562,N_484,N_215);
nor U4563 (N_4563,N_1868,N_1683);
or U4564 (N_4564,N_1621,N_784);
and U4565 (N_4565,N_2533,N_1817);
nand U4566 (N_4566,N_545,N_76);
nand U4567 (N_4567,N_1504,N_863);
nand U4568 (N_4568,N_2914,N_2699);
nor U4569 (N_4569,N_1223,N_1476);
nand U4570 (N_4570,N_1432,N_2523);
nor U4571 (N_4571,N_1627,N_1359);
nor U4572 (N_4572,N_2940,N_717);
nand U4573 (N_4573,N_2727,N_2635);
or U4574 (N_4574,N_1941,N_2771);
nor U4575 (N_4575,N_1414,N_1010);
or U4576 (N_4576,N_1973,N_2759);
or U4577 (N_4577,N_704,N_1659);
or U4578 (N_4578,N_310,N_90);
nand U4579 (N_4579,N_2063,N_321);
nor U4580 (N_4580,N_978,N_2244);
xnor U4581 (N_4581,N_207,N_1512);
xor U4582 (N_4582,N_1666,N_2827);
nand U4583 (N_4583,N_1355,N_188);
nor U4584 (N_4584,N_917,N_2253);
and U4585 (N_4585,N_1010,N_2751);
or U4586 (N_4586,N_405,N_783);
nor U4587 (N_4587,N_2153,N_1180);
nand U4588 (N_4588,N_2162,N_2725);
xnor U4589 (N_4589,N_2874,N_2686);
nor U4590 (N_4590,N_418,N_2110);
nand U4591 (N_4591,N_2382,N_53);
nand U4592 (N_4592,N_2864,N_454);
or U4593 (N_4593,N_2085,N_2771);
xnor U4594 (N_4594,N_802,N_1405);
xnor U4595 (N_4595,N_2861,N_1718);
or U4596 (N_4596,N_1451,N_36);
nand U4597 (N_4597,N_976,N_622);
or U4598 (N_4598,N_1284,N_329);
nor U4599 (N_4599,N_2254,N_756);
and U4600 (N_4600,N_2841,N_530);
and U4601 (N_4601,N_2213,N_1227);
xor U4602 (N_4602,N_790,N_1175);
and U4603 (N_4603,N_838,N_1017);
nand U4604 (N_4604,N_2683,N_2092);
nor U4605 (N_4605,N_2707,N_726);
xnor U4606 (N_4606,N_2160,N_2887);
xor U4607 (N_4607,N_529,N_2972);
nor U4608 (N_4608,N_829,N_806);
nor U4609 (N_4609,N_2240,N_1798);
and U4610 (N_4610,N_137,N_2788);
nand U4611 (N_4611,N_1807,N_2973);
or U4612 (N_4612,N_1550,N_115);
nand U4613 (N_4613,N_51,N_2452);
nand U4614 (N_4614,N_1626,N_1730);
nor U4615 (N_4615,N_192,N_1773);
nand U4616 (N_4616,N_2994,N_892);
nand U4617 (N_4617,N_646,N_2087);
nand U4618 (N_4618,N_176,N_1127);
nand U4619 (N_4619,N_1099,N_2143);
xnor U4620 (N_4620,N_1400,N_950);
or U4621 (N_4621,N_362,N_2014);
nand U4622 (N_4622,N_586,N_170);
nor U4623 (N_4623,N_1405,N_1126);
and U4624 (N_4624,N_791,N_1585);
nor U4625 (N_4625,N_1420,N_893);
nand U4626 (N_4626,N_1178,N_738);
or U4627 (N_4627,N_1864,N_2492);
or U4628 (N_4628,N_2521,N_2693);
nand U4629 (N_4629,N_640,N_2053);
nor U4630 (N_4630,N_1548,N_1352);
nand U4631 (N_4631,N_57,N_2038);
and U4632 (N_4632,N_442,N_1277);
and U4633 (N_4633,N_385,N_1669);
nand U4634 (N_4634,N_234,N_2819);
or U4635 (N_4635,N_186,N_2789);
nand U4636 (N_4636,N_1632,N_1823);
nand U4637 (N_4637,N_1761,N_382);
or U4638 (N_4638,N_2920,N_1167);
nor U4639 (N_4639,N_1127,N_2356);
nand U4640 (N_4640,N_849,N_1804);
nand U4641 (N_4641,N_1546,N_259);
or U4642 (N_4642,N_2110,N_618);
nand U4643 (N_4643,N_2252,N_2213);
or U4644 (N_4644,N_1276,N_21);
and U4645 (N_4645,N_2584,N_1728);
xor U4646 (N_4646,N_1805,N_325);
or U4647 (N_4647,N_2109,N_675);
nand U4648 (N_4648,N_2466,N_118);
xnor U4649 (N_4649,N_851,N_2329);
nand U4650 (N_4650,N_875,N_1383);
nor U4651 (N_4651,N_2231,N_1300);
nor U4652 (N_4652,N_2136,N_1318);
or U4653 (N_4653,N_1970,N_605);
and U4654 (N_4654,N_1627,N_2889);
and U4655 (N_4655,N_1847,N_2141);
xnor U4656 (N_4656,N_2246,N_2162);
nand U4657 (N_4657,N_2485,N_2642);
or U4658 (N_4658,N_1512,N_487);
nor U4659 (N_4659,N_876,N_1749);
nor U4660 (N_4660,N_1030,N_182);
and U4661 (N_4661,N_1262,N_628);
nand U4662 (N_4662,N_573,N_2816);
or U4663 (N_4663,N_2082,N_1508);
or U4664 (N_4664,N_2969,N_62);
nor U4665 (N_4665,N_2344,N_121);
xnor U4666 (N_4666,N_482,N_983);
nand U4667 (N_4667,N_673,N_353);
xor U4668 (N_4668,N_1222,N_377);
nand U4669 (N_4669,N_1194,N_307);
or U4670 (N_4670,N_1113,N_17);
nand U4671 (N_4671,N_232,N_2717);
and U4672 (N_4672,N_545,N_1975);
or U4673 (N_4673,N_1485,N_1101);
or U4674 (N_4674,N_2497,N_396);
nand U4675 (N_4675,N_828,N_1253);
and U4676 (N_4676,N_1494,N_843);
xor U4677 (N_4677,N_625,N_568);
nand U4678 (N_4678,N_802,N_1384);
nor U4679 (N_4679,N_2015,N_103);
nand U4680 (N_4680,N_1757,N_1686);
and U4681 (N_4681,N_8,N_693);
nand U4682 (N_4682,N_765,N_595);
nand U4683 (N_4683,N_2280,N_1290);
nand U4684 (N_4684,N_2373,N_1231);
nor U4685 (N_4685,N_248,N_229);
xnor U4686 (N_4686,N_2225,N_2845);
nor U4687 (N_4687,N_1235,N_1155);
or U4688 (N_4688,N_2331,N_1253);
or U4689 (N_4689,N_697,N_655);
or U4690 (N_4690,N_1008,N_2606);
or U4691 (N_4691,N_1459,N_1557);
nor U4692 (N_4692,N_1947,N_1712);
and U4693 (N_4693,N_1326,N_2466);
or U4694 (N_4694,N_2501,N_1034);
nand U4695 (N_4695,N_742,N_1879);
nor U4696 (N_4696,N_1163,N_340);
nand U4697 (N_4697,N_1820,N_2092);
nor U4698 (N_4698,N_1271,N_1189);
and U4699 (N_4699,N_1463,N_366);
nor U4700 (N_4700,N_785,N_1049);
nor U4701 (N_4701,N_2847,N_630);
and U4702 (N_4702,N_158,N_630);
and U4703 (N_4703,N_1582,N_2194);
nor U4704 (N_4704,N_2843,N_655);
and U4705 (N_4705,N_2533,N_992);
or U4706 (N_4706,N_629,N_1580);
nor U4707 (N_4707,N_1127,N_32);
nor U4708 (N_4708,N_2250,N_455);
nand U4709 (N_4709,N_2066,N_976);
nor U4710 (N_4710,N_392,N_2245);
nand U4711 (N_4711,N_1065,N_2260);
or U4712 (N_4712,N_1654,N_881);
and U4713 (N_4713,N_1299,N_1641);
and U4714 (N_4714,N_336,N_2670);
and U4715 (N_4715,N_1523,N_1873);
or U4716 (N_4716,N_958,N_1257);
xnor U4717 (N_4717,N_167,N_1381);
nor U4718 (N_4718,N_852,N_470);
and U4719 (N_4719,N_1018,N_2296);
nor U4720 (N_4720,N_1176,N_825);
or U4721 (N_4721,N_2547,N_1654);
nor U4722 (N_4722,N_1130,N_1184);
nand U4723 (N_4723,N_1079,N_1305);
xor U4724 (N_4724,N_683,N_464);
nor U4725 (N_4725,N_130,N_960);
or U4726 (N_4726,N_2596,N_2407);
or U4727 (N_4727,N_1962,N_2071);
and U4728 (N_4728,N_2653,N_723);
or U4729 (N_4729,N_231,N_469);
and U4730 (N_4730,N_628,N_2996);
and U4731 (N_4731,N_890,N_2447);
nand U4732 (N_4732,N_203,N_626);
or U4733 (N_4733,N_2222,N_1636);
and U4734 (N_4734,N_1985,N_172);
nor U4735 (N_4735,N_596,N_2734);
nand U4736 (N_4736,N_700,N_247);
nand U4737 (N_4737,N_1349,N_1975);
nand U4738 (N_4738,N_1662,N_1566);
nand U4739 (N_4739,N_742,N_71);
nor U4740 (N_4740,N_435,N_808);
nor U4741 (N_4741,N_1261,N_2074);
nor U4742 (N_4742,N_2559,N_648);
and U4743 (N_4743,N_1533,N_2893);
or U4744 (N_4744,N_387,N_1914);
xnor U4745 (N_4745,N_2910,N_60);
nor U4746 (N_4746,N_1859,N_282);
or U4747 (N_4747,N_2440,N_218);
or U4748 (N_4748,N_2454,N_2221);
and U4749 (N_4749,N_823,N_1818);
or U4750 (N_4750,N_1234,N_2410);
or U4751 (N_4751,N_407,N_2307);
nor U4752 (N_4752,N_1634,N_1314);
nor U4753 (N_4753,N_900,N_2284);
nor U4754 (N_4754,N_978,N_2048);
nand U4755 (N_4755,N_2536,N_581);
or U4756 (N_4756,N_243,N_720);
or U4757 (N_4757,N_1264,N_2093);
or U4758 (N_4758,N_1533,N_2084);
and U4759 (N_4759,N_2547,N_1628);
nor U4760 (N_4760,N_58,N_468);
or U4761 (N_4761,N_2225,N_1028);
nor U4762 (N_4762,N_182,N_381);
or U4763 (N_4763,N_1353,N_2997);
nor U4764 (N_4764,N_965,N_1390);
or U4765 (N_4765,N_1957,N_627);
xnor U4766 (N_4766,N_72,N_517);
and U4767 (N_4767,N_1329,N_992);
nor U4768 (N_4768,N_1331,N_723);
and U4769 (N_4769,N_2074,N_1352);
and U4770 (N_4770,N_454,N_1244);
nor U4771 (N_4771,N_1359,N_1261);
and U4772 (N_4772,N_1768,N_2268);
nand U4773 (N_4773,N_859,N_1911);
and U4774 (N_4774,N_1569,N_1270);
or U4775 (N_4775,N_2512,N_2265);
xnor U4776 (N_4776,N_648,N_2528);
nor U4777 (N_4777,N_1869,N_278);
or U4778 (N_4778,N_1190,N_887);
or U4779 (N_4779,N_2110,N_1435);
nor U4780 (N_4780,N_1702,N_2311);
and U4781 (N_4781,N_2100,N_424);
nand U4782 (N_4782,N_1092,N_1935);
or U4783 (N_4783,N_1855,N_2753);
and U4784 (N_4784,N_447,N_2753);
and U4785 (N_4785,N_1261,N_136);
and U4786 (N_4786,N_855,N_1469);
or U4787 (N_4787,N_1735,N_2010);
or U4788 (N_4788,N_1136,N_585);
nor U4789 (N_4789,N_1081,N_1796);
and U4790 (N_4790,N_2776,N_2259);
xnor U4791 (N_4791,N_375,N_2501);
and U4792 (N_4792,N_1622,N_139);
nand U4793 (N_4793,N_1157,N_698);
nand U4794 (N_4794,N_2977,N_155);
and U4795 (N_4795,N_2957,N_2382);
nand U4796 (N_4796,N_2984,N_406);
nand U4797 (N_4797,N_2727,N_1962);
or U4798 (N_4798,N_69,N_735);
and U4799 (N_4799,N_2814,N_2167);
and U4800 (N_4800,N_4,N_1200);
nand U4801 (N_4801,N_1428,N_1557);
nand U4802 (N_4802,N_1885,N_2519);
nor U4803 (N_4803,N_2277,N_2264);
nand U4804 (N_4804,N_1546,N_766);
nor U4805 (N_4805,N_1776,N_2477);
nand U4806 (N_4806,N_2028,N_2952);
or U4807 (N_4807,N_1906,N_2476);
xnor U4808 (N_4808,N_1052,N_1693);
and U4809 (N_4809,N_1898,N_1619);
nor U4810 (N_4810,N_2308,N_1984);
or U4811 (N_4811,N_2754,N_510);
or U4812 (N_4812,N_1182,N_1275);
or U4813 (N_4813,N_1845,N_2202);
nand U4814 (N_4814,N_2253,N_1719);
nand U4815 (N_4815,N_1751,N_2628);
or U4816 (N_4816,N_1290,N_16);
nor U4817 (N_4817,N_1987,N_1348);
nand U4818 (N_4818,N_1934,N_1104);
and U4819 (N_4819,N_1595,N_1740);
nand U4820 (N_4820,N_2200,N_946);
and U4821 (N_4821,N_1912,N_1963);
nor U4822 (N_4822,N_858,N_2319);
nand U4823 (N_4823,N_2881,N_2747);
nor U4824 (N_4824,N_1329,N_893);
or U4825 (N_4825,N_1708,N_1221);
or U4826 (N_4826,N_912,N_2386);
nand U4827 (N_4827,N_817,N_277);
or U4828 (N_4828,N_195,N_217);
and U4829 (N_4829,N_1730,N_2502);
or U4830 (N_4830,N_965,N_2838);
or U4831 (N_4831,N_1372,N_774);
or U4832 (N_4832,N_2127,N_1996);
nand U4833 (N_4833,N_874,N_1230);
nor U4834 (N_4834,N_1064,N_2048);
or U4835 (N_4835,N_1138,N_1699);
xnor U4836 (N_4836,N_1954,N_2574);
nor U4837 (N_4837,N_929,N_8);
and U4838 (N_4838,N_352,N_2446);
nand U4839 (N_4839,N_294,N_1873);
or U4840 (N_4840,N_1603,N_2627);
nand U4841 (N_4841,N_1012,N_1458);
nand U4842 (N_4842,N_1106,N_2997);
nand U4843 (N_4843,N_651,N_630);
and U4844 (N_4844,N_2635,N_2342);
or U4845 (N_4845,N_1307,N_1277);
and U4846 (N_4846,N_2143,N_1267);
nand U4847 (N_4847,N_1189,N_286);
nand U4848 (N_4848,N_1069,N_2339);
and U4849 (N_4849,N_2592,N_1840);
nor U4850 (N_4850,N_431,N_673);
and U4851 (N_4851,N_1502,N_2147);
and U4852 (N_4852,N_308,N_2297);
or U4853 (N_4853,N_965,N_2037);
xnor U4854 (N_4854,N_1435,N_1555);
nor U4855 (N_4855,N_2865,N_1567);
nand U4856 (N_4856,N_2802,N_49);
nor U4857 (N_4857,N_273,N_1365);
nor U4858 (N_4858,N_2303,N_2004);
and U4859 (N_4859,N_1714,N_2094);
nand U4860 (N_4860,N_2586,N_2538);
nand U4861 (N_4861,N_1348,N_1184);
and U4862 (N_4862,N_71,N_1915);
nor U4863 (N_4863,N_465,N_313);
nor U4864 (N_4864,N_2445,N_1148);
or U4865 (N_4865,N_170,N_1230);
and U4866 (N_4866,N_1886,N_2072);
nand U4867 (N_4867,N_183,N_2742);
nand U4868 (N_4868,N_832,N_2367);
xnor U4869 (N_4869,N_1825,N_857);
or U4870 (N_4870,N_1160,N_534);
nand U4871 (N_4871,N_689,N_2182);
or U4872 (N_4872,N_447,N_63);
nor U4873 (N_4873,N_241,N_82);
nand U4874 (N_4874,N_2981,N_407);
nor U4875 (N_4875,N_1928,N_1243);
nor U4876 (N_4876,N_970,N_2515);
nor U4877 (N_4877,N_241,N_2348);
or U4878 (N_4878,N_343,N_1164);
xnor U4879 (N_4879,N_714,N_2695);
and U4880 (N_4880,N_1861,N_1239);
or U4881 (N_4881,N_225,N_2334);
xnor U4882 (N_4882,N_1914,N_682);
nand U4883 (N_4883,N_2957,N_1470);
and U4884 (N_4884,N_1592,N_1923);
or U4885 (N_4885,N_599,N_1178);
and U4886 (N_4886,N_2914,N_2208);
nand U4887 (N_4887,N_2902,N_1138);
nand U4888 (N_4888,N_2333,N_1941);
or U4889 (N_4889,N_1258,N_2044);
nor U4890 (N_4890,N_116,N_414);
or U4891 (N_4891,N_1238,N_2831);
and U4892 (N_4892,N_1506,N_2744);
and U4893 (N_4893,N_514,N_330);
nor U4894 (N_4894,N_1115,N_1821);
or U4895 (N_4895,N_1386,N_1400);
nand U4896 (N_4896,N_1109,N_255);
nand U4897 (N_4897,N_729,N_1112);
nor U4898 (N_4898,N_1364,N_2777);
or U4899 (N_4899,N_164,N_1763);
nor U4900 (N_4900,N_2496,N_561);
nor U4901 (N_4901,N_1702,N_1275);
nor U4902 (N_4902,N_88,N_1700);
nor U4903 (N_4903,N_422,N_714);
or U4904 (N_4904,N_1085,N_1893);
xor U4905 (N_4905,N_1271,N_1487);
or U4906 (N_4906,N_1207,N_2872);
or U4907 (N_4907,N_361,N_1770);
nand U4908 (N_4908,N_1324,N_2808);
or U4909 (N_4909,N_2320,N_1163);
nand U4910 (N_4910,N_1510,N_362);
and U4911 (N_4911,N_1472,N_43);
or U4912 (N_4912,N_2237,N_613);
xor U4913 (N_4913,N_160,N_515);
xor U4914 (N_4914,N_1809,N_35);
or U4915 (N_4915,N_2778,N_133);
or U4916 (N_4916,N_2266,N_1964);
xnor U4917 (N_4917,N_1839,N_1109);
nor U4918 (N_4918,N_461,N_58);
or U4919 (N_4919,N_969,N_640);
and U4920 (N_4920,N_2356,N_644);
and U4921 (N_4921,N_2168,N_953);
nand U4922 (N_4922,N_261,N_807);
nor U4923 (N_4923,N_1933,N_652);
and U4924 (N_4924,N_209,N_868);
nor U4925 (N_4925,N_1652,N_306);
nand U4926 (N_4926,N_1561,N_2803);
nor U4927 (N_4927,N_1240,N_1518);
xnor U4928 (N_4928,N_1457,N_807);
or U4929 (N_4929,N_412,N_2587);
nand U4930 (N_4930,N_2904,N_2348);
or U4931 (N_4931,N_1487,N_2948);
or U4932 (N_4932,N_2957,N_1437);
nor U4933 (N_4933,N_1809,N_1285);
and U4934 (N_4934,N_1907,N_1210);
nor U4935 (N_4935,N_932,N_881);
nor U4936 (N_4936,N_692,N_1518);
nand U4937 (N_4937,N_1200,N_2452);
or U4938 (N_4938,N_190,N_307);
and U4939 (N_4939,N_1545,N_1795);
or U4940 (N_4940,N_2862,N_1712);
nand U4941 (N_4941,N_1833,N_2060);
and U4942 (N_4942,N_1790,N_412);
nand U4943 (N_4943,N_901,N_170);
nor U4944 (N_4944,N_2556,N_1835);
xor U4945 (N_4945,N_1392,N_1219);
or U4946 (N_4946,N_1325,N_2516);
nand U4947 (N_4947,N_1985,N_2471);
nand U4948 (N_4948,N_2132,N_2259);
or U4949 (N_4949,N_523,N_985);
nor U4950 (N_4950,N_1067,N_1501);
nand U4951 (N_4951,N_1970,N_176);
nor U4952 (N_4952,N_1916,N_777);
nand U4953 (N_4953,N_1541,N_2292);
nor U4954 (N_4954,N_215,N_1413);
or U4955 (N_4955,N_2299,N_2204);
nor U4956 (N_4956,N_89,N_594);
or U4957 (N_4957,N_164,N_125);
xnor U4958 (N_4958,N_1538,N_307);
or U4959 (N_4959,N_2497,N_2837);
nor U4960 (N_4960,N_2628,N_2547);
nand U4961 (N_4961,N_942,N_2771);
and U4962 (N_4962,N_2726,N_1243);
and U4963 (N_4963,N_2006,N_2425);
nor U4964 (N_4964,N_1218,N_1364);
nand U4965 (N_4965,N_893,N_2769);
nor U4966 (N_4966,N_1410,N_1162);
nand U4967 (N_4967,N_1459,N_2916);
or U4968 (N_4968,N_2707,N_1975);
nor U4969 (N_4969,N_2532,N_499);
nand U4970 (N_4970,N_2222,N_1283);
xor U4971 (N_4971,N_2724,N_651);
xor U4972 (N_4972,N_194,N_213);
or U4973 (N_4973,N_1989,N_2502);
and U4974 (N_4974,N_880,N_256);
and U4975 (N_4975,N_1078,N_2150);
or U4976 (N_4976,N_1651,N_1555);
or U4977 (N_4977,N_2562,N_2399);
or U4978 (N_4978,N_499,N_2051);
nand U4979 (N_4979,N_2158,N_832);
xnor U4980 (N_4980,N_1036,N_660);
and U4981 (N_4981,N_499,N_998);
nor U4982 (N_4982,N_492,N_2789);
or U4983 (N_4983,N_925,N_275);
nand U4984 (N_4984,N_2755,N_992);
nor U4985 (N_4985,N_2679,N_2773);
or U4986 (N_4986,N_2873,N_2526);
xor U4987 (N_4987,N_1527,N_2173);
nand U4988 (N_4988,N_227,N_766);
and U4989 (N_4989,N_58,N_321);
nand U4990 (N_4990,N_1027,N_1586);
or U4991 (N_4991,N_2961,N_1941);
or U4992 (N_4992,N_1824,N_745);
and U4993 (N_4993,N_1487,N_2999);
or U4994 (N_4994,N_2093,N_2750);
nand U4995 (N_4995,N_948,N_664);
xor U4996 (N_4996,N_898,N_651);
nand U4997 (N_4997,N_2683,N_2978);
nand U4998 (N_4998,N_1812,N_1808);
and U4999 (N_4999,N_833,N_2202);
nand U5000 (N_5000,N_2613,N_2893);
or U5001 (N_5001,N_1671,N_2992);
nor U5002 (N_5002,N_576,N_887);
or U5003 (N_5003,N_2674,N_618);
nand U5004 (N_5004,N_2064,N_2075);
nand U5005 (N_5005,N_281,N_2827);
and U5006 (N_5006,N_2920,N_1244);
or U5007 (N_5007,N_1287,N_881);
xor U5008 (N_5008,N_1207,N_2657);
and U5009 (N_5009,N_1695,N_1730);
nand U5010 (N_5010,N_2857,N_2475);
or U5011 (N_5011,N_1815,N_2937);
nand U5012 (N_5012,N_1596,N_2157);
xor U5013 (N_5013,N_1340,N_25);
or U5014 (N_5014,N_2493,N_906);
and U5015 (N_5015,N_2336,N_600);
nor U5016 (N_5016,N_1903,N_1645);
nor U5017 (N_5017,N_1161,N_2477);
nor U5018 (N_5018,N_1842,N_1981);
xor U5019 (N_5019,N_2211,N_708);
or U5020 (N_5020,N_2406,N_1898);
nor U5021 (N_5021,N_47,N_561);
nor U5022 (N_5022,N_1335,N_1036);
or U5023 (N_5023,N_850,N_332);
or U5024 (N_5024,N_1552,N_2201);
nor U5025 (N_5025,N_1296,N_1374);
nor U5026 (N_5026,N_135,N_536);
nand U5027 (N_5027,N_1176,N_1418);
nor U5028 (N_5028,N_2302,N_122);
nand U5029 (N_5029,N_2994,N_920);
or U5030 (N_5030,N_1490,N_677);
nor U5031 (N_5031,N_2336,N_1663);
or U5032 (N_5032,N_1384,N_2912);
or U5033 (N_5033,N_2986,N_2099);
or U5034 (N_5034,N_1297,N_1419);
or U5035 (N_5035,N_40,N_206);
nor U5036 (N_5036,N_1859,N_2364);
nor U5037 (N_5037,N_2818,N_1504);
and U5038 (N_5038,N_986,N_115);
xnor U5039 (N_5039,N_2517,N_1859);
and U5040 (N_5040,N_1962,N_140);
xor U5041 (N_5041,N_610,N_657);
and U5042 (N_5042,N_1646,N_134);
nand U5043 (N_5043,N_588,N_2295);
nand U5044 (N_5044,N_876,N_2896);
and U5045 (N_5045,N_513,N_2467);
or U5046 (N_5046,N_2699,N_647);
nor U5047 (N_5047,N_115,N_2665);
and U5048 (N_5048,N_841,N_811);
nor U5049 (N_5049,N_1414,N_16);
and U5050 (N_5050,N_2375,N_2366);
nor U5051 (N_5051,N_2824,N_2339);
or U5052 (N_5052,N_1355,N_1270);
nand U5053 (N_5053,N_2876,N_2943);
nor U5054 (N_5054,N_450,N_2358);
nor U5055 (N_5055,N_1588,N_1473);
and U5056 (N_5056,N_988,N_824);
and U5057 (N_5057,N_2295,N_212);
nand U5058 (N_5058,N_2668,N_2637);
or U5059 (N_5059,N_2230,N_1272);
and U5060 (N_5060,N_1083,N_547);
xnor U5061 (N_5061,N_1368,N_895);
nor U5062 (N_5062,N_1474,N_2960);
and U5063 (N_5063,N_1331,N_2827);
nand U5064 (N_5064,N_429,N_2691);
nor U5065 (N_5065,N_2734,N_1214);
nand U5066 (N_5066,N_1422,N_1745);
nand U5067 (N_5067,N_2807,N_2936);
or U5068 (N_5068,N_1136,N_2791);
xor U5069 (N_5069,N_691,N_184);
nand U5070 (N_5070,N_1863,N_2293);
or U5071 (N_5071,N_685,N_12);
and U5072 (N_5072,N_1372,N_131);
nand U5073 (N_5073,N_79,N_1735);
nand U5074 (N_5074,N_2105,N_2119);
nor U5075 (N_5075,N_2711,N_138);
or U5076 (N_5076,N_1044,N_1791);
nand U5077 (N_5077,N_107,N_1452);
nand U5078 (N_5078,N_289,N_673);
nor U5079 (N_5079,N_2060,N_596);
xor U5080 (N_5080,N_1,N_1554);
and U5081 (N_5081,N_2018,N_2632);
nor U5082 (N_5082,N_23,N_2124);
xor U5083 (N_5083,N_1960,N_1686);
and U5084 (N_5084,N_1727,N_517);
and U5085 (N_5085,N_423,N_1751);
nand U5086 (N_5086,N_156,N_2454);
and U5087 (N_5087,N_332,N_291);
and U5088 (N_5088,N_1627,N_269);
or U5089 (N_5089,N_1711,N_151);
and U5090 (N_5090,N_2059,N_1830);
and U5091 (N_5091,N_1504,N_1361);
nor U5092 (N_5092,N_2105,N_2766);
xor U5093 (N_5093,N_1104,N_2935);
and U5094 (N_5094,N_1931,N_1654);
nor U5095 (N_5095,N_2470,N_2387);
or U5096 (N_5096,N_2697,N_1536);
and U5097 (N_5097,N_2967,N_1308);
and U5098 (N_5098,N_1441,N_174);
and U5099 (N_5099,N_2794,N_2913);
or U5100 (N_5100,N_88,N_228);
nor U5101 (N_5101,N_965,N_1957);
or U5102 (N_5102,N_558,N_551);
and U5103 (N_5103,N_1073,N_1763);
nor U5104 (N_5104,N_64,N_152);
or U5105 (N_5105,N_2870,N_1361);
or U5106 (N_5106,N_974,N_1008);
or U5107 (N_5107,N_1796,N_312);
and U5108 (N_5108,N_2611,N_2502);
nor U5109 (N_5109,N_2155,N_2188);
nor U5110 (N_5110,N_1960,N_2993);
or U5111 (N_5111,N_2533,N_1117);
nor U5112 (N_5112,N_2339,N_4);
nand U5113 (N_5113,N_634,N_2881);
and U5114 (N_5114,N_772,N_315);
nor U5115 (N_5115,N_1572,N_562);
or U5116 (N_5116,N_1194,N_296);
and U5117 (N_5117,N_66,N_2950);
and U5118 (N_5118,N_2778,N_2505);
nand U5119 (N_5119,N_1813,N_328);
nor U5120 (N_5120,N_2105,N_1331);
or U5121 (N_5121,N_1791,N_497);
and U5122 (N_5122,N_1,N_2657);
nor U5123 (N_5123,N_1748,N_2757);
or U5124 (N_5124,N_1223,N_1173);
nand U5125 (N_5125,N_439,N_1759);
nand U5126 (N_5126,N_2096,N_1219);
or U5127 (N_5127,N_1013,N_1912);
nor U5128 (N_5128,N_2853,N_2513);
xnor U5129 (N_5129,N_1033,N_2528);
nand U5130 (N_5130,N_1247,N_2290);
nand U5131 (N_5131,N_298,N_211);
or U5132 (N_5132,N_1667,N_53);
nand U5133 (N_5133,N_1778,N_1964);
and U5134 (N_5134,N_2078,N_464);
nand U5135 (N_5135,N_51,N_2045);
and U5136 (N_5136,N_1110,N_376);
nand U5137 (N_5137,N_74,N_2472);
or U5138 (N_5138,N_1715,N_459);
and U5139 (N_5139,N_88,N_1563);
or U5140 (N_5140,N_1503,N_562);
and U5141 (N_5141,N_2919,N_872);
and U5142 (N_5142,N_434,N_2976);
nand U5143 (N_5143,N_85,N_1212);
xor U5144 (N_5144,N_2399,N_2527);
nand U5145 (N_5145,N_559,N_1977);
nand U5146 (N_5146,N_1456,N_2975);
nor U5147 (N_5147,N_1846,N_1978);
and U5148 (N_5148,N_1643,N_1584);
nand U5149 (N_5149,N_356,N_496);
nand U5150 (N_5150,N_1511,N_1786);
xnor U5151 (N_5151,N_1156,N_704);
nor U5152 (N_5152,N_508,N_1784);
nor U5153 (N_5153,N_1669,N_966);
and U5154 (N_5154,N_1601,N_2079);
or U5155 (N_5155,N_2233,N_1079);
and U5156 (N_5156,N_78,N_2691);
nor U5157 (N_5157,N_1957,N_2487);
or U5158 (N_5158,N_162,N_96);
and U5159 (N_5159,N_2250,N_1627);
and U5160 (N_5160,N_770,N_1704);
or U5161 (N_5161,N_2165,N_2563);
or U5162 (N_5162,N_1327,N_1588);
and U5163 (N_5163,N_2937,N_1428);
nand U5164 (N_5164,N_1370,N_2718);
nor U5165 (N_5165,N_582,N_881);
and U5166 (N_5166,N_1273,N_1818);
or U5167 (N_5167,N_564,N_1295);
and U5168 (N_5168,N_507,N_680);
nand U5169 (N_5169,N_2352,N_2949);
or U5170 (N_5170,N_459,N_2731);
and U5171 (N_5171,N_2202,N_503);
xor U5172 (N_5172,N_802,N_2207);
or U5173 (N_5173,N_2606,N_757);
or U5174 (N_5174,N_2760,N_2331);
or U5175 (N_5175,N_2049,N_1085);
nor U5176 (N_5176,N_951,N_2694);
or U5177 (N_5177,N_2929,N_2749);
nor U5178 (N_5178,N_2762,N_1179);
nor U5179 (N_5179,N_1287,N_436);
or U5180 (N_5180,N_1307,N_1356);
and U5181 (N_5181,N_369,N_1407);
or U5182 (N_5182,N_1796,N_2639);
nand U5183 (N_5183,N_533,N_2544);
nor U5184 (N_5184,N_955,N_1210);
or U5185 (N_5185,N_1717,N_1009);
nand U5186 (N_5186,N_1319,N_2500);
or U5187 (N_5187,N_1393,N_2914);
or U5188 (N_5188,N_928,N_1773);
xnor U5189 (N_5189,N_321,N_803);
and U5190 (N_5190,N_2028,N_2355);
xor U5191 (N_5191,N_1686,N_2996);
xnor U5192 (N_5192,N_584,N_2921);
xnor U5193 (N_5193,N_357,N_1161);
nor U5194 (N_5194,N_2709,N_1020);
xnor U5195 (N_5195,N_540,N_121);
nand U5196 (N_5196,N_337,N_2402);
nand U5197 (N_5197,N_2317,N_1978);
nand U5198 (N_5198,N_1092,N_2715);
nand U5199 (N_5199,N_1651,N_2791);
nand U5200 (N_5200,N_32,N_2932);
nor U5201 (N_5201,N_945,N_82);
nor U5202 (N_5202,N_878,N_2957);
or U5203 (N_5203,N_2569,N_2885);
or U5204 (N_5204,N_1047,N_537);
nor U5205 (N_5205,N_208,N_1748);
xor U5206 (N_5206,N_764,N_1974);
nor U5207 (N_5207,N_585,N_2280);
nor U5208 (N_5208,N_2705,N_2102);
nand U5209 (N_5209,N_551,N_79);
and U5210 (N_5210,N_2048,N_973);
nor U5211 (N_5211,N_1302,N_1433);
xnor U5212 (N_5212,N_1241,N_1613);
nand U5213 (N_5213,N_626,N_2829);
or U5214 (N_5214,N_213,N_2312);
or U5215 (N_5215,N_1849,N_2758);
or U5216 (N_5216,N_836,N_1224);
nand U5217 (N_5217,N_2365,N_387);
nor U5218 (N_5218,N_1213,N_2811);
and U5219 (N_5219,N_1992,N_2668);
and U5220 (N_5220,N_1921,N_1439);
and U5221 (N_5221,N_86,N_1754);
or U5222 (N_5222,N_2405,N_145);
or U5223 (N_5223,N_229,N_2582);
and U5224 (N_5224,N_1944,N_2550);
or U5225 (N_5225,N_2406,N_2419);
and U5226 (N_5226,N_2652,N_2252);
or U5227 (N_5227,N_2009,N_1985);
nor U5228 (N_5228,N_420,N_563);
and U5229 (N_5229,N_329,N_722);
or U5230 (N_5230,N_2367,N_560);
nand U5231 (N_5231,N_21,N_618);
and U5232 (N_5232,N_2014,N_2479);
and U5233 (N_5233,N_1795,N_2899);
or U5234 (N_5234,N_1425,N_592);
and U5235 (N_5235,N_255,N_711);
nor U5236 (N_5236,N_505,N_2494);
and U5237 (N_5237,N_368,N_1462);
nor U5238 (N_5238,N_1447,N_2093);
or U5239 (N_5239,N_262,N_305);
or U5240 (N_5240,N_1368,N_553);
and U5241 (N_5241,N_1760,N_2551);
nand U5242 (N_5242,N_2591,N_592);
nor U5243 (N_5243,N_2596,N_46);
nand U5244 (N_5244,N_1372,N_616);
nand U5245 (N_5245,N_1038,N_2169);
nand U5246 (N_5246,N_1170,N_138);
and U5247 (N_5247,N_1747,N_1917);
nor U5248 (N_5248,N_2902,N_2508);
and U5249 (N_5249,N_1537,N_749);
and U5250 (N_5250,N_6,N_1716);
nand U5251 (N_5251,N_2607,N_2013);
nand U5252 (N_5252,N_286,N_388);
or U5253 (N_5253,N_2089,N_1589);
and U5254 (N_5254,N_2092,N_871);
nor U5255 (N_5255,N_952,N_1945);
or U5256 (N_5256,N_77,N_998);
and U5257 (N_5257,N_1114,N_437);
nand U5258 (N_5258,N_2253,N_946);
nor U5259 (N_5259,N_1339,N_2265);
xnor U5260 (N_5260,N_1214,N_2006);
xor U5261 (N_5261,N_804,N_1902);
nand U5262 (N_5262,N_201,N_39);
and U5263 (N_5263,N_2113,N_999);
nand U5264 (N_5264,N_2495,N_2553);
nor U5265 (N_5265,N_2312,N_1787);
or U5266 (N_5266,N_2139,N_2666);
and U5267 (N_5267,N_2686,N_640);
or U5268 (N_5268,N_2386,N_1785);
nor U5269 (N_5269,N_2163,N_59);
or U5270 (N_5270,N_838,N_2236);
nor U5271 (N_5271,N_2930,N_2319);
nand U5272 (N_5272,N_2596,N_676);
nor U5273 (N_5273,N_2734,N_1370);
xor U5274 (N_5274,N_634,N_846);
nand U5275 (N_5275,N_180,N_1769);
nor U5276 (N_5276,N_1229,N_2096);
nor U5277 (N_5277,N_2675,N_2190);
and U5278 (N_5278,N_2751,N_1381);
nor U5279 (N_5279,N_1791,N_1803);
or U5280 (N_5280,N_1698,N_1761);
xnor U5281 (N_5281,N_1288,N_198);
nand U5282 (N_5282,N_305,N_1115);
and U5283 (N_5283,N_2184,N_2772);
or U5284 (N_5284,N_1152,N_2069);
nand U5285 (N_5285,N_1249,N_2429);
and U5286 (N_5286,N_807,N_1636);
and U5287 (N_5287,N_2842,N_1936);
and U5288 (N_5288,N_2122,N_1910);
and U5289 (N_5289,N_782,N_2218);
and U5290 (N_5290,N_559,N_823);
xor U5291 (N_5291,N_2968,N_2158);
nand U5292 (N_5292,N_120,N_392);
or U5293 (N_5293,N_1237,N_155);
or U5294 (N_5294,N_390,N_992);
and U5295 (N_5295,N_2017,N_1289);
nand U5296 (N_5296,N_2107,N_479);
nor U5297 (N_5297,N_2081,N_1449);
nand U5298 (N_5298,N_2853,N_1234);
nand U5299 (N_5299,N_2628,N_2447);
or U5300 (N_5300,N_1639,N_1216);
nor U5301 (N_5301,N_1233,N_193);
nor U5302 (N_5302,N_2867,N_1118);
nor U5303 (N_5303,N_2076,N_934);
nand U5304 (N_5304,N_474,N_950);
nor U5305 (N_5305,N_1936,N_2057);
nand U5306 (N_5306,N_648,N_290);
nor U5307 (N_5307,N_1503,N_2214);
or U5308 (N_5308,N_2270,N_1149);
or U5309 (N_5309,N_2018,N_1704);
nor U5310 (N_5310,N_414,N_2005);
and U5311 (N_5311,N_469,N_2556);
nand U5312 (N_5312,N_2047,N_2631);
and U5313 (N_5313,N_167,N_1273);
nand U5314 (N_5314,N_998,N_53);
nor U5315 (N_5315,N_2075,N_707);
nor U5316 (N_5316,N_1477,N_1475);
xor U5317 (N_5317,N_458,N_980);
and U5318 (N_5318,N_559,N_1173);
nand U5319 (N_5319,N_1554,N_375);
nor U5320 (N_5320,N_1327,N_464);
nor U5321 (N_5321,N_1267,N_2315);
nor U5322 (N_5322,N_2236,N_605);
nand U5323 (N_5323,N_1086,N_1936);
nor U5324 (N_5324,N_2625,N_92);
and U5325 (N_5325,N_2523,N_2899);
or U5326 (N_5326,N_1452,N_700);
nand U5327 (N_5327,N_2994,N_2217);
xor U5328 (N_5328,N_2220,N_1535);
nand U5329 (N_5329,N_2329,N_1011);
or U5330 (N_5330,N_92,N_254);
nor U5331 (N_5331,N_381,N_2931);
and U5332 (N_5332,N_1232,N_2856);
xnor U5333 (N_5333,N_2271,N_1181);
or U5334 (N_5334,N_583,N_1011);
nor U5335 (N_5335,N_2862,N_2171);
and U5336 (N_5336,N_150,N_2788);
and U5337 (N_5337,N_1009,N_2781);
or U5338 (N_5338,N_1532,N_87);
and U5339 (N_5339,N_2719,N_67);
nand U5340 (N_5340,N_1050,N_2141);
and U5341 (N_5341,N_2765,N_1670);
nor U5342 (N_5342,N_1988,N_2868);
and U5343 (N_5343,N_1865,N_1375);
xor U5344 (N_5344,N_1796,N_1355);
nand U5345 (N_5345,N_620,N_416);
and U5346 (N_5346,N_2666,N_722);
xnor U5347 (N_5347,N_404,N_964);
nand U5348 (N_5348,N_1765,N_1743);
or U5349 (N_5349,N_1033,N_678);
and U5350 (N_5350,N_627,N_2573);
and U5351 (N_5351,N_1866,N_1981);
nand U5352 (N_5352,N_2819,N_2544);
nand U5353 (N_5353,N_151,N_1357);
nor U5354 (N_5354,N_2899,N_2320);
and U5355 (N_5355,N_2309,N_1732);
or U5356 (N_5356,N_629,N_2797);
and U5357 (N_5357,N_2698,N_2001);
nand U5358 (N_5358,N_442,N_1863);
nand U5359 (N_5359,N_2596,N_2580);
or U5360 (N_5360,N_193,N_1273);
nor U5361 (N_5361,N_2593,N_222);
or U5362 (N_5362,N_2366,N_208);
nor U5363 (N_5363,N_1826,N_1536);
or U5364 (N_5364,N_698,N_544);
and U5365 (N_5365,N_1048,N_2939);
nor U5366 (N_5366,N_875,N_687);
nand U5367 (N_5367,N_907,N_2073);
nor U5368 (N_5368,N_802,N_2718);
nor U5369 (N_5369,N_463,N_1984);
nand U5370 (N_5370,N_743,N_752);
and U5371 (N_5371,N_897,N_2386);
xnor U5372 (N_5372,N_1428,N_595);
nand U5373 (N_5373,N_649,N_1423);
nor U5374 (N_5374,N_1038,N_1008);
nand U5375 (N_5375,N_1759,N_1415);
nand U5376 (N_5376,N_990,N_338);
xnor U5377 (N_5377,N_1611,N_247);
and U5378 (N_5378,N_2700,N_1331);
xnor U5379 (N_5379,N_1193,N_772);
nand U5380 (N_5380,N_2953,N_1061);
and U5381 (N_5381,N_2038,N_734);
nor U5382 (N_5382,N_1064,N_70);
nor U5383 (N_5383,N_287,N_1549);
nand U5384 (N_5384,N_122,N_1139);
or U5385 (N_5385,N_1966,N_2841);
and U5386 (N_5386,N_1394,N_778);
or U5387 (N_5387,N_429,N_782);
and U5388 (N_5388,N_2582,N_2250);
nand U5389 (N_5389,N_2990,N_1330);
nand U5390 (N_5390,N_711,N_1802);
nor U5391 (N_5391,N_1356,N_2517);
and U5392 (N_5392,N_1727,N_2058);
or U5393 (N_5393,N_2398,N_1013);
and U5394 (N_5394,N_2469,N_94);
nand U5395 (N_5395,N_2348,N_2236);
and U5396 (N_5396,N_2544,N_2627);
and U5397 (N_5397,N_2729,N_2563);
nand U5398 (N_5398,N_1203,N_1107);
nand U5399 (N_5399,N_528,N_917);
xor U5400 (N_5400,N_2136,N_1399);
nor U5401 (N_5401,N_1038,N_1768);
nor U5402 (N_5402,N_1605,N_1419);
nor U5403 (N_5403,N_1046,N_2475);
nand U5404 (N_5404,N_439,N_1140);
xor U5405 (N_5405,N_2447,N_880);
nor U5406 (N_5406,N_959,N_1459);
nor U5407 (N_5407,N_407,N_1205);
and U5408 (N_5408,N_2174,N_914);
nor U5409 (N_5409,N_2668,N_2198);
or U5410 (N_5410,N_1264,N_14);
nor U5411 (N_5411,N_2140,N_1916);
nor U5412 (N_5412,N_1174,N_259);
nand U5413 (N_5413,N_755,N_2029);
nand U5414 (N_5414,N_970,N_1138);
nand U5415 (N_5415,N_163,N_155);
nor U5416 (N_5416,N_1981,N_994);
or U5417 (N_5417,N_2114,N_836);
nand U5418 (N_5418,N_2318,N_937);
nand U5419 (N_5419,N_2564,N_1941);
nor U5420 (N_5420,N_88,N_1853);
and U5421 (N_5421,N_1274,N_942);
or U5422 (N_5422,N_1964,N_457);
or U5423 (N_5423,N_1962,N_1354);
xor U5424 (N_5424,N_2604,N_2559);
nand U5425 (N_5425,N_743,N_849);
or U5426 (N_5426,N_564,N_1643);
nand U5427 (N_5427,N_2708,N_1820);
nor U5428 (N_5428,N_2539,N_1816);
xnor U5429 (N_5429,N_562,N_1184);
and U5430 (N_5430,N_566,N_1035);
nor U5431 (N_5431,N_2801,N_1101);
or U5432 (N_5432,N_2161,N_2497);
or U5433 (N_5433,N_1517,N_86);
nand U5434 (N_5434,N_500,N_2000);
or U5435 (N_5435,N_379,N_1660);
nor U5436 (N_5436,N_2761,N_1201);
or U5437 (N_5437,N_1644,N_2401);
nor U5438 (N_5438,N_295,N_2820);
or U5439 (N_5439,N_901,N_1419);
xor U5440 (N_5440,N_208,N_2911);
and U5441 (N_5441,N_862,N_2359);
xor U5442 (N_5442,N_2021,N_1169);
xnor U5443 (N_5443,N_2617,N_1436);
and U5444 (N_5444,N_2169,N_1752);
or U5445 (N_5445,N_802,N_630);
and U5446 (N_5446,N_919,N_1814);
and U5447 (N_5447,N_45,N_2454);
nor U5448 (N_5448,N_1556,N_2734);
or U5449 (N_5449,N_270,N_670);
and U5450 (N_5450,N_2904,N_2311);
nor U5451 (N_5451,N_146,N_1956);
and U5452 (N_5452,N_813,N_271);
and U5453 (N_5453,N_656,N_1579);
or U5454 (N_5454,N_1566,N_601);
or U5455 (N_5455,N_2444,N_1789);
or U5456 (N_5456,N_165,N_1792);
and U5457 (N_5457,N_1962,N_727);
nand U5458 (N_5458,N_637,N_791);
or U5459 (N_5459,N_2125,N_1070);
nor U5460 (N_5460,N_57,N_897);
or U5461 (N_5461,N_1472,N_367);
or U5462 (N_5462,N_417,N_991);
or U5463 (N_5463,N_2945,N_1843);
nand U5464 (N_5464,N_2003,N_665);
and U5465 (N_5465,N_798,N_836);
nand U5466 (N_5466,N_2179,N_765);
and U5467 (N_5467,N_2124,N_2405);
xor U5468 (N_5468,N_1978,N_541);
or U5469 (N_5469,N_1170,N_2163);
and U5470 (N_5470,N_1011,N_1417);
or U5471 (N_5471,N_1261,N_2727);
nand U5472 (N_5472,N_1812,N_2372);
nand U5473 (N_5473,N_2788,N_1750);
or U5474 (N_5474,N_1575,N_142);
nand U5475 (N_5475,N_407,N_88);
and U5476 (N_5476,N_2592,N_715);
or U5477 (N_5477,N_86,N_2834);
nor U5478 (N_5478,N_1477,N_2030);
or U5479 (N_5479,N_1490,N_1489);
nand U5480 (N_5480,N_2452,N_712);
nor U5481 (N_5481,N_2094,N_676);
nand U5482 (N_5482,N_1655,N_353);
or U5483 (N_5483,N_2360,N_2803);
or U5484 (N_5484,N_1237,N_446);
and U5485 (N_5485,N_120,N_2915);
and U5486 (N_5486,N_1351,N_567);
and U5487 (N_5487,N_1015,N_770);
and U5488 (N_5488,N_129,N_959);
and U5489 (N_5489,N_2011,N_743);
or U5490 (N_5490,N_1095,N_2153);
nand U5491 (N_5491,N_153,N_466);
nor U5492 (N_5492,N_2077,N_2730);
nand U5493 (N_5493,N_116,N_123);
nor U5494 (N_5494,N_2810,N_148);
nor U5495 (N_5495,N_1027,N_948);
or U5496 (N_5496,N_2557,N_2550);
nand U5497 (N_5497,N_2371,N_2235);
nor U5498 (N_5498,N_1374,N_591);
nand U5499 (N_5499,N_1528,N_1853);
or U5500 (N_5500,N_1802,N_2420);
xor U5501 (N_5501,N_1115,N_62);
xnor U5502 (N_5502,N_2246,N_1819);
nor U5503 (N_5503,N_1969,N_1395);
or U5504 (N_5504,N_2895,N_2551);
and U5505 (N_5505,N_594,N_1112);
and U5506 (N_5506,N_163,N_397);
and U5507 (N_5507,N_66,N_405);
nor U5508 (N_5508,N_238,N_866);
nor U5509 (N_5509,N_2879,N_2142);
nand U5510 (N_5510,N_2256,N_2078);
nor U5511 (N_5511,N_360,N_808);
nand U5512 (N_5512,N_1482,N_1639);
nand U5513 (N_5513,N_1870,N_2105);
nor U5514 (N_5514,N_2211,N_1531);
nor U5515 (N_5515,N_2618,N_2487);
and U5516 (N_5516,N_2481,N_312);
xnor U5517 (N_5517,N_428,N_248);
or U5518 (N_5518,N_2469,N_750);
nor U5519 (N_5519,N_368,N_313);
and U5520 (N_5520,N_2319,N_913);
nor U5521 (N_5521,N_1133,N_244);
nor U5522 (N_5522,N_2639,N_165);
nor U5523 (N_5523,N_1146,N_701);
nand U5524 (N_5524,N_649,N_488);
or U5525 (N_5525,N_2588,N_1109);
nor U5526 (N_5526,N_1067,N_1036);
or U5527 (N_5527,N_2213,N_1635);
and U5528 (N_5528,N_1693,N_1390);
nor U5529 (N_5529,N_2782,N_104);
and U5530 (N_5530,N_2248,N_1881);
nor U5531 (N_5531,N_2475,N_716);
nor U5532 (N_5532,N_315,N_1689);
or U5533 (N_5533,N_1596,N_1537);
nor U5534 (N_5534,N_2141,N_2363);
nand U5535 (N_5535,N_2102,N_2407);
and U5536 (N_5536,N_1320,N_1403);
or U5537 (N_5537,N_2673,N_1735);
or U5538 (N_5538,N_412,N_1959);
nand U5539 (N_5539,N_947,N_2005);
and U5540 (N_5540,N_2016,N_358);
xor U5541 (N_5541,N_2597,N_1044);
nand U5542 (N_5542,N_1561,N_2616);
and U5543 (N_5543,N_1134,N_2503);
nor U5544 (N_5544,N_1585,N_1888);
and U5545 (N_5545,N_1878,N_838);
nand U5546 (N_5546,N_2511,N_1008);
and U5547 (N_5547,N_992,N_1367);
nor U5548 (N_5548,N_248,N_2341);
or U5549 (N_5549,N_2373,N_2585);
nor U5550 (N_5550,N_1039,N_692);
nor U5551 (N_5551,N_4,N_1349);
or U5552 (N_5552,N_316,N_1246);
and U5553 (N_5553,N_123,N_2494);
nand U5554 (N_5554,N_1120,N_2391);
and U5555 (N_5555,N_378,N_1665);
xor U5556 (N_5556,N_54,N_1879);
nor U5557 (N_5557,N_2506,N_1986);
and U5558 (N_5558,N_262,N_1536);
nor U5559 (N_5559,N_802,N_334);
nor U5560 (N_5560,N_2753,N_1038);
nor U5561 (N_5561,N_2060,N_224);
and U5562 (N_5562,N_742,N_2562);
or U5563 (N_5563,N_258,N_1909);
and U5564 (N_5564,N_2576,N_1818);
xor U5565 (N_5565,N_1988,N_1633);
and U5566 (N_5566,N_2872,N_2360);
nor U5567 (N_5567,N_719,N_1172);
nand U5568 (N_5568,N_38,N_116);
xnor U5569 (N_5569,N_2746,N_1121);
and U5570 (N_5570,N_2669,N_1529);
and U5571 (N_5571,N_926,N_2663);
nand U5572 (N_5572,N_1148,N_449);
and U5573 (N_5573,N_1254,N_2997);
and U5574 (N_5574,N_812,N_2993);
nor U5575 (N_5575,N_715,N_2394);
nand U5576 (N_5576,N_1061,N_2485);
nand U5577 (N_5577,N_2712,N_498);
or U5578 (N_5578,N_1516,N_2467);
or U5579 (N_5579,N_2015,N_236);
nor U5580 (N_5580,N_2643,N_56);
and U5581 (N_5581,N_964,N_591);
and U5582 (N_5582,N_805,N_732);
or U5583 (N_5583,N_1237,N_2832);
or U5584 (N_5584,N_1979,N_602);
or U5585 (N_5585,N_1600,N_1359);
and U5586 (N_5586,N_626,N_187);
nand U5587 (N_5587,N_914,N_2671);
nand U5588 (N_5588,N_1015,N_2793);
nor U5589 (N_5589,N_174,N_2106);
and U5590 (N_5590,N_2484,N_1866);
and U5591 (N_5591,N_2907,N_20);
nor U5592 (N_5592,N_1336,N_128);
nor U5593 (N_5593,N_118,N_1678);
nor U5594 (N_5594,N_434,N_923);
nor U5595 (N_5595,N_2958,N_840);
or U5596 (N_5596,N_1416,N_2903);
and U5597 (N_5597,N_2980,N_2730);
and U5598 (N_5598,N_1748,N_2896);
nand U5599 (N_5599,N_1553,N_253);
xor U5600 (N_5600,N_1226,N_83);
and U5601 (N_5601,N_1550,N_1989);
nand U5602 (N_5602,N_971,N_255);
or U5603 (N_5603,N_1167,N_2815);
nand U5604 (N_5604,N_1523,N_1126);
nand U5605 (N_5605,N_1850,N_62);
and U5606 (N_5606,N_129,N_2250);
xnor U5607 (N_5607,N_2119,N_873);
nand U5608 (N_5608,N_2534,N_1046);
and U5609 (N_5609,N_1738,N_1444);
nand U5610 (N_5610,N_134,N_1989);
nand U5611 (N_5611,N_402,N_2162);
nand U5612 (N_5612,N_544,N_2275);
or U5613 (N_5613,N_2811,N_1);
or U5614 (N_5614,N_400,N_1417);
nand U5615 (N_5615,N_2330,N_1089);
nor U5616 (N_5616,N_2498,N_1121);
nand U5617 (N_5617,N_2692,N_1818);
or U5618 (N_5618,N_1888,N_1494);
nand U5619 (N_5619,N_41,N_818);
nor U5620 (N_5620,N_1576,N_140);
xor U5621 (N_5621,N_1759,N_2289);
xor U5622 (N_5622,N_1586,N_2539);
or U5623 (N_5623,N_30,N_1373);
xnor U5624 (N_5624,N_241,N_2481);
nor U5625 (N_5625,N_2878,N_2643);
or U5626 (N_5626,N_2537,N_750);
nor U5627 (N_5627,N_376,N_1525);
nand U5628 (N_5628,N_493,N_2048);
or U5629 (N_5629,N_2551,N_246);
nor U5630 (N_5630,N_1410,N_1880);
and U5631 (N_5631,N_1928,N_623);
xor U5632 (N_5632,N_2382,N_2129);
and U5633 (N_5633,N_2791,N_843);
nand U5634 (N_5634,N_1868,N_814);
nand U5635 (N_5635,N_1402,N_2911);
nor U5636 (N_5636,N_2616,N_2086);
nor U5637 (N_5637,N_2969,N_1045);
or U5638 (N_5638,N_549,N_578);
nand U5639 (N_5639,N_371,N_1015);
xor U5640 (N_5640,N_1314,N_2061);
nand U5641 (N_5641,N_1777,N_1772);
nor U5642 (N_5642,N_2812,N_1127);
nand U5643 (N_5643,N_1167,N_2049);
or U5644 (N_5644,N_2284,N_2053);
nor U5645 (N_5645,N_2572,N_1654);
xnor U5646 (N_5646,N_2802,N_923);
or U5647 (N_5647,N_1257,N_1723);
or U5648 (N_5648,N_1765,N_2450);
nor U5649 (N_5649,N_2152,N_1368);
nor U5650 (N_5650,N_1952,N_530);
and U5651 (N_5651,N_54,N_473);
and U5652 (N_5652,N_2124,N_1139);
and U5653 (N_5653,N_1090,N_549);
or U5654 (N_5654,N_1472,N_2215);
nor U5655 (N_5655,N_1234,N_1635);
xnor U5656 (N_5656,N_1470,N_1729);
nand U5657 (N_5657,N_898,N_1724);
or U5658 (N_5658,N_667,N_2690);
nor U5659 (N_5659,N_330,N_2198);
xnor U5660 (N_5660,N_264,N_1416);
or U5661 (N_5661,N_2416,N_14);
nor U5662 (N_5662,N_1874,N_879);
xnor U5663 (N_5663,N_1232,N_2042);
and U5664 (N_5664,N_1677,N_1789);
and U5665 (N_5665,N_981,N_1654);
xnor U5666 (N_5666,N_821,N_2507);
and U5667 (N_5667,N_1743,N_896);
nand U5668 (N_5668,N_718,N_2342);
nor U5669 (N_5669,N_2469,N_1912);
nand U5670 (N_5670,N_162,N_2885);
nand U5671 (N_5671,N_1709,N_400);
nor U5672 (N_5672,N_247,N_1247);
nor U5673 (N_5673,N_1354,N_1699);
nand U5674 (N_5674,N_2187,N_662);
and U5675 (N_5675,N_2992,N_737);
nor U5676 (N_5676,N_466,N_2845);
nand U5677 (N_5677,N_484,N_375);
and U5678 (N_5678,N_2966,N_2290);
nor U5679 (N_5679,N_2638,N_680);
nand U5680 (N_5680,N_2589,N_1923);
nand U5681 (N_5681,N_2268,N_347);
xnor U5682 (N_5682,N_732,N_1909);
nand U5683 (N_5683,N_958,N_1123);
nor U5684 (N_5684,N_253,N_1361);
and U5685 (N_5685,N_2534,N_2057);
nor U5686 (N_5686,N_2559,N_1289);
nor U5687 (N_5687,N_135,N_724);
nor U5688 (N_5688,N_930,N_2451);
nand U5689 (N_5689,N_1400,N_1848);
and U5690 (N_5690,N_100,N_1710);
nor U5691 (N_5691,N_46,N_564);
nand U5692 (N_5692,N_472,N_388);
or U5693 (N_5693,N_2073,N_2421);
nand U5694 (N_5694,N_270,N_785);
nand U5695 (N_5695,N_1564,N_151);
and U5696 (N_5696,N_1120,N_2610);
nor U5697 (N_5697,N_1902,N_200);
or U5698 (N_5698,N_1129,N_1027);
or U5699 (N_5699,N_1252,N_1199);
nor U5700 (N_5700,N_40,N_483);
or U5701 (N_5701,N_1784,N_1928);
or U5702 (N_5702,N_25,N_975);
and U5703 (N_5703,N_2609,N_645);
or U5704 (N_5704,N_568,N_1339);
or U5705 (N_5705,N_990,N_2311);
nor U5706 (N_5706,N_1247,N_395);
nor U5707 (N_5707,N_999,N_1138);
nand U5708 (N_5708,N_2393,N_1139);
nand U5709 (N_5709,N_2435,N_1193);
nor U5710 (N_5710,N_1170,N_486);
or U5711 (N_5711,N_1872,N_2574);
nand U5712 (N_5712,N_726,N_221);
or U5713 (N_5713,N_595,N_466);
and U5714 (N_5714,N_1044,N_1148);
and U5715 (N_5715,N_2549,N_2373);
and U5716 (N_5716,N_1049,N_570);
nand U5717 (N_5717,N_2100,N_1315);
nor U5718 (N_5718,N_336,N_2189);
nor U5719 (N_5719,N_681,N_836);
or U5720 (N_5720,N_2089,N_182);
nor U5721 (N_5721,N_2076,N_1609);
xnor U5722 (N_5722,N_896,N_643);
nand U5723 (N_5723,N_2660,N_40);
nor U5724 (N_5724,N_2266,N_431);
nand U5725 (N_5725,N_1985,N_903);
nor U5726 (N_5726,N_2795,N_2042);
nand U5727 (N_5727,N_903,N_1030);
or U5728 (N_5728,N_266,N_2967);
and U5729 (N_5729,N_359,N_2441);
xnor U5730 (N_5730,N_2495,N_2685);
nand U5731 (N_5731,N_2285,N_743);
nand U5732 (N_5732,N_1703,N_2615);
nor U5733 (N_5733,N_1485,N_893);
nor U5734 (N_5734,N_574,N_2499);
or U5735 (N_5735,N_2703,N_1852);
and U5736 (N_5736,N_887,N_235);
nand U5737 (N_5737,N_2129,N_760);
nand U5738 (N_5738,N_1676,N_1365);
or U5739 (N_5739,N_977,N_1140);
or U5740 (N_5740,N_2620,N_1436);
and U5741 (N_5741,N_165,N_713);
nand U5742 (N_5742,N_2998,N_445);
xor U5743 (N_5743,N_2468,N_494);
and U5744 (N_5744,N_2568,N_2383);
nor U5745 (N_5745,N_987,N_1801);
nand U5746 (N_5746,N_1467,N_823);
or U5747 (N_5747,N_985,N_223);
nand U5748 (N_5748,N_25,N_1492);
and U5749 (N_5749,N_141,N_2090);
nor U5750 (N_5750,N_1810,N_810);
nor U5751 (N_5751,N_2568,N_266);
nor U5752 (N_5752,N_666,N_544);
nand U5753 (N_5753,N_1537,N_2421);
or U5754 (N_5754,N_866,N_840);
or U5755 (N_5755,N_832,N_188);
nand U5756 (N_5756,N_1990,N_138);
nand U5757 (N_5757,N_1540,N_1552);
and U5758 (N_5758,N_1180,N_2371);
and U5759 (N_5759,N_1788,N_1596);
nand U5760 (N_5760,N_1177,N_1579);
nor U5761 (N_5761,N_2991,N_1484);
nor U5762 (N_5762,N_1850,N_404);
nor U5763 (N_5763,N_473,N_607);
or U5764 (N_5764,N_2353,N_2681);
nand U5765 (N_5765,N_89,N_432);
or U5766 (N_5766,N_1836,N_1391);
or U5767 (N_5767,N_1860,N_2246);
and U5768 (N_5768,N_2510,N_675);
and U5769 (N_5769,N_143,N_2127);
nor U5770 (N_5770,N_2970,N_365);
xnor U5771 (N_5771,N_1473,N_2637);
nor U5772 (N_5772,N_468,N_214);
or U5773 (N_5773,N_2859,N_1083);
and U5774 (N_5774,N_1470,N_620);
or U5775 (N_5775,N_192,N_2373);
nor U5776 (N_5776,N_312,N_2070);
and U5777 (N_5777,N_350,N_1677);
nand U5778 (N_5778,N_2461,N_1672);
nor U5779 (N_5779,N_2359,N_2519);
and U5780 (N_5780,N_2217,N_1522);
nand U5781 (N_5781,N_1362,N_475);
and U5782 (N_5782,N_968,N_2832);
nor U5783 (N_5783,N_810,N_2632);
or U5784 (N_5784,N_2489,N_1578);
and U5785 (N_5785,N_12,N_793);
and U5786 (N_5786,N_2896,N_1514);
or U5787 (N_5787,N_903,N_901);
or U5788 (N_5788,N_913,N_2341);
or U5789 (N_5789,N_2462,N_1874);
nand U5790 (N_5790,N_1757,N_404);
or U5791 (N_5791,N_1060,N_972);
nor U5792 (N_5792,N_1018,N_1713);
xnor U5793 (N_5793,N_1075,N_2304);
or U5794 (N_5794,N_550,N_1941);
and U5795 (N_5795,N_2753,N_2679);
and U5796 (N_5796,N_2646,N_1604);
or U5797 (N_5797,N_164,N_275);
or U5798 (N_5798,N_683,N_392);
nand U5799 (N_5799,N_110,N_2420);
and U5800 (N_5800,N_2444,N_816);
nand U5801 (N_5801,N_997,N_2927);
and U5802 (N_5802,N_1560,N_1299);
nand U5803 (N_5803,N_1203,N_1891);
and U5804 (N_5804,N_1189,N_2555);
xnor U5805 (N_5805,N_777,N_2766);
xor U5806 (N_5806,N_2311,N_2582);
nand U5807 (N_5807,N_688,N_1091);
or U5808 (N_5808,N_1141,N_2373);
or U5809 (N_5809,N_2691,N_16);
nor U5810 (N_5810,N_1154,N_1842);
xnor U5811 (N_5811,N_2645,N_404);
nor U5812 (N_5812,N_2273,N_1675);
nand U5813 (N_5813,N_877,N_470);
or U5814 (N_5814,N_2655,N_2665);
and U5815 (N_5815,N_141,N_2342);
nor U5816 (N_5816,N_672,N_1264);
nand U5817 (N_5817,N_752,N_2236);
and U5818 (N_5818,N_703,N_231);
xnor U5819 (N_5819,N_1036,N_1607);
and U5820 (N_5820,N_2684,N_1228);
nor U5821 (N_5821,N_145,N_2971);
or U5822 (N_5822,N_99,N_687);
xor U5823 (N_5823,N_28,N_2335);
or U5824 (N_5824,N_2051,N_2310);
xnor U5825 (N_5825,N_2596,N_1106);
or U5826 (N_5826,N_2296,N_2532);
nand U5827 (N_5827,N_1850,N_2049);
or U5828 (N_5828,N_1418,N_1207);
or U5829 (N_5829,N_1224,N_2180);
and U5830 (N_5830,N_2269,N_2563);
or U5831 (N_5831,N_2820,N_1242);
and U5832 (N_5832,N_1138,N_2721);
xnor U5833 (N_5833,N_896,N_884);
and U5834 (N_5834,N_1546,N_2702);
and U5835 (N_5835,N_2787,N_2581);
or U5836 (N_5836,N_117,N_1060);
nand U5837 (N_5837,N_1828,N_568);
or U5838 (N_5838,N_950,N_2520);
and U5839 (N_5839,N_2977,N_1455);
nor U5840 (N_5840,N_610,N_2911);
nand U5841 (N_5841,N_2250,N_476);
nor U5842 (N_5842,N_1014,N_1207);
or U5843 (N_5843,N_1325,N_1095);
and U5844 (N_5844,N_292,N_195);
nand U5845 (N_5845,N_2849,N_1725);
and U5846 (N_5846,N_542,N_747);
and U5847 (N_5847,N_2700,N_759);
and U5848 (N_5848,N_984,N_660);
nand U5849 (N_5849,N_2029,N_2979);
nand U5850 (N_5850,N_2010,N_582);
or U5851 (N_5851,N_818,N_1570);
and U5852 (N_5852,N_1020,N_2286);
or U5853 (N_5853,N_1195,N_1730);
and U5854 (N_5854,N_1980,N_2777);
nand U5855 (N_5855,N_1541,N_1795);
or U5856 (N_5856,N_1034,N_1335);
nor U5857 (N_5857,N_2888,N_1704);
or U5858 (N_5858,N_949,N_2918);
and U5859 (N_5859,N_2193,N_2137);
and U5860 (N_5860,N_2635,N_1680);
nand U5861 (N_5861,N_1501,N_2245);
nor U5862 (N_5862,N_1829,N_2100);
nor U5863 (N_5863,N_1518,N_2297);
nor U5864 (N_5864,N_2512,N_167);
or U5865 (N_5865,N_1504,N_1376);
and U5866 (N_5866,N_49,N_2365);
or U5867 (N_5867,N_2665,N_926);
nand U5868 (N_5868,N_1930,N_1138);
nor U5869 (N_5869,N_800,N_1861);
and U5870 (N_5870,N_1505,N_2318);
nand U5871 (N_5871,N_1303,N_905);
or U5872 (N_5872,N_527,N_756);
or U5873 (N_5873,N_422,N_2425);
nor U5874 (N_5874,N_1499,N_2163);
nand U5875 (N_5875,N_2635,N_432);
nor U5876 (N_5876,N_2787,N_1697);
and U5877 (N_5877,N_257,N_2854);
or U5878 (N_5878,N_935,N_1506);
nand U5879 (N_5879,N_1249,N_1866);
and U5880 (N_5880,N_1574,N_1815);
xnor U5881 (N_5881,N_541,N_2938);
or U5882 (N_5882,N_2594,N_2117);
and U5883 (N_5883,N_1055,N_1304);
or U5884 (N_5884,N_212,N_2424);
or U5885 (N_5885,N_890,N_1776);
and U5886 (N_5886,N_82,N_277);
nand U5887 (N_5887,N_2285,N_1688);
nand U5888 (N_5888,N_2058,N_2844);
or U5889 (N_5889,N_1767,N_2475);
nand U5890 (N_5890,N_215,N_403);
or U5891 (N_5891,N_2277,N_2971);
nand U5892 (N_5892,N_2127,N_952);
nand U5893 (N_5893,N_956,N_339);
nand U5894 (N_5894,N_2790,N_1299);
or U5895 (N_5895,N_294,N_723);
and U5896 (N_5896,N_2508,N_2771);
and U5897 (N_5897,N_1026,N_991);
or U5898 (N_5898,N_1126,N_134);
nor U5899 (N_5899,N_671,N_824);
and U5900 (N_5900,N_1655,N_1037);
or U5901 (N_5901,N_2060,N_2305);
nand U5902 (N_5902,N_1505,N_1850);
and U5903 (N_5903,N_1707,N_719);
or U5904 (N_5904,N_2832,N_2661);
nand U5905 (N_5905,N_1103,N_422);
xor U5906 (N_5906,N_942,N_127);
nor U5907 (N_5907,N_1801,N_1011);
nor U5908 (N_5908,N_666,N_502);
xor U5909 (N_5909,N_2809,N_1199);
nand U5910 (N_5910,N_1339,N_1746);
nand U5911 (N_5911,N_199,N_1869);
xor U5912 (N_5912,N_2969,N_2170);
nor U5913 (N_5913,N_804,N_879);
nand U5914 (N_5914,N_2507,N_2513);
xnor U5915 (N_5915,N_1071,N_782);
nand U5916 (N_5916,N_517,N_841);
xnor U5917 (N_5917,N_1206,N_2563);
or U5918 (N_5918,N_1593,N_15);
or U5919 (N_5919,N_1479,N_196);
or U5920 (N_5920,N_2912,N_1474);
and U5921 (N_5921,N_464,N_1289);
nand U5922 (N_5922,N_224,N_354);
and U5923 (N_5923,N_2040,N_2286);
or U5924 (N_5924,N_2408,N_106);
and U5925 (N_5925,N_2390,N_1858);
nor U5926 (N_5926,N_669,N_1574);
xor U5927 (N_5927,N_2553,N_310);
xor U5928 (N_5928,N_1817,N_2895);
nand U5929 (N_5929,N_394,N_250);
nand U5930 (N_5930,N_1112,N_589);
or U5931 (N_5931,N_538,N_735);
or U5932 (N_5932,N_365,N_2154);
nand U5933 (N_5933,N_310,N_1046);
nand U5934 (N_5934,N_986,N_1059);
or U5935 (N_5935,N_841,N_2389);
xnor U5936 (N_5936,N_2591,N_1809);
or U5937 (N_5937,N_2599,N_979);
nor U5938 (N_5938,N_936,N_1426);
nand U5939 (N_5939,N_2411,N_745);
nand U5940 (N_5940,N_183,N_659);
nor U5941 (N_5941,N_1993,N_1382);
and U5942 (N_5942,N_197,N_1157);
nand U5943 (N_5943,N_2707,N_954);
or U5944 (N_5944,N_911,N_2660);
nand U5945 (N_5945,N_852,N_1400);
nand U5946 (N_5946,N_2446,N_1857);
nor U5947 (N_5947,N_1558,N_279);
xor U5948 (N_5948,N_125,N_19);
nor U5949 (N_5949,N_1462,N_282);
nand U5950 (N_5950,N_784,N_2549);
nand U5951 (N_5951,N_932,N_1563);
or U5952 (N_5952,N_2721,N_2589);
or U5953 (N_5953,N_1122,N_1722);
and U5954 (N_5954,N_733,N_988);
nand U5955 (N_5955,N_761,N_570);
nor U5956 (N_5956,N_2571,N_540);
nand U5957 (N_5957,N_344,N_1943);
xor U5958 (N_5958,N_2000,N_742);
nor U5959 (N_5959,N_990,N_43);
and U5960 (N_5960,N_2939,N_2933);
and U5961 (N_5961,N_1621,N_268);
nor U5962 (N_5962,N_339,N_2260);
and U5963 (N_5963,N_543,N_2505);
and U5964 (N_5964,N_1777,N_415);
and U5965 (N_5965,N_1530,N_1480);
and U5966 (N_5966,N_2448,N_1384);
nand U5967 (N_5967,N_2422,N_527);
and U5968 (N_5968,N_234,N_1583);
nor U5969 (N_5969,N_188,N_957);
nand U5970 (N_5970,N_643,N_2478);
nor U5971 (N_5971,N_1250,N_2647);
and U5972 (N_5972,N_2916,N_2109);
and U5973 (N_5973,N_1671,N_2018);
nor U5974 (N_5974,N_690,N_696);
and U5975 (N_5975,N_909,N_198);
nand U5976 (N_5976,N_1843,N_2797);
nor U5977 (N_5977,N_2902,N_2555);
nand U5978 (N_5978,N_1648,N_372);
nor U5979 (N_5979,N_1931,N_1209);
or U5980 (N_5980,N_256,N_1481);
and U5981 (N_5981,N_2918,N_308);
nand U5982 (N_5982,N_1617,N_925);
and U5983 (N_5983,N_1852,N_2917);
nor U5984 (N_5984,N_1671,N_1486);
or U5985 (N_5985,N_188,N_2473);
nand U5986 (N_5986,N_158,N_1813);
and U5987 (N_5987,N_2394,N_1363);
and U5988 (N_5988,N_442,N_1189);
nand U5989 (N_5989,N_550,N_2002);
nor U5990 (N_5990,N_2109,N_1897);
or U5991 (N_5991,N_767,N_25);
and U5992 (N_5992,N_2563,N_40);
nor U5993 (N_5993,N_2942,N_2223);
nor U5994 (N_5994,N_1710,N_1255);
or U5995 (N_5995,N_964,N_2510);
nand U5996 (N_5996,N_2857,N_126);
nand U5997 (N_5997,N_2790,N_1677);
nor U5998 (N_5998,N_718,N_2927);
xnor U5999 (N_5999,N_2375,N_2806);
and U6000 (N_6000,N_3810,N_4474);
or U6001 (N_6001,N_3583,N_5028);
and U6002 (N_6002,N_5523,N_5215);
nand U6003 (N_6003,N_5204,N_5533);
or U6004 (N_6004,N_4224,N_4262);
or U6005 (N_6005,N_3112,N_5192);
nand U6006 (N_6006,N_5304,N_4562);
or U6007 (N_6007,N_5267,N_5394);
or U6008 (N_6008,N_4628,N_4795);
nor U6009 (N_6009,N_4433,N_4554);
nand U6010 (N_6010,N_5881,N_3631);
or U6011 (N_6011,N_5236,N_3005);
and U6012 (N_6012,N_5769,N_5067);
and U6013 (N_6013,N_4134,N_5144);
nor U6014 (N_6014,N_3272,N_5126);
nor U6015 (N_6015,N_5366,N_4201);
and U6016 (N_6016,N_3694,N_4106);
nor U6017 (N_6017,N_4338,N_3687);
and U6018 (N_6018,N_3813,N_3315);
or U6019 (N_6019,N_4049,N_5805);
nand U6020 (N_6020,N_5275,N_3513);
nor U6021 (N_6021,N_4571,N_4863);
or U6022 (N_6022,N_3178,N_4990);
nand U6023 (N_6023,N_3650,N_5337);
or U6024 (N_6024,N_5750,N_3353);
and U6025 (N_6025,N_3267,N_3461);
xor U6026 (N_6026,N_4001,N_3798);
nand U6027 (N_6027,N_4721,N_3531);
and U6028 (N_6028,N_4384,N_4075);
and U6029 (N_6029,N_3479,N_4036);
nor U6030 (N_6030,N_5602,N_5447);
nand U6031 (N_6031,N_3724,N_4889);
nor U6032 (N_6032,N_5690,N_5564);
nand U6033 (N_6033,N_4362,N_5214);
nand U6034 (N_6034,N_3812,N_5831);
nor U6035 (N_6035,N_3638,N_3447);
or U6036 (N_6036,N_3982,N_4765);
nand U6037 (N_6037,N_3301,N_3207);
and U6038 (N_6038,N_5980,N_4963);
and U6039 (N_6039,N_5520,N_5677);
or U6040 (N_6040,N_4725,N_4425);
nor U6041 (N_6041,N_3264,N_4417);
nand U6042 (N_6042,N_5694,N_4724);
or U6043 (N_6043,N_3254,N_4412);
and U6044 (N_6044,N_4938,N_5551);
nand U6045 (N_6045,N_3951,N_3708);
nor U6046 (N_6046,N_3168,N_3403);
nand U6047 (N_6047,N_4778,N_3457);
nand U6048 (N_6048,N_4408,N_5614);
or U6049 (N_6049,N_3079,N_5092);
or U6050 (N_6050,N_3374,N_4824);
or U6051 (N_6051,N_3892,N_3429);
or U6052 (N_6052,N_3743,N_5175);
and U6053 (N_6053,N_3700,N_3030);
and U6054 (N_6054,N_5473,N_3647);
nand U6055 (N_6055,N_4798,N_5790);
or U6056 (N_6056,N_5024,N_3197);
or U6057 (N_6057,N_5507,N_5591);
nor U6058 (N_6058,N_5847,N_4089);
nand U6059 (N_6059,N_3815,N_4306);
or U6060 (N_6060,N_5370,N_4897);
and U6061 (N_6061,N_5432,N_4916);
and U6062 (N_6062,N_4368,N_5912);
nand U6063 (N_6063,N_4861,N_5997);
nor U6064 (N_6064,N_4788,N_4299);
and U6065 (N_6065,N_3418,N_4665);
nand U6066 (N_6066,N_5829,N_3009);
nor U6067 (N_6067,N_5102,N_3794);
nand U6068 (N_6068,N_3472,N_4409);
nor U6069 (N_6069,N_5451,N_5163);
nand U6070 (N_6070,N_4991,N_4742);
or U6071 (N_6071,N_4928,N_5334);
and U6072 (N_6072,N_3099,N_5566);
and U6073 (N_6073,N_3397,N_4222);
xor U6074 (N_6074,N_3507,N_5240);
nor U6075 (N_6075,N_4213,N_4214);
or U6076 (N_6076,N_5177,N_3784);
or U6077 (N_6077,N_3714,N_3106);
nor U6078 (N_6078,N_4559,N_5048);
nand U6079 (N_6079,N_5587,N_5721);
and U6080 (N_6080,N_4260,N_4290);
and U6081 (N_6081,N_4553,N_5408);
and U6082 (N_6082,N_4206,N_5913);
nand U6083 (N_6083,N_5804,N_3808);
nor U6084 (N_6084,N_3801,N_5521);
nand U6085 (N_6085,N_5524,N_3899);
or U6086 (N_6086,N_4601,N_5436);
or U6087 (N_6087,N_3477,N_4052);
and U6088 (N_6088,N_3059,N_3963);
or U6089 (N_6089,N_5468,N_3114);
and U6090 (N_6090,N_4870,N_5395);
nand U6091 (N_6091,N_5181,N_5187);
or U6092 (N_6092,N_3485,N_3535);
nor U6093 (N_6093,N_4613,N_5885);
xnor U6094 (N_6094,N_5469,N_5426);
and U6095 (N_6095,N_4178,N_5570);
and U6096 (N_6096,N_3887,N_5379);
nand U6097 (N_6097,N_3764,N_3920);
nand U6098 (N_6098,N_5149,N_5630);
or U6099 (N_6099,N_5044,N_4387);
nand U6100 (N_6100,N_5556,N_3065);
and U6101 (N_6101,N_4495,N_3048);
nand U6102 (N_6102,N_4268,N_4173);
nand U6103 (N_6103,N_3719,N_5316);
and U6104 (N_6104,N_4239,N_3824);
and U6105 (N_6105,N_5397,N_5617);
nand U6106 (N_6106,N_4092,N_4492);
nor U6107 (N_6107,N_5380,N_5061);
nor U6108 (N_6108,N_3837,N_3475);
nand U6109 (N_6109,N_4083,N_5688);
nand U6110 (N_6110,N_3860,N_3672);
or U6111 (N_6111,N_3186,N_5327);
nor U6112 (N_6112,N_5069,N_3959);
xnor U6113 (N_6113,N_3536,N_3143);
nor U6114 (N_6114,N_3589,N_4681);
and U6115 (N_6115,N_3659,N_5902);
nor U6116 (N_6116,N_5990,N_3234);
or U6117 (N_6117,N_5388,N_3093);
nand U6118 (N_6118,N_5534,N_5080);
xnor U6119 (N_6119,N_4316,N_5223);
and U6120 (N_6120,N_3149,N_5216);
or U6121 (N_6121,N_5697,N_3710);
and U6122 (N_6122,N_5636,N_4398);
nor U6123 (N_6123,N_4662,N_3725);
nor U6124 (N_6124,N_5445,N_3966);
nand U6125 (N_6125,N_4920,N_5441);
nor U6126 (N_6126,N_4834,N_5384);
nor U6127 (N_6127,N_5031,N_3242);
nand U6128 (N_6128,N_5479,N_5708);
nor U6129 (N_6129,N_5935,N_4403);
and U6130 (N_6130,N_5001,N_4210);
nand U6131 (N_6131,N_5577,N_3929);
xor U6132 (N_6132,N_5233,N_4586);
nand U6133 (N_6133,N_3804,N_5908);
xnor U6134 (N_6134,N_3741,N_4892);
nor U6135 (N_6135,N_5243,N_5017);
nand U6136 (N_6136,N_4321,N_5284);
and U6137 (N_6137,N_5321,N_3739);
and U6138 (N_6138,N_4568,N_3590);
nand U6139 (N_6139,N_4658,N_3407);
nand U6140 (N_6140,N_4774,N_5153);
and U6141 (N_6141,N_3751,N_4097);
and U6142 (N_6142,N_5136,N_4955);
and U6143 (N_6143,N_4564,N_4978);
and U6144 (N_6144,N_5221,N_4718);
nand U6145 (N_6145,N_3709,N_3574);
nand U6146 (N_6146,N_5869,N_3451);
and U6147 (N_6147,N_4904,N_5903);
nor U6148 (N_6148,N_5907,N_5484);
nand U6149 (N_6149,N_5002,N_5797);
and U6150 (N_6150,N_3555,N_3426);
nand U6151 (N_6151,N_3282,N_3597);
and U6152 (N_6152,N_3104,N_4779);
and U6153 (N_6153,N_5856,N_3593);
and U6154 (N_6154,N_3090,N_3329);
and U6155 (N_6155,N_5817,N_5665);
nor U6156 (N_6156,N_4069,N_5634);
and U6157 (N_6157,N_5825,N_4740);
nor U6158 (N_6158,N_5383,N_5867);
or U6159 (N_6159,N_3934,N_4827);
nand U6160 (N_6160,N_4274,N_3139);
and U6161 (N_6161,N_4982,N_4814);
xnor U6162 (N_6162,N_5578,N_5363);
and U6163 (N_6163,N_4701,N_4256);
and U6164 (N_6164,N_3303,N_4805);
nand U6165 (N_6165,N_3493,N_3399);
or U6166 (N_6166,N_5607,N_4790);
nand U6167 (N_6167,N_3690,N_5117);
nor U6168 (N_6168,N_4657,N_5501);
and U6169 (N_6169,N_3446,N_5405);
and U6170 (N_6170,N_4062,N_3110);
or U6171 (N_6171,N_4797,N_5631);
nor U6172 (N_6172,N_5234,N_3086);
nand U6173 (N_6173,N_3692,N_3545);
and U6174 (N_6174,N_3428,N_3806);
and U6175 (N_6175,N_3842,N_5411);
or U6176 (N_6176,N_5763,N_5495);
nor U6177 (N_6177,N_5043,N_3533);
nand U6178 (N_6178,N_4843,N_3703);
or U6179 (N_6179,N_4249,N_3733);
nand U6180 (N_6180,N_4741,N_4782);
xor U6181 (N_6181,N_4190,N_3134);
xor U6182 (N_6182,N_4308,N_3338);
nand U6183 (N_6183,N_5116,N_4633);
nor U6184 (N_6184,N_5344,N_5088);
nand U6185 (N_6185,N_5399,N_4828);
nor U6186 (N_6186,N_3828,N_5960);
nor U6187 (N_6187,N_4370,N_3420);
nor U6188 (N_6188,N_4703,N_3283);
or U6189 (N_6189,N_3623,N_3877);
xnor U6190 (N_6190,N_3989,N_5816);
xor U6191 (N_6191,N_5669,N_4102);
or U6192 (N_6192,N_3482,N_5716);
xor U6193 (N_6193,N_3383,N_3003);
or U6194 (N_6194,N_3586,N_4737);
nand U6195 (N_6195,N_3787,N_3939);
or U6196 (N_6196,N_4654,N_5986);
and U6197 (N_6197,N_3408,N_3393);
or U6198 (N_6198,N_4896,N_4046);
nor U6199 (N_6199,N_3381,N_5936);
and U6200 (N_6200,N_3715,N_5349);
nor U6201 (N_6201,N_3871,N_3746);
nand U6202 (N_6202,N_3101,N_3384);
nor U6203 (N_6203,N_4612,N_4549);
and U6204 (N_6204,N_4527,N_5278);
nor U6205 (N_6205,N_3083,N_3632);
xnor U6206 (N_6206,N_5004,N_3067);
nand U6207 (N_6207,N_5815,N_5416);
nor U6208 (N_6208,N_3246,N_5844);
nand U6209 (N_6209,N_5635,N_4029);
nor U6210 (N_6210,N_3553,N_3052);
nor U6211 (N_6211,N_5619,N_4195);
nand U6212 (N_6212,N_4873,N_3753);
xnor U6213 (N_6213,N_3612,N_5073);
and U6214 (N_6214,N_5406,N_5325);
nor U6215 (N_6215,N_4819,N_4915);
nor U6216 (N_6216,N_4357,N_5212);
nand U6217 (N_6217,N_4627,N_3859);
nor U6218 (N_6218,N_5466,N_4908);
or U6219 (N_6219,N_4063,N_4161);
nor U6220 (N_6220,N_4678,N_3732);
nand U6221 (N_6221,N_5667,N_4676);
nand U6222 (N_6222,N_3167,N_5282);
or U6223 (N_6223,N_5601,N_5542);
nand U6224 (N_6224,N_5417,N_3915);
and U6225 (N_6225,N_4526,N_5306);
nand U6226 (N_6226,N_3085,N_3833);
xor U6227 (N_6227,N_3095,N_3102);
or U6228 (N_6228,N_4674,N_5746);
or U6229 (N_6229,N_5323,N_3772);
nand U6230 (N_6230,N_5717,N_5803);
nor U6231 (N_6231,N_4958,N_4642);
and U6232 (N_6232,N_3161,N_3922);
nor U6233 (N_6233,N_3268,N_3789);
nand U6234 (N_6234,N_5637,N_5165);
or U6235 (N_6235,N_4793,N_3941);
or U6236 (N_6236,N_5166,N_5753);
nor U6237 (N_6237,N_4380,N_5748);
or U6238 (N_6238,N_5703,N_4269);
and U6239 (N_6239,N_4525,N_3174);
or U6240 (N_6240,N_5606,N_3988);
nand U6241 (N_6241,N_4539,N_4939);
and U6242 (N_6242,N_4242,N_4661);
and U6243 (N_6243,N_3195,N_4739);
nor U6244 (N_6244,N_3856,N_4248);
and U6245 (N_6245,N_5013,N_3500);
or U6246 (N_6246,N_5872,N_5821);
and U6247 (N_6247,N_3217,N_4589);
nand U6248 (N_6248,N_4135,N_3904);
and U6249 (N_6249,N_4883,N_3498);
nor U6250 (N_6250,N_5588,N_4961);
nor U6251 (N_6251,N_5120,N_3550);
and U6252 (N_6252,N_4111,N_5218);
nand U6253 (N_6253,N_4405,N_5164);
or U6254 (N_6254,N_5137,N_4365);
xor U6255 (N_6255,N_4512,N_4708);
xnor U6256 (N_6256,N_3441,N_4026);
xor U6257 (N_6257,N_4085,N_3109);
nand U6258 (N_6258,N_5288,N_5329);
or U6259 (N_6259,N_3296,N_5303);
xnor U6260 (N_6260,N_5442,N_5579);
xor U6261 (N_6261,N_4881,N_4126);
nand U6262 (N_6262,N_3999,N_4020);
nand U6263 (N_6263,N_3449,N_4530);
nand U6264 (N_6264,N_3280,N_5726);
nor U6265 (N_6265,N_3544,N_3861);
and U6266 (N_6266,N_4878,N_4257);
or U6267 (N_6267,N_3519,N_3524);
or U6268 (N_6268,N_4558,N_4022);
xnor U6269 (N_6269,N_5193,N_3832);
and U6270 (N_6270,N_3950,N_4451);
nor U6271 (N_6271,N_4054,N_5128);
or U6272 (N_6272,N_3644,N_4537);
nand U6273 (N_6273,N_4070,N_3678);
or U6274 (N_6274,N_5851,N_5747);
nor U6275 (N_6275,N_5706,N_5318);
nand U6276 (N_6276,N_4643,N_4799);
xor U6277 (N_6277,N_5202,N_4670);
and U6278 (N_6278,N_5308,N_4098);
nor U6279 (N_6279,N_3907,N_3117);
or U6280 (N_6280,N_4127,N_4108);
nand U6281 (N_6281,N_4951,N_3598);
or U6282 (N_6282,N_3335,N_5265);
and U6283 (N_6283,N_5951,N_4956);
nor U6284 (N_6284,N_5826,N_4597);
nand U6285 (N_6285,N_5958,N_4595);
nand U6286 (N_6286,N_3229,N_4479);
or U6287 (N_6287,N_5527,N_3115);
and U6288 (N_6288,N_4902,N_4501);
nand U6289 (N_6289,N_5553,N_5955);
or U6290 (N_6290,N_5709,N_5921);
or U6291 (N_6291,N_5889,N_3875);
or U6292 (N_6292,N_5194,N_3967);
or U6293 (N_6293,N_3554,N_4686);
nand U6294 (N_6294,N_5108,N_3184);
xnor U6295 (N_6295,N_3573,N_3113);
nor U6296 (N_6296,N_5271,N_3413);
nor U6297 (N_6297,N_5970,N_3294);
nand U6298 (N_6298,N_5324,N_3629);
nand U6299 (N_6299,N_3034,N_5361);
nor U6300 (N_6300,N_4952,N_5727);
or U6301 (N_6301,N_5387,N_4252);
xor U6302 (N_6302,N_4270,N_4569);
nand U6303 (N_6303,N_3853,N_5155);
nor U6304 (N_6304,N_4682,N_3776);
and U6305 (N_6305,N_4728,N_4519);
and U6306 (N_6306,N_4509,N_3993);
and U6307 (N_6307,N_4906,N_5414);
nand U6308 (N_6308,N_4552,N_4604);
and U6309 (N_6309,N_5857,N_4281);
xor U6310 (N_6310,N_5899,N_5824);
nor U6311 (N_6311,N_5609,N_5160);
and U6312 (N_6312,N_3570,N_5643);
or U6313 (N_6313,N_3293,N_3673);
nor U6314 (N_6314,N_3504,N_5326);
nand U6315 (N_6315,N_4692,N_4780);
xnor U6316 (N_6316,N_4862,N_5161);
nor U6317 (N_6317,N_5298,N_3525);
or U6318 (N_6318,N_3033,N_5828);
nand U6319 (N_6319,N_3701,N_4051);
and U6320 (N_6320,N_3865,N_4748);
and U6321 (N_6321,N_3394,N_3767);
or U6322 (N_6322,N_4375,N_4444);
or U6323 (N_6323,N_5819,N_4716);
and U6324 (N_6324,N_5691,N_3088);
and U6325 (N_6325,N_3474,N_3971);
or U6326 (N_6326,N_5622,N_4940);
nor U6327 (N_6327,N_3058,N_5478);
or U6328 (N_6328,N_3225,N_3809);
nand U6329 (N_6329,N_5532,N_3818);
nand U6330 (N_6330,N_5084,N_3285);
and U6331 (N_6331,N_5079,N_4985);
nor U6332 (N_6332,N_3416,N_4261);
nand U6333 (N_6333,N_5294,N_5794);
and U6334 (N_6334,N_4023,N_3992);
and U6335 (N_6335,N_3721,N_4844);
and U6336 (N_6336,N_3863,N_5754);
nor U6337 (N_6337,N_4067,N_4285);
and U6338 (N_6338,N_3157,N_3170);
xor U6339 (N_6339,N_4599,N_5793);
nand U6340 (N_6340,N_4304,N_4998);
nor U6341 (N_6341,N_4557,N_5528);
and U6342 (N_6342,N_3923,N_4124);
and U6343 (N_6343,N_3062,N_3556);
and U6344 (N_6344,N_3082,N_5890);
xor U6345 (N_6345,N_3053,N_3193);
and U6346 (N_6346,N_5642,N_5232);
or U6347 (N_6347,N_3541,N_4399);
nand U6348 (N_6348,N_5771,N_4867);
and U6349 (N_6349,N_3938,N_3452);
nor U6350 (N_6350,N_4625,N_4719);
nor U6351 (N_6351,N_5046,N_3945);
or U6352 (N_6352,N_3979,N_3502);
nand U6353 (N_6353,N_4523,N_3046);
nand U6354 (N_6354,N_4091,N_4473);
or U6355 (N_6355,N_4651,N_3518);
and U6356 (N_6356,N_3903,N_4443);
nor U6357 (N_6357,N_5206,N_5015);
nor U6358 (N_6358,N_3440,N_3857);
and U6359 (N_6359,N_4969,N_5977);
nor U6360 (N_6360,N_4637,N_3406);
or U6361 (N_6361,N_4645,N_4540);
nor U6362 (N_6362,N_5320,N_5742);
nor U6363 (N_6363,N_4033,N_5229);
nand U6364 (N_6364,N_5672,N_5503);
nand U6365 (N_6365,N_3654,N_5608);
nor U6366 (N_6366,N_5456,N_4061);
and U6367 (N_6367,N_3037,N_3747);
nor U6368 (N_6368,N_4855,N_5254);
or U6369 (N_6369,N_5693,N_5178);
nor U6370 (N_6370,N_5089,N_4872);
and U6371 (N_6371,N_3284,N_3497);
and U6372 (N_6372,N_4228,N_3649);
nor U6373 (N_6373,N_4730,N_5180);
nand U6374 (N_6374,N_5376,N_5281);
and U6375 (N_6375,N_4406,N_5262);
nand U6376 (N_6376,N_4818,N_4112);
xnor U6377 (N_6377,N_3147,N_3377);
or U6378 (N_6378,N_4141,N_4264);
and U6379 (N_6379,N_4864,N_3445);
and U6380 (N_6380,N_5719,N_4917);
or U6381 (N_6381,N_3491,N_3879);
or U6382 (N_6382,N_5791,N_3022);
or U6383 (N_6383,N_5250,N_5685);
nand U6384 (N_6384,N_3470,N_5778);
or U6385 (N_6385,N_5841,N_3214);
xor U6386 (N_6386,N_5743,N_4008);
or U6387 (N_6387,N_5858,N_3239);
and U6388 (N_6388,N_4749,N_3918);
nand U6389 (N_6389,N_5745,N_5657);
or U6390 (N_6390,N_3852,N_3674);
nor U6391 (N_6391,N_4673,N_3713);
nor U6392 (N_6392,N_4310,N_4900);
nor U6393 (N_6393,N_4103,N_5260);
or U6394 (N_6394,N_5560,N_4416);
and U6395 (N_6395,N_3218,N_4690);
nand U6396 (N_6396,N_5603,N_5652);
nor U6397 (N_6397,N_5513,N_5953);
or U6398 (N_6398,N_3409,N_5530);
nand U6399 (N_6399,N_4047,N_3858);
xnor U6400 (N_6400,N_4689,N_5973);
nand U6401 (N_6401,N_5345,N_3237);
nand U6402 (N_6402,N_3306,N_4305);
xor U6403 (N_6403,N_3961,N_3780);
and U6404 (N_6404,N_5364,N_5139);
nand U6405 (N_6405,N_5335,N_3205);
xnor U6406 (N_6406,N_4731,N_5488);
nor U6407 (N_6407,N_4351,N_3360);
nand U6408 (N_6408,N_5241,N_3671);
nand U6409 (N_6409,N_3466,N_5944);
and U6410 (N_6410,N_3323,N_3213);
or U6411 (N_6411,N_4396,N_3969);
and U6412 (N_6412,N_5425,N_5809);
nand U6413 (N_6413,N_4429,N_4456);
nand U6414 (N_6414,N_5845,N_3578);
nor U6415 (N_6415,N_5836,N_4079);
nor U6416 (N_6416,N_3089,N_4954);
and U6417 (N_6417,N_4837,N_3805);
and U6418 (N_6418,N_5531,N_5252);
nor U6419 (N_6419,N_4194,N_4042);
nor U6420 (N_6420,N_4439,N_5396);
and U6421 (N_6421,N_5620,N_4932);
nand U6422 (N_6422,N_3116,N_5550);
nand U6423 (N_6423,N_4332,N_3092);
and U6424 (N_6424,N_3027,N_3069);
and U6425 (N_6425,N_4803,N_5839);
or U6426 (N_6426,N_3434,N_5276);
nor U6427 (N_6427,N_5700,N_4496);
and U6428 (N_6428,N_4747,N_5317);
or U6429 (N_6429,N_5732,N_3811);
xnor U6430 (N_6430,N_3585,N_3221);
and U6431 (N_6431,N_3361,N_4469);
nor U6432 (N_6432,N_3001,N_4197);
xor U6433 (N_6433,N_4435,N_4055);
xor U6434 (N_6434,N_5033,N_3995);
or U6435 (N_6435,N_4346,N_3252);
or U6436 (N_6436,N_5993,N_3224);
nor U6437 (N_6437,N_5768,N_5401);
or U6438 (N_6438,N_3888,N_3984);
nand U6439 (N_6439,N_3977,N_3476);
nor U6440 (N_6440,N_5471,N_4838);
xor U6441 (N_6441,N_5348,N_3896);
or U6442 (N_6442,N_5744,N_5535);
or U6443 (N_6443,N_4034,N_5076);
or U6444 (N_6444,N_3281,N_3921);
or U6445 (N_6445,N_3681,N_5115);
nor U6446 (N_6446,N_5689,N_4971);
nand U6447 (N_6447,N_3129,N_3869);
nor U6448 (N_6448,N_4572,N_3722);
xnor U6449 (N_6449,N_3595,N_4813);
or U6450 (N_6450,N_3362,N_4983);
nand U6451 (N_6451,N_4035,N_3260);
nand U6452 (N_6452,N_5684,N_5118);
nor U6453 (N_6453,N_4183,N_3777);
and U6454 (N_6454,N_4841,N_4039);
and U6455 (N_6455,N_3799,N_3177);
nand U6456 (N_6456,N_3473,N_5671);
or U6457 (N_6457,N_3287,N_5151);
nand U6458 (N_6458,N_3210,N_5998);
and U6459 (N_6459,N_3986,N_3564);
nor U6460 (N_6460,N_4964,N_3825);
nand U6461 (N_6461,N_4136,N_4221);
and U6462 (N_6462,N_3230,N_4484);
nor U6463 (N_6463,N_5755,N_3571);
and U6464 (N_6464,N_3797,N_3501);
and U6465 (N_6465,N_5248,N_3467);
nor U6466 (N_6466,N_4723,N_3685);
nor U6467 (N_6467,N_4936,N_4041);
nand U6468 (N_6468,N_4354,N_4358);
or U6469 (N_6469,N_3094,N_3508);
or U6470 (N_6470,N_3049,N_5975);
or U6471 (N_6471,N_3289,N_5592);
or U6472 (N_6472,N_3744,N_4415);
and U6473 (N_6473,N_4198,N_5461);
and U6474 (N_6474,N_3146,N_5311);
and U6475 (N_6475,N_5779,N_4428);
nand U6476 (N_6476,N_5292,N_5668);
and U6477 (N_6477,N_5525,N_5492);
nor U6478 (N_6478,N_4717,N_4073);
xnor U6479 (N_6479,N_3270,N_3054);
xor U6480 (N_6480,N_5597,N_4411);
and U6481 (N_6481,N_3130,N_3854);
nand U6482 (N_6482,N_4542,N_3738);
nor U6483 (N_6483,N_3697,N_5096);
xnor U6484 (N_6484,N_5367,N_4199);
nand U6485 (N_6485,N_5259,N_3346);
and U6486 (N_6486,N_3304,N_3873);
or U6487 (N_6487,N_4816,N_3641);
nor U6488 (N_6488,N_4736,N_4935);
and U6489 (N_6489,N_3762,N_3581);
or U6490 (N_6490,N_3412,N_3994);
nor U6491 (N_6491,N_5185,N_4436);
nand U6492 (N_6492,N_5059,N_3081);
nand U6493 (N_6493,N_3019,N_3734);
and U6494 (N_6494,N_4082,N_3886);
nor U6495 (N_6495,N_5083,N_5111);
and U6496 (N_6496,N_5230,N_4850);
nor U6497 (N_6497,N_3509,N_3029);
nor U6498 (N_6498,N_4187,N_4040);
and U6499 (N_6499,N_4158,N_4060);
and U6500 (N_6500,N_3665,N_5511);
nand U6501 (N_6501,N_4447,N_5526);
nand U6502 (N_6502,N_5100,N_4133);
nand U6503 (N_6503,N_5658,N_5095);
or U6504 (N_6504,N_5598,N_5571);
and U6505 (N_6505,N_4705,N_3070);
or U6506 (N_6506,N_4154,N_4327);
nor U6507 (N_6507,N_5911,N_3791);
or U6508 (N_6508,N_5720,N_5981);
and U6509 (N_6509,N_4699,N_5453);
nor U6510 (N_6510,N_5464,N_3220);
or U6511 (N_6511,N_5751,N_4675);
nand U6512 (N_6512,N_3582,N_3996);
nor U6513 (N_6513,N_4390,N_5315);
and U6514 (N_6514,N_3495,N_5782);
nand U6515 (N_6515,N_3868,N_3527);
or U6516 (N_6516,N_4857,N_4996);
and U6517 (N_6517,N_3368,N_5737);
and U6518 (N_6518,N_4929,N_3552);
and U6519 (N_6519,N_3247,N_4829);
nor U6520 (N_6520,N_3579,N_4566);
nor U6521 (N_6521,N_4648,N_4267);
and U6522 (N_6522,N_3758,N_3201);
nand U6523 (N_6523,N_4574,N_3729);
nor U6524 (N_6524,N_3537,N_5849);
nand U6525 (N_6525,N_5496,N_4209);
and U6526 (N_6526,N_3964,N_3295);
nand U6527 (N_6527,N_5430,N_5167);
nor U6528 (N_6528,N_5891,N_5901);
or U6529 (N_6529,N_4712,N_3292);
or U6530 (N_6530,N_5444,N_5071);
nor U6531 (N_6531,N_5457,N_5554);
xnor U6532 (N_6532,N_3897,N_3973);
and U6533 (N_6533,N_5974,N_4948);
and U6534 (N_6534,N_3529,N_3244);
nor U6535 (N_6535,N_4095,N_3136);
and U6536 (N_6536,N_5301,N_3845);
and U6537 (N_6537,N_4140,N_5741);
and U6538 (N_6538,N_4353,N_3651);
nand U6539 (N_6539,N_3816,N_4962);
or U6540 (N_6540,N_4044,N_3870);
nand U6541 (N_6541,N_4548,N_5567);
or U6542 (N_6542,N_3388,N_5025);
and U6543 (N_6543,N_3334,N_4700);
or U6544 (N_6544,N_5860,N_3520);
or U6545 (N_6545,N_4710,N_3291);
or U6546 (N_6546,N_5280,N_4325);
nor U6547 (N_6547,N_4934,N_4784);
or U6548 (N_6548,N_4204,N_5625);
nor U6549 (N_6549,N_3142,N_3297);
nor U6550 (N_6550,N_5517,N_3044);
nor U6551 (N_6551,N_3290,N_3188);
nand U6552 (N_6552,N_5626,N_4766);
and U6553 (N_6553,N_5130,N_5659);
nand U6554 (N_6554,N_4515,N_3263);
nand U6555 (N_6555,N_4340,N_4392);
and U6556 (N_6556,N_5147,N_5670);
or U6557 (N_6557,N_3551,N_4440);
or U6558 (N_6558,N_5353,N_4099);
and U6559 (N_6559,N_3192,N_5736);
xor U6560 (N_6560,N_4250,N_3991);
or U6561 (N_6561,N_5003,N_5010);
nor U6562 (N_6562,N_5522,N_5680);
nor U6563 (N_6563,N_4272,N_3792);
xor U6564 (N_6564,N_5075,N_5702);
nand U6565 (N_6565,N_4804,N_4757);
nor U6566 (N_6566,N_3121,N_4967);
and U6567 (N_6567,N_4984,N_5418);
nor U6568 (N_6568,N_3442,N_5909);
nor U6569 (N_6569,N_5045,N_4225);
nor U6570 (N_6570,N_4812,N_4735);
and U6571 (N_6571,N_3432,N_5309);
nor U6572 (N_6572,N_3179,N_3455);
nor U6573 (N_6573,N_4498,N_5360);
nor U6574 (N_6574,N_4755,N_3517);
nand U6575 (N_6575,N_4776,N_4946);
nor U6576 (N_6576,N_4196,N_5465);
nand U6577 (N_6577,N_3611,N_5713);
or U6578 (N_6578,N_3919,N_4016);
or U6579 (N_6579,N_5386,N_5228);
nor U6580 (N_6580,N_5107,N_3949);
or U6581 (N_6581,N_5701,N_4833);
nor U6582 (N_6582,N_4809,N_3790);
nand U6583 (N_6583,N_4068,N_4711);
nand U6584 (N_6584,N_3312,N_4842);
nor U6585 (N_6585,N_5382,N_4848);
nand U6586 (N_6586,N_3983,N_4426);
nand U6587 (N_6587,N_3779,N_5833);
nand U6588 (N_6588,N_3761,N_5971);
or U6589 (N_6589,N_3013,N_4149);
nand U6590 (N_6590,N_4815,N_5786);
nor U6591 (N_6591,N_5235,N_5956);
and U6592 (N_6592,N_5342,N_4110);
nor U6593 (N_6593,N_4822,N_4300);
or U6594 (N_6594,N_4852,N_3402);
nand U6595 (N_6595,N_5949,N_3496);
and U6596 (N_6596,N_3118,N_5371);
and U6597 (N_6597,N_4663,N_3411);
or U6598 (N_6598,N_5113,N_4800);
or U6599 (N_6599,N_5470,N_4606);
nand U6600 (N_6600,N_4907,N_4679);
nand U6601 (N_6601,N_3901,N_3439);
and U6602 (N_6602,N_4517,N_4871);
and U6603 (N_6603,N_3636,N_5289);
nand U6604 (N_6604,N_3515,N_5176);
or U6605 (N_6605,N_3358,N_3365);
and U6606 (N_6606,N_4808,N_5573);
or U6607 (N_6607,N_4533,N_3389);
nor U6608 (N_6608,N_4620,N_4382);
xnor U6609 (N_6609,N_4374,N_5519);
nand U6610 (N_6610,N_3909,N_4631);
nor U6611 (N_6611,N_5056,N_3028);
or U6612 (N_6612,N_5864,N_5226);
or U6613 (N_6613,N_3444,N_4400);
or U6614 (N_6614,N_4845,N_5783);
or U6615 (N_6615,N_3591,N_3542);
nand U6616 (N_6616,N_3404,N_3460);
and U6617 (N_6617,N_5359,N_4282);
or U6618 (N_6618,N_4487,N_5880);
nor U6619 (N_6619,N_4746,N_3516);
and U6620 (N_6620,N_4388,N_3176);
xnor U6621 (N_6621,N_4002,N_4510);
or U6622 (N_6622,N_4185,N_4372);
nor U6623 (N_6623,N_5012,N_3187);
or U6624 (N_6624,N_5066,N_3051);
nand U6625 (N_6625,N_5094,N_5879);
nor U6626 (N_6626,N_5925,N_3337);
or U6627 (N_6627,N_5332,N_5812);
nor U6628 (N_6628,N_5286,N_3233);
or U6629 (N_6629,N_3666,N_4579);
nand U6630 (N_6630,N_3004,N_3530);
or U6631 (N_6631,N_3124,N_5018);
nor U6632 (N_6632,N_4989,N_5623);
or U6633 (N_6633,N_5253,N_4671);
nand U6634 (N_6634,N_5020,N_3313);
and U6635 (N_6635,N_5219,N_3152);
or U6636 (N_6636,N_3155,N_3538);
and U6637 (N_6637,N_3890,N_4817);
nor U6638 (N_6638,N_5296,N_4122);
nor U6639 (N_6639,N_3012,N_3073);
nor U6640 (N_6640,N_4339,N_4117);
nand U6641 (N_6641,N_5287,N_5735);
and U6642 (N_6642,N_4421,N_3712);
or U6643 (N_6643,N_5338,N_4660);
or U6644 (N_6644,N_4003,N_3259);
and U6645 (N_6645,N_4015,N_5290);
nor U6646 (N_6646,N_4301,N_5112);
and U6647 (N_6647,N_5068,N_3249);
and U6648 (N_6648,N_5410,N_5295);
xor U6649 (N_6649,N_3874,N_4298);
nand U6650 (N_6650,N_4379,N_5840);
and U6651 (N_6651,N_3340,N_5963);
nand U6652 (N_6652,N_3342,N_4649);
or U6653 (N_6653,N_5874,N_3718);
xor U6654 (N_6654,N_4471,N_4756);
nand U6655 (N_6655,N_5946,N_3930);
nand U6656 (N_6656,N_4933,N_3047);
and U6657 (N_6657,N_4999,N_4970);
and U6658 (N_6658,N_4578,N_3819);
nand U6659 (N_6659,N_5774,N_5687);
nor U6660 (N_6660,N_4313,N_3622);
nand U6661 (N_6661,N_5242,N_3584);
and U6662 (N_6662,N_5231,N_4006);
nand U6663 (N_6663,N_5150,N_5933);
nand U6664 (N_6664,N_4216,N_4284);
nor U6665 (N_6665,N_5389,N_4875);
or U6666 (N_6666,N_5506,N_5208);
or U6667 (N_6667,N_5052,N_5699);
xnor U6668 (N_6668,N_4707,N_3068);
nand U6669 (N_6669,N_5972,N_4065);
nor U6670 (N_6670,N_4422,N_5413);
nor U6671 (N_6671,N_4105,N_3042);
or U6672 (N_6672,N_4182,N_5158);
and U6673 (N_6673,N_5191,N_5244);
or U6674 (N_6674,N_5900,N_5247);
nor U6675 (N_6675,N_4959,N_4189);
or U6676 (N_6676,N_4887,N_5655);
xor U6677 (N_6677,N_4614,N_3663);
or U6678 (N_6678,N_3248,N_4156);
nor U6679 (N_6679,N_3618,N_5293);
nor U6680 (N_6680,N_3363,N_3424);
nand U6681 (N_6681,N_5129,N_5624);
nor U6682 (N_6682,N_3577,N_4465);
nor U6683 (N_6683,N_3330,N_5093);
xor U6684 (N_6684,N_3974,N_3607);
and U6685 (N_6685,N_3726,N_3215);
nor U6686 (N_6686,N_3990,N_4888);
and U6687 (N_6687,N_4342,N_3844);
or U6688 (N_6688,N_5238,N_4789);
nor U6689 (N_6689,N_4455,N_3640);
nand U6690 (N_6690,N_5799,N_3895);
or U6691 (N_6691,N_4672,N_5948);
nor U6692 (N_6692,N_3898,N_3077);
or U6693 (N_6693,N_4516,N_5450);
nand U6694 (N_6694,N_3014,N_5199);
nor U6695 (N_6695,N_5696,N_4483);
and U6696 (N_6696,N_5853,N_4493);
and U6697 (N_6697,N_3752,N_3375);
and U6698 (N_6698,N_3100,N_4702);
xor U6699 (N_6699,N_5541,N_3341);
nand U6700 (N_6700,N_4835,N_4148);
and U6701 (N_6701,N_3369,N_3605);
and U6702 (N_6702,N_3814,N_5640);
nor U6703 (N_6703,N_5547,N_4997);
and U6704 (N_6704,N_4807,N_4840);
nand U6705 (N_6705,N_5728,N_3275);
and U6706 (N_6706,N_4950,N_4212);
nand U6707 (N_6707,N_3199,N_5171);
nor U6708 (N_6708,N_4100,N_4616);
nor U6709 (N_6709,N_5510,N_4596);
and U6710 (N_6710,N_5969,N_5504);
and U6711 (N_6711,N_3039,N_4116);
xor U6712 (N_6712,N_4074,N_5548);
xor U6713 (N_6713,N_3706,N_5463);
nand U6714 (N_6714,N_5227,N_4096);
or U6715 (N_6715,N_5322,N_5483);
nand U6716 (N_6716,N_3425,N_4420);
or U6717 (N_6717,N_5629,N_5792);
nor U6718 (N_6718,N_4919,N_4981);
nor U6719 (N_6719,N_5611,N_4477);
nand U6720 (N_6720,N_3781,N_4090);
nor U6721 (N_6721,N_3023,N_3646);
or U6722 (N_6722,N_3940,N_5307);
and U6723 (N_6723,N_5644,N_4449);
nand U6724 (N_6724,N_3664,N_5683);
and U6725 (N_6725,N_4927,N_3894);
and U6726 (N_6726,N_4640,N_5285);
nand U6727 (N_6727,N_3223,N_4169);
or U6728 (N_6728,N_3987,N_3097);
nand U6729 (N_6729,N_5589,N_5203);
nor U6730 (N_6730,N_3534,N_3450);
or U6731 (N_6731,N_4466,N_3357);
or U6732 (N_6732,N_5448,N_4937);
and U6733 (N_6733,N_5133,N_3040);
or U6734 (N_6734,N_5211,N_3469);
or U6735 (N_6735,N_3271,N_3981);
and U6736 (N_6736,N_4292,N_4753);
and U6737 (N_6737,N_5105,N_5369);
and U6738 (N_6738,N_3126,N_3560);
nor U6739 (N_6739,N_3774,N_5827);
and U6740 (N_6740,N_4485,N_3608);
nor U6741 (N_6741,N_4972,N_5639);
nor U6742 (N_6742,N_4028,N_3928);
or U6743 (N_6743,N_4078,N_3592);
and U6744 (N_6744,N_3351,N_3944);
or U6745 (N_6745,N_4885,N_5035);
nand U6746 (N_6746,N_5649,N_3135);
or U6747 (N_6747,N_3717,N_4629);
or U6748 (N_6748,N_5940,N_4164);
and U6749 (N_6749,N_5310,N_4513);
and U6750 (N_6750,N_3565,N_4311);
nor U6751 (N_6751,N_5711,N_3838);
xnor U6752 (N_6752,N_4000,N_3775);
or U6753 (N_6753,N_3691,N_4617);
and U6754 (N_6754,N_3937,N_3698);
or U6755 (N_6755,N_4511,N_5170);
nand U6756 (N_6756,N_3619,N_4364);
or U6757 (N_6757,N_5749,N_4745);
or U6758 (N_6758,N_4953,N_3882);
nor U6759 (N_6759,N_5054,N_3795);
nand U6760 (N_6760,N_3893,N_4450);
nand U6761 (N_6761,N_5552,N_4794);
or U6762 (N_6762,N_4275,N_5916);
nand U6763 (N_6763,N_4738,N_4772);
nand U6764 (N_6764,N_5498,N_4220);
nor U6765 (N_6765,N_3968,N_5435);
xor U6766 (N_6766,N_5784,N_5679);
nand U6767 (N_6767,N_5945,N_4754);
nand U6768 (N_6768,N_5283,N_5057);
or U6769 (N_6769,N_4475,N_3667);
and U6770 (N_6770,N_5460,N_3198);
or U6771 (N_6771,N_3021,N_3367);
nor U6772 (N_6772,N_4157,N_4234);
xnor U6773 (N_6773,N_4180,N_5957);
nor U6774 (N_6774,N_5272,N_4144);
and U6775 (N_6775,N_4622,N_4630);
nor U6776 (N_6776,N_3914,N_4905);
nor U6777 (N_6777,N_4431,N_5101);
and U6778 (N_6778,N_3333,N_5565);
and U6779 (N_6779,N_5795,N_3415);
and U6780 (N_6780,N_3933,N_3122);
and U6781 (N_6781,N_5255,N_3347);
nand U6782 (N_6782,N_5818,N_3601);
nand U6783 (N_6783,N_3151,N_5540);
or U6784 (N_6784,N_5264,N_3604);
or U6785 (N_6785,N_4334,N_3523);
or U6786 (N_6786,N_4005,N_4294);
or U6787 (N_6787,N_3002,N_5351);
nor U6788 (N_6788,N_5581,N_4605);
and U6789 (N_6789,N_5731,N_3066);
or U6790 (N_6790,N_3906,N_4319);
nor U6791 (N_6791,N_5739,N_4626);
and U6792 (N_6792,N_3318,N_4704);
xor U6793 (N_6793,N_3288,N_4893);
nor U6794 (N_6794,N_4879,N_4464);
or U6795 (N_6795,N_3613,N_3172);
nor U6796 (N_6796,N_4752,N_4709);
or U6797 (N_6797,N_3972,N_3720);
nor U6798 (N_6798,N_5557,N_3015);
nand U6799 (N_6799,N_4610,N_3947);
and U6800 (N_6800,N_5246,N_5569);
or U6801 (N_6801,N_3386,N_3309);
and U6802 (N_6802,N_5539,N_3807);
nand U6803 (N_6803,N_5452,N_3038);
nor U6804 (N_6804,N_3140,N_4193);
nand U6805 (N_6805,N_5065,N_4811);
and U6806 (N_6806,N_4247,N_4345);
or U6807 (N_6807,N_3954,N_4229);
nand U6808 (N_6808,N_4366,N_4418);
xnor U6809 (N_6809,N_3379,N_4012);
and U6810 (N_6810,N_4750,N_3768);
or U6811 (N_6811,N_4181,N_5852);
nand U6812 (N_6812,N_3778,N_5950);
and U6813 (N_6813,N_3737,N_4773);
xor U6814 (N_6814,N_3727,N_3336);
nand U6815 (N_6815,N_3162,N_4168);
nor U6816 (N_6816,N_4177,N_5336);
nand U6817 (N_6817,N_5583,N_4980);
or U6818 (N_6818,N_4427,N_3596);
and U6819 (N_6819,N_4395,N_5174);
nand U6820 (N_6820,N_5486,N_4528);
nor U6821 (N_6821,N_4820,N_4030);
nand U6822 (N_6822,N_4531,N_3503);
nand U6823 (N_6823,N_5673,N_4592);
nor U6824 (N_6824,N_5437,N_4452);
nand U6825 (N_6825,N_5224,N_5789);
nor U6826 (N_6826,N_3422,N_4166);
or U6827 (N_6827,N_4874,N_4810);
or U6828 (N_6828,N_3878,N_3785);
and U6829 (N_6829,N_5796,N_4071);
nor U6830 (N_6830,N_4128,N_4541);
or U6831 (N_6831,N_5559,N_4058);
xor U6832 (N_6832,N_3946,N_3266);
nor U6833 (N_6833,N_4391,N_3707);
nor U6834 (N_6834,N_3238,N_5661);
nor U6835 (N_6835,N_3154,N_5145);
xor U6836 (N_6836,N_5429,N_4356);
nand U6837 (N_6837,N_4866,N_5428);
nor U6838 (N_6838,N_3060,N_5368);
nand U6839 (N_6839,N_3316,N_5016);
nand U6840 (N_6840,N_3373,N_5740);
xnor U6841 (N_6841,N_5072,N_3063);
and U6842 (N_6842,N_5568,N_3600);
nand U6843 (N_6843,N_5654,N_4322);
or U6844 (N_6844,N_4460,N_3822);
nand U6845 (N_6845,N_3072,N_5777);
or U6846 (N_6846,N_3735,N_4925);
xor U6847 (N_6847,N_3209,N_5220);
xor U6848 (N_6848,N_3325,N_4550);
nor U6849 (N_6849,N_5838,N_4289);
nand U6850 (N_6850,N_4445,N_3376);
and U6851 (N_6851,N_3699,N_4577);
nand U6852 (N_6852,N_3817,N_4901);
or U6853 (N_6853,N_3000,N_4534);
nor U6854 (N_6854,N_4659,N_3936);
nor U6855 (N_6855,N_4115,N_5976);
or U6856 (N_6856,N_5767,N_3277);
nand U6857 (N_6857,N_4373,N_3486);
nand U6858 (N_6858,N_5188,N_4481);
or U6859 (N_6859,N_4491,N_3594);
or U6860 (N_6860,N_4394,N_4323);
or U6861 (N_6861,N_4205,N_3696);
or U6862 (N_6862,N_5663,N_4966);
nor U6863 (N_6863,N_3423,N_5766);
nand U6864 (N_6864,N_3834,N_5011);
nor U6865 (N_6865,N_3782,N_3243);
and U6866 (N_6866,N_4635,N_3431);
and U6867 (N_6867,N_4618,N_5961);
xor U6868 (N_6868,N_5143,N_3830);
or U6869 (N_6869,N_5995,N_3900);
nor U6870 (N_6870,N_3016,N_4836);
or U6871 (N_6871,N_3400,N_3658);
or U6872 (N_6872,N_5582,N_4532);
or U6873 (N_6873,N_3148,N_5647);
and U6874 (N_6874,N_3257,N_3499);
nand U6875 (N_6875,N_3314,N_5027);
and U6876 (N_6876,N_4960,N_4072);
xnor U6877 (N_6877,N_3165,N_3736);
nand U6878 (N_6878,N_4995,N_5772);
nor U6879 (N_6879,N_3965,N_4768);
or U6880 (N_6880,N_4297,N_4004);
nor U6881 (N_6881,N_4508,N_4238);
nand U6882 (N_6882,N_4245,N_5705);
nand U6883 (N_6883,N_4744,N_5381);
and U6884 (N_6884,N_3226,N_3740);
nor U6885 (N_6885,N_5404,N_5109);
nand U6886 (N_6886,N_3683,N_4462);
nor U6887 (N_6887,N_4974,N_3343);
or U6888 (N_6888,N_4666,N_4547);
nor U6889 (N_6889,N_4424,N_5964);
nand U6890 (N_6890,N_5561,N_3025);
and U6891 (N_6891,N_4066,N_5914);
and U6892 (N_6892,N_3931,N_3250);
nor U6893 (N_6893,N_3849,N_3693);
nand U6894 (N_6894,N_4343,N_4293);
or U6895 (N_6895,N_4430,N_4575);
nand U6896 (N_6896,N_4949,N_4987);
nor U6897 (N_6897,N_4088,N_4505);
or U6898 (N_6898,N_5832,N_4324);
nor U6899 (N_6899,N_4265,N_4170);
xnor U6900 (N_6900,N_4713,N_3557);
or U6901 (N_6901,N_3222,N_5785);
or U6902 (N_6902,N_3748,N_3302);
or U6903 (N_6903,N_3855,N_4802);
or U6904 (N_6904,N_4404,N_5042);
and U6905 (N_6905,N_5110,N_4360);
and U6906 (N_6906,N_5196,N_5656);
and U6907 (N_6907,N_5007,N_3208);
xnor U6908 (N_6908,N_5681,N_4142);
or U6909 (N_6909,N_5886,N_3355);
nand U6910 (N_6910,N_5403,N_3757);
or U6911 (N_6911,N_5341,N_3026);
and U6912 (N_6912,N_3156,N_4385);
or U6913 (N_6913,N_4184,N_4854);
nand U6914 (N_6914,N_3352,N_4407);
nand U6915 (N_6915,N_5374,N_4202);
nand U6916 (N_6916,N_3417,N_4646);
and U6917 (N_6917,N_3419,N_5865);
nand U6918 (N_6918,N_4331,N_3041);
nor U6919 (N_6919,N_5494,N_3031);
nand U6920 (N_6920,N_3344,N_3107);
nor U6921 (N_6921,N_5596,N_5558);
nand U6922 (N_6922,N_5585,N_4697);
and U6923 (N_6923,N_4120,N_5760);
nand U6924 (N_6924,N_5131,N_3255);
xnor U6925 (N_6925,N_3175,N_5929);
or U6926 (N_6926,N_5866,N_4726);
xor U6927 (N_6927,N_4317,N_4506);
and U6928 (N_6928,N_3310,N_3181);
nand U6929 (N_6929,N_3036,N_5124);
and U6930 (N_6930,N_4957,N_3943);
xnor U6931 (N_6931,N_4638,N_5761);
or U6932 (N_6932,N_5146,N_5978);
nand U6933 (N_6933,N_3345,N_3253);
nand U6934 (N_6934,N_5455,N_5924);
or U6935 (N_6935,N_5114,N_3750);
nor U6936 (N_6936,N_5141,N_3459);
and U6937 (N_6937,N_4280,N_3625);
nor U6938 (N_6938,N_4913,N_5385);
and U6939 (N_6939,N_3235,N_4764);
nor U6940 (N_6940,N_4080,N_5628);
xor U6941 (N_6941,N_4172,N_3615);
nor U6942 (N_6942,N_5493,N_4457);
nor U6943 (N_6943,N_3912,N_5040);
nand U6944 (N_6944,N_3203,N_4188);
nand U6945 (N_6945,N_5086,N_3823);
and U6946 (N_6946,N_5882,N_5132);
xor U6947 (N_6947,N_3478,N_3061);
nand U6948 (N_6948,N_5600,N_4330);
and U6949 (N_6949,N_3141,N_3273);
or U6950 (N_6950,N_4018,N_3670);
or U6951 (N_6951,N_5339,N_4847);
and U6952 (N_6952,N_3653,N_4335);
or U6953 (N_6953,N_4243,N_3276);
nand U6954 (N_6954,N_3561,N_3153);
and U6955 (N_6955,N_4580,N_3864);
or U6956 (N_6956,N_5305,N_5605);
nand U6957 (N_6957,N_3018,N_5173);
nor U6958 (N_6958,N_4478,N_5099);
and U6959 (N_6959,N_5302,N_5538);
xnor U6960 (N_6960,N_5883,N_4868);
or U6961 (N_6961,N_4573,N_5356);
nor U6962 (N_6962,N_4147,N_4488);
and U6963 (N_6963,N_5932,N_4101);
and U6964 (N_6964,N_5443,N_5999);
nand U6965 (N_6965,N_3096,N_4732);
nor U6966 (N_6966,N_3463,N_4698);
nor U6967 (N_6967,N_3826,N_5627);
nor U6968 (N_6968,N_3371,N_4895);
xor U6969 (N_6969,N_4608,N_3158);
and U6970 (N_6970,N_5848,N_4988);
and U6971 (N_6971,N_4053,N_4922);
and U6972 (N_6972,N_3138,N_4529);
nor U6973 (N_6973,N_4639,N_5811);
xor U6974 (N_6974,N_3677,N_5053);
nand U6975 (N_6975,N_5407,N_5314);
nand U6976 (N_6976,N_3880,N_4655);
nor U6977 (N_6977,N_3228,N_4434);
nand U6978 (N_6978,N_3045,N_5034);
and U6979 (N_6979,N_3074,N_4413);
nor U6980 (N_6980,N_5168,N_5449);
or U6981 (N_6981,N_3558,N_5169);
and U6982 (N_6982,N_3145,N_5261);
or U6983 (N_6983,N_4603,N_4696);
or U6984 (N_6984,N_5480,N_4320);
nor U6985 (N_6985,N_4591,N_5050);
or U6986 (N_6986,N_4179,N_4877);
nor U6987 (N_6987,N_3843,N_5968);
nand U6988 (N_6988,N_5876,N_5477);
and U6989 (N_6989,N_5752,N_3311);
nand U6990 (N_6990,N_5729,N_4792);
and U6991 (N_6991,N_4636,N_3055);
or U6992 (N_6992,N_5299,N_4151);
or U6993 (N_6993,N_4414,N_3511);
nand U6994 (N_6994,N_4200,N_3071);
or U6995 (N_6995,N_3364,N_3128);
and U6996 (N_6996,N_4472,N_4137);
or U6997 (N_6997,N_5422,N_4632);
nor U6998 (N_6998,N_4386,N_5835);
nor U6999 (N_6999,N_5546,N_4146);
nand U7000 (N_7000,N_3241,N_4315);
or U7001 (N_7001,N_3396,N_5781);
nand U7002 (N_7002,N_4944,N_3883);
and U7003 (N_7003,N_3392,N_4056);
nand U7004 (N_7004,N_4232,N_3105);
nor U7005 (N_7005,N_4683,N_3755);
and U7006 (N_7006,N_5277,N_3587);
nand U7007 (N_7007,N_5575,N_3827);
nor U7008 (N_7008,N_4024,N_5555);
nand U7009 (N_7009,N_4163,N_5032);
nor U7010 (N_7010,N_4760,N_5140);
or U7011 (N_7011,N_3274,N_4467);
or U7012 (N_7012,N_3256,N_3387);
or U7013 (N_7013,N_4361,N_5842);
or U7014 (N_7014,N_5675,N_5482);
or U7015 (N_7015,N_4770,N_4993);
nand U7016 (N_7016,N_3688,N_5650);
or U7017 (N_7017,N_3676,N_3159);
nand U7018 (N_7018,N_5545,N_4729);
and U7019 (N_7019,N_5920,N_4367);
nor U7020 (N_7020,N_5952,N_5355);
xnor U7021 (N_7021,N_3862,N_4383);
nor U7022 (N_7022,N_5878,N_5186);
xnor U7023 (N_7023,N_5722,N_3240);
nor U7024 (N_7024,N_3164,N_3786);
xor U7025 (N_7025,N_5632,N_4143);
xnor U7026 (N_7026,N_3682,N_4751);
and U7027 (N_7027,N_3648,N_4909);
or U7028 (N_7028,N_5509,N_4556);
or U7029 (N_7029,N_5438,N_4882);
nand U7030 (N_7030,N_5458,N_3621);
nor U7031 (N_7031,N_5563,N_5319);
nor U7032 (N_7032,N_5590,N_5487);
and U7033 (N_7033,N_4227,N_4255);
nor U7034 (N_7034,N_3802,N_4393);
and U7035 (N_7035,N_3189,N_3540);
and U7036 (N_7036,N_4186,N_3236);
or U7037 (N_7037,N_5938,N_4576);
and U7038 (N_7038,N_3328,N_5423);
or U7039 (N_7039,N_5892,N_5764);
or U7040 (N_7040,N_3307,N_3532);
nand U7041 (N_7041,N_4976,N_5104);
and U7042 (N_7042,N_3262,N_5269);
or U7043 (N_7043,N_3978,N_4832);
nor U7044 (N_7044,N_3024,N_5499);
and U7045 (N_7045,N_4208,N_5331);
and U7046 (N_7046,N_3035,N_4680);
nand U7047 (N_7047,N_4734,N_3390);
nand U7048 (N_7048,N_3510,N_3169);
or U7049 (N_7049,N_5947,N_5029);
nand U7050 (N_7050,N_4114,N_5822);
or U7051 (N_7051,N_4437,N_5979);
nand U7052 (N_7052,N_4226,N_4762);
and U7053 (N_7053,N_3382,N_4992);
or U7054 (N_7054,N_3111,N_4743);
or U7055 (N_7055,N_4551,N_5103);
xor U7056 (N_7056,N_3348,N_4191);
nand U7057 (N_7057,N_5362,N_3087);
xor U7058 (N_7058,N_5820,N_3836);
and U7059 (N_7059,N_3962,N_4880);
nor U7060 (N_7060,N_5198,N_5459);
xnor U7061 (N_7061,N_3620,N_5268);
nor U7062 (N_7062,N_4215,N_4621);
nand U7063 (N_7063,N_3326,N_3905);
and U7064 (N_7064,N_5850,N_5266);
or U7065 (N_7065,N_4045,N_5718);
nor U7066 (N_7066,N_5930,N_3349);
nor U7067 (N_7067,N_3723,N_3662);
xor U7068 (N_7068,N_5917,N_4521);
and U7069 (N_7069,N_3796,N_4341);
and U7070 (N_7070,N_4806,N_3232);
nand U7071 (N_7071,N_4441,N_3227);
nor U7072 (N_7072,N_5350,N_4536);
xnor U7073 (N_7073,N_5863,N_3976);
nor U7074 (N_7074,N_3885,N_5312);
nor U7075 (N_7075,N_4514,N_3840);
and U7076 (N_7076,N_5871,N_3952);
xor U7077 (N_7077,N_5063,N_4884);
xor U7078 (N_7078,N_4624,N_5134);
or U7079 (N_7079,N_5162,N_5877);
xnor U7080 (N_7080,N_4783,N_5047);
and U7081 (N_7081,N_4107,N_4086);
nand U7082 (N_7082,N_3771,N_4125);
nor U7083 (N_7083,N_4011,N_3265);
nor U7084 (N_7084,N_4910,N_3567);
and U7085 (N_7085,N_3916,N_3075);
nor U7086 (N_7086,N_5039,N_4463);
nand U7087 (N_7087,N_3078,N_3471);
nor U7088 (N_7088,N_4207,N_5270);
xnor U7089 (N_7089,N_5106,N_5707);
and U7090 (N_7090,N_3191,N_4942);
or U7091 (N_7091,N_5992,N_4359);
nor U7092 (N_7092,N_5431,N_5440);
nor U7093 (N_7093,N_4656,N_4266);
xor U7094 (N_7094,N_4584,N_4014);
nor U7095 (N_7095,N_5896,N_4786);
nand U7096 (N_7096,N_3366,N_4397);
nor U7097 (N_7097,N_3829,N_3998);
or U7098 (N_7098,N_3675,N_4767);
or U7099 (N_7099,N_4979,N_3588);
or U7100 (N_7100,N_4715,N_4865);
and U7101 (N_7101,N_4653,N_3547);
nand U7102 (N_7102,N_5514,N_5420);
nand U7103 (N_7103,N_4087,N_5122);
or U7104 (N_7104,N_4973,N_3955);
nor U7105 (N_7105,N_4503,N_5873);
nand U7106 (N_7106,N_3926,N_5653);
nor U7107 (N_7107,N_4602,N_5586);
or U7108 (N_7108,N_5894,N_4233);
nor U7109 (N_7109,N_3660,N_3851);
and U7110 (N_7110,N_5943,N_4013);
nor U7111 (N_7111,N_5041,N_4858);
nor U7112 (N_7112,N_5190,N_3549);
and U7113 (N_7113,N_3910,N_3202);
or U7114 (N_7114,N_5328,N_4499);
or U7115 (N_7115,N_4371,N_3730);
and U7116 (N_7116,N_5928,N_4230);
or U7117 (N_7117,N_3872,N_4775);
nand U7118 (N_7118,N_5810,N_5926);
or U7119 (N_7119,N_3076,N_5965);
and U7120 (N_7120,N_4287,N_4031);
or U7121 (N_7121,N_4563,N_4497);
or U7122 (N_7122,N_4378,N_5249);
nand U7123 (N_7123,N_4518,N_3884);
or U7124 (N_7124,N_4522,N_4057);
nor U7125 (N_7125,N_3925,N_5415);
nand U7126 (N_7126,N_4312,N_4389);
and U7127 (N_7127,N_4898,N_3391);
nor U7128 (N_7128,N_4667,N_4860);
nor U7129 (N_7129,N_3020,N_4027);
and U7130 (N_7130,N_3848,N_3300);
xnor U7131 (N_7131,N_3427,N_5474);
or U7132 (N_7132,N_5051,N_3639);
and U7133 (N_7133,N_4500,N_4377);
or U7134 (N_7134,N_3769,N_3120);
or U7135 (N_7135,N_3032,N_5373);
or U7136 (N_7136,N_5472,N_5273);
nand U7137 (N_7137,N_5923,N_5087);
and U7138 (N_7138,N_4856,N_3630);
and U7139 (N_7139,N_5686,N_5476);
and U7140 (N_7140,N_5987,N_4240);
nand U7141 (N_7141,N_5009,N_3339);
xnor U7142 (N_7142,N_5788,N_3405);
nor U7143 (N_7143,N_4468,N_4259);
and U7144 (N_7144,N_3711,N_4830);
nor U7145 (N_7145,N_4758,N_4337);
nor U7146 (N_7146,N_4174,N_4546);
nor U7147 (N_7147,N_5612,N_5257);
nand U7148 (N_7148,N_3773,N_5674);
xnor U7149 (N_7149,N_3960,N_4759);
nand U7150 (N_7150,N_5148,N_3219);
or U7151 (N_7151,N_5695,N_4994);
and U7152 (N_7152,N_3007,N_3745);
or U7153 (N_7153,N_4600,N_5082);
or U7154 (N_7154,N_3448,N_3783);
and U7155 (N_7155,N_5184,N_5159);
nor U7156 (N_7156,N_5922,N_5939);
or U7157 (N_7157,N_5446,N_4355);
nor U7158 (N_7158,N_5036,N_3435);
or U7159 (N_7159,N_5757,N_4869);
or U7160 (N_7160,N_3891,N_5770);
xor U7161 (N_7161,N_4461,N_5991);
or U7162 (N_7162,N_5375,N_5152);
nand U7163 (N_7163,N_3841,N_3522);
xnor U7164 (N_7164,N_3462,N_3456);
and U7165 (N_7165,N_5000,N_3803);
nand U7166 (N_7166,N_4271,N_3258);
or U7167 (N_7167,N_4009,N_5393);
or U7168 (N_7168,N_4470,N_3204);
nand U7169 (N_7169,N_3749,N_4263);
nor U7170 (N_7170,N_3610,N_5201);
and U7171 (N_7171,N_4258,N_4921);
xnor U7172 (N_7172,N_4459,N_5723);
or U7173 (N_7173,N_4918,N_5098);
nand U7174 (N_7174,N_3514,N_3380);
nor U7175 (N_7175,N_4442,N_3182);
xor U7176 (N_7176,N_4968,N_5775);
or U7177 (N_7177,N_4943,N_5125);
nor U7178 (N_7178,N_4714,N_3652);
or U7179 (N_7179,N_5910,N_3846);
or U7180 (N_7180,N_4545,N_4504);
and U7181 (N_7181,N_4150,N_4831);
and U7182 (N_7182,N_3200,N_4594);
nand U7183 (N_7183,N_3354,N_4344);
xnor U7184 (N_7184,N_5439,N_4160);
xnor U7185 (N_7185,N_5419,N_3902);
and U7186 (N_7186,N_3150,N_3043);
and U7187 (N_7187,N_3484,N_5172);
or U7188 (N_7188,N_3617,N_4823);
or U7189 (N_7189,N_5934,N_4021);
and U7190 (N_7190,N_3637,N_4890);
and U7191 (N_7191,N_4695,N_5801);
and U7192 (N_7192,N_3831,N_3957);
nor U7193 (N_7193,N_5988,N_5692);
and U7194 (N_7194,N_4241,N_5698);
xnor U7195 (N_7195,N_4288,N_3760);
nand U7196 (N_7196,N_4291,N_5006);
or U7197 (N_7197,N_4965,N_5424);
nand U7198 (N_7198,N_3645,N_4283);
nand U7199 (N_7199,N_3098,N_5544);
and U7200 (N_7200,N_5135,N_3206);
and U7201 (N_7201,N_4192,N_4476);
nand U7202 (N_7202,N_3765,N_4796);
nor U7203 (N_7203,N_4218,N_3702);
nor U7204 (N_7204,N_4025,N_3453);
nand U7205 (N_7205,N_3684,N_3528);
and U7206 (N_7206,N_5121,N_4203);
xor U7207 (N_7207,N_3575,N_3231);
and U7208 (N_7208,N_5906,N_5014);
or U7209 (N_7209,N_4923,N_3378);
or U7210 (N_7210,N_4318,N_5142);
nor U7211 (N_7211,N_4945,N_3103);
and U7212 (N_7212,N_5904,N_3728);
or U7213 (N_7213,N_4277,N_3319);
nor U7214 (N_7214,N_5377,N_5279);
or U7215 (N_7215,N_4132,N_5195);
or U7216 (N_7216,N_5983,N_3091);
nor U7217 (N_7217,N_4453,N_4891);
and U7218 (N_7218,N_4336,N_5733);
nand U7219 (N_7219,N_3481,N_5433);
nand U7220 (N_7220,N_4886,N_4401);
and U7221 (N_7221,N_4423,N_4876);
nand U7222 (N_7222,N_5251,N_4329);
nor U7223 (N_7223,N_5776,N_3526);
xor U7224 (N_7224,N_3788,N_3763);
xor U7225 (N_7225,N_3298,N_4236);
nor U7226 (N_7226,N_5762,N_5154);
nand U7227 (N_7227,N_4911,N_5942);
and U7228 (N_7228,N_5064,N_4145);
or U7229 (N_7229,N_4165,N_3010);
or U7230 (N_7230,N_4644,N_3850);
or U7231 (N_7231,N_3793,N_5576);
nand U7232 (N_7232,N_5802,N_5837);
or U7233 (N_7233,N_5756,N_3881);
or U7234 (N_7234,N_5421,N_4903);
nand U7235 (N_7235,N_5962,N_5651);
nand U7236 (N_7236,N_3433,N_5664);
and U7237 (N_7237,N_4846,N_5209);
and U7238 (N_7238,N_3137,N_3050);
and U7239 (N_7239,N_5927,N_5807);
or U7240 (N_7240,N_3669,N_5937);
nand U7241 (N_7241,N_4017,N_5985);
nand U7242 (N_7242,N_3847,N_3657);
and U7243 (N_7243,N_4139,N_4652);
and U7244 (N_7244,N_3866,N_4582);
nor U7245 (N_7245,N_3464,N_5138);
or U7246 (N_7246,N_3332,N_5502);
and U7247 (N_7247,N_3245,N_4851);
or U7248 (N_7248,N_4130,N_4722);
and U7249 (N_7249,N_4129,N_3194);
nor U7250 (N_7250,N_3144,N_4419);
nand U7251 (N_7251,N_4785,N_3488);
xnor U7252 (N_7252,N_5931,N_5021);
or U7253 (N_7253,N_4231,N_4480);
nand U7254 (N_7254,N_4650,N_3458);
or U7255 (N_7255,N_5898,N_5843);
or U7256 (N_7256,N_4352,N_3913);
or U7257 (N_7257,N_5515,N_5467);
and U7258 (N_7258,N_3668,N_5333);
nand U7259 (N_7259,N_4914,N_5989);
and U7260 (N_7260,N_3190,N_5682);
nor U7261 (N_7261,N_5222,N_3562);
and U7262 (N_7262,N_3820,N_3614);
and U7263 (N_7263,N_3559,N_3643);
nand U7264 (N_7264,N_3278,N_3770);
nand U7265 (N_7265,N_4131,N_3704);
or U7266 (N_7266,N_4664,N_3211);
nor U7267 (N_7267,N_3716,N_4543);
nand U7268 (N_7268,N_5019,N_3468);
nand U7269 (N_7269,N_4273,N_3492);
nand U7270 (N_7270,N_4524,N_5887);
and U7271 (N_7271,N_3430,N_4350);
nor U7272 (N_7272,N_5870,N_5516);
nand U7273 (N_7273,N_5862,N_4677);
or U7274 (N_7274,N_3867,N_5562);
and U7275 (N_7275,N_3064,N_5179);
and U7276 (N_7276,N_5005,N_4314);
or U7277 (N_7277,N_3494,N_4007);
nand U7278 (N_7278,N_5616,N_4763);
nand U7279 (N_7279,N_3490,N_3171);
and U7280 (N_7280,N_4668,N_3437);
nand U7281 (N_7281,N_3321,N_3935);
nor U7282 (N_7282,N_5967,N_5518);
or U7283 (N_7283,N_5895,N_5022);
nor U7284 (N_7284,N_3017,N_3251);
and U7285 (N_7285,N_5549,N_5217);
or U7286 (N_7286,N_4010,N_5712);
or U7287 (N_7287,N_5391,N_3958);
nor U7288 (N_7288,N_4244,N_4781);
and U7289 (N_7289,N_5966,N_5330);
or U7290 (N_7290,N_5300,N_5357);
nor U7291 (N_7291,N_4853,N_3566);
xor U7292 (N_7292,N_3953,N_4076);
and U7293 (N_7293,N_5263,N_4162);
nand U7294 (N_7294,N_5959,N_3320);
xnor U7295 (N_7295,N_3350,N_3635);
xnor U7296 (N_7296,N_5372,N_4691);
and U7297 (N_7297,N_5941,N_5427);
or U7298 (N_7298,N_4494,N_4894);
xnor U7299 (N_7299,N_4733,N_5758);
nand U7300 (N_7300,N_5481,N_4121);
nand U7301 (N_7301,N_5123,N_4825);
and U7302 (N_7302,N_3216,N_3759);
and U7303 (N_7303,N_5434,N_5049);
nand U7304 (N_7304,N_3599,N_3634);
nor U7305 (N_7305,N_5905,N_4849);
nor U7306 (N_7306,N_5352,N_4986);
xor U7307 (N_7307,N_5823,N_5537);
or U7308 (N_7308,N_4926,N_4585);
xor U7309 (N_7309,N_3572,N_4685);
or U7310 (N_7310,N_3766,N_3173);
nor U7311 (N_7311,N_3539,N_3997);
and U7312 (N_7312,N_3308,N_4155);
nand U7313 (N_7313,N_4727,N_5340);
nor U7314 (N_7314,N_5454,N_3008);
nor U7315 (N_7315,N_4769,N_5038);
nand U7316 (N_7316,N_5645,N_3512);
or U7317 (N_7317,N_3414,N_3506);
nand U7318 (N_7318,N_3756,N_5830);
or U7319 (N_7319,N_4611,N_3212);
nand U7320 (N_7320,N_5489,N_4561);
or U7321 (N_7321,N_3356,N_3395);
nand U7322 (N_7322,N_4048,N_4050);
or U7323 (N_7323,N_4159,N_4947);
nor U7324 (N_7324,N_3421,N_3924);
nor U7325 (N_7325,N_5081,N_5676);
and U7326 (N_7326,N_5884,N_4432);
and U7327 (N_7327,N_4223,N_3132);
nor U7328 (N_7328,N_5580,N_3286);
nand U7329 (N_7329,N_3372,N_4931);
or U7330 (N_7330,N_3580,N_3322);
and U7331 (N_7331,N_5734,N_3119);
and U7332 (N_7332,N_4538,N_3569);
or U7333 (N_7333,N_3661,N_3606);
nor U7334 (N_7334,N_4520,N_3932);
or U7335 (N_7335,N_4246,N_5861);
nand U7336 (N_7336,N_5074,N_5813);
or U7337 (N_7337,N_4777,N_3603);
or U7338 (N_7338,N_3731,N_4482);
nor U7339 (N_7339,N_4363,N_4043);
nor U7340 (N_7340,N_3985,N_4839);
nand U7341 (N_7341,N_4217,N_3800);
xnor U7342 (N_7342,N_4093,N_3821);
nand U7343 (N_7343,N_4211,N_3911);
xnor U7344 (N_7344,N_5704,N_5297);
nor U7345 (N_7345,N_5814,N_5584);
xor U7346 (N_7346,N_4609,N_4295);
nand U7347 (N_7347,N_5354,N_3133);
nand U7348 (N_7348,N_3689,N_4376);
nand U7349 (N_7349,N_3742,N_5365);
nor U7350 (N_7350,N_5023,N_4924);
or U7351 (N_7351,N_4251,N_5759);
xor U7352 (N_7352,N_3006,N_5638);
or U7353 (N_7353,N_4381,N_4941);
nor U7354 (N_7354,N_4593,N_5291);
or U7355 (N_7355,N_3123,N_4064);
and U7356 (N_7356,N_4235,N_4038);
nor U7357 (N_7357,N_4175,N_4555);
and U7358 (N_7358,N_4059,N_5714);
nor U7359 (N_7359,N_5213,N_3754);
nand U7360 (N_7360,N_3975,N_5893);
nor U7361 (N_7361,N_5621,N_3080);
nand U7362 (N_7362,N_4402,N_3927);
and U7363 (N_7363,N_4619,N_5646);
nand U7364 (N_7364,N_4583,N_5529);
or U7365 (N_7365,N_4438,N_5996);
nor U7366 (N_7366,N_3908,N_5787);
nor U7367 (N_7367,N_5641,N_4279);
nor U7368 (N_7368,N_4826,N_3160);
nand U7369 (N_7369,N_4171,N_3279);
xor U7370 (N_7370,N_5715,N_4975);
nor U7371 (N_7371,N_5239,N_4565);
xnor U7372 (N_7372,N_5662,N_4607);
nor U7373 (N_7373,N_4502,N_4567);
or U7374 (N_7374,N_5543,N_3835);
nor U7375 (N_7375,N_5613,N_4912);
or U7376 (N_7376,N_4507,N_5207);
nor U7377 (N_7377,N_4219,N_4032);
or U7378 (N_7378,N_5055,N_4254);
nor U7379 (N_7379,N_5205,N_5182);
nor U7380 (N_7380,N_5347,N_3948);
nand U7381 (N_7381,N_3370,N_4623);
xor U7382 (N_7382,N_4647,N_3505);
nand U7383 (N_7383,N_4118,N_5508);
or U7384 (N_7384,N_4333,N_4693);
and U7385 (N_7385,N_5197,N_4490);
or U7386 (N_7386,N_5008,N_4084);
xnor U7387 (N_7387,N_3633,N_3839);
or U7388 (N_7388,N_4152,N_5725);
nand U7389 (N_7389,N_3602,N_4369);
nor U7390 (N_7390,N_3084,N_3695);
xor U7391 (N_7391,N_5402,N_5274);
and U7392 (N_7392,N_5710,N_4787);
nor U7393 (N_7393,N_4615,N_5800);
nand U7394 (N_7394,N_5512,N_5412);
nor U7395 (N_7395,N_5855,N_5313);
or U7396 (N_7396,N_5572,N_5030);
nor U7397 (N_7397,N_4153,N_5859);
nor U7398 (N_7398,N_4899,N_5599);
nand U7399 (N_7399,N_5062,N_4821);
or U7400 (N_7400,N_5392,N_5485);
and U7401 (N_7401,N_5026,N_5037);
and U7402 (N_7402,N_3942,N_3680);
or U7403 (N_7403,N_5400,N_5200);
or U7404 (N_7404,N_5090,N_5536);
and U7405 (N_7405,N_5500,N_5398);
or U7406 (N_7406,N_4859,N_4598);
and U7407 (N_7407,N_3305,N_4123);
and U7408 (N_7408,N_5773,N_4348);
or U7409 (N_7409,N_3196,N_5660);
nor U7410 (N_7410,N_5189,N_5256);
xnor U7411 (N_7411,N_4326,N_5724);
xnor U7412 (N_7412,N_4458,N_5595);
nor U7413 (N_7413,N_5780,N_5808);
and U7414 (N_7414,N_3889,N_5505);
or U7415 (N_7415,N_5854,N_4278);
and U7416 (N_7416,N_3686,N_3465);
nor U7417 (N_7417,N_5730,N_4694);
or U7418 (N_7418,N_5868,N_3398);
or U7419 (N_7419,N_5834,N_4081);
or U7420 (N_7420,N_5058,N_5806);
nor U7421 (N_7421,N_3876,N_5409);
or U7422 (N_7422,N_5633,N_4544);
and U7423 (N_7423,N_3324,N_4791);
nand U7424 (N_7424,N_3317,N_4347);
nand U7425 (N_7425,N_5915,N_4138);
xor U7426 (N_7426,N_4176,N_4570);
and U7427 (N_7427,N_4761,N_3543);
nor U7428 (N_7428,N_4486,N_5604);
nor U7429 (N_7429,N_5490,N_3628);
nand U7430 (N_7430,N_5574,N_5875);
or U7431 (N_7431,N_5919,N_5077);
and U7432 (N_7432,N_5497,N_5245);
nor U7433 (N_7433,N_3163,N_3269);
and U7434 (N_7434,N_5157,N_5648);
xnor U7435 (N_7435,N_4706,N_5070);
nand U7436 (N_7436,N_5127,N_3401);
and U7437 (N_7437,N_4687,N_5678);
nor U7438 (N_7438,N_3656,N_3489);
or U7439 (N_7439,N_3679,N_3568);
nor U7440 (N_7440,N_3185,N_3546);
nor U7441 (N_7441,N_4801,N_4590);
or U7442 (N_7442,N_5225,N_5982);
and U7443 (N_7443,N_5846,N_5078);
xor U7444 (N_7444,N_4581,N_3483);
nand U7445 (N_7445,N_4119,N_4446);
nor U7446 (N_7446,N_4634,N_4448);
and U7447 (N_7447,N_3626,N_3480);
or U7448 (N_7448,N_4489,N_5918);
nand U7449 (N_7449,N_5593,N_4587);
and U7450 (N_7450,N_5462,N_3436);
nor U7451 (N_7451,N_5210,N_4454);
or U7452 (N_7452,N_5156,N_4930);
or U7453 (N_7453,N_3108,N_3563);
xnor U7454 (N_7454,N_3980,N_3183);
or U7455 (N_7455,N_5897,N_3970);
or U7456 (N_7456,N_4077,N_4588);
or U7457 (N_7457,N_3180,N_3616);
and U7458 (N_7458,N_4669,N_5060);
nor U7459 (N_7459,N_4113,N_3624);
or U7460 (N_7460,N_4094,N_4019);
nand U7461 (N_7461,N_3131,N_4307);
nand U7462 (N_7462,N_3548,N_4771);
or U7463 (N_7463,N_4167,N_4535);
nand U7464 (N_7464,N_3327,N_5475);
nand U7465 (N_7465,N_5798,N_3299);
and U7466 (N_7466,N_5666,N_5258);
or U7467 (N_7467,N_3261,N_3655);
or U7468 (N_7468,N_3443,N_4977);
and U7469 (N_7469,N_4684,N_4237);
and U7470 (N_7470,N_4286,N_3705);
and U7471 (N_7471,N_4109,N_4296);
and U7472 (N_7472,N_4303,N_3385);
or U7473 (N_7473,N_5119,N_5738);
or U7474 (N_7474,N_5343,N_3917);
and U7475 (N_7475,N_4641,N_3487);
and U7476 (N_7476,N_4328,N_4037);
or U7477 (N_7477,N_3359,N_5346);
or U7478 (N_7478,N_4560,N_5378);
or U7479 (N_7479,N_3576,N_3642);
nor U7480 (N_7480,N_4309,N_5594);
and U7481 (N_7481,N_5888,N_3125);
nand U7482 (N_7482,N_5091,N_5237);
nand U7483 (N_7483,N_5615,N_5610);
and U7484 (N_7484,N_4410,N_3438);
or U7485 (N_7485,N_4253,N_5994);
and U7486 (N_7486,N_5618,N_3454);
or U7487 (N_7487,N_3609,N_5765);
nand U7488 (N_7488,N_3011,N_3331);
and U7489 (N_7489,N_3956,N_4302);
nor U7490 (N_7490,N_4276,N_5984);
and U7491 (N_7491,N_3521,N_4104);
nor U7492 (N_7492,N_3057,N_5390);
or U7493 (N_7493,N_3166,N_4720);
and U7494 (N_7494,N_4349,N_5358);
nand U7495 (N_7495,N_3127,N_5491);
and U7496 (N_7496,N_5097,N_3627);
and U7497 (N_7497,N_5085,N_3410);
and U7498 (N_7498,N_4688,N_5183);
nor U7499 (N_7499,N_3056,N_5954);
nor U7500 (N_7500,N_3881,N_5480);
xnor U7501 (N_7501,N_5997,N_5844);
nand U7502 (N_7502,N_4687,N_3897);
nor U7503 (N_7503,N_4981,N_3575);
or U7504 (N_7504,N_4353,N_3805);
xnor U7505 (N_7505,N_3519,N_4505);
nor U7506 (N_7506,N_3896,N_3503);
or U7507 (N_7507,N_4503,N_5639);
and U7508 (N_7508,N_3404,N_3366);
or U7509 (N_7509,N_3606,N_5537);
nor U7510 (N_7510,N_3542,N_5258);
nor U7511 (N_7511,N_4542,N_4838);
and U7512 (N_7512,N_3878,N_4744);
or U7513 (N_7513,N_5137,N_4582);
or U7514 (N_7514,N_4732,N_3298);
xnor U7515 (N_7515,N_3333,N_4835);
xnor U7516 (N_7516,N_4935,N_3731);
nand U7517 (N_7517,N_3798,N_5813);
nor U7518 (N_7518,N_5521,N_5200);
or U7519 (N_7519,N_3481,N_4381);
nand U7520 (N_7520,N_5157,N_4375);
nand U7521 (N_7521,N_4349,N_4953);
nor U7522 (N_7522,N_5634,N_3295);
nand U7523 (N_7523,N_4583,N_4625);
and U7524 (N_7524,N_4634,N_5514);
or U7525 (N_7525,N_5728,N_3708);
nor U7526 (N_7526,N_4082,N_4249);
and U7527 (N_7527,N_3194,N_3090);
nor U7528 (N_7528,N_4516,N_3227);
nor U7529 (N_7529,N_3899,N_3377);
or U7530 (N_7530,N_5420,N_4714);
nand U7531 (N_7531,N_5521,N_3319);
nor U7532 (N_7532,N_3461,N_4831);
and U7533 (N_7533,N_3548,N_3990);
nand U7534 (N_7534,N_4588,N_3598);
nor U7535 (N_7535,N_5516,N_4747);
or U7536 (N_7536,N_5729,N_5488);
and U7537 (N_7537,N_5814,N_5459);
nor U7538 (N_7538,N_5663,N_5770);
nor U7539 (N_7539,N_4665,N_4792);
and U7540 (N_7540,N_4200,N_3926);
and U7541 (N_7541,N_5562,N_3066);
xnor U7542 (N_7542,N_4955,N_3036);
and U7543 (N_7543,N_3528,N_4228);
nand U7544 (N_7544,N_5935,N_4058);
or U7545 (N_7545,N_3088,N_4220);
and U7546 (N_7546,N_3293,N_3481);
and U7547 (N_7547,N_4932,N_5854);
or U7548 (N_7548,N_3419,N_4059);
nor U7549 (N_7549,N_5749,N_5192);
nand U7550 (N_7550,N_4498,N_5692);
nor U7551 (N_7551,N_5731,N_3385);
nand U7552 (N_7552,N_3018,N_5709);
and U7553 (N_7553,N_3256,N_4931);
or U7554 (N_7554,N_5357,N_5803);
and U7555 (N_7555,N_4815,N_4170);
nand U7556 (N_7556,N_4993,N_4617);
xnor U7557 (N_7557,N_4590,N_4011);
or U7558 (N_7558,N_3037,N_3516);
nor U7559 (N_7559,N_3789,N_4132);
xnor U7560 (N_7560,N_4967,N_5181);
or U7561 (N_7561,N_5050,N_5031);
and U7562 (N_7562,N_4150,N_5115);
and U7563 (N_7563,N_5551,N_4654);
or U7564 (N_7564,N_4559,N_4729);
or U7565 (N_7565,N_5341,N_4249);
and U7566 (N_7566,N_4395,N_5306);
nor U7567 (N_7567,N_3660,N_4423);
or U7568 (N_7568,N_3594,N_4872);
or U7569 (N_7569,N_3595,N_5213);
nor U7570 (N_7570,N_3001,N_4125);
nor U7571 (N_7571,N_5173,N_5484);
xnor U7572 (N_7572,N_5925,N_5240);
or U7573 (N_7573,N_5084,N_4646);
nand U7574 (N_7574,N_3503,N_4667);
or U7575 (N_7575,N_3077,N_4108);
nor U7576 (N_7576,N_3587,N_5648);
nor U7577 (N_7577,N_4462,N_3032);
or U7578 (N_7578,N_3392,N_3199);
nand U7579 (N_7579,N_4791,N_3800);
xnor U7580 (N_7580,N_5871,N_5915);
and U7581 (N_7581,N_3927,N_3403);
nand U7582 (N_7582,N_4244,N_3343);
or U7583 (N_7583,N_3677,N_5570);
or U7584 (N_7584,N_4467,N_3114);
nor U7585 (N_7585,N_4084,N_3309);
and U7586 (N_7586,N_3775,N_4063);
or U7587 (N_7587,N_5386,N_3399);
or U7588 (N_7588,N_4195,N_3989);
nand U7589 (N_7589,N_4839,N_5424);
nor U7590 (N_7590,N_4459,N_4397);
or U7591 (N_7591,N_3422,N_4026);
and U7592 (N_7592,N_5554,N_3254);
nor U7593 (N_7593,N_3156,N_5954);
and U7594 (N_7594,N_5533,N_3841);
or U7595 (N_7595,N_4433,N_5907);
and U7596 (N_7596,N_5301,N_3531);
nand U7597 (N_7597,N_5495,N_5038);
nand U7598 (N_7598,N_3627,N_3505);
nand U7599 (N_7599,N_3240,N_3034);
nand U7600 (N_7600,N_4624,N_3852);
xnor U7601 (N_7601,N_4274,N_3500);
nor U7602 (N_7602,N_4273,N_3453);
and U7603 (N_7603,N_4339,N_5531);
or U7604 (N_7604,N_4657,N_3766);
nand U7605 (N_7605,N_5246,N_5395);
nand U7606 (N_7606,N_4745,N_4489);
and U7607 (N_7607,N_3548,N_5006);
and U7608 (N_7608,N_4703,N_5326);
and U7609 (N_7609,N_4706,N_5101);
nor U7610 (N_7610,N_5320,N_3762);
or U7611 (N_7611,N_5361,N_5743);
nor U7612 (N_7612,N_5477,N_3993);
nor U7613 (N_7613,N_4961,N_4909);
nor U7614 (N_7614,N_3446,N_4767);
or U7615 (N_7615,N_3661,N_4277);
and U7616 (N_7616,N_5133,N_4021);
and U7617 (N_7617,N_5133,N_3995);
nor U7618 (N_7618,N_3999,N_4176);
nor U7619 (N_7619,N_4526,N_4674);
and U7620 (N_7620,N_4235,N_4817);
or U7621 (N_7621,N_3785,N_5368);
or U7622 (N_7622,N_5628,N_3904);
or U7623 (N_7623,N_5820,N_4458);
nand U7624 (N_7624,N_4371,N_3188);
nor U7625 (N_7625,N_5548,N_4370);
nand U7626 (N_7626,N_5747,N_3889);
nand U7627 (N_7627,N_4468,N_4179);
or U7628 (N_7628,N_4796,N_3175);
xor U7629 (N_7629,N_3260,N_4123);
and U7630 (N_7630,N_5543,N_3531);
and U7631 (N_7631,N_3760,N_4398);
and U7632 (N_7632,N_5959,N_3231);
xor U7633 (N_7633,N_5254,N_3021);
xor U7634 (N_7634,N_3222,N_4945);
nand U7635 (N_7635,N_5642,N_5962);
and U7636 (N_7636,N_4985,N_5354);
or U7637 (N_7637,N_3507,N_4972);
nand U7638 (N_7638,N_4578,N_5875);
or U7639 (N_7639,N_5265,N_4280);
nor U7640 (N_7640,N_4343,N_5728);
nand U7641 (N_7641,N_3400,N_5261);
nor U7642 (N_7642,N_4338,N_5312);
nor U7643 (N_7643,N_5226,N_3218);
or U7644 (N_7644,N_5742,N_5273);
and U7645 (N_7645,N_3182,N_3325);
or U7646 (N_7646,N_5619,N_4213);
nor U7647 (N_7647,N_3481,N_3387);
xnor U7648 (N_7648,N_5138,N_4904);
and U7649 (N_7649,N_3952,N_3828);
nand U7650 (N_7650,N_4801,N_4272);
nand U7651 (N_7651,N_3190,N_4044);
nand U7652 (N_7652,N_5488,N_3517);
nor U7653 (N_7653,N_4221,N_4022);
or U7654 (N_7654,N_5655,N_4933);
and U7655 (N_7655,N_3900,N_5533);
or U7656 (N_7656,N_3922,N_4474);
nand U7657 (N_7657,N_4054,N_5350);
nor U7658 (N_7658,N_5420,N_4905);
nor U7659 (N_7659,N_3685,N_4098);
or U7660 (N_7660,N_4569,N_4724);
xnor U7661 (N_7661,N_4932,N_4150);
nor U7662 (N_7662,N_3166,N_4320);
nor U7663 (N_7663,N_3692,N_4706);
or U7664 (N_7664,N_3735,N_5104);
nor U7665 (N_7665,N_3624,N_5949);
nor U7666 (N_7666,N_3653,N_4770);
nand U7667 (N_7667,N_3311,N_5283);
nand U7668 (N_7668,N_5151,N_4932);
or U7669 (N_7669,N_4349,N_5939);
and U7670 (N_7670,N_3277,N_3289);
nor U7671 (N_7671,N_3510,N_5253);
and U7672 (N_7672,N_5417,N_4462);
or U7673 (N_7673,N_5726,N_5418);
nor U7674 (N_7674,N_3039,N_3443);
or U7675 (N_7675,N_5226,N_3328);
and U7676 (N_7676,N_4703,N_5172);
nor U7677 (N_7677,N_3595,N_3252);
and U7678 (N_7678,N_3175,N_3924);
or U7679 (N_7679,N_5261,N_3612);
or U7680 (N_7680,N_5802,N_5554);
and U7681 (N_7681,N_4573,N_5328);
and U7682 (N_7682,N_5893,N_4216);
xor U7683 (N_7683,N_5028,N_3117);
nor U7684 (N_7684,N_3218,N_5900);
and U7685 (N_7685,N_5367,N_5805);
or U7686 (N_7686,N_3915,N_3447);
or U7687 (N_7687,N_5040,N_5576);
nand U7688 (N_7688,N_5592,N_3799);
and U7689 (N_7689,N_3782,N_5745);
or U7690 (N_7690,N_3744,N_3100);
nand U7691 (N_7691,N_3580,N_4186);
or U7692 (N_7692,N_4255,N_3683);
or U7693 (N_7693,N_4992,N_5922);
or U7694 (N_7694,N_3487,N_3011);
xnor U7695 (N_7695,N_4430,N_3993);
xor U7696 (N_7696,N_5462,N_3220);
or U7697 (N_7697,N_3646,N_3642);
nand U7698 (N_7698,N_5113,N_4298);
nor U7699 (N_7699,N_4261,N_4759);
nand U7700 (N_7700,N_3175,N_3131);
and U7701 (N_7701,N_5518,N_4609);
and U7702 (N_7702,N_4136,N_4161);
or U7703 (N_7703,N_4821,N_4867);
nor U7704 (N_7704,N_4272,N_4038);
nand U7705 (N_7705,N_5051,N_3767);
or U7706 (N_7706,N_5414,N_5177);
xor U7707 (N_7707,N_3686,N_5768);
nor U7708 (N_7708,N_4280,N_5131);
or U7709 (N_7709,N_4503,N_5079);
or U7710 (N_7710,N_4265,N_3287);
nand U7711 (N_7711,N_4876,N_4251);
or U7712 (N_7712,N_3717,N_3154);
nand U7713 (N_7713,N_5954,N_3323);
nand U7714 (N_7714,N_4660,N_4173);
nand U7715 (N_7715,N_4440,N_4984);
or U7716 (N_7716,N_3508,N_3837);
nand U7717 (N_7717,N_3904,N_5553);
and U7718 (N_7718,N_4963,N_4430);
or U7719 (N_7719,N_5249,N_5072);
nor U7720 (N_7720,N_5817,N_3196);
nand U7721 (N_7721,N_3974,N_4383);
nor U7722 (N_7722,N_4840,N_3892);
xor U7723 (N_7723,N_5156,N_3992);
or U7724 (N_7724,N_3235,N_3317);
or U7725 (N_7725,N_3769,N_5512);
or U7726 (N_7726,N_4338,N_4584);
or U7727 (N_7727,N_3406,N_3556);
or U7728 (N_7728,N_3185,N_3711);
or U7729 (N_7729,N_4369,N_4746);
and U7730 (N_7730,N_3100,N_5068);
and U7731 (N_7731,N_3138,N_3777);
or U7732 (N_7732,N_4989,N_3695);
nor U7733 (N_7733,N_5585,N_3435);
xor U7734 (N_7734,N_3809,N_5506);
or U7735 (N_7735,N_5664,N_4910);
nand U7736 (N_7736,N_3568,N_4240);
or U7737 (N_7737,N_4438,N_3591);
or U7738 (N_7738,N_3082,N_5663);
nor U7739 (N_7739,N_4579,N_5744);
and U7740 (N_7740,N_4924,N_3587);
or U7741 (N_7741,N_5587,N_5692);
and U7742 (N_7742,N_4767,N_5807);
nand U7743 (N_7743,N_5948,N_3698);
or U7744 (N_7744,N_4767,N_5044);
nor U7745 (N_7745,N_5216,N_4799);
and U7746 (N_7746,N_4374,N_4684);
and U7747 (N_7747,N_3554,N_3060);
nor U7748 (N_7748,N_3152,N_3483);
xnor U7749 (N_7749,N_3077,N_5852);
or U7750 (N_7750,N_5182,N_4538);
and U7751 (N_7751,N_3770,N_4181);
xor U7752 (N_7752,N_5310,N_5407);
and U7753 (N_7753,N_3114,N_4651);
and U7754 (N_7754,N_5854,N_3116);
and U7755 (N_7755,N_3326,N_3396);
nor U7756 (N_7756,N_5066,N_4088);
nand U7757 (N_7757,N_4251,N_5420);
or U7758 (N_7758,N_5819,N_5495);
or U7759 (N_7759,N_5146,N_3124);
and U7760 (N_7760,N_4025,N_5546);
or U7761 (N_7761,N_3225,N_4240);
nand U7762 (N_7762,N_3739,N_5957);
and U7763 (N_7763,N_4883,N_5864);
nor U7764 (N_7764,N_3287,N_4428);
or U7765 (N_7765,N_4222,N_5329);
xor U7766 (N_7766,N_3464,N_5147);
nor U7767 (N_7767,N_4053,N_4299);
xnor U7768 (N_7768,N_3939,N_4229);
or U7769 (N_7769,N_4498,N_5568);
or U7770 (N_7770,N_4487,N_5356);
nand U7771 (N_7771,N_5200,N_5575);
xor U7772 (N_7772,N_5115,N_3733);
nor U7773 (N_7773,N_5693,N_3256);
and U7774 (N_7774,N_4278,N_4006);
and U7775 (N_7775,N_3413,N_5765);
and U7776 (N_7776,N_3397,N_4874);
nor U7777 (N_7777,N_5673,N_4731);
nor U7778 (N_7778,N_3016,N_3539);
nor U7779 (N_7779,N_4485,N_5060);
and U7780 (N_7780,N_5978,N_4652);
nor U7781 (N_7781,N_3578,N_5657);
and U7782 (N_7782,N_5746,N_4106);
or U7783 (N_7783,N_5931,N_5554);
xor U7784 (N_7784,N_3375,N_5523);
xor U7785 (N_7785,N_5578,N_3604);
and U7786 (N_7786,N_4868,N_5315);
and U7787 (N_7787,N_5104,N_5999);
nand U7788 (N_7788,N_5684,N_4568);
or U7789 (N_7789,N_4814,N_3562);
nor U7790 (N_7790,N_3210,N_3881);
nand U7791 (N_7791,N_4092,N_5744);
and U7792 (N_7792,N_4409,N_4151);
and U7793 (N_7793,N_5106,N_3146);
and U7794 (N_7794,N_4994,N_3326);
xor U7795 (N_7795,N_5359,N_4134);
nor U7796 (N_7796,N_4337,N_4660);
and U7797 (N_7797,N_4680,N_4375);
and U7798 (N_7798,N_4620,N_4520);
nand U7799 (N_7799,N_4481,N_5475);
or U7800 (N_7800,N_5381,N_4157);
nor U7801 (N_7801,N_4000,N_3064);
and U7802 (N_7802,N_5934,N_5641);
nand U7803 (N_7803,N_3436,N_5950);
nor U7804 (N_7804,N_4491,N_4333);
or U7805 (N_7805,N_4790,N_3293);
and U7806 (N_7806,N_3273,N_5264);
xnor U7807 (N_7807,N_5092,N_5567);
and U7808 (N_7808,N_4767,N_3010);
or U7809 (N_7809,N_5969,N_5721);
and U7810 (N_7810,N_4044,N_4123);
or U7811 (N_7811,N_4549,N_3467);
xor U7812 (N_7812,N_5811,N_5507);
nor U7813 (N_7813,N_4585,N_5894);
or U7814 (N_7814,N_5978,N_3280);
and U7815 (N_7815,N_3102,N_3964);
or U7816 (N_7816,N_3542,N_4585);
nand U7817 (N_7817,N_5374,N_3954);
or U7818 (N_7818,N_4823,N_4109);
nand U7819 (N_7819,N_3922,N_3893);
or U7820 (N_7820,N_5263,N_4937);
nor U7821 (N_7821,N_5010,N_3391);
and U7822 (N_7822,N_5015,N_4994);
and U7823 (N_7823,N_4534,N_3554);
and U7824 (N_7824,N_5413,N_3909);
xor U7825 (N_7825,N_4078,N_4208);
nand U7826 (N_7826,N_3089,N_5930);
nor U7827 (N_7827,N_4604,N_4823);
and U7828 (N_7828,N_5188,N_4794);
and U7829 (N_7829,N_5211,N_3480);
nor U7830 (N_7830,N_5438,N_4717);
or U7831 (N_7831,N_3460,N_3025);
nand U7832 (N_7832,N_4095,N_4872);
nand U7833 (N_7833,N_5076,N_4185);
xnor U7834 (N_7834,N_3687,N_4497);
nand U7835 (N_7835,N_4292,N_4882);
and U7836 (N_7836,N_4165,N_5769);
nor U7837 (N_7837,N_5517,N_3860);
nand U7838 (N_7838,N_5867,N_4526);
or U7839 (N_7839,N_3514,N_3275);
and U7840 (N_7840,N_3279,N_5518);
nor U7841 (N_7841,N_5205,N_4340);
or U7842 (N_7842,N_3735,N_4194);
nor U7843 (N_7843,N_3983,N_3395);
xnor U7844 (N_7844,N_4174,N_3200);
nand U7845 (N_7845,N_5929,N_4680);
nor U7846 (N_7846,N_3224,N_4602);
nand U7847 (N_7847,N_3791,N_3091);
nor U7848 (N_7848,N_3825,N_3536);
nor U7849 (N_7849,N_5253,N_5317);
or U7850 (N_7850,N_4134,N_4937);
xor U7851 (N_7851,N_5971,N_4515);
nand U7852 (N_7852,N_5866,N_3338);
xor U7853 (N_7853,N_4117,N_4923);
nand U7854 (N_7854,N_3186,N_4163);
nor U7855 (N_7855,N_3989,N_5649);
xor U7856 (N_7856,N_3629,N_3229);
nor U7857 (N_7857,N_4458,N_5752);
xnor U7858 (N_7858,N_4286,N_5978);
or U7859 (N_7859,N_5046,N_5332);
nor U7860 (N_7860,N_3953,N_5777);
and U7861 (N_7861,N_3305,N_4212);
and U7862 (N_7862,N_5677,N_5597);
or U7863 (N_7863,N_5457,N_3174);
and U7864 (N_7864,N_5265,N_4433);
nor U7865 (N_7865,N_4782,N_5954);
or U7866 (N_7866,N_5701,N_3290);
nor U7867 (N_7867,N_4652,N_3132);
nand U7868 (N_7868,N_5662,N_3406);
and U7869 (N_7869,N_3916,N_3057);
or U7870 (N_7870,N_3468,N_5417);
nand U7871 (N_7871,N_3980,N_3858);
nand U7872 (N_7872,N_3680,N_5870);
or U7873 (N_7873,N_3103,N_4061);
nand U7874 (N_7874,N_5877,N_5193);
xnor U7875 (N_7875,N_5659,N_5571);
nor U7876 (N_7876,N_4135,N_4477);
and U7877 (N_7877,N_4631,N_5870);
nand U7878 (N_7878,N_3595,N_5312);
or U7879 (N_7879,N_3256,N_5120);
xnor U7880 (N_7880,N_4600,N_4736);
nand U7881 (N_7881,N_5456,N_4970);
nand U7882 (N_7882,N_5525,N_3743);
or U7883 (N_7883,N_3833,N_3997);
and U7884 (N_7884,N_4783,N_3062);
nand U7885 (N_7885,N_4624,N_5474);
nor U7886 (N_7886,N_3980,N_4696);
or U7887 (N_7887,N_5304,N_3369);
and U7888 (N_7888,N_5100,N_3293);
nor U7889 (N_7889,N_3008,N_3720);
nor U7890 (N_7890,N_3300,N_3522);
nand U7891 (N_7891,N_4398,N_5039);
nor U7892 (N_7892,N_3723,N_4627);
nor U7893 (N_7893,N_4350,N_3800);
or U7894 (N_7894,N_4795,N_3570);
and U7895 (N_7895,N_4506,N_3638);
nand U7896 (N_7896,N_4905,N_4454);
nand U7897 (N_7897,N_4433,N_3570);
and U7898 (N_7898,N_5583,N_4673);
nand U7899 (N_7899,N_5873,N_3293);
and U7900 (N_7900,N_4587,N_4437);
nor U7901 (N_7901,N_3063,N_4459);
or U7902 (N_7902,N_5861,N_4978);
nor U7903 (N_7903,N_3024,N_4673);
nor U7904 (N_7904,N_5155,N_4451);
xor U7905 (N_7905,N_4263,N_4722);
nor U7906 (N_7906,N_4138,N_5402);
and U7907 (N_7907,N_5796,N_4969);
and U7908 (N_7908,N_3202,N_4064);
nor U7909 (N_7909,N_3260,N_5820);
or U7910 (N_7910,N_3127,N_3393);
nor U7911 (N_7911,N_3511,N_4318);
and U7912 (N_7912,N_3599,N_3863);
and U7913 (N_7913,N_5325,N_3725);
nand U7914 (N_7914,N_5720,N_5226);
and U7915 (N_7915,N_4186,N_4091);
or U7916 (N_7916,N_4889,N_5446);
and U7917 (N_7917,N_5283,N_3309);
and U7918 (N_7918,N_3832,N_3759);
xnor U7919 (N_7919,N_3857,N_4425);
or U7920 (N_7920,N_3018,N_5263);
and U7921 (N_7921,N_3390,N_4709);
nand U7922 (N_7922,N_3362,N_4647);
nor U7923 (N_7923,N_4224,N_3119);
and U7924 (N_7924,N_3402,N_4591);
nor U7925 (N_7925,N_3365,N_3257);
nand U7926 (N_7926,N_3561,N_5812);
nor U7927 (N_7927,N_5030,N_5376);
nor U7928 (N_7928,N_4682,N_5837);
nor U7929 (N_7929,N_3400,N_3804);
nand U7930 (N_7930,N_3777,N_4083);
or U7931 (N_7931,N_4952,N_3858);
nor U7932 (N_7932,N_5354,N_5048);
nor U7933 (N_7933,N_4737,N_4817);
nor U7934 (N_7934,N_5828,N_3561);
xnor U7935 (N_7935,N_4733,N_4830);
and U7936 (N_7936,N_4276,N_3156);
nand U7937 (N_7937,N_5439,N_4554);
or U7938 (N_7938,N_3575,N_5835);
nand U7939 (N_7939,N_5731,N_5525);
and U7940 (N_7940,N_5974,N_4212);
nor U7941 (N_7941,N_3710,N_5933);
nand U7942 (N_7942,N_4534,N_4593);
nor U7943 (N_7943,N_3890,N_3279);
nor U7944 (N_7944,N_3843,N_5783);
nand U7945 (N_7945,N_5483,N_5121);
or U7946 (N_7946,N_5748,N_3195);
nor U7947 (N_7947,N_4732,N_5849);
and U7948 (N_7948,N_3031,N_5312);
and U7949 (N_7949,N_4966,N_4327);
nor U7950 (N_7950,N_3705,N_4293);
nor U7951 (N_7951,N_5668,N_3016);
and U7952 (N_7952,N_5710,N_4213);
nand U7953 (N_7953,N_5285,N_3888);
xor U7954 (N_7954,N_3289,N_4737);
nor U7955 (N_7955,N_5908,N_4874);
nand U7956 (N_7956,N_4072,N_4765);
xor U7957 (N_7957,N_3837,N_5300);
or U7958 (N_7958,N_5305,N_5939);
nor U7959 (N_7959,N_4142,N_3073);
nand U7960 (N_7960,N_5192,N_5333);
and U7961 (N_7961,N_3117,N_3551);
and U7962 (N_7962,N_4209,N_4541);
or U7963 (N_7963,N_5446,N_5043);
and U7964 (N_7964,N_4205,N_3730);
nor U7965 (N_7965,N_5746,N_5951);
or U7966 (N_7966,N_5782,N_4690);
and U7967 (N_7967,N_4424,N_5379);
or U7968 (N_7968,N_5072,N_5300);
or U7969 (N_7969,N_5911,N_5917);
nor U7970 (N_7970,N_3782,N_5988);
nand U7971 (N_7971,N_4242,N_3432);
nor U7972 (N_7972,N_4284,N_4391);
and U7973 (N_7973,N_3949,N_4432);
or U7974 (N_7974,N_4543,N_4183);
or U7975 (N_7975,N_4694,N_5297);
nor U7976 (N_7976,N_4404,N_3304);
nand U7977 (N_7977,N_4006,N_3997);
nand U7978 (N_7978,N_3020,N_5054);
nand U7979 (N_7979,N_3462,N_4321);
and U7980 (N_7980,N_5026,N_4687);
or U7981 (N_7981,N_5146,N_4350);
nand U7982 (N_7982,N_4746,N_3102);
xor U7983 (N_7983,N_4031,N_3748);
and U7984 (N_7984,N_5285,N_3871);
or U7985 (N_7985,N_4882,N_5231);
and U7986 (N_7986,N_5147,N_3033);
nand U7987 (N_7987,N_3576,N_3285);
xor U7988 (N_7988,N_3158,N_4803);
nand U7989 (N_7989,N_5643,N_3751);
nor U7990 (N_7990,N_3758,N_4439);
nand U7991 (N_7991,N_3279,N_5333);
nor U7992 (N_7992,N_4676,N_3719);
and U7993 (N_7993,N_3200,N_5384);
nand U7994 (N_7994,N_4562,N_5425);
nor U7995 (N_7995,N_4514,N_4591);
and U7996 (N_7996,N_5009,N_3967);
nand U7997 (N_7997,N_4696,N_3910);
nor U7998 (N_7998,N_3944,N_3283);
and U7999 (N_7999,N_5713,N_4577);
and U8000 (N_8000,N_4859,N_3469);
or U8001 (N_8001,N_4601,N_5901);
and U8002 (N_8002,N_5772,N_3149);
nand U8003 (N_8003,N_3138,N_3225);
nor U8004 (N_8004,N_3426,N_5038);
nand U8005 (N_8005,N_4249,N_3884);
and U8006 (N_8006,N_3290,N_4175);
nand U8007 (N_8007,N_5778,N_3906);
or U8008 (N_8008,N_3385,N_4015);
or U8009 (N_8009,N_3657,N_3426);
nand U8010 (N_8010,N_4922,N_4270);
and U8011 (N_8011,N_5337,N_5425);
and U8012 (N_8012,N_4116,N_5849);
nor U8013 (N_8013,N_4249,N_4757);
and U8014 (N_8014,N_5001,N_5842);
nand U8015 (N_8015,N_5100,N_4293);
nor U8016 (N_8016,N_5996,N_4869);
nor U8017 (N_8017,N_5985,N_4232);
nand U8018 (N_8018,N_5147,N_4517);
or U8019 (N_8019,N_5946,N_5378);
nor U8020 (N_8020,N_3848,N_5556);
nor U8021 (N_8021,N_4584,N_5018);
xor U8022 (N_8022,N_3167,N_5064);
nand U8023 (N_8023,N_5300,N_5902);
xnor U8024 (N_8024,N_5317,N_4928);
nor U8025 (N_8025,N_3899,N_5373);
or U8026 (N_8026,N_3472,N_4343);
nor U8027 (N_8027,N_5138,N_3316);
xor U8028 (N_8028,N_5766,N_3182);
nand U8029 (N_8029,N_5547,N_4872);
or U8030 (N_8030,N_5118,N_5319);
nand U8031 (N_8031,N_3865,N_5660);
or U8032 (N_8032,N_5376,N_4614);
and U8033 (N_8033,N_5997,N_4807);
nand U8034 (N_8034,N_3050,N_5071);
nand U8035 (N_8035,N_4707,N_4524);
and U8036 (N_8036,N_3169,N_4193);
and U8037 (N_8037,N_5285,N_4211);
nor U8038 (N_8038,N_3267,N_4282);
nor U8039 (N_8039,N_3813,N_3740);
and U8040 (N_8040,N_3686,N_5191);
xor U8041 (N_8041,N_5340,N_5443);
nor U8042 (N_8042,N_5198,N_4261);
or U8043 (N_8043,N_3559,N_5613);
and U8044 (N_8044,N_3028,N_3851);
or U8045 (N_8045,N_3901,N_3333);
nand U8046 (N_8046,N_5421,N_4520);
nand U8047 (N_8047,N_3836,N_5125);
xor U8048 (N_8048,N_5384,N_5913);
xnor U8049 (N_8049,N_5794,N_4860);
or U8050 (N_8050,N_3009,N_4613);
xnor U8051 (N_8051,N_4966,N_3121);
nor U8052 (N_8052,N_5409,N_5081);
nand U8053 (N_8053,N_5727,N_4649);
or U8054 (N_8054,N_3189,N_4810);
nor U8055 (N_8055,N_3959,N_5477);
or U8056 (N_8056,N_4863,N_5866);
nor U8057 (N_8057,N_3162,N_3831);
nor U8058 (N_8058,N_4854,N_3708);
nand U8059 (N_8059,N_4718,N_3776);
nor U8060 (N_8060,N_3529,N_4747);
nor U8061 (N_8061,N_4334,N_5815);
nor U8062 (N_8062,N_5288,N_5198);
nor U8063 (N_8063,N_5133,N_4983);
or U8064 (N_8064,N_5204,N_5977);
and U8065 (N_8065,N_4008,N_4005);
or U8066 (N_8066,N_4386,N_5078);
and U8067 (N_8067,N_4748,N_5856);
nand U8068 (N_8068,N_5029,N_5766);
nand U8069 (N_8069,N_5910,N_3125);
or U8070 (N_8070,N_5232,N_5865);
nand U8071 (N_8071,N_4998,N_4850);
or U8072 (N_8072,N_4682,N_4646);
nand U8073 (N_8073,N_5838,N_4974);
nor U8074 (N_8074,N_5940,N_4396);
nor U8075 (N_8075,N_3257,N_5022);
nor U8076 (N_8076,N_3045,N_3439);
nor U8077 (N_8077,N_3691,N_5660);
nand U8078 (N_8078,N_4843,N_5311);
nor U8079 (N_8079,N_3750,N_5989);
nor U8080 (N_8080,N_3410,N_5841);
xnor U8081 (N_8081,N_5258,N_3920);
and U8082 (N_8082,N_3967,N_3932);
nor U8083 (N_8083,N_4665,N_5340);
nor U8084 (N_8084,N_4993,N_3077);
nor U8085 (N_8085,N_4038,N_5533);
or U8086 (N_8086,N_5327,N_4145);
nor U8087 (N_8087,N_3538,N_3087);
or U8088 (N_8088,N_4744,N_3694);
nor U8089 (N_8089,N_4491,N_5856);
and U8090 (N_8090,N_4821,N_4271);
or U8091 (N_8091,N_5332,N_5162);
nor U8092 (N_8092,N_3811,N_3401);
or U8093 (N_8093,N_4697,N_5552);
or U8094 (N_8094,N_5485,N_3492);
nor U8095 (N_8095,N_4238,N_4726);
and U8096 (N_8096,N_3693,N_3536);
nor U8097 (N_8097,N_5894,N_3860);
nor U8098 (N_8098,N_4330,N_5342);
and U8099 (N_8099,N_5949,N_5546);
nand U8100 (N_8100,N_4699,N_5775);
nand U8101 (N_8101,N_3849,N_3833);
nor U8102 (N_8102,N_4043,N_5530);
or U8103 (N_8103,N_5853,N_3913);
xor U8104 (N_8104,N_5308,N_3513);
or U8105 (N_8105,N_4148,N_4205);
and U8106 (N_8106,N_4654,N_5118);
or U8107 (N_8107,N_5332,N_4161);
and U8108 (N_8108,N_3201,N_3980);
and U8109 (N_8109,N_3567,N_4884);
xor U8110 (N_8110,N_4143,N_5806);
nand U8111 (N_8111,N_5167,N_3180);
or U8112 (N_8112,N_3746,N_4345);
nand U8113 (N_8113,N_3823,N_4331);
nand U8114 (N_8114,N_3286,N_5961);
xor U8115 (N_8115,N_4687,N_4408);
and U8116 (N_8116,N_4887,N_5989);
or U8117 (N_8117,N_4870,N_3611);
nand U8118 (N_8118,N_4906,N_3784);
or U8119 (N_8119,N_3401,N_5705);
nand U8120 (N_8120,N_5588,N_3810);
nor U8121 (N_8121,N_3872,N_5299);
nor U8122 (N_8122,N_3585,N_3321);
nor U8123 (N_8123,N_3970,N_4454);
or U8124 (N_8124,N_5461,N_5571);
or U8125 (N_8125,N_5826,N_5533);
or U8126 (N_8126,N_3906,N_3008);
and U8127 (N_8127,N_4028,N_5433);
or U8128 (N_8128,N_3247,N_5301);
or U8129 (N_8129,N_4671,N_3590);
nand U8130 (N_8130,N_5313,N_4823);
nand U8131 (N_8131,N_4368,N_5035);
nor U8132 (N_8132,N_5883,N_4812);
and U8133 (N_8133,N_5661,N_5973);
and U8134 (N_8134,N_3561,N_5408);
nand U8135 (N_8135,N_5575,N_5973);
nand U8136 (N_8136,N_3243,N_3042);
or U8137 (N_8137,N_4048,N_4084);
and U8138 (N_8138,N_5169,N_4169);
nor U8139 (N_8139,N_5095,N_3453);
or U8140 (N_8140,N_5376,N_5469);
nor U8141 (N_8141,N_5128,N_3353);
and U8142 (N_8142,N_5675,N_3027);
or U8143 (N_8143,N_5471,N_4409);
or U8144 (N_8144,N_3167,N_5164);
or U8145 (N_8145,N_5346,N_3675);
and U8146 (N_8146,N_3702,N_4461);
nand U8147 (N_8147,N_3645,N_3466);
nand U8148 (N_8148,N_5877,N_4594);
nand U8149 (N_8149,N_4594,N_3667);
and U8150 (N_8150,N_4617,N_5632);
nor U8151 (N_8151,N_5016,N_5783);
nand U8152 (N_8152,N_5235,N_3479);
nand U8153 (N_8153,N_3632,N_4851);
or U8154 (N_8154,N_4176,N_4739);
and U8155 (N_8155,N_5095,N_5854);
and U8156 (N_8156,N_4491,N_4298);
nor U8157 (N_8157,N_3710,N_5949);
and U8158 (N_8158,N_3028,N_3804);
and U8159 (N_8159,N_4743,N_4492);
nor U8160 (N_8160,N_5028,N_3068);
or U8161 (N_8161,N_3406,N_3976);
nor U8162 (N_8162,N_4987,N_5783);
nor U8163 (N_8163,N_5106,N_3445);
nor U8164 (N_8164,N_4324,N_3769);
or U8165 (N_8165,N_4797,N_4988);
or U8166 (N_8166,N_5788,N_5197);
and U8167 (N_8167,N_5529,N_3632);
or U8168 (N_8168,N_5598,N_5200);
nor U8169 (N_8169,N_4641,N_5642);
or U8170 (N_8170,N_5287,N_3436);
nor U8171 (N_8171,N_3272,N_5482);
or U8172 (N_8172,N_4745,N_4637);
nand U8173 (N_8173,N_4523,N_3104);
nor U8174 (N_8174,N_4928,N_5525);
nor U8175 (N_8175,N_5924,N_4106);
or U8176 (N_8176,N_4708,N_4559);
or U8177 (N_8177,N_3874,N_4779);
nor U8178 (N_8178,N_3900,N_4419);
nor U8179 (N_8179,N_4544,N_4546);
and U8180 (N_8180,N_5895,N_3580);
or U8181 (N_8181,N_4855,N_4846);
or U8182 (N_8182,N_5939,N_3555);
or U8183 (N_8183,N_4351,N_5106);
nor U8184 (N_8184,N_5904,N_4731);
xnor U8185 (N_8185,N_4578,N_5754);
nor U8186 (N_8186,N_5752,N_5312);
nand U8187 (N_8187,N_4762,N_4620);
nor U8188 (N_8188,N_5439,N_5793);
and U8189 (N_8189,N_4681,N_4256);
or U8190 (N_8190,N_5981,N_3586);
nor U8191 (N_8191,N_4080,N_5767);
nor U8192 (N_8192,N_4093,N_4397);
nand U8193 (N_8193,N_5937,N_3870);
nand U8194 (N_8194,N_4192,N_4892);
and U8195 (N_8195,N_5707,N_4656);
nor U8196 (N_8196,N_4175,N_4575);
and U8197 (N_8197,N_3861,N_4005);
nor U8198 (N_8198,N_5663,N_5058);
xor U8199 (N_8199,N_5780,N_4716);
or U8200 (N_8200,N_4268,N_5963);
nand U8201 (N_8201,N_5291,N_5063);
or U8202 (N_8202,N_3470,N_5281);
and U8203 (N_8203,N_3733,N_3883);
and U8204 (N_8204,N_4803,N_5117);
nor U8205 (N_8205,N_5970,N_5992);
xnor U8206 (N_8206,N_3865,N_3663);
nor U8207 (N_8207,N_5437,N_3747);
nor U8208 (N_8208,N_3968,N_4170);
xnor U8209 (N_8209,N_4295,N_4159);
nand U8210 (N_8210,N_4329,N_3291);
nand U8211 (N_8211,N_5426,N_3057);
and U8212 (N_8212,N_3143,N_5258);
nor U8213 (N_8213,N_4016,N_3654);
or U8214 (N_8214,N_5178,N_5442);
nand U8215 (N_8215,N_4448,N_4318);
nand U8216 (N_8216,N_4254,N_5064);
nand U8217 (N_8217,N_4194,N_3767);
and U8218 (N_8218,N_5523,N_5824);
and U8219 (N_8219,N_3662,N_3103);
or U8220 (N_8220,N_3510,N_5305);
and U8221 (N_8221,N_4457,N_4786);
or U8222 (N_8222,N_4743,N_4262);
or U8223 (N_8223,N_5334,N_5941);
xnor U8224 (N_8224,N_3455,N_3281);
and U8225 (N_8225,N_4352,N_3722);
nand U8226 (N_8226,N_3057,N_4369);
nand U8227 (N_8227,N_5563,N_3277);
or U8228 (N_8228,N_4817,N_5743);
nand U8229 (N_8229,N_3379,N_5911);
and U8230 (N_8230,N_3459,N_3489);
or U8231 (N_8231,N_4060,N_5762);
nand U8232 (N_8232,N_4757,N_3075);
or U8233 (N_8233,N_3250,N_5670);
nand U8234 (N_8234,N_5529,N_3805);
nand U8235 (N_8235,N_5620,N_4594);
xor U8236 (N_8236,N_3656,N_5036);
and U8237 (N_8237,N_3681,N_4316);
nor U8238 (N_8238,N_5348,N_5504);
xor U8239 (N_8239,N_4163,N_5189);
nor U8240 (N_8240,N_3562,N_3216);
and U8241 (N_8241,N_3967,N_5668);
or U8242 (N_8242,N_3751,N_3814);
and U8243 (N_8243,N_4046,N_5784);
xnor U8244 (N_8244,N_5930,N_3942);
xnor U8245 (N_8245,N_4343,N_3575);
nor U8246 (N_8246,N_4770,N_5095);
and U8247 (N_8247,N_3117,N_5320);
and U8248 (N_8248,N_3629,N_4869);
xor U8249 (N_8249,N_3117,N_5527);
or U8250 (N_8250,N_3022,N_4081);
xnor U8251 (N_8251,N_4800,N_4352);
nor U8252 (N_8252,N_5512,N_3288);
nand U8253 (N_8253,N_3649,N_4000);
or U8254 (N_8254,N_3941,N_3036);
nand U8255 (N_8255,N_4729,N_4717);
and U8256 (N_8256,N_3896,N_5195);
nand U8257 (N_8257,N_5590,N_3897);
nor U8258 (N_8258,N_3224,N_3851);
nor U8259 (N_8259,N_3529,N_5640);
nand U8260 (N_8260,N_3587,N_3239);
and U8261 (N_8261,N_4099,N_4013);
nand U8262 (N_8262,N_5665,N_5536);
nand U8263 (N_8263,N_4866,N_4960);
nand U8264 (N_8264,N_3737,N_5062);
nor U8265 (N_8265,N_5369,N_4370);
xor U8266 (N_8266,N_3416,N_5562);
nor U8267 (N_8267,N_5661,N_5279);
nor U8268 (N_8268,N_5069,N_3221);
or U8269 (N_8269,N_5677,N_5862);
nor U8270 (N_8270,N_4613,N_3510);
nand U8271 (N_8271,N_3835,N_5190);
nand U8272 (N_8272,N_5692,N_5287);
nand U8273 (N_8273,N_3293,N_3579);
and U8274 (N_8274,N_5804,N_3654);
and U8275 (N_8275,N_5986,N_3553);
xor U8276 (N_8276,N_3258,N_5100);
or U8277 (N_8277,N_3409,N_4735);
and U8278 (N_8278,N_5617,N_4994);
or U8279 (N_8279,N_5887,N_3888);
and U8280 (N_8280,N_3131,N_5028);
or U8281 (N_8281,N_5000,N_5989);
nand U8282 (N_8282,N_4536,N_3754);
and U8283 (N_8283,N_4015,N_3802);
and U8284 (N_8284,N_3263,N_4121);
nor U8285 (N_8285,N_4253,N_5630);
and U8286 (N_8286,N_3118,N_3262);
or U8287 (N_8287,N_3184,N_3523);
nor U8288 (N_8288,N_4553,N_5981);
nor U8289 (N_8289,N_5823,N_4040);
xnor U8290 (N_8290,N_4733,N_4013);
nand U8291 (N_8291,N_5611,N_3812);
xor U8292 (N_8292,N_4006,N_5687);
and U8293 (N_8293,N_5272,N_3227);
or U8294 (N_8294,N_3621,N_3120);
nor U8295 (N_8295,N_4430,N_3682);
or U8296 (N_8296,N_3289,N_5483);
and U8297 (N_8297,N_3153,N_5406);
nor U8298 (N_8298,N_3783,N_5795);
and U8299 (N_8299,N_5009,N_4440);
and U8300 (N_8300,N_4551,N_3463);
xor U8301 (N_8301,N_3062,N_5746);
nand U8302 (N_8302,N_4155,N_4407);
nand U8303 (N_8303,N_3112,N_3901);
xnor U8304 (N_8304,N_3576,N_3556);
nor U8305 (N_8305,N_5338,N_5035);
nand U8306 (N_8306,N_4997,N_5784);
nor U8307 (N_8307,N_4755,N_3225);
or U8308 (N_8308,N_3793,N_4330);
or U8309 (N_8309,N_4004,N_4840);
or U8310 (N_8310,N_5972,N_3835);
nor U8311 (N_8311,N_4793,N_5268);
nor U8312 (N_8312,N_3159,N_4803);
xnor U8313 (N_8313,N_5529,N_4751);
or U8314 (N_8314,N_4032,N_5474);
nand U8315 (N_8315,N_3961,N_4356);
and U8316 (N_8316,N_3596,N_4581);
nand U8317 (N_8317,N_4678,N_3268);
and U8318 (N_8318,N_4219,N_3932);
nor U8319 (N_8319,N_4568,N_4988);
nor U8320 (N_8320,N_3719,N_3117);
nor U8321 (N_8321,N_5100,N_4471);
nor U8322 (N_8322,N_4507,N_4246);
nor U8323 (N_8323,N_4931,N_5337);
and U8324 (N_8324,N_3029,N_3491);
and U8325 (N_8325,N_4220,N_4982);
or U8326 (N_8326,N_4590,N_5066);
nand U8327 (N_8327,N_5921,N_4309);
nor U8328 (N_8328,N_5028,N_4502);
nor U8329 (N_8329,N_4735,N_5560);
or U8330 (N_8330,N_4463,N_3865);
or U8331 (N_8331,N_5411,N_4604);
and U8332 (N_8332,N_3950,N_5590);
and U8333 (N_8333,N_4099,N_5817);
or U8334 (N_8334,N_4843,N_4557);
or U8335 (N_8335,N_4005,N_4728);
nand U8336 (N_8336,N_5196,N_4856);
and U8337 (N_8337,N_3196,N_4761);
xnor U8338 (N_8338,N_4677,N_3216);
nand U8339 (N_8339,N_3430,N_4302);
xor U8340 (N_8340,N_3471,N_3988);
nor U8341 (N_8341,N_5201,N_5785);
or U8342 (N_8342,N_4696,N_3387);
and U8343 (N_8343,N_3190,N_5325);
and U8344 (N_8344,N_5536,N_5383);
xor U8345 (N_8345,N_4605,N_3720);
or U8346 (N_8346,N_4940,N_4309);
and U8347 (N_8347,N_5744,N_4510);
nand U8348 (N_8348,N_5154,N_3735);
or U8349 (N_8349,N_4485,N_5419);
xor U8350 (N_8350,N_4221,N_4929);
nand U8351 (N_8351,N_4432,N_4048);
nand U8352 (N_8352,N_4566,N_4797);
or U8353 (N_8353,N_3683,N_5105);
or U8354 (N_8354,N_4426,N_4838);
nand U8355 (N_8355,N_3052,N_4167);
nand U8356 (N_8356,N_3180,N_4420);
and U8357 (N_8357,N_5218,N_4560);
or U8358 (N_8358,N_4686,N_5301);
or U8359 (N_8359,N_5907,N_4253);
or U8360 (N_8360,N_4948,N_5353);
and U8361 (N_8361,N_3074,N_5418);
nor U8362 (N_8362,N_4051,N_3689);
nand U8363 (N_8363,N_4476,N_3879);
nand U8364 (N_8364,N_3703,N_5974);
or U8365 (N_8365,N_5281,N_4838);
nand U8366 (N_8366,N_5327,N_4864);
nand U8367 (N_8367,N_4388,N_4418);
nor U8368 (N_8368,N_3919,N_4224);
or U8369 (N_8369,N_5213,N_5671);
nand U8370 (N_8370,N_4524,N_4587);
or U8371 (N_8371,N_3249,N_3460);
nand U8372 (N_8372,N_3636,N_5043);
and U8373 (N_8373,N_5049,N_4917);
and U8374 (N_8374,N_3641,N_4773);
nand U8375 (N_8375,N_5287,N_3092);
and U8376 (N_8376,N_4323,N_3319);
nor U8377 (N_8377,N_5278,N_4427);
nor U8378 (N_8378,N_4209,N_3562);
nand U8379 (N_8379,N_4148,N_3003);
and U8380 (N_8380,N_3186,N_5725);
nand U8381 (N_8381,N_5333,N_4856);
or U8382 (N_8382,N_4401,N_5858);
or U8383 (N_8383,N_4697,N_3554);
or U8384 (N_8384,N_4342,N_3000);
and U8385 (N_8385,N_3068,N_3476);
or U8386 (N_8386,N_4503,N_4208);
and U8387 (N_8387,N_5601,N_3667);
or U8388 (N_8388,N_4804,N_3401);
and U8389 (N_8389,N_3258,N_3426);
or U8390 (N_8390,N_4155,N_5473);
nand U8391 (N_8391,N_3182,N_3882);
xnor U8392 (N_8392,N_3972,N_3472);
or U8393 (N_8393,N_3438,N_5281);
and U8394 (N_8394,N_5810,N_3594);
nor U8395 (N_8395,N_4543,N_4954);
xor U8396 (N_8396,N_3384,N_4547);
nor U8397 (N_8397,N_5051,N_3970);
or U8398 (N_8398,N_5060,N_5434);
nor U8399 (N_8399,N_4833,N_3411);
nor U8400 (N_8400,N_3876,N_5141);
and U8401 (N_8401,N_4386,N_4823);
and U8402 (N_8402,N_5142,N_3325);
xor U8403 (N_8403,N_3285,N_3073);
nor U8404 (N_8404,N_5064,N_4258);
or U8405 (N_8405,N_5281,N_4101);
and U8406 (N_8406,N_4845,N_4763);
and U8407 (N_8407,N_4404,N_5415);
xor U8408 (N_8408,N_5236,N_4667);
or U8409 (N_8409,N_5138,N_3258);
or U8410 (N_8410,N_5149,N_5096);
xnor U8411 (N_8411,N_4359,N_5042);
nand U8412 (N_8412,N_4331,N_5975);
or U8413 (N_8413,N_5170,N_3896);
or U8414 (N_8414,N_4402,N_4644);
nand U8415 (N_8415,N_5158,N_4203);
and U8416 (N_8416,N_3430,N_5351);
nor U8417 (N_8417,N_4534,N_4999);
nor U8418 (N_8418,N_3279,N_5071);
or U8419 (N_8419,N_3388,N_5535);
nand U8420 (N_8420,N_3875,N_5762);
nand U8421 (N_8421,N_4177,N_4596);
or U8422 (N_8422,N_3570,N_5329);
and U8423 (N_8423,N_3282,N_5749);
and U8424 (N_8424,N_3360,N_4814);
nand U8425 (N_8425,N_5994,N_4533);
xnor U8426 (N_8426,N_4519,N_5907);
and U8427 (N_8427,N_5734,N_5404);
nor U8428 (N_8428,N_3408,N_3601);
xor U8429 (N_8429,N_5572,N_4027);
nor U8430 (N_8430,N_3612,N_3437);
and U8431 (N_8431,N_5956,N_4084);
nand U8432 (N_8432,N_5457,N_4602);
nor U8433 (N_8433,N_4893,N_3095);
nor U8434 (N_8434,N_3734,N_3042);
or U8435 (N_8435,N_4925,N_5359);
and U8436 (N_8436,N_5022,N_4994);
nor U8437 (N_8437,N_5606,N_5160);
or U8438 (N_8438,N_5590,N_5604);
nand U8439 (N_8439,N_4081,N_4880);
nor U8440 (N_8440,N_4651,N_3426);
and U8441 (N_8441,N_4366,N_5771);
and U8442 (N_8442,N_5761,N_5852);
xnor U8443 (N_8443,N_4212,N_4353);
or U8444 (N_8444,N_3759,N_4682);
nand U8445 (N_8445,N_5452,N_4436);
or U8446 (N_8446,N_5946,N_3365);
nor U8447 (N_8447,N_3201,N_5551);
nand U8448 (N_8448,N_5902,N_3902);
nand U8449 (N_8449,N_3287,N_5554);
and U8450 (N_8450,N_4432,N_4316);
and U8451 (N_8451,N_4185,N_4127);
or U8452 (N_8452,N_5851,N_5359);
nand U8453 (N_8453,N_5197,N_3391);
or U8454 (N_8454,N_4232,N_5713);
xnor U8455 (N_8455,N_5298,N_5471);
and U8456 (N_8456,N_5748,N_5298);
nand U8457 (N_8457,N_5555,N_3590);
and U8458 (N_8458,N_3402,N_5426);
xor U8459 (N_8459,N_5269,N_3021);
and U8460 (N_8460,N_3028,N_3013);
nor U8461 (N_8461,N_5172,N_3317);
and U8462 (N_8462,N_4931,N_5664);
nand U8463 (N_8463,N_4566,N_4735);
xor U8464 (N_8464,N_4233,N_3408);
xnor U8465 (N_8465,N_3687,N_5854);
nor U8466 (N_8466,N_3261,N_3995);
and U8467 (N_8467,N_5535,N_4783);
or U8468 (N_8468,N_4820,N_5742);
nand U8469 (N_8469,N_5126,N_3869);
xor U8470 (N_8470,N_5415,N_5593);
and U8471 (N_8471,N_3722,N_3830);
xor U8472 (N_8472,N_5755,N_4063);
nor U8473 (N_8473,N_4271,N_4527);
nor U8474 (N_8474,N_3001,N_4490);
or U8475 (N_8475,N_5721,N_3817);
nor U8476 (N_8476,N_4797,N_5345);
nand U8477 (N_8477,N_5175,N_3290);
or U8478 (N_8478,N_4840,N_5229);
nor U8479 (N_8479,N_5989,N_5474);
or U8480 (N_8480,N_3264,N_4774);
nor U8481 (N_8481,N_4304,N_3756);
xor U8482 (N_8482,N_3185,N_5739);
nor U8483 (N_8483,N_5823,N_5339);
and U8484 (N_8484,N_5833,N_5143);
nor U8485 (N_8485,N_4456,N_5741);
and U8486 (N_8486,N_5122,N_3020);
or U8487 (N_8487,N_4663,N_4492);
nand U8488 (N_8488,N_5758,N_4043);
and U8489 (N_8489,N_3192,N_5596);
and U8490 (N_8490,N_5577,N_4718);
and U8491 (N_8491,N_3528,N_3086);
nand U8492 (N_8492,N_4942,N_4083);
or U8493 (N_8493,N_4291,N_5528);
or U8494 (N_8494,N_4070,N_4686);
nor U8495 (N_8495,N_3198,N_4586);
or U8496 (N_8496,N_5955,N_4763);
or U8497 (N_8497,N_4042,N_3293);
nand U8498 (N_8498,N_5016,N_5872);
xor U8499 (N_8499,N_3917,N_5958);
nand U8500 (N_8500,N_5148,N_5074);
nand U8501 (N_8501,N_5897,N_5902);
xnor U8502 (N_8502,N_3883,N_3350);
xor U8503 (N_8503,N_4351,N_3127);
or U8504 (N_8504,N_4065,N_5278);
nand U8505 (N_8505,N_4850,N_5033);
and U8506 (N_8506,N_3373,N_4113);
and U8507 (N_8507,N_3700,N_5079);
and U8508 (N_8508,N_4286,N_3874);
nor U8509 (N_8509,N_5356,N_5941);
or U8510 (N_8510,N_4742,N_3285);
or U8511 (N_8511,N_5940,N_5950);
nand U8512 (N_8512,N_4224,N_5571);
and U8513 (N_8513,N_5716,N_4072);
nor U8514 (N_8514,N_5983,N_4158);
nor U8515 (N_8515,N_4993,N_5621);
and U8516 (N_8516,N_5052,N_5482);
nor U8517 (N_8517,N_5200,N_3010);
and U8518 (N_8518,N_5646,N_3149);
or U8519 (N_8519,N_3025,N_5542);
nor U8520 (N_8520,N_3012,N_4696);
or U8521 (N_8521,N_3232,N_4486);
or U8522 (N_8522,N_3272,N_4321);
and U8523 (N_8523,N_5486,N_5818);
xor U8524 (N_8524,N_5659,N_3880);
or U8525 (N_8525,N_5362,N_3281);
nand U8526 (N_8526,N_4474,N_4084);
nand U8527 (N_8527,N_4767,N_3216);
and U8528 (N_8528,N_4170,N_5008);
nand U8529 (N_8529,N_3259,N_4574);
or U8530 (N_8530,N_4202,N_4347);
nor U8531 (N_8531,N_3319,N_4985);
and U8532 (N_8532,N_4522,N_3094);
or U8533 (N_8533,N_5895,N_3496);
or U8534 (N_8534,N_5571,N_5602);
nand U8535 (N_8535,N_3839,N_4993);
nand U8536 (N_8536,N_3349,N_5642);
nor U8537 (N_8537,N_4916,N_4764);
and U8538 (N_8538,N_5365,N_4371);
nand U8539 (N_8539,N_4257,N_4745);
or U8540 (N_8540,N_4467,N_4585);
nor U8541 (N_8541,N_4292,N_3266);
nand U8542 (N_8542,N_3272,N_5795);
nor U8543 (N_8543,N_5810,N_5157);
nand U8544 (N_8544,N_4923,N_3674);
xor U8545 (N_8545,N_4004,N_3208);
and U8546 (N_8546,N_3095,N_3749);
and U8547 (N_8547,N_5562,N_5475);
and U8548 (N_8548,N_3037,N_5067);
nand U8549 (N_8549,N_3948,N_3022);
xnor U8550 (N_8550,N_5081,N_3079);
or U8551 (N_8551,N_4580,N_5127);
or U8552 (N_8552,N_3905,N_3713);
nor U8553 (N_8553,N_4471,N_3071);
or U8554 (N_8554,N_4014,N_4363);
nand U8555 (N_8555,N_4325,N_3644);
nand U8556 (N_8556,N_3189,N_3351);
nor U8557 (N_8557,N_3983,N_3732);
nand U8558 (N_8558,N_5296,N_5889);
nor U8559 (N_8559,N_3241,N_3851);
nor U8560 (N_8560,N_3548,N_3528);
nand U8561 (N_8561,N_5451,N_5740);
and U8562 (N_8562,N_3027,N_4342);
and U8563 (N_8563,N_3421,N_4279);
and U8564 (N_8564,N_5397,N_5496);
and U8565 (N_8565,N_3697,N_5208);
or U8566 (N_8566,N_3759,N_5919);
nand U8567 (N_8567,N_3456,N_4019);
and U8568 (N_8568,N_3625,N_3737);
xnor U8569 (N_8569,N_3677,N_5178);
nor U8570 (N_8570,N_4528,N_5054);
and U8571 (N_8571,N_4150,N_5570);
nor U8572 (N_8572,N_4519,N_5029);
and U8573 (N_8573,N_5583,N_4177);
or U8574 (N_8574,N_5693,N_4193);
and U8575 (N_8575,N_5885,N_3954);
or U8576 (N_8576,N_4169,N_3829);
or U8577 (N_8577,N_5416,N_3774);
xnor U8578 (N_8578,N_5958,N_3366);
nand U8579 (N_8579,N_4821,N_3793);
nor U8580 (N_8580,N_3393,N_4737);
or U8581 (N_8581,N_4163,N_5385);
nand U8582 (N_8582,N_5148,N_5828);
and U8583 (N_8583,N_5995,N_3924);
and U8584 (N_8584,N_4557,N_5015);
nand U8585 (N_8585,N_3671,N_5157);
nor U8586 (N_8586,N_3146,N_3395);
and U8587 (N_8587,N_4061,N_4011);
nor U8588 (N_8588,N_4139,N_4374);
or U8589 (N_8589,N_5446,N_5756);
nor U8590 (N_8590,N_3341,N_5039);
and U8591 (N_8591,N_4308,N_4103);
nor U8592 (N_8592,N_3158,N_3555);
xnor U8593 (N_8593,N_3463,N_5080);
or U8594 (N_8594,N_3278,N_3999);
xnor U8595 (N_8595,N_5312,N_5916);
and U8596 (N_8596,N_3757,N_5632);
nand U8597 (N_8597,N_4599,N_5703);
and U8598 (N_8598,N_4733,N_3440);
or U8599 (N_8599,N_4896,N_4452);
nor U8600 (N_8600,N_4604,N_3402);
and U8601 (N_8601,N_3382,N_4997);
or U8602 (N_8602,N_3999,N_5714);
or U8603 (N_8603,N_3793,N_5264);
nand U8604 (N_8604,N_4074,N_4658);
nor U8605 (N_8605,N_4044,N_4752);
and U8606 (N_8606,N_5300,N_4303);
xor U8607 (N_8607,N_5497,N_5566);
and U8608 (N_8608,N_4150,N_4745);
nor U8609 (N_8609,N_4713,N_4192);
nor U8610 (N_8610,N_5003,N_3214);
or U8611 (N_8611,N_5111,N_4624);
or U8612 (N_8612,N_5950,N_3741);
and U8613 (N_8613,N_5481,N_5222);
or U8614 (N_8614,N_5680,N_4571);
nand U8615 (N_8615,N_5258,N_4996);
or U8616 (N_8616,N_5685,N_4303);
nor U8617 (N_8617,N_5723,N_4148);
nor U8618 (N_8618,N_3270,N_5873);
xor U8619 (N_8619,N_5598,N_5297);
nand U8620 (N_8620,N_5011,N_3979);
xnor U8621 (N_8621,N_4475,N_5367);
xor U8622 (N_8622,N_5230,N_3509);
or U8623 (N_8623,N_5880,N_3238);
nor U8624 (N_8624,N_4434,N_5220);
nand U8625 (N_8625,N_5873,N_4121);
or U8626 (N_8626,N_3541,N_3963);
or U8627 (N_8627,N_5902,N_3430);
and U8628 (N_8628,N_5302,N_4535);
nand U8629 (N_8629,N_4088,N_5271);
and U8630 (N_8630,N_4886,N_5106);
xor U8631 (N_8631,N_3887,N_5444);
nor U8632 (N_8632,N_3039,N_4835);
nand U8633 (N_8633,N_3765,N_3991);
or U8634 (N_8634,N_4497,N_5839);
nor U8635 (N_8635,N_5736,N_5216);
or U8636 (N_8636,N_4540,N_3927);
nand U8637 (N_8637,N_3264,N_5183);
and U8638 (N_8638,N_5354,N_5585);
nor U8639 (N_8639,N_4731,N_5876);
nor U8640 (N_8640,N_4885,N_4634);
nor U8641 (N_8641,N_4831,N_4520);
or U8642 (N_8642,N_5049,N_5462);
nor U8643 (N_8643,N_3488,N_4871);
and U8644 (N_8644,N_4860,N_4770);
nor U8645 (N_8645,N_4203,N_3113);
and U8646 (N_8646,N_3897,N_5828);
and U8647 (N_8647,N_5053,N_3239);
and U8648 (N_8648,N_3977,N_3374);
and U8649 (N_8649,N_5393,N_4717);
and U8650 (N_8650,N_4567,N_4185);
nand U8651 (N_8651,N_3765,N_4751);
and U8652 (N_8652,N_4261,N_4336);
and U8653 (N_8653,N_5535,N_3769);
nor U8654 (N_8654,N_5074,N_4279);
nand U8655 (N_8655,N_4612,N_4723);
nand U8656 (N_8656,N_4407,N_5289);
nor U8657 (N_8657,N_5527,N_3473);
nand U8658 (N_8658,N_4388,N_3333);
and U8659 (N_8659,N_3800,N_3763);
nand U8660 (N_8660,N_3471,N_4774);
nor U8661 (N_8661,N_3983,N_5892);
and U8662 (N_8662,N_4754,N_3076);
nor U8663 (N_8663,N_3137,N_3683);
or U8664 (N_8664,N_4781,N_4846);
nor U8665 (N_8665,N_5293,N_5393);
and U8666 (N_8666,N_3193,N_3106);
nor U8667 (N_8667,N_4561,N_5788);
nand U8668 (N_8668,N_3299,N_5197);
and U8669 (N_8669,N_5855,N_3383);
nand U8670 (N_8670,N_4709,N_4556);
nand U8671 (N_8671,N_4829,N_4006);
and U8672 (N_8672,N_3569,N_3860);
nor U8673 (N_8673,N_4843,N_4336);
and U8674 (N_8674,N_3471,N_5263);
and U8675 (N_8675,N_4746,N_5818);
and U8676 (N_8676,N_3933,N_5370);
and U8677 (N_8677,N_4472,N_5709);
and U8678 (N_8678,N_5047,N_4578);
and U8679 (N_8679,N_3695,N_4611);
nand U8680 (N_8680,N_3801,N_5411);
nand U8681 (N_8681,N_3016,N_4471);
xnor U8682 (N_8682,N_5296,N_3434);
and U8683 (N_8683,N_5753,N_4881);
and U8684 (N_8684,N_4161,N_3443);
nand U8685 (N_8685,N_4104,N_4175);
nor U8686 (N_8686,N_3645,N_4081);
xnor U8687 (N_8687,N_4398,N_4167);
nand U8688 (N_8688,N_4050,N_4693);
and U8689 (N_8689,N_5284,N_5299);
nand U8690 (N_8690,N_3111,N_4158);
nand U8691 (N_8691,N_3158,N_3191);
or U8692 (N_8692,N_4657,N_4904);
nor U8693 (N_8693,N_3407,N_4519);
or U8694 (N_8694,N_3759,N_5679);
nor U8695 (N_8695,N_5041,N_3206);
and U8696 (N_8696,N_5651,N_4899);
nand U8697 (N_8697,N_4938,N_4172);
nor U8698 (N_8698,N_3915,N_5704);
and U8699 (N_8699,N_3842,N_3109);
and U8700 (N_8700,N_4077,N_5037);
and U8701 (N_8701,N_5036,N_4273);
and U8702 (N_8702,N_4250,N_4970);
xnor U8703 (N_8703,N_5096,N_5679);
nand U8704 (N_8704,N_4821,N_5667);
and U8705 (N_8705,N_5880,N_4106);
xor U8706 (N_8706,N_5607,N_4775);
and U8707 (N_8707,N_4482,N_4692);
or U8708 (N_8708,N_3497,N_5493);
or U8709 (N_8709,N_5628,N_4917);
or U8710 (N_8710,N_4099,N_4237);
nor U8711 (N_8711,N_4221,N_3774);
nor U8712 (N_8712,N_4366,N_3844);
nand U8713 (N_8713,N_4223,N_3874);
nand U8714 (N_8714,N_3768,N_4670);
nand U8715 (N_8715,N_4884,N_3634);
and U8716 (N_8716,N_5517,N_5707);
nor U8717 (N_8717,N_3920,N_4718);
or U8718 (N_8718,N_3178,N_5809);
and U8719 (N_8719,N_5857,N_3657);
or U8720 (N_8720,N_3682,N_5323);
or U8721 (N_8721,N_3055,N_3914);
xor U8722 (N_8722,N_3186,N_3848);
nand U8723 (N_8723,N_3404,N_4564);
xor U8724 (N_8724,N_4995,N_3535);
nand U8725 (N_8725,N_3764,N_5681);
or U8726 (N_8726,N_4102,N_3097);
nor U8727 (N_8727,N_3494,N_5974);
xor U8728 (N_8728,N_4315,N_4462);
and U8729 (N_8729,N_3190,N_5997);
and U8730 (N_8730,N_5412,N_3488);
nand U8731 (N_8731,N_4261,N_5005);
and U8732 (N_8732,N_3477,N_4594);
nand U8733 (N_8733,N_3080,N_3348);
nand U8734 (N_8734,N_5386,N_3104);
nand U8735 (N_8735,N_4151,N_4740);
and U8736 (N_8736,N_5687,N_4181);
nor U8737 (N_8737,N_3788,N_3109);
xor U8738 (N_8738,N_4090,N_3057);
nor U8739 (N_8739,N_4407,N_3374);
or U8740 (N_8740,N_3263,N_4061);
xor U8741 (N_8741,N_3470,N_3376);
xor U8742 (N_8742,N_5193,N_4098);
or U8743 (N_8743,N_3132,N_5313);
and U8744 (N_8744,N_4928,N_4424);
nor U8745 (N_8745,N_3635,N_5115);
and U8746 (N_8746,N_3630,N_4731);
nor U8747 (N_8747,N_5754,N_3027);
or U8748 (N_8748,N_3506,N_3049);
nor U8749 (N_8749,N_5453,N_5311);
and U8750 (N_8750,N_4535,N_5749);
and U8751 (N_8751,N_5562,N_5481);
nand U8752 (N_8752,N_3465,N_5864);
or U8753 (N_8753,N_4131,N_3672);
or U8754 (N_8754,N_4012,N_3662);
nand U8755 (N_8755,N_4269,N_3004);
nor U8756 (N_8756,N_3293,N_5551);
and U8757 (N_8757,N_5838,N_3006);
xor U8758 (N_8758,N_5164,N_3643);
nor U8759 (N_8759,N_4446,N_4340);
nand U8760 (N_8760,N_3236,N_4837);
nand U8761 (N_8761,N_3246,N_5566);
xor U8762 (N_8762,N_5627,N_5202);
and U8763 (N_8763,N_3087,N_5671);
nand U8764 (N_8764,N_3172,N_5896);
and U8765 (N_8765,N_5000,N_5732);
and U8766 (N_8766,N_4939,N_4034);
or U8767 (N_8767,N_5458,N_4490);
and U8768 (N_8768,N_4948,N_4859);
or U8769 (N_8769,N_4252,N_5973);
and U8770 (N_8770,N_3868,N_5002);
nand U8771 (N_8771,N_3235,N_3115);
or U8772 (N_8772,N_4920,N_5964);
nand U8773 (N_8773,N_5684,N_5872);
and U8774 (N_8774,N_4984,N_4049);
nand U8775 (N_8775,N_4643,N_4010);
nand U8776 (N_8776,N_5301,N_5716);
or U8777 (N_8777,N_5451,N_3780);
nand U8778 (N_8778,N_5081,N_3353);
and U8779 (N_8779,N_5233,N_4877);
or U8780 (N_8780,N_5951,N_4003);
or U8781 (N_8781,N_3461,N_4719);
or U8782 (N_8782,N_3791,N_4375);
or U8783 (N_8783,N_5559,N_4307);
xor U8784 (N_8784,N_3315,N_4191);
nor U8785 (N_8785,N_3406,N_5865);
nor U8786 (N_8786,N_4609,N_4544);
and U8787 (N_8787,N_4089,N_3938);
and U8788 (N_8788,N_3325,N_3856);
nor U8789 (N_8789,N_3513,N_3237);
nand U8790 (N_8790,N_3336,N_4813);
nor U8791 (N_8791,N_5011,N_4348);
and U8792 (N_8792,N_5452,N_3719);
nor U8793 (N_8793,N_3797,N_4175);
nor U8794 (N_8794,N_4399,N_4559);
or U8795 (N_8795,N_5282,N_4948);
and U8796 (N_8796,N_4462,N_3578);
nor U8797 (N_8797,N_3062,N_5321);
and U8798 (N_8798,N_4129,N_3783);
and U8799 (N_8799,N_4334,N_4603);
and U8800 (N_8800,N_3895,N_3084);
and U8801 (N_8801,N_4627,N_5833);
and U8802 (N_8802,N_4967,N_4425);
or U8803 (N_8803,N_3273,N_5714);
nand U8804 (N_8804,N_4481,N_4557);
nand U8805 (N_8805,N_4980,N_3000);
nand U8806 (N_8806,N_4731,N_5136);
nand U8807 (N_8807,N_3614,N_4741);
nor U8808 (N_8808,N_4092,N_3631);
nand U8809 (N_8809,N_3747,N_3256);
and U8810 (N_8810,N_5894,N_3039);
or U8811 (N_8811,N_3230,N_4736);
nor U8812 (N_8812,N_3341,N_4149);
or U8813 (N_8813,N_3399,N_5766);
and U8814 (N_8814,N_3675,N_4027);
nand U8815 (N_8815,N_5897,N_5564);
nor U8816 (N_8816,N_4415,N_4989);
and U8817 (N_8817,N_3746,N_3005);
nand U8818 (N_8818,N_4259,N_4655);
or U8819 (N_8819,N_5785,N_3774);
and U8820 (N_8820,N_4112,N_5874);
or U8821 (N_8821,N_5142,N_5732);
nor U8822 (N_8822,N_3267,N_5101);
or U8823 (N_8823,N_4201,N_3317);
nor U8824 (N_8824,N_3909,N_4223);
or U8825 (N_8825,N_3909,N_5272);
nand U8826 (N_8826,N_3434,N_5474);
and U8827 (N_8827,N_3688,N_5350);
and U8828 (N_8828,N_5645,N_4759);
or U8829 (N_8829,N_5061,N_3233);
nor U8830 (N_8830,N_4157,N_5763);
or U8831 (N_8831,N_4905,N_5735);
xor U8832 (N_8832,N_4386,N_4202);
nor U8833 (N_8833,N_4012,N_3757);
nor U8834 (N_8834,N_5943,N_3228);
nand U8835 (N_8835,N_4657,N_5778);
or U8836 (N_8836,N_4825,N_5224);
or U8837 (N_8837,N_5974,N_3452);
or U8838 (N_8838,N_4127,N_4176);
nor U8839 (N_8839,N_4529,N_4953);
nand U8840 (N_8840,N_5647,N_4779);
nor U8841 (N_8841,N_5370,N_4709);
xor U8842 (N_8842,N_3638,N_4166);
and U8843 (N_8843,N_5589,N_5166);
or U8844 (N_8844,N_5379,N_5188);
xor U8845 (N_8845,N_3817,N_4149);
nand U8846 (N_8846,N_4941,N_3908);
or U8847 (N_8847,N_5625,N_5807);
nor U8848 (N_8848,N_4414,N_3360);
nand U8849 (N_8849,N_3653,N_5976);
xor U8850 (N_8850,N_5771,N_3415);
nor U8851 (N_8851,N_4993,N_3216);
or U8852 (N_8852,N_5019,N_5729);
or U8853 (N_8853,N_5701,N_5095);
and U8854 (N_8854,N_3664,N_5083);
or U8855 (N_8855,N_3105,N_5539);
or U8856 (N_8856,N_3329,N_3138);
or U8857 (N_8857,N_3095,N_3262);
nand U8858 (N_8858,N_5872,N_3069);
xor U8859 (N_8859,N_5843,N_5784);
and U8860 (N_8860,N_3287,N_3608);
nand U8861 (N_8861,N_4306,N_5795);
or U8862 (N_8862,N_3211,N_3539);
nand U8863 (N_8863,N_3225,N_4949);
or U8864 (N_8864,N_5412,N_3169);
or U8865 (N_8865,N_3538,N_4231);
nor U8866 (N_8866,N_4666,N_4538);
nand U8867 (N_8867,N_4739,N_4880);
and U8868 (N_8868,N_3229,N_5619);
or U8869 (N_8869,N_5640,N_4637);
and U8870 (N_8870,N_5040,N_5284);
and U8871 (N_8871,N_4229,N_4207);
and U8872 (N_8872,N_5476,N_3649);
and U8873 (N_8873,N_4364,N_4954);
xor U8874 (N_8874,N_3947,N_5040);
nand U8875 (N_8875,N_3374,N_4385);
nand U8876 (N_8876,N_5354,N_4681);
or U8877 (N_8877,N_4615,N_5645);
xor U8878 (N_8878,N_4862,N_3478);
or U8879 (N_8879,N_4727,N_5158);
or U8880 (N_8880,N_5601,N_3210);
nor U8881 (N_8881,N_5639,N_4992);
xor U8882 (N_8882,N_4156,N_3402);
xnor U8883 (N_8883,N_5605,N_3488);
nor U8884 (N_8884,N_3779,N_5805);
nand U8885 (N_8885,N_4795,N_3950);
and U8886 (N_8886,N_3275,N_5068);
or U8887 (N_8887,N_3262,N_5842);
or U8888 (N_8888,N_3397,N_3875);
nor U8889 (N_8889,N_3889,N_5586);
or U8890 (N_8890,N_4793,N_3076);
nor U8891 (N_8891,N_5330,N_4383);
or U8892 (N_8892,N_4195,N_3846);
or U8893 (N_8893,N_3635,N_5866);
nand U8894 (N_8894,N_3202,N_4296);
nand U8895 (N_8895,N_4094,N_5297);
nand U8896 (N_8896,N_3938,N_5510);
or U8897 (N_8897,N_3252,N_4183);
or U8898 (N_8898,N_3198,N_3088);
or U8899 (N_8899,N_5797,N_4998);
and U8900 (N_8900,N_4385,N_3301);
or U8901 (N_8901,N_3784,N_3499);
or U8902 (N_8902,N_4316,N_3430);
nand U8903 (N_8903,N_4897,N_5451);
and U8904 (N_8904,N_3967,N_5464);
or U8905 (N_8905,N_3463,N_5475);
and U8906 (N_8906,N_4424,N_5944);
nand U8907 (N_8907,N_4018,N_4342);
or U8908 (N_8908,N_5984,N_3655);
and U8909 (N_8909,N_5794,N_3343);
and U8910 (N_8910,N_4622,N_4750);
xor U8911 (N_8911,N_5409,N_4545);
xor U8912 (N_8912,N_3308,N_5761);
nand U8913 (N_8913,N_3652,N_4115);
and U8914 (N_8914,N_4636,N_4159);
nand U8915 (N_8915,N_4334,N_3652);
and U8916 (N_8916,N_5130,N_3678);
nand U8917 (N_8917,N_3138,N_3931);
or U8918 (N_8918,N_5706,N_3762);
nor U8919 (N_8919,N_3016,N_3870);
nor U8920 (N_8920,N_3318,N_5987);
and U8921 (N_8921,N_5633,N_3218);
and U8922 (N_8922,N_3817,N_4988);
and U8923 (N_8923,N_5998,N_4907);
nand U8924 (N_8924,N_4149,N_5401);
and U8925 (N_8925,N_4523,N_4563);
and U8926 (N_8926,N_5893,N_3019);
and U8927 (N_8927,N_4214,N_5165);
or U8928 (N_8928,N_3125,N_3676);
nor U8929 (N_8929,N_3087,N_3602);
nor U8930 (N_8930,N_3067,N_5909);
xor U8931 (N_8931,N_4275,N_5616);
or U8932 (N_8932,N_3499,N_3878);
nor U8933 (N_8933,N_3435,N_3742);
xnor U8934 (N_8934,N_4525,N_4355);
nor U8935 (N_8935,N_3428,N_4154);
and U8936 (N_8936,N_4388,N_3668);
and U8937 (N_8937,N_4914,N_4238);
nor U8938 (N_8938,N_3525,N_5246);
nor U8939 (N_8939,N_5987,N_5136);
and U8940 (N_8940,N_4901,N_3194);
and U8941 (N_8941,N_3150,N_5952);
nand U8942 (N_8942,N_4941,N_5079);
or U8943 (N_8943,N_3397,N_5005);
and U8944 (N_8944,N_3452,N_4946);
nand U8945 (N_8945,N_4804,N_3884);
xnor U8946 (N_8946,N_3841,N_3057);
nand U8947 (N_8947,N_4539,N_4252);
or U8948 (N_8948,N_3506,N_5424);
nor U8949 (N_8949,N_3836,N_4075);
or U8950 (N_8950,N_4381,N_3876);
and U8951 (N_8951,N_3779,N_3737);
and U8952 (N_8952,N_5259,N_3416);
or U8953 (N_8953,N_3424,N_4838);
or U8954 (N_8954,N_3601,N_5983);
nand U8955 (N_8955,N_3567,N_4349);
nand U8956 (N_8956,N_5090,N_4113);
or U8957 (N_8957,N_3674,N_4820);
or U8958 (N_8958,N_5074,N_3175);
nand U8959 (N_8959,N_4031,N_3393);
nand U8960 (N_8960,N_5013,N_4684);
and U8961 (N_8961,N_3589,N_5152);
nor U8962 (N_8962,N_3981,N_5552);
xnor U8963 (N_8963,N_5812,N_4041);
nand U8964 (N_8964,N_5703,N_3655);
and U8965 (N_8965,N_3287,N_3396);
nor U8966 (N_8966,N_4909,N_3472);
nand U8967 (N_8967,N_4152,N_3601);
and U8968 (N_8968,N_4045,N_3948);
or U8969 (N_8969,N_4317,N_5662);
nor U8970 (N_8970,N_5539,N_4850);
or U8971 (N_8971,N_3404,N_4870);
and U8972 (N_8972,N_5733,N_3583);
or U8973 (N_8973,N_5303,N_3740);
nand U8974 (N_8974,N_5778,N_3504);
nand U8975 (N_8975,N_5740,N_3726);
nand U8976 (N_8976,N_3552,N_3661);
or U8977 (N_8977,N_5740,N_4006);
or U8978 (N_8978,N_3804,N_4144);
nand U8979 (N_8979,N_5276,N_5889);
nand U8980 (N_8980,N_5437,N_3602);
nand U8981 (N_8981,N_5890,N_5996);
nand U8982 (N_8982,N_3693,N_3587);
and U8983 (N_8983,N_5426,N_4662);
nor U8984 (N_8984,N_4001,N_3409);
nand U8985 (N_8985,N_3521,N_5760);
nand U8986 (N_8986,N_5556,N_5593);
and U8987 (N_8987,N_3997,N_5486);
nor U8988 (N_8988,N_4223,N_4281);
nor U8989 (N_8989,N_3753,N_4707);
and U8990 (N_8990,N_4638,N_4596);
nor U8991 (N_8991,N_5412,N_4379);
nor U8992 (N_8992,N_3848,N_3424);
nand U8993 (N_8993,N_4577,N_5289);
nor U8994 (N_8994,N_3670,N_3644);
nand U8995 (N_8995,N_4224,N_4072);
or U8996 (N_8996,N_4426,N_4233);
xnor U8997 (N_8997,N_4053,N_5851);
nor U8998 (N_8998,N_3949,N_5136);
or U8999 (N_8999,N_4138,N_5327);
or U9000 (N_9000,N_7704,N_6089);
nand U9001 (N_9001,N_6642,N_8402);
nand U9002 (N_9002,N_6180,N_6674);
or U9003 (N_9003,N_8354,N_7083);
and U9004 (N_9004,N_7631,N_7254);
and U9005 (N_9005,N_8740,N_8092);
and U9006 (N_9006,N_7817,N_6799);
or U9007 (N_9007,N_7085,N_8657);
or U9008 (N_9008,N_6067,N_8477);
xor U9009 (N_9009,N_8855,N_7033);
and U9010 (N_9010,N_8864,N_7217);
and U9011 (N_9011,N_8704,N_6195);
nor U9012 (N_9012,N_6033,N_6850);
and U9013 (N_9013,N_7000,N_6316);
nor U9014 (N_9014,N_6554,N_8427);
nand U9015 (N_9015,N_7749,N_6958);
and U9016 (N_9016,N_7393,N_8062);
and U9017 (N_9017,N_8885,N_8533);
nand U9018 (N_9018,N_6189,N_7331);
and U9019 (N_9019,N_7663,N_7606);
xor U9020 (N_9020,N_7414,N_7781);
and U9021 (N_9021,N_8504,N_8975);
nand U9022 (N_9022,N_8482,N_6348);
or U9023 (N_9023,N_8136,N_8023);
or U9024 (N_9024,N_8996,N_6226);
nand U9025 (N_9025,N_6061,N_8626);
xnor U9026 (N_9026,N_8033,N_7601);
or U9027 (N_9027,N_7994,N_8258);
nand U9028 (N_9028,N_8526,N_7947);
or U9029 (N_9029,N_6974,N_6950);
or U9030 (N_9030,N_6599,N_6752);
nand U9031 (N_9031,N_6279,N_7437);
nor U9032 (N_9032,N_8237,N_8946);
nand U9033 (N_9033,N_7482,N_7481);
xor U9034 (N_9034,N_8254,N_8791);
nor U9035 (N_9035,N_7826,N_8490);
nand U9036 (N_9036,N_6526,N_6838);
or U9037 (N_9037,N_6987,N_6614);
or U9038 (N_9038,N_6429,N_7005);
or U9039 (N_9039,N_7539,N_6314);
nand U9040 (N_9040,N_7181,N_8038);
or U9041 (N_9041,N_6182,N_7889);
nor U9042 (N_9042,N_7777,N_7304);
nand U9043 (N_9043,N_6567,N_6106);
nand U9044 (N_9044,N_7291,N_7837);
or U9045 (N_9045,N_8350,N_6294);
and U9046 (N_9046,N_7792,N_8901);
and U9047 (N_9047,N_8164,N_8966);
nor U9048 (N_9048,N_6233,N_7941);
nand U9049 (N_9049,N_7712,N_6703);
nand U9050 (N_9050,N_8824,N_8424);
xnor U9051 (N_9051,N_6630,N_6946);
nand U9052 (N_9052,N_8681,N_6980);
and U9053 (N_9053,N_6051,N_6865);
xnor U9054 (N_9054,N_8257,N_8869);
nand U9055 (N_9055,N_6737,N_8381);
or U9056 (N_9056,N_6011,N_6345);
xnor U9057 (N_9057,N_7988,N_7840);
or U9058 (N_9058,N_7132,N_7533);
nor U9059 (N_9059,N_6172,N_8884);
nand U9060 (N_9060,N_8573,N_8319);
or U9061 (N_9061,N_6660,N_6307);
or U9062 (N_9062,N_6343,N_7557);
xnor U9063 (N_9063,N_7963,N_8637);
xor U9064 (N_9064,N_7905,N_8069);
nand U9065 (N_9065,N_8801,N_7330);
nor U9066 (N_9066,N_8478,N_6449);
or U9067 (N_9067,N_8135,N_7850);
and U9068 (N_9068,N_7469,N_6286);
and U9069 (N_9069,N_6517,N_7411);
nor U9070 (N_9070,N_8588,N_6330);
xnor U9071 (N_9071,N_6009,N_8882);
nand U9072 (N_9072,N_7268,N_8090);
or U9073 (N_9073,N_7412,N_7078);
or U9074 (N_9074,N_7435,N_8894);
nor U9075 (N_9075,N_8779,N_6112);
nand U9076 (N_9076,N_7324,N_8611);
nor U9077 (N_9077,N_8969,N_7667);
or U9078 (N_9078,N_8234,N_6891);
or U9079 (N_9079,N_6717,N_8925);
nand U9080 (N_9080,N_6159,N_8857);
or U9081 (N_9081,N_8875,N_7306);
or U9082 (N_9082,N_7483,N_8302);
xor U9083 (N_9083,N_8455,N_7086);
xnor U9084 (N_9084,N_7782,N_7389);
nor U9085 (N_9085,N_6149,N_7733);
nand U9086 (N_9086,N_6275,N_6028);
xnor U9087 (N_9087,N_8182,N_7114);
nor U9088 (N_9088,N_6693,N_8728);
xor U9089 (N_9089,N_6131,N_6624);
and U9090 (N_9090,N_8244,N_6486);
or U9091 (N_9091,N_8191,N_7929);
nand U9092 (N_9092,N_8432,N_7658);
nor U9093 (N_9093,N_8229,N_8660);
or U9094 (N_9094,N_6967,N_8685);
and U9095 (N_9095,N_8199,N_8390);
nor U9096 (N_9096,N_6218,N_7462);
or U9097 (N_9097,N_6476,N_8138);
and U9098 (N_9098,N_8070,N_6601);
or U9099 (N_9099,N_7346,N_6962);
or U9100 (N_9100,N_8224,N_7451);
and U9101 (N_9101,N_6473,N_7368);
nand U9102 (N_9102,N_7496,N_8297);
nor U9103 (N_9103,N_7099,N_6368);
nand U9104 (N_9104,N_7823,N_7727);
and U9105 (N_9105,N_7651,N_6075);
nand U9106 (N_9106,N_7904,N_6653);
or U9107 (N_9107,N_8389,N_6474);
and U9108 (N_9108,N_8643,N_8718);
or U9109 (N_9109,N_8453,N_8775);
or U9110 (N_9110,N_7380,N_7997);
nor U9111 (N_9111,N_7774,N_6032);
nor U9112 (N_9112,N_6750,N_8345);
and U9113 (N_9113,N_7731,N_7550);
or U9114 (N_9114,N_7418,N_8896);
nor U9115 (N_9115,N_6446,N_8930);
nand U9116 (N_9116,N_8145,N_7366);
xnor U9117 (N_9117,N_8418,N_7476);
or U9118 (N_9118,N_7685,N_8113);
nor U9119 (N_9119,N_8711,N_6856);
nor U9120 (N_9120,N_8906,N_8167);
or U9121 (N_9121,N_6467,N_6217);
nor U9122 (N_9122,N_8835,N_6022);
xor U9123 (N_9123,N_6543,N_7620);
or U9124 (N_9124,N_6827,N_7864);
nor U9125 (N_9125,N_7130,N_6125);
nor U9126 (N_9126,N_7416,N_6049);
or U9127 (N_9127,N_6949,N_7137);
xnor U9128 (N_9128,N_6768,N_6230);
nand U9129 (N_9129,N_8570,N_7543);
nor U9130 (N_9130,N_6825,N_7236);
or U9131 (N_9131,N_6315,N_7421);
nor U9132 (N_9132,N_6214,N_6928);
nand U9133 (N_9133,N_8587,N_6966);
xnor U9134 (N_9134,N_8359,N_6886);
xor U9135 (N_9135,N_7926,N_8408);
xnor U9136 (N_9136,N_7135,N_6899);
nor U9137 (N_9137,N_8933,N_6727);
nor U9138 (N_9138,N_6686,N_7394);
xnor U9139 (N_9139,N_7068,N_8115);
nor U9140 (N_9140,N_7711,N_6885);
xor U9141 (N_9141,N_8180,N_8619);
nand U9142 (N_9142,N_8541,N_8509);
nor U9143 (N_9143,N_6124,N_6138);
and U9144 (N_9144,N_8238,N_6837);
nor U9145 (N_9145,N_6421,N_8093);
nor U9146 (N_9146,N_7252,N_7795);
nand U9147 (N_9147,N_7095,N_6143);
or U9148 (N_9148,N_7800,N_6789);
nor U9149 (N_9149,N_6834,N_8014);
and U9150 (N_9150,N_8656,N_6568);
or U9151 (N_9151,N_7454,N_6258);
and U9152 (N_9152,N_8365,N_7742);
or U9153 (N_9153,N_8442,N_7398);
and U9154 (N_9154,N_6297,N_8688);
nand U9155 (N_9155,N_8374,N_8571);
nand U9156 (N_9156,N_7561,N_7503);
and U9157 (N_9157,N_8220,N_7057);
nand U9158 (N_9158,N_8591,N_6097);
or U9159 (N_9159,N_6764,N_8963);
or U9160 (N_9160,N_8039,N_6020);
nor U9161 (N_9161,N_7653,N_7403);
xor U9162 (N_9162,N_6540,N_8780);
and U9163 (N_9163,N_7261,N_8843);
nand U9164 (N_9164,N_8705,N_8452);
nand U9165 (N_9165,N_6362,N_7447);
and U9166 (N_9166,N_6785,N_6771);
and U9167 (N_9167,N_6809,N_7419);
nand U9168 (N_9168,N_7689,N_7635);
nand U9169 (N_9169,N_8753,N_6426);
or U9170 (N_9170,N_7626,N_6744);
xnor U9171 (N_9171,N_7449,N_7359);
or U9172 (N_9172,N_8123,N_7450);
or U9173 (N_9173,N_6623,N_8841);
and U9174 (N_9174,N_7344,N_7280);
nor U9175 (N_9175,N_8461,N_8269);
nor U9176 (N_9176,N_7713,N_6448);
nand U9177 (N_9177,N_6773,N_7211);
nand U9178 (N_9178,N_6171,N_6493);
and U9179 (N_9179,N_6321,N_6581);
and U9180 (N_9180,N_8814,N_7783);
nand U9181 (N_9181,N_8782,N_6589);
nor U9182 (N_9182,N_7453,N_8179);
and U9183 (N_9183,N_8472,N_8595);
xnor U9184 (N_9184,N_6821,N_7102);
nand U9185 (N_9185,N_8513,N_7319);
nor U9186 (N_9186,N_7479,N_7071);
and U9187 (N_9187,N_6290,N_7004);
nor U9188 (N_9188,N_7231,N_6205);
or U9189 (N_9189,N_6973,N_8967);
and U9190 (N_9190,N_8076,N_8936);
and U9191 (N_9191,N_6084,N_8306);
or U9192 (N_9192,N_7870,N_8948);
and U9193 (N_9193,N_7722,N_7410);
xor U9194 (N_9194,N_8264,N_8926);
xor U9195 (N_9195,N_8360,N_8883);
or U9196 (N_9196,N_8808,N_6369);
nand U9197 (N_9197,N_7015,N_7556);
nand U9198 (N_9198,N_6453,N_6519);
or U9199 (N_9199,N_7846,N_7311);
or U9200 (N_9200,N_8233,N_8682);
nand U9201 (N_9201,N_7659,N_6720);
nor U9202 (N_9202,N_6266,N_8899);
or U9203 (N_9203,N_6298,N_6847);
or U9204 (N_9204,N_6144,N_8734);
and U9205 (N_9205,N_7853,N_8912);
and U9206 (N_9206,N_7661,N_7180);
xnor U9207 (N_9207,N_6137,N_8805);
xor U9208 (N_9208,N_8056,N_8828);
nand U9209 (N_9209,N_8804,N_6168);
nor U9210 (N_9210,N_6541,N_6129);
nor U9211 (N_9211,N_8286,N_8386);
and U9212 (N_9212,N_6603,N_7519);
nor U9213 (N_9213,N_8772,N_7644);
or U9214 (N_9214,N_7420,N_7726);
and U9215 (N_9215,N_8543,N_7176);
nand U9216 (N_9216,N_8836,N_8152);
and U9217 (N_9217,N_6412,N_7750);
nor U9218 (N_9218,N_7467,N_7505);
or U9219 (N_9219,N_8760,N_6238);
and U9220 (N_9220,N_8289,N_8583);
nand U9221 (N_9221,N_6695,N_8677);
nand U9222 (N_9222,N_6547,N_6350);
nor U9223 (N_9223,N_7353,N_7526);
nand U9224 (N_9224,N_7401,N_8582);
or U9225 (N_9225,N_7300,N_6497);
and U9226 (N_9226,N_7248,N_8029);
or U9227 (N_9227,N_6518,N_7002);
xor U9228 (N_9228,N_6659,N_7232);
and U9229 (N_9229,N_8341,N_7347);
or U9230 (N_9230,N_7212,N_8785);
xnor U9231 (N_9231,N_7869,N_8003);
nor U9232 (N_9232,N_7725,N_6701);
nor U9233 (N_9233,N_7534,N_7513);
or U9234 (N_9234,N_6783,N_6499);
or U9235 (N_9235,N_7547,N_7703);
or U9236 (N_9236,N_7955,N_8781);
or U9237 (N_9237,N_6360,N_7954);
nand U9238 (N_9238,N_6329,N_8880);
and U9239 (N_9239,N_7422,N_7919);
nor U9240 (N_9240,N_6078,N_6188);
or U9241 (N_9241,N_6611,N_8539);
or U9242 (N_9242,N_8126,N_8377);
nand U9243 (N_9243,N_7912,N_7832);
nor U9244 (N_9244,N_7719,N_6573);
nor U9245 (N_9245,N_7396,N_6048);
and U9246 (N_9246,N_8125,N_8046);
and U9247 (N_9247,N_6787,N_8200);
and U9248 (N_9248,N_8714,N_8535);
xnor U9249 (N_9249,N_6139,N_7569);
nand U9250 (N_9250,N_6811,N_7686);
xnor U9251 (N_9251,N_8428,N_7318);
xnor U9252 (N_9252,N_7812,N_7174);
and U9253 (N_9253,N_7738,N_7303);
nand U9254 (N_9254,N_6372,N_6835);
xor U9255 (N_9255,N_6181,N_6242);
or U9256 (N_9256,N_8903,N_7351);
nand U9257 (N_9257,N_6248,N_6714);
and U9258 (N_9258,N_6110,N_8053);
or U9259 (N_9259,N_7830,N_8520);
and U9260 (N_9260,N_8633,N_6496);
nor U9261 (N_9261,N_6118,N_8147);
nand U9262 (N_9262,N_8833,N_8529);
and U9263 (N_9263,N_7821,N_7743);
nor U9264 (N_9264,N_6400,N_8988);
or U9265 (N_9265,N_7171,N_6732);
nand U9266 (N_9266,N_6957,N_6481);
nand U9267 (N_9267,N_6012,N_7073);
and U9268 (N_9268,N_8048,N_6583);
and U9269 (N_9269,N_7332,N_8187);
or U9270 (N_9270,N_6937,N_6651);
or U9271 (N_9271,N_8347,N_8096);
nand U9272 (N_9272,N_7754,N_6463);
nor U9273 (N_9273,N_6044,N_6709);
nand U9274 (N_9274,N_6031,N_7859);
and U9275 (N_9275,N_7956,N_8777);
nor U9276 (N_9276,N_8887,N_7056);
nand U9277 (N_9277,N_8944,N_6101);
or U9278 (N_9278,N_7699,N_7247);
and U9279 (N_9279,N_8653,N_7751);
or U9280 (N_9280,N_7582,N_8021);
nand U9281 (N_9281,N_8989,N_7983);
or U9282 (N_9282,N_8502,N_7982);
and U9283 (N_9283,N_6801,N_7509);
nor U9284 (N_9284,N_8079,N_7977);
nor U9285 (N_9285,N_6841,N_8255);
nand U9286 (N_9286,N_8786,N_6951);
and U9287 (N_9287,N_7094,N_6665);
nand U9288 (N_9288,N_7442,N_6428);
nor U9289 (N_9289,N_7234,N_8223);
and U9290 (N_9290,N_8197,N_8666);
nor U9291 (N_9291,N_8008,N_6193);
nor U9292 (N_9292,N_7555,N_6741);
and U9293 (N_9293,N_6207,N_6490);
or U9294 (N_9294,N_8958,N_8101);
and U9295 (N_9295,N_7500,N_6502);
or U9296 (N_9296,N_6961,N_7493);
nor U9297 (N_9297,N_6970,N_7737);
nor U9298 (N_9298,N_8285,N_7278);
nor U9299 (N_9299,N_8028,N_8108);
nand U9300 (N_9300,N_8324,N_8613);
and U9301 (N_9301,N_6860,N_8252);
nand U9302 (N_9302,N_6346,N_6705);
nor U9303 (N_9303,N_8361,N_6052);
and U9304 (N_9304,N_8045,N_6025);
or U9305 (N_9305,N_8487,N_7018);
nor U9306 (N_9306,N_7400,N_8132);
and U9307 (N_9307,N_6539,N_7196);
and U9308 (N_9308,N_8937,N_6152);
xor U9309 (N_9309,N_8983,N_7066);
nor U9310 (N_9310,N_7136,N_7946);
and U9311 (N_9311,N_6262,N_8031);
or U9312 (N_9312,N_6639,N_8175);
nor U9313 (N_9313,N_8217,N_8391);
and U9314 (N_9314,N_7824,N_6954);
or U9315 (N_9315,N_7770,N_7991);
nor U9316 (N_9316,N_6743,N_7046);
or U9317 (N_9317,N_6246,N_7588);
or U9318 (N_9318,N_7720,N_6797);
nor U9319 (N_9319,N_7537,N_6923);
and U9320 (N_9320,N_8236,N_8993);
and U9321 (N_9321,N_8456,N_7577);
or U9322 (N_9322,N_8431,N_6609);
nand U9323 (N_9323,N_7138,N_7913);
nor U9324 (N_9324,N_6320,N_7141);
nor U9325 (N_9325,N_8776,N_8144);
or U9326 (N_9326,N_8109,N_8940);
xor U9327 (N_9327,N_8403,N_6508);
nor U9328 (N_9328,N_6645,N_6672);
nand U9329 (N_9329,N_6939,N_8450);
xor U9330 (N_9330,N_7921,N_7803);
nand U9331 (N_9331,N_6223,N_8834);
nand U9332 (N_9332,N_8140,N_7460);
or U9333 (N_9333,N_7295,N_7544);
nor U9334 (N_9334,N_8041,N_8505);
or U9335 (N_9335,N_8204,N_7901);
and U9336 (N_9336,N_8066,N_6887);
nand U9337 (N_9337,N_7896,N_7219);
nor U9338 (N_9338,N_8054,N_7198);
nand U9339 (N_9339,N_8343,N_6688);
xnor U9340 (N_9340,N_7063,N_6439);
nand U9341 (N_9341,N_8004,N_8877);
or U9342 (N_9342,N_6014,N_7814);
nand U9343 (N_9343,N_7321,N_7809);
or U9344 (N_9344,N_8454,N_6933);
and U9345 (N_9345,N_7805,N_7061);
nand U9346 (N_9346,N_8328,N_6255);
nand U9347 (N_9347,N_6045,N_7191);
or U9348 (N_9348,N_7164,N_8852);
nand U9349 (N_9349,N_7273,N_6515);
and U9350 (N_9350,N_8909,N_6796);
and U9351 (N_9351,N_7275,N_8886);
and U9352 (N_9352,N_7377,N_7111);
nand U9353 (N_9353,N_6074,N_6489);
or U9354 (N_9354,N_8614,N_7801);
and U9355 (N_9355,N_6965,N_7144);
or U9356 (N_9356,N_6240,N_7225);
xor U9357 (N_9357,N_7104,N_8344);
and U9358 (N_9358,N_7251,N_8463);
xnor U9359 (N_9359,N_8349,N_6006);
nor U9360 (N_9360,N_6495,N_7314);
nor U9361 (N_9361,N_7958,N_8537);
nor U9362 (N_9362,N_7657,N_6790);
or U9363 (N_9363,N_6935,N_8521);
xnor U9364 (N_9364,N_6964,N_8568);
nand U9365 (N_9365,N_6324,N_8304);
nor U9366 (N_9366,N_8250,N_8928);
nand U9367 (N_9367,N_7966,N_8796);
and U9368 (N_9368,N_6706,N_8837);
and U9369 (N_9369,N_6237,N_8610);
nand U9370 (N_9370,N_8327,N_6930);
or U9371 (N_9371,N_6668,N_6409);
or U9372 (N_9372,N_6460,N_8679);
nand U9373 (N_9373,N_7843,N_6981);
nand U9374 (N_9374,N_6817,N_6812);
nor U9375 (N_9375,N_7489,N_6563);
and U9376 (N_9376,N_8184,N_6215);
nand U9377 (N_9377,N_6212,N_6803);
or U9378 (N_9378,N_7034,N_8476);
nor U9379 (N_9379,N_6085,N_7647);
and U9380 (N_9380,N_6745,N_7634);
or U9381 (N_9381,N_6304,N_6558);
nand U9382 (N_9382,N_6135,N_8670);
nand U9383 (N_9383,N_8815,N_6487);
and U9384 (N_9384,N_8429,N_8577);
and U9385 (N_9385,N_8488,N_8052);
or U9386 (N_9386,N_8542,N_7884);
xnor U9387 (N_9387,N_7862,N_6736);
xnor U9388 (N_9388,N_7927,N_6786);
nor U9389 (N_9389,N_8865,N_6179);
nor U9390 (N_9390,N_8661,N_7611);
and U9391 (N_9391,N_6806,N_8331);
and U9392 (N_9392,N_7706,N_6272);
or U9393 (N_9393,N_8914,N_8676);
nand U9394 (N_9394,N_8689,N_8932);
nor U9395 (N_9395,N_6361,N_7554);
and U9396 (N_9396,N_7260,N_6612);
or U9397 (N_9397,N_6302,N_6396);
xnor U9398 (N_9398,N_8557,N_6919);
nor U9399 (N_9399,N_6281,N_8658);
or U9400 (N_9400,N_7798,N_6236);
or U9401 (N_9401,N_8272,N_6424);
xor U9402 (N_9402,N_7957,N_6986);
nand U9403 (N_9403,N_7852,N_7811);
and U9404 (N_9404,N_8321,N_8318);
nand U9405 (N_9405,N_6384,N_8230);
and U9406 (N_9406,N_8648,N_8771);
and U9407 (N_9407,N_7655,N_6929);
nand U9408 (N_9408,N_7408,N_6832);
nand U9409 (N_9409,N_6571,N_8881);
or U9410 (N_9410,N_8956,N_8957);
and U9411 (N_9411,N_8270,N_6284);
nand U9412 (N_9412,N_8392,N_7666);
nor U9413 (N_9413,N_6332,N_7501);
or U9414 (N_9414,N_6585,N_8916);
nand U9415 (N_9415,N_6952,N_6667);
and U9416 (N_9416,N_7335,N_7125);
nor U9417 (N_9417,N_6059,N_7806);
nor U9418 (N_9418,N_6017,N_6784);
or U9419 (N_9419,N_6083,N_8443);
and U9420 (N_9420,N_6158,N_7692);
nand U9421 (N_9421,N_7333,N_6523);
nor U9422 (N_9422,N_8009,N_7761);
and U9423 (N_9423,N_8609,N_7494);
nand U9424 (N_9424,N_6572,N_6437);
xnor U9425 (N_9425,N_7267,N_8949);
xor U9426 (N_9426,N_6909,N_6578);
nand U9427 (N_9427,N_8995,N_7326);
xor U9428 (N_9428,N_6823,N_6358);
and U9429 (N_9429,N_8671,N_6922);
or U9430 (N_9430,N_8508,N_6605);
nand U9431 (N_9431,N_6140,N_6733);
nor U9432 (N_9432,N_7025,N_8111);
nor U9433 (N_9433,N_8083,N_7150);
and U9434 (N_9434,N_7887,N_6874);
xnor U9435 (N_9435,N_7652,N_8767);
nor U9436 (N_9436,N_7802,N_7027);
nor U9437 (N_9437,N_8919,N_8171);
and U9438 (N_9438,N_6510,N_6387);
or U9439 (N_9439,N_7014,N_6096);
or U9440 (N_9440,N_8050,N_8495);
nor U9441 (N_9441,N_7230,N_8485);
and U9442 (N_9442,N_6157,N_6819);
nor U9443 (N_9443,N_8606,N_8065);
or U9444 (N_9444,N_6288,N_6162);
nor U9445 (N_9445,N_8300,N_8231);
or U9446 (N_9446,N_8524,N_7881);
or U9447 (N_9447,N_8961,N_6826);
nor U9448 (N_9448,N_6092,N_6708);
and U9449 (N_9449,N_8575,N_8178);
nor U9450 (N_9450,N_6003,N_6698);
xor U9451 (N_9451,N_6274,N_8799);
or U9452 (N_9452,N_6710,N_7789);
or U9453 (N_9453,N_6596,N_7299);
and U9454 (N_9454,N_6920,N_8690);
and U9455 (N_9455,N_7928,N_6586);
nor U9456 (N_9456,N_8523,N_6146);
and U9457 (N_9457,N_8817,N_7356);
xnor U9458 (N_9458,N_8710,N_6985);
nand U9459 (N_9459,N_8669,N_8985);
nand U9460 (N_9460,N_7178,N_7724);
and U9461 (N_9461,N_8675,N_6378);
or U9462 (N_9462,N_7337,N_8228);
nand U9463 (N_9463,N_6451,N_7842);
or U9464 (N_9464,N_6969,N_6730);
or U9465 (N_9465,N_7502,N_6760);
and U9466 (N_9466,N_6388,N_8554);
or U9467 (N_9467,N_8134,N_6050);
and U9468 (N_9468,N_8118,N_8787);
and U9469 (N_9469,N_7213,N_6715);
nand U9470 (N_9470,N_7316,N_8744);
and U9471 (N_9471,N_8712,N_7939);
xnor U9472 (N_9472,N_7224,N_7807);
and U9473 (N_9473,N_6895,N_8694);
nor U9474 (N_9474,N_8460,N_8947);
or U9475 (N_9475,N_7117,N_8260);
and U9476 (N_9476,N_7495,N_6203);
nor U9477 (N_9477,N_7361,N_8629);
nand U9478 (N_9478,N_7548,N_8839);
and U9479 (N_9479,N_7159,N_8516);
or U9480 (N_9480,N_8726,N_6024);
xnor U9481 (N_9481,N_8122,N_6443);
nor U9482 (N_9482,N_8942,N_6511);
nand U9483 (N_9483,N_7374,N_6725);
nor U9484 (N_9484,N_7820,N_6793);
nor U9485 (N_9485,N_7031,N_8420);
or U9486 (N_9486,N_8263,N_7143);
or U9487 (N_9487,N_6778,N_6882);
and U9488 (N_9488,N_7087,N_6150);
or U9489 (N_9489,N_8256,N_8183);
and U9490 (N_9490,N_6333,N_6114);
nor U9491 (N_9491,N_6491,N_7490);
nand U9492 (N_9492,N_6076,N_8642);
nand U9493 (N_9493,N_8051,N_6010);
nor U9494 (N_9494,N_8202,N_8756);
and U9495 (N_9495,N_8018,N_6917);
or U9496 (N_9496,N_8729,N_6444);
nor U9497 (N_9497,N_7257,N_8545);
nand U9498 (N_9498,N_8974,N_8596);
and U9499 (N_9499,N_8405,N_6459);
nand U9500 (N_9500,N_8830,N_6382);
and U9501 (N_9501,N_7604,N_7709);
nor U9502 (N_9502,N_7907,N_8645);
xnor U9503 (N_9503,N_8829,N_8421);
xnor U9504 (N_9504,N_8737,N_8735);
or U9505 (N_9505,N_6173,N_6300);
or U9506 (N_9506,N_7976,N_8385);
and U9507 (N_9507,N_7701,N_6331);
and U9508 (N_9508,N_7521,N_6979);
and U9509 (N_9509,N_7863,N_6054);
and U9510 (N_9510,N_6607,N_7683);
or U9511 (N_9511,N_8586,N_6175);
and U9512 (N_9512,N_7608,N_7128);
and U9513 (N_9513,N_8507,N_7432);
xnor U9514 (N_9514,N_7679,N_7161);
or U9515 (N_9515,N_6676,N_8888);
nor U9516 (N_9516,N_6311,N_6690);
or U9517 (N_9517,N_8308,N_6419);
nand U9518 (N_9518,N_8020,N_6127);
or U9519 (N_9519,N_8222,N_7200);
or U9520 (N_9520,N_8567,N_7008);
and U9521 (N_9521,N_8470,N_7916);
or U9522 (N_9522,N_8706,N_7404);
or U9523 (N_9523,N_7465,N_8481);
nand U9524 (N_9524,N_6728,N_7478);
and U9525 (N_9525,N_7172,N_8623);
nand U9526 (N_9526,N_6512,N_8742);
and U9527 (N_9527,N_8266,N_7387);
or U9528 (N_9528,N_6533,N_6220);
nor U9529 (N_9529,N_7458,N_8743);
nand U9530 (N_9530,N_8840,N_7734);
nand U9531 (N_9531,N_6627,N_6640);
and U9532 (N_9532,N_7384,N_8578);
or U9533 (N_9533,N_7153,N_7900);
and U9534 (N_9534,N_8559,N_7097);
nor U9535 (N_9535,N_6893,N_7633);
nor U9536 (N_9536,N_8063,N_8962);
and U9537 (N_9537,N_6682,N_7480);
nand U9538 (N_9538,N_8209,N_8602);
and U9539 (N_9539,N_7309,N_7902);
nand U9540 (N_9540,N_7160,N_7974);
or U9541 (N_9541,N_7345,N_6620);
and U9542 (N_9542,N_6132,N_8773);
or U9543 (N_9543,N_7839,N_7184);
and U9544 (N_9544,N_6145,N_7284);
nand U9545 (N_9545,N_6684,N_6638);
or U9546 (N_9546,N_7336,N_6848);
and U9547 (N_9547,N_7506,N_6751);
nand U9548 (N_9548,N_6047,N_6046);
and U9549 (N_9549,N_6066,N_7274);
nand U9550 (N_9550,N_7879,N_6818);
or U9551 (N_9551,N_7531,N_8362);
nor U9552 (N_9552,N_8934,N_7517);
and U9553 (N_9553,N_6295,N_6846);
nand U9554 (N_9554,N_8594,N_7108);
xor U9555 (N_9555,N_8720,N_7662);
nand U9556 (N_9556,N_8186,N_6404);
or U9557 (N_9557,N_7948,N_7854);
or U9558 (N_9558,N_6610,N_8338);
xor U9559 (N_9559,N_8271,N_7768);
and U9560 (N_9560,N_8968,N_8576);
nand U9561 (N_9561,N_7990,N_8275);
xor U9562 (N_9562,N_7152,N_8001);
and U9563 (N_9563,N_6628,N_6662);
and U9564 (N_9564,N_8862,N_6244);
and U9565 (N_9565,N_8299,N_8847);
xnor U9566 (N_9566,N_7438,N_6643);
nor U9567 (N_9567,N_6527,N_6911);
or U9568 (N_9568,N_7660,N_6004);
nor U9569 (N_9569,N_8802,N_6077);
nor U9570 (N_9570,N_6829,N_6142);
and U9571 (N_9571,N_7216,N_7691);
xor U9572 (N_9572,N_8225,N_7834);
or U9573 (N_9573,N_8097,N_8754);
nor U9574 (N_9574,N_7518,N_7047);
nor U9575 (N_9575,N_7603,N_8156);
and U9576 (N_9576,N_7625,N_8525);
nand U9577 (N_9577,N_6019,N_8556);
nor U9578 (N_9578,N_6317,N_8784);
and U9579 (N_9579,N_8764,N_6183);
nor U9580 (N_9580,N_7283,N_7147);
or U9581 (N_9581,N_8953,N_6340);
nand U9582 (N_9582,N_8783,N_7717);
nand U9583 (N_9583,N_8905,N_8316);
xnor U9584 (N_9584,N_7922,N_7204);
and U9585 (N_9585,N_6813,N_8240);
or U9586 (N_9586,N_8859,N_6622);
or U9587 (N_9587,N_6209,N_8169);
nor U9588 (N_9588,N_6761,N_7020);
nor U9589 (N_9589,N_6654,N_6683);
or U9590 (N_9590,N_6239,N_8986);
or U9591 (N_9591,N_6503,N_6757);
nor U9592 (N_9592,N_7741,N_7044);
or U9593 (N_9593,N_6041,N_6312);
or U9594 (N_9594,N_7037,N_6983);
or U9595 (N_9595,N_8624,N_8697);
nor U9596 (N_9596,N_6397,N_6398);
xor U9597 (N_9597,N_7600,N_8005);
nand U9598 (N_9598,N_8047,N_7700);
nor U9599 (N_9599,N_7908,N_7357);
or U9600 (N_9600,N_7987,N_7787);
nand U9601 (N_9601,N_8298,N_8212);
nor U9602 (N_9602,N_6206,N_7223);
xor U9603 (N_9603,N_6065,N_7522);
or U9604 (N_9604,N_8457,N_7082);
and U9605 (N_9605,N_8411,N_8310);
nor U9606 (N_9606,N_7228,N_7290);
or U9607 (N_9607,N_7006,N_7732);
and U9608 (N_9608,N_8011,N_8528);
and U9609 (N_9609,N_6808,N_6088);
and U9610 (N_9610,N_6136,N_6866);
xnor U9611 (N_9611,N_7338,N_8026);
and U9612 (N_9612,N_8854,N_7856);
or U9613 (N_9613,N_6501,N_7425);
or U9614 (N_9614,N_7113,N_6507);
nor U9615 (N_9615,N_7950,N_8439);
and U9616 (N_9616,N_7177,N_8288);
nand U9617 (N_9617,N_7233,N_8168);
nand U9618 (N_9618,N_7355,N_7288);
nand U9619 (N_9619,N_7857,N_7621);
nor U9620 (N_9620,N_7767,N_7865);
or U9621 (N_9621,N_7484,N_6270);
nand U9622 (N_9622,N_7845,N_7665);
nor U9623 (N_9623,N_8492,N_8084);
and U9624 (N_9624,N_8352,N_8900);
and U9625 (N_9625,N_7431,N_8698);
nor U9626 (N_9626,N_7586,N_7329);
and U9627 (N_9627,N_6504,N_6494);
xor U9628 (N_9628,N_8444,N_7485);
nor U9629 (N_9629,N_6323,N_6121);
and U9630 (N_9630,N_7112,N_6905);
and U9631 (N_9631,N_7584,N_7838);
nor U9632 (N_9632,N_6861,N_6881);
xnor U9633 (N_9633,N_8550,N_6855);
nor U9634 (N_9634,N_6367,N_7581);
nor U9635 (N_9635,N_6222,N_8043);
nand U9636 (N_9636,N_8412,N_8155);
nand U9637 (N_9637,N_6291,N_6178);
nand U9638 (N_9638,N_7090,N_7639);
nor U9639 (N_9639,N_7549,N_7360);
nor U9640 (N_9640,N_6308,N_6679);
or U9641 (N_9641,N_6364,N_6549);
or U9642 (N_9642,N_7936,N_6184);
and U9643 (N_9643,N_8547,N_7443);
nand U9644 (N_9644,N_7197,N_6174);
and U9645 (N_9645,N_7003,N_8378);
xor U9646 (N_9646,N_7906,N_7334);
nand U9647 (N_9647,N_7121,N_8034);
and U9648 (N_9648,N_7017,N_8496);
and U9649 (N_9649,N_7226,N_8207);
or U9650 (N_9650,N_8752,N_6098);
and U9651 (N_9651,N_7861,N_7362);
or U9652 (N_9652,N_8356,N_8294);
or U9653 (N_9653,N_8089,N_7434);
or U9654 (N_9654,N_6402,N_8863);
nand U9655 (N_9655,N_7825,N_6673);
or U9656 (N_9656,N_8683,N_6644);
or U9657 (N_9657,N_8499,N_8721);
xor U9658 (N_9658,N_8709,N_7263);
and U9659 (N_9659,N_8466,N_7716);
or U9660 (N_9660,N_6349,N_7618);
nand U9661 (N_9661,N_6550,N_6250);
and U9662 (N_9662,N_6590,N_7256);
nor U9663 (N_9663,N_6313,N_7486);
nand U9664 (N_9664,N_6342,N_7613);
or U9665 (N_9665,N_6072,N_8668);
xnor U9666 (N_9666,N_7320,N_7886);
or U9667 (N_9667,N_8649,N_6774);
nor U9668 (N_9668,N_7898,N_8827);
nand U9669 (N_9669,N_7512,N_6754);
or U9670 (N_9670,N_7455,N_7769);
or U9671 (N_9671,N_8994,N_8433);
nand U9672 (N_9672,N_6959,N_7038);
nand U9673 (N_9673,N_7835,N_7131);
xnor U9674 (N_9674,N_8205,N_6445);
nand U9675 (N_9675,N_7429,N_8406);
and U9676 (N_9676,N_6574,N_8722);
xnor U9677 (N_9677,N_6155,N_7592);
xnor U9678 (N_9678,N_6671,N_6769);
nor U9679 (N_9679,N_7698,N_6726);
and U9680 (N_9680,N_7790,N_6254);
xor U9681 (N_9681,N_8651,N_8923);
or U9682 (N_9682,N_6901,N_6299);
nor U9683 (N_9683,N_8129,N_6219);
nor U9684 (N_9684,N_6735,N_6247);
nor U9685 (N_9685,N_7693,N_7560);
nor U9686 (N_9686,N_8110,N_7671);
nand U9687 (N_9687,N_6399,N_7327);
and U9688 (N_9688,N_6661,N_8372);
xor U9689 (N_9689,N_6411,N_6147);
and U9690 (N_9690,N_7289,N_7866);
xnor U9691 (N_9691,N_8959,N_7109);
or U9692 (N_9692,N_7142,N_7202);
or U9693 (N_9693,N_7715,N_8518);
and U9694 (N_9694,N_8080,N_7165);
or U9695 (N_9695,N_6781,N_6766);
nand U9696 (N_9696,N_7123,N_7218);
and U9697 (N_9697,N_8592,N_7100);
nor U9698 (N_9698,N_7092,N_6927);
or U9699 (N_9699,N_8303,N_6666);
nor U9700 (N_9700,N_7969,N_6553);
nand U9701 (N_9701,N_7785,N_8617);
nand U9702 (N_9702,N_8173,N_7786);
xor U9703 (N_9703,N_6341,N_7690);
xor U9704 (N_9704,N_6753,N_8278);
or U9705 (N_9705,N_8908,N_8873);
and U9706 (N_9706,N_8440,N_6894);
nor U9707 (N_9707,N_8691,N_6842);
or U9708 (N_9708,N_7705,N_6390);
and U9709 (N_9709,N_8346,N_6351);
or U9710 (N_9710,N_7841,N_7973);
nor U9711 (N_9711,N_8816,N_6765);
or U9712 (N_9712,N_7562,N_8999);
or U9713 (N_9713,N_8162,N_8100);
and U9714 (N_9714,N_7563,N_8652);
nand U9715 (N_9715,N_8534,N_6636);
or U9716 (N_9716,N_8295,N_8640);
or U9717 (N_9717,N_6691,N_6466);
or U9718 (N_9718,N_8560,N_8239);
xor U9719 (N_9719,N_8503,N_7022);
nor U9720 (N_9720,N_8196,N_6151);
nand U9721 (N_9721,N_7060,N_7423);
nand U9722 (N_9722,N_7784,N_7933);
and U9723 (N_9723,N_6423,N_6839);
xor U9724 (N_9724,N_8635,N_7587);
and U9725 (N_9725,N_8336,N_8544);
nand U9726 (N_9726,N_8449,N_8572);
or U9727 (N_9727,N_6021,N_7298);
or U9728 (N_9728,N_8663,N_7026);
and U9729 (N_9729,N_6161,N_7446);
nor U9730 (N_9730,N_8077,N_7757);
nand U9731 (N_9731,N_7681,N_8639);
nand U9732 (N_9732,N_8831,N_7406);
nand U9733 (N_9733,N_7669,N_6431);
and U9734 (N_9734,N_7893,N_8013);
or U9735 (N_9735,N_8647,N_7996);
or U9736 (N_9736,N_8511,N_6256);
nand U9737 (N_9737,N_8790,N_6000);
nand U9738 (N_9738,N_6278,N_6822);
and U9739 (N_9739,N_8732,N_8119);
nand U9740 (N_9740,N_8630,N_6176);
nand U9741 (N_9741,N_7897,N_6530);
nor U9742 (N_9742,N_8404,N_6902);
nor U9743 (N_9743,N_7179,N_6309);
nor U9744 (N_9744,N_7827,N_8104);
or U9745 (N_9745,N_6621,N_7167);
nand U9746 (N_9746,N_6433,N_8818);
nor U9747 (N_9747,N_8589,N_6857);
or U9748 (N_9748,N_7978,N_7468);
or U9749 (N_9749,N_7773,N_7011);
nand U9750 (N_9750,N_7058,N_6655);
nand U9751 (N_9751,N_7910,N_6921);
nand U9752 (N_9752,N_6115,N_8291);
nand U9753 (N_9753,N_7747,N_6505);
or U9754 (N_9754,N_6945,N_6117);
nor U9755 (N_9755,N_8279,N_7594);
nand U9756 (N_9756,N_7262,N_8469);
nand U9757 (N_9757,N_6613,N_7778);
and U9758 (N_9758,N_7407,N_6984);
nand U9759 (N_9759,N_6196,N_7215);
or U9760 (N_9760,N_8027,N_8131);
and U9761 (N_9761,N_6377,N_8176);
nand U9762 (N_9762,N_6575,N_7649);
or U9763 (N_9763,N_8845,N_6267);
or U9764 (N_9764,N_6436,N_7473);
or U9765 (N_9765,N_8190,N_8292);
nand U9766 (N_9766,N_8044,N_6593);
or U9767 (N_9767,N_7729,N_7255);
and U9768 (N_9768,N_6908,N_8713);
nand U9769 (N_9769,N_7540,N_7708);
or U9770 (N_9770,N_7118,N_6652);
and U9771 (N_9771,N_8770,N_7810);
and U9772 (N_9772,N_7098,N_6198);
or U9773 (N_9773,N_8317,N_8032);
nand U9774 (N_9774,N_8654,N_7242);
nor U9775 (N_9775,N_7032,N_7746);
and U9776 (N_9776,N_7186,N_7855);
nor U9777 (N_9777,N_6190,N_7391);
nor U9778 (N_9778,N_8437,N_7595);
and U9779 (N_9779,N_8363,N_6148);
and U9780 (N_9780,N_6748,N_6723);
or U9781 (N_9781,N_7190,N_8581);
and U9782 (N_9782,N_6303,N_6259);
nand U9783 (N_9783,N_7139,N_6462);
or U9784 (N_9784,N_6221,N_6542);
nand U9785 (N_9785,N_6016,N_6030);
xnor U9786 (N_9786,N_6509,N_8927);
or U9787 (N_9787,N_6128,N_6213);
or U9788 (N_9788,N_8935,N_7545);
nor U9789 (N_9789,N_6792,N_6354);
nand U9790 (N_9790,N_8128,N_6169);
nor U9791 (N_9791,N_6363,N_8284);
nor U9792 (N_9792,N_8977,N_6366);
or U9793 (N_9793,N_6854,N_7890);
or U9794 (N_9794,N_6039,N_6301);
nand U9795 (N_9795,N_8856,N_7642);
and U9796 (N_9796,N_8064,N_7598);
or U9797 (N_9797,N_7258,N_8954);
nor U9798 (N_9798,N_6287,N_7873);
nor U9799 (N_9799,N_7195,N_6738);
or U9800 (N_9800,N_7794,N_7209);
nor U9801 (N_9801,N_6485,N_6976);
nand U9802 (N_9802,N_7249,N_7456);
nand U9803 (N_9803,N_6227,N_6767);
or U9804 (N_9804,N_6104,N_7461);
or U9805 (N_9805,N_7375,N_6062);
and U9806 (N_9806,N_8902,N_8215);
nor U9807 (N_9807,N_6156,N_8307);
xnor U9808 (N_9808,N_6836,N_7492);
nor U9809 (N_9809,N_6564,N_6334);
nor U9810 (N_9810,N_7246,N_6971);
nor U9811 (N_9811,N_8615,N_6001);
nand U9812 (N_9812,N_7385,N_7080);
nor U9813 (N_9813,N_6594,N_7122);
nand U9814 (N_9814,N_7464,N_8858);
or U9815 (N_9815,N_6658,N_6931);
or U9816 (N_9816,N_7899,N_8702);
or U9817 (N_9817,N_8232,N_6231);
nor U9818 (N_9818,N_8150,N_7740);
nand U9819 (N_9819,N_8751,N_6456);
or U9820 (N_9820,N_7877,N_6253);
and U9821 (N_9821,N_7612,N_8312);
and U9822 (N_9822,N_8358,N_8072);
nor U9823 (N_9823,N_8965,N_7040);
nand U9824 (N_9824,N_6955,N_6664);
xor U9825 (N_9825,N_6532,N_8422);
and U9826 (N_9826,N_7917,N_7430);
nor U9827 (N_9827,N_8320,N_6026);
nand U9828 (N_9828,N_6815,N_7187);
and U9829 (N_9829,N_8159,N_6747);
and U9830 (N_9830,N_8563,N_7390);
xor U9831 (N_9831,N_8620,N_8489);
nand U9832 (N_9832,N_8325,N_6982);
nand U9833 (N_9833,N_8616,N_7428);
and U9834 (N_9834,N_7684,N_7016);
xnor U9835 (N_9835,N_6677,N_6941);
nand U9836 (N_9836,N_7129,N_6249);
nand U9837 (N_9837,N_7301,N_7682);
nand U9838 (N_9838,N_6940,N_7170);
nand U9839 (N_9839,N_6408,N_8793);
and U9840 (N_9840,N_6177,N_7436);
and U9841 (N_9841,N_8010,N_7676);
nand U9842 (N_9842,N_6853,N_8514);
nand U9843 (N_9843,N_6276,N_8512);
xor U9844 (N_9844,N_8099,N_8153);
or U9845 (N_9845,N_7819,N_7892);
nor U9846 (N_9846,N_8579,N_7710);
nand U9847 (N_9847,N_7589,N_8293);
or U9848 (N_9848,N_7221,N_7297);
or U9849 (N_9849,N_8368,N_6876);
or U9850 (N_9850,N_6700,N_6170);
and U9851 (N_9851,N_6619,N_8074);
nor U9852 (N_9852,N_8939,N_7903);
or U9853 (N_9853,N_8467,N_8448);
xor U9854 (N_9854,N_7565,N_6528);
nand U9855 (N_9855,N_7417,N_7619);
or U9856 (N_9856,N_8979,N_6915);
or U9857 (N_9857,N_8030,N_8253);
nand U9858 (N_9858,N_7564,N_8407);
nand U9859 (N_9859,N_6872,N_6814);
or U9860 (N_9860,N_8561,N_8917);
xor U9861 (N_9861,N_6699,N_6410);
nand U9862 (N_9862,N_6868,N_6153);
nand U9863 (N_9863,N_7622,N_7934);
nor U9864 (N_9864,N_7452,N_8904);
nand U9865 (N_9865,N_8311,N_6450);
and U9866 (N_9866,N_6777,N_7804);
or U9867 (N_9867,N_8017,N_8114);
nor U9868 (N_9868,N_7084,N_6385);
xor U9869 (N_9869,N_7599,N_8267);
xor U9870 (N_9870,N_8248,N_7093);
and U9871 (N_9871,N_7343,N_7636);
xor U9872 (N_9872,N_8120,N_6210);
nand U9873 (N_9873,N_7688,N_7967);
or U9874 (N_9874,N_8872,N_6108);
and U9875 (N_9875,N_7146,N_7972);
or U9876 (N_9876,N_6353,N_6465);
nor U9877 (N_9877,N_8867,N_7286);
nand U9878 (N_9878,N_8794,N_7372);
nand U9879 (N_9879,N_8715,N_7210);
or U9880 (N_9880,N_8910,N_8792);
xor U9881 (N_9881,N_7220,N_7024);
and U9882 (N_9882,N_6296,N_6896);
nor U9883 (N_9883,N_7076,N_7953);
or U9884 (N_9884,N_7585,N_7779);
and U9885 (N_9885,N_8569,N_6461);
nand U9886 (N_9886,N_7053,N_6713);
nor U9887 (N_9887,N_7448,N_6995);
xnor U9888 (N_9888,N_8763,N_6458);
or U9889 (N_9889,N_7007,N_8259);
xor U9890 (N_9890,N_7940,N_8553);
nand U9891 (N_9891,N_6641,N_7822);
xnor U9892 (N_9892,N_7580,N_7148);
and U9893 (N_9893,N_6993,N_8015);
nor U9894 (N_9894,N_6718,N_6595);
and U9895 (N_9895,N_6994,N_6015);
and U9896 (N_9896,N_7664,N_6245);
nor U9897 (N_9897,N_6201,N_6005);
xor U9898 (N_9898,N_7036,N_6251);
nor U9899 (N_9899,N_8800,N_6211);
or U9900 (N_9900,N_7188,N_8636);
or U9901 (N_9901,N_6435,N_6252);
nand U9902 (N_9902,N_6029,N_7415);
or U9903 (N_9903,N_7678,N_7192);
xor U9904 (N_9904,N_8952,N_7514);
or U9905 (N_9905,N_6037,N_6626);
or U9906 (N_9906,N_8861,N_8078);
nand U9907 (N_9907,N_8826,N_6898);
and U9908 (N_9908,N_7739,N_8139);
nand U9909 (N_9909,N_8479,N_8446);
or U9910 (N_9910,N_7341,N_6916);
xnor U9911 (N_9911,N_7874,N_7885);
xor U9912 (N_9912,N_8494,N_7993);
nor U9913 (N_9913,N_6186,N_8340);
or U9914 (N_9914,N_6998,N_7088);
or U9915 (N_9915,N_8984,N_7497);
or U9916 (N_9916,N_6432,N_8738);
nand U9917 (N_9917,N_7116,N_8326);
nand U9918 (N_9918,N_6057,N_6166);
or U9919 (N_9919,N_8059,N_8436);
or U9920 (N_9920,N_7816,N_7317);
nor U9921 (N_9921,N_7567,N_8211);
nor U9922 (N_9922,N_8314,N_7880);
or U9923 (N_9923,N_6631,N_8701);
nor U9924 (N_9924,N_8960,N_7472);
nor U9925 (N_9925,N_8061,N_7352);
nor U9926 (N_9926,N_6795,N_8201);
nor U9927 (N_9927,N_7145,N_6265);
nor U9928 (N_9928,N_8329,N_8414);
or U9929 (N_9929,N_7119,N_6663);
or U9930 (N_9930,N_7516,N_8491);
and U9931 (N_9931,N_8538,N_6326);
or U9932 (N_9932,N_8811,N_7105);
xor U9933 (N_9933,N_7369,N_7775);
and U9934 (N_9934,N_8376,N_7630);
nor U9935 (N_9935,N_8551,N_7532);
or U9936 (N_9936,N_8193,N_6888);
nor U9937 (N_9937,N_6406,N_8393);
and U9938 (N_9938,N_8747,N_7340);
xor U9939 (N_9939,N_7579,N_7089);
and U9940 (N_9940,N_6820,N_8251);
nor U9941 (N_9941,N_8876,N_6403);
nor U9942 (N_9942,N_6926,N_7815);
or U9943 (N_9943,N_6438,N_8493);
xnor U9944 (N_9944,N_6216,N_7388);
nand U9945 (N_9945,N_6430,N_6734);
nor U9946 (N_9946,N_7339,N_8382);
xnor U9947 (N_9947,N_6875,N_6191);
and U9948 (N_9948,N_7558,N_8650);
xnor U9949 (N_9949,N_7271,N_7882);
or U9950 (N_9950,N_6960,N_6711);
or U9951 (N_9951,N_6988,N_6694);
and U9952 (N_9952,N_8214,N_8945);
and U9953 (N_9953,N_8366,N_7096);
or U9954 (N_9954,N_7163,N_8203);
nand U9955 (N_9955,N_7062,N_6625);
nand U9956 (N_9956,N_7593,N_6791);
xor U9957 (N_9957,N_8387,N_8208);
and U9958 (N_9958,N_6008,N_7952);
nand U9959 (N_9959,N_6689,N_6721);
nand U9960 (N_9960,N_7222,N_6580);
or U9961 (N_9961,N_7364,N_8604);
nor U9962 (N_9962,N_6413,N_7610);
nor U9963 (N_9963,N_7459,N_7030);
and U9964 (N_9964,N_7285,N_6914);
nand U9965 (N_9965,N_8621,N_6126);
nor U9966 (N_9966,N_6670,N_6798);
nand U9967 (N_9967,N_8860,N_7474);
or U9968 (N_9968,N_6592,N_8667);
nand U9969 (N_9969,N_8664,N_6696);
and U9970 (N_9970,N_6851,N_8458);
nand U9971 (N_9971,N_8095,N_7559);
nand U9972 (N_9972,N_6477,N_7227);
nor U9973 (N_9973,N_6910,N_8580);
or U9974 (N_9974,N_7107,N_6165);
nand U9975 (N_9975,N_7766,N_8332);
nor U9976 (N_9976,N_8552,N_7624);
xnor U9977 (N_9977,N_7091,N_7951);
xor U9978 (N_9978,N_7245,N_6678);
xor U9979 (N_9979,N_8415,N_8601);
or U9980 (N_9980,N_6833,N_8868);
nor U9981 (N_9981,N_7860,N_8997);
nor U9982 (N_9982,N_7238,N_6687);
nor U9983 (N_9983,N_6794,N_7602);
nor U9984 (N_9984,N_7043,N_6943);
nand U9985 (N_9985,N_8081,N_8605);
nand U9986 (N_9986,N_8438,N_7760);
and U9987 (N_9987,N_7402,N_7596);
or U9988 (N_9988,N_6879,N_6417);
nand U9989 (N_9989,N_8662,N_6440);
or U9990 (N_9990,N_6729,N_7718);
and U9991 (N_9991,N_8395,N_7637);
and U9992 (N_9992,N_6918,N_6830);
or U9993 (N_9993,N_8277,N_8305);
nor U9994 (N_9994,N_7551,N_8235);
nor U9995 (N_9995,N_8117,N_7915);
and U9996 (N_9996,N_8607,N_6134);
or U9997 (N_9997,N_7162,N_8445);
and U9998 (N_9998,N_6685,N_6119);
and U9999 (N_9999,N_8245,N_8716);
xnor U10000 (N_10000,N_6130,N_7891);
xnor U10001 (N_10001,N_6060,N_8500);
nand U10002 (N_10002,N_6560,N_6344);
nand U10003 (N_10003,N_7771,N_7848);
nand U10004 (N_10004,N_7001,N_7645);
nor U10005 (N_10005,N_6185,N_7654);
nand U10006 (N_10006,N_8972,N_7694);
nor U10007 (N_10007,N_6991,N_8717);
nand U10008 (N_10008,N_6932,N_8590);
nand U10009 (N_10009,N_7048,N_7376);
nand U10010 (N_10010,N_7173,N_7851);
and U10011 (N_10011,N_6948,N_8788);
xnor U10012 (N_10012,N_7680,N_7039);
and U10013 (N_10013,N_6657,N_7413);
nor U10014 (N_10014,N_7386,N_6749);
xnor U10015 (N_10015,N_8584,N_8177);
and U10016 (N_10016,N_6053,N_7570);
or U10017 (N_10017,N_8795,N_6978);
nand U10018 (N_10018,N_8821,N_8820);
and U10019 (N_10019,N_6762,N_8628);
nand U10020 (N_10020,N_7986,N_6365);
and U10021 (N_10021,N_7833,N_8127);
xor U10022 (N_10022,N_8262,N_6634);
and U10023 (N_10023,N_8762,N_8646);
xor U10024 (N_10024,N_7444,N_6069);
xor U10025 (N_10025,N_8562,N_8848);
nand U10026 (N_10026,N_7294,N_8674);
nand U10027 (N_10027,N_7313,N_6637);
and U10028 (N_10028,N_8879,N_8941);
nor U10029 (N_10029,N_7012,N_6697);
nand U10030 (N_10030,N_6035,N_6849);
or U10031 (N_10031,N_7797,N_6434);
or U10032 (N_10032,N_8273,N_6018);
and U10033 (N_10033,N_8210,N_6925);
xor U10034 (N_10034,N_7793,N_7572);
xnor U10035 (N_10035,N_7072,N_7511);
nor U10036 (N_10036,N_6282,N_8441);
or U10037 (N_10037,N_7189,N_7149);
xnor U10038 (N_10038,N_6099,N_7932);
xnor U10039 (N_10039,N_7373,N_6040);
nand U10040 (N_10040,N_6702,N_7134);
and U10041 (N_10041,N_6569,N_6319);
xor U10042 (N_10042,N_6187,N_8468);
nand U10043 (N_10043,N_6405,N_6828);
nor U10044 (N_10044,N_7847,N_8599);
nand U10045 (N_10045,N_6538,N_7925);
or U10046 (N_10046,N_7296,N_7064);
and U10047 (N_10047,N_6055,N_8483);
nand U10048 (N_10048,N_8249,N_7894);
xnor U10049 (N_10049,N_6565,N_7103);
xor U10050 (N_10050,N_6776,N_8546);
nor U10051 (N_10051,N_6391,N_8759);
xnor U10052 (N_10052,N_7183,N_8842);
xor U10053 (N_10053,N_7302,N_6339);
or U10054 (N_10054,N_6731,N_8758);
nor U10055 (N_10055,N_8161,N_7627);
and U10056 (N_10056,N_8851,N_7818);
and U10057 (N_10057,N_7470,N_6452);
xnor U10058 (N_10058,N_6269,N_8068);
and U10059 (N_10059,N_7583,N_6427);
or U10060 (N_10060,N_8322,N_7538);
nor U10061 (N_10061,N_6805,N_8219);
or U10062 (N_10062,N_8281,N_7541);
nand U10063 (N_10063,N_8964,N_6468);
nor U10064 (N_10064,N_6420,N_7477);
xor U10065 (N_10065,N_7721,N_7305);
nand U10066 (N_10066,N_7962,N_6604);
or U10067 (N_10067,N_8803,N_8419);
nor U10068 (N_10068,N_8655,N_6534);
nand U10069 (N_10069,N_8339,N_7253);
and U10070 (N_10070,N_6414,N_6782);
and U10071 (N_10071,N_7735,N_8143);
or U10072 (N_10072,N_8558,N_8137);
or U10073 (N_10073,N_8086,N_7989);
nor U10074 (N_10074,N_7515,N_8276);
and U10075 (N_10075,N_6079,N_7277);
nor U10076 (N_10076,N_7575,N_7266);
xor U10077 (N_10077,N_6873,N_6478);
and U10078 (N_10078,N_7203,N_6883);
nand U10079 (N_10079,N_8736,N_7392);
nor U10080 (N_10080,N_8330,N_7959);
nor U10081 (N_10081,N_8394,N_6722);
nor U10082 (N_10082,N_6113,N_6963);
nor U10083 (N_10083,N_8823,N_7844);
nand U10084 (N_10084,N_7762,N_6357);
xor U10085 (N_10085,N_7378,N_7695);
and U10086 (N_10086,N_7566,N_6356);
xnor U10087 (N_10087,N_8243,N_8768);
nor U10088 (N_10088,N_7250,N_8342);
xor U10089 (N_10089,N_8416,N_8430);
nor U10090 (N_10090,N_8246,N_7965);
and U10091 (N_10091,N_6924,N_7523);
or U10092 (N_10092,N_8644,N_8172);
and U10093 (N_10093,N_8367,N_8618);
and U10094 (N_10094,N_8274,N_6870);
and U10095 (N_10095,N_7487,N_6310);
or U10096 (N_10096,N_7381,N_6498);
nand U10097 (N_10097,N_6858,N_6649);
nand U10098 (N_10098,N_8810,N_8425);
nor U10099 (N_10099,N_7208,N_7282);
nor U10100 (N_10100,N_7829,N_6264);
or U10101 (N_10101,N_7553,N_6257);
nand U10102 (N_10102,N_8730,N_8838);
nor U10103 (N_10103,N_7240,N_7791);
nor U10104 (N_10104,N_8739,N_7867);
nand U10105 (N_10105,N_7441,N_6788);
nand U10106 (N_10106,N_6355,N_6975);
nor U10107 (N_10107,N_7571,N_7696);
nor U10108 (N_10108,N_8315,N_7409);
xnor U10109 (N_10109,N_7574,N_6043);
nand U10110 (N_10110,N_8049,N_8920);
nand U10111 (N_10111,N_8075,N_8597);
nor U10112 (N_10112,N_6648,N_8778);
nor U10113 (N_10113,N_6680,N_6335);
and U10114 (N_10114,N_8924,N_6442);
nand U10115 (N_10115,N_7028,N_7010);
nor U10116 (N_10116,N_8060,N_8333);
nor U10117 (N_10117,N_6824,N_7828);
or U10118 (N_10118,N_8151,N_8192);
nor U10119 (N_10119,N_8955,N_8931);
nor U10120 (N_10120,N_6889,N_8695);
nor U10121 (N_10121,N_7182,N_6544);
xor U10122 (N_10122,N_8067,N_6845);
and U10123 (N_10123,N_7042,N_7875);
nand U10124 (N_10124,N_8464,N_8992);
nor U10125 (N_10125,N_8913,N_8798);
and U10126 (N_10126,N_6376,N_8227);
nor U10127 (N_10127,N_6869,N_6013);
nand U10128 (N_10128,N_6906,N_8625);
nand U10129 (N_10129,N_7744,N_6576);
nor U10130 (N_10130,N_7591,N_7930);
and U10131 (N_10131,N_8921,N_6742);
or U10132 (N_10132,N_6234,N_8185);
xnor U10133 (N_10133,N_8130,N_8612);
and U10134 (N_10134,N_7687,N_6968);
or U10135 (N_10135,N_7772,N_6561);
and U10136 (N_10136,N_6073,N_6475);
nor U10137 (N_10137,N_6068,N_8384);
or U10138 (N_10138,N_6577,N_6816);
or U10139 (N_10139,N_7504,N_7168);
nor U10140 (N_10140,N_8943,N_6164);
xnor U10141 (N_10141,N_7397,N_8218);
or U10142 (N_10142,N_7937,N_7041);
nor U10143 (N_10143,N_8723,N_8515);
nor U10144 (N_10144,N_7269,N_7127);
or U10145 (N_10145,N_7244,N_6007);
nor U10146 (N_10146,N_7281,N_6229);
nand U10147 (N_10147,N_7979,N_6457);
or U10148 (N_10148,N_7140,N_8486);
xnor U10149 (N_10149,N_6602,N_7615);
nand U10150 (N_10150,N_7052,N_6163);
nand U10151 (N_10151,N_6194,N_6633);
or U10152 (N_10152,N_6283,N_8098);
nand U10153 (N_10153,N_6516,N_7365);
and U10154 (N_10154,N_6395,N_6615);
and U10155 (N_10155,N_7752,N_7672);
nor U10156 (N_10156,N_6202,N_8970);
and U10157 (N_10157,N_6864,N_6483);
xor U10158 (N_10158,N_6904,N_8750);
xor U10159 (N_10159,N_7310,N_8684);
and U10160 (N_10160,N_6337,N_8103);
nand U10161 (N_10161,N_6759,N_8731);
nor U10162 (N_10162,N_6070,N_7367);
nor U10163 (N_10163,N_7970,N_7552);
and U10164 (N_10164,N_8133,N_6650);
nor U10165 (N_10165,N_6036,N_8632);
and U10166 (N_10166,N_6352,N_7942);
or U10167 (N_10167,N_6632,N_7307);
xor U10168 (N_10168,N_8915,N_7780);
or U10169 (N_10169,N_7895,N_8035);
and U10170 (N_10170,N_8435,N_6482);
nand U10171 (N_10171,N_6082,N_6802);
nand U10172 (N_10172,N_7463,N_8825);
nand U10173 (N_10173,N_8746,N_8141);
xor U10174 (N_10174,N_7745,N_6545);
nor U10175 (N_10175,N_6897,N_7055);
nor U10176 (N_10176,N_8585,N_6447);
xor U10177 (N_10177,N_7883,N_6780);
nor U10178 (N_10178,N_8091,N_6383);
nor U10179 (N_10179,N_8166,N_8699);
nor U10180 (N_10180,N_8761,N_6380);
nor U10181 (N_10181,N_8895,N_8398);
nor U10182 (N_10182,N_8846,N_8409);
or U10183 (N_10183,N_6584,N_6506);
nand U10184 (N_10184,N_6514,N_6675);
xor U10185 (N_10185,N_7035,N_6109);
nand U10186 (N_10186,N_6522,N_7714);
nand U10187 (N_10187,N_8142,N_8369);
nor U10188 (N_10188,N_6635,N_6002);
nor U10189 (N_10189,N_7350,N_6862);
nand U10190 (N_10190,N_6656,N_6154);
and U10191 (N_10191,N_8188,N_8198);
nand U10192 (N_10192,N_6160,N_6086);
nand U10193 (N_10193,N_7763,N_6739);
or U10194 (N_10194,N_7508,N_8174);
nor U10195 (N_10195,N_7021,N_8990);
nor U10196 (N_10196,N_7590,N_8058);
and U10197 (N_10197,N_6277,N_6081);
or U10198 (N_10198,N_8548,N_8918);
or U10199 (N_10199,N_8216,N_7201);
or U10200 (N_10200,N_7638,N_6386);
nand U10201 (N_10201,N_7293,N_7279);
and U10202 (N_10202,N_8040,N_8019);
xor U10203 (N_10203,N_8399,N_8106);
and U10204 (N_10204,N_8980,N_6758);
nor U10205 (N_10205,N_8410,N_8893);
and U10206 (N_10206,N_6763,N_8000);
nor U10207 (N_10207,N_8396,N_6877);
and U10208 (N_10208,N_6401,N_6263);
or U10209 (N_10209,N_6285,N_6373);
nand U10210 (N_10210,N_6772,N_6608);
nand U10211 (N_10211,N_8870,N_6770);
or U10212 (N_10212,N_7265,N_7924);
nor U10213 (N_10213,N_7126,N_6102);
nand U10214 (N_10214,N_7529,N_7405);
or U10215 (N_10215,N_7009,N_7650);
and U10216 (N_10216,N_6027,N_6095);
and U10217 (N_10217,N_8462,N_6600);
and U10218 (N_10218,N_7609,N_8085);
and U10219 (N_10219,N_7945,N_8423);
or U10220 (N_10220,N_6105,N_8163);
and U10221 (N_10221,N_7629,N_8866);
nand U10222 (N_10222,N_7237,N_7349);
nand U10223 (N_10223,N_6422,N_7054);
nor U10224 (N_10224,N_8071,N_6997);
nor U10225 (N_10225,N_7999,N_8154);
nand U10226 (N_10226,N_8522,N_7379);
nor U10227 (N_10227,N_6704,N_8774);
and U10228 (N_10228,N_8686,N_6197);
xnor U10229 (N_10229,N_7264,N_7081);
or U10230 (N_10230,N_6884,N_6235);
nand U10231 (N_10231,N_8678,N_8981);
or U10232 (N_10232,N_7788,N_7110);
xor U10233 (N_10233,N_7961,N_7205);
xor U10234 (N_10234,N_8749,N_7259);
nor U10235 (N_10235,N_8745,N_7199);
xor U10236 (N_10236,N_8181,N_6454);
nand U10237 (N_10237,N_8094,N_7154);
nand U10238 (N_10238,N_7949,N_8971);
nand U10239 (N_10239,N_7440,N_6111);
and U10240 (N_10240,N_6167,N_7229);
nor U10241 (N_10241,N_8348,N_6280);
nand U10242 (N_10242,N_6555,N_8510);
or U10243 (N_10243,N_8708,N_8447);
nand U10244 (N_10244,N_8337,N_8727);
and U10245 (N_10245,N_6521,N_7528);
nor U10246 (N_10246,N_8375,N_8242);
or U10247 (N_10247,N_8370,N_7019);
xnor U10248 (N_10248,N_6322,N_7510);
and U10249 (N_10249,N_8189,N_8025);
or U10250 (N_10250,N_7849,N_7998);
and U10251 (N_10251,N_6535,N_8598);
nor U10252 (N_10252,N_6479,N_6755);
nand U10253 (N_10253,N_7158,N_7270);
nand U10254 (N_10254,N_8950,N_8938);
xor U10255 (N_10255,N_7981,N_8809);
nor U10256 (N_10256,N_6724,N_6415);
or U10257 (N_10257,N_8401,N_7325);
nand U10258 (N_10258,N_7736,N_7214);
and U10259 (N_10259,N_8006,N_7535);
nand U10260 (N_10260,N_8268,N_8353);
or U10261 (N_10261,N_6852,N_6807);
and U10262 (N_10262,N_8226,N_6141);
nand U10263 (N_10263,N_7471,N_7079);
or U10264 (N_10264,N_6394,N_6719);
xnor U10265 (N_10265,N_8105,N_6551);
and U10266 (N_10266,N_8357,N_8832);
nand U10267 (N_10267,N_6570,N_8290);
nand U10268 (N_10268,N_7120,N_8976);
or U10269 (N_10269,N_8696,N_6318);
xnor U10270 (N_10270,N_8638,N_8849);
nand U10271 (N_10271,N_7984,N_7272);
and U10272 (N_10272,N_6972,N_7520);
nand U10273 (N_10273,N_8388,N_8484);
or U10274 (N_10274,N_8850,N_8891);
or U10275 (N_10275,N_7985,N_8160);
nor U10276 (N_10276,N_6913,N_7426);
nand U10277 (N_10277,N_7909,N_7756);
or U10278 (N_10278,N_6938,N_7674);
nand U10279 (N_10279,N_6347,N_6381);
and U10280 (N_10280,N_8892,N_7169);
or U10281 (N_10281,N_6912,N_8608);
or U10282 (N_10282,N_6562,N_6588);
nand U10283 (N_10283,N_7157,N_8165);
or U10284 (N_10284,N_6775,N_6305);
nor U10285 (N_10285,N_8241,N_7395);
or U10286 (N_10286,N_8555,N_8002);
and U10287 (N_10287,N_6579,N_6232);
and U10288 (N_10288,N_6804,N_8480);
nor U10289 (N_10289,N_8532,N_8465);
or U10290 (N_10290,N_8373,N_7241);
nand U10291 (N_10291,N_7992,N_8951);
or U10292 (N_10292,N_7185,N_7427);
xor U10293 (N_10293,N_7858,N_8283);
nand U10294 (N_10294,N_8323,N_7641);
or U10295 (N_10295,N_7399,N_7067);
and U10296 (N_10296,N_8593,N_6859);
and U10297 (N_10297,N_8121,N_8022);
and U10298 (N_10298,N_6261,N_8335);
nand U10299 (N_10299,N_6292,N_8687);
xnor U10300 (N_10300,N_7616,N_8889);
nand U10301 (N_10301,N_6990,N_6224);
nand U10302 (N_10302,N_7433,N_6546);
nand U10303 (N_10303,N_6880,N_6617);
nor U10304 (N_10304,N_8213,N_6903);
and U10305 (N_10305,N_8693,N_8703);
nand U10306 (N_10306,N_6524,N_6520);
nand U10307 (N_10307,N_7070,N_6587);
nor U10308 (N_10308,N_7628,N_8898);
nor U10309 (N_10309,N_6844,N_7292);
nand U10310 (N_10310,N_7935,N_8400);
xnor U10311 (N_10311,N_6707,N_7322);
and U10312 (N_10312,N_6464,N_6090);
nand U10313 (N_10313,N_6071,N_8055);
or U10314 (N_10314,N_8673,N_8634);
nor U10315 (N_10315,N_7975,N_7878);
nand U10316 (N_10316,N_7075,N_6370);
nor U10317 (N_10317,N_6556,N_7960);
and U10318 (N_10318,N_7524,N_6469);
nor U10319 (N_10319,N_6716,N_8042);
or U10320 (N_10320,N_8631,N_7943);
nand U10321 (N_10321,N_8725,N_6999);
or U10322 (N_10322,N_6058,N_8564);
nand U10323 (N_10323,N_8531,N_7348);
and U10324 (N_10324,N_8765,N_6472);
or U10325 (N_10325,N_7315,N_8692);
nand U10326 (N_10326,N_7632,N_6034);
or U10327 (N_10327,N_8672,N_7156);
nor U10328 (N_10328,N_6557,N_7527);
or U10329 (N_10329,N_6944,N_7640);
nand U10330 (N_10330,N_6120,N_7546);
nand U10331 (N_10331,N_7755,N_7466);
xor U10332 (N_10332,N_8309,N_8282);
and U10333 (N_10333,N_8680,N_7931);
nand U10334 (N_10334,N_6756,N_7617);
or U10335 (N_10335,N_7308,N_6480);
and U10336 (N_10336,N_7106,N_8016);
and U10337 (N_10337,N_8741,N_6056);
nand U10338 (N_10338,N_8313,N_7457);
nand U10339 (N_10339,N_7872,N_6379);
nand U10340 (N_10340,N_8498,N_8540);
nand U10341 (N_10341,N_6692,N_7646);
and U10342 (N_10342,N_7723,N_7813);
and U10343 (N_10343,N_7920,N_6992);
or U10344 (N_10344,N_8146,N_8057);
or U10345 (N_10345,N_8124,N_6359);
or U10346 (N_10346,N_8364,N_6289);
nand U10347 (N_10347,N_8265,N_8280);
or U10348 (N_10348,N_8112,N_7475);
nor U10349 (N_10349,N_6063,N_8890);
and U10350 (N_10350,N_6843,N_6271);
and U10351 (N_10351,N_8874,N_7576);
nand U10352 (N_10352,N_7065,N_7836);
and U10353 (N_10353,N_7342,N_8102);
or U10354 (N_10354,N_6389,N_8527);
nor U10355 (N_10355,N_6325,N_8806);
or U10356 (N_10356,N_7748,N_6513);
xor U10357 (N_10357,N_8813,N_6094);
nand U10358 (N_10358,N_7918,N_7643);
or U10359 (N_10359,N_7051,N_6293);
xnor U10360 (N_10360,N_6942,N_6746);
nand U10361 (N_10361,N_6484,N_7069);
nor U10362 (N_10362,N_8036,N_8844);
nand U10363 (N_10363,N_6934,N_6531);
xor U10364 (N_10364,N_7536,N_7911);
nor U10365 (N_10365,N_7675,N_6425);
nor U10366 (N_10366,N_7124,N_8497);
nor U10367 (N_10367,N_8978,N_6996);
and U10368 (N_10368,N_7876,N_8929);
or U10369 (N_10369,N_8797,N_7808);
or U10370 (N_10370,N_6023,N_7439);
or U10371 (N_10371,N_7730,N_8748);
and U10372 (N_10372,N_7656,N_8700);
nand U10373 (N_10373,N_7614,N_7424);
and U10374 (N_10374,N_8757,N_7914);
and U10375 (N_10375,N_7358,N_6375);
nand U10376 (N_10376,N_6393,N_6371);
and U10377 (N_10377,N_7371,N_7702);
nand U10378 (N_10378,N_6407,N_8158);
nand U10379 (N_10379,N_7995,N_7155);
or U10380 (N_10380,N_8475,N_6548);
nand U10381 (N_10381,N_7871,N_7578);
nor U10382 (N_10382,N_7077,N_7968);
nand U10383 (N_10383,N_6907,N_8724);
nor U10384 (N_10384,N_8600,N_6525);
nor U10385 (N_10385,N_6740,N_6455);
or U10386 (N_10386,N_6989,N_6228);
or U10387 (N_10387,N_7445,N_8719);
nor U10388 (N_10388,N_8380,N_7607);
nor U10389 (N_10389,N_7573,N_6116);
or U10390 (N_10390,N_8426,N_6338);
or U10391 (N_10391,N_6268,N_7074);
nand U10392 (N_10392,N_6093,N_6441);
and U10393 (N_10393,N_8149,N_6591);
nor U10394 (N_10394,N_7759,N_7568);
nand U10395 (N_10395,N_8565,N_6947);
nand U10396 (N_10396,N_7276,N_6225);
nand U10397 (N_10397,N_6681,N_7059);
or U10398 (N_10398,N_8073,N_7133);
or U10399 (N_10399,N_8379,N_7799);
and U10400 (N_10400,N_7542,N_7623);
nor U10401 (N_10401,N_6892,N_6328);
or U10402 (N_10402,N_8549,N_6133);
nor U10403 (N_10403,N_8982,N_6629);
or U10404 (N_10404,N_8355,N_8506);
or U10405 (N_10405,N_7964,N_7507);
nor U10406 (N_10406,N_8194,N_7888);
and U10407 (N_10407,N_7938,N_8334);
or U10408 (N_10408,N_6597,N_6080);
nor U10409 (N_10409,N_6470,N_8987);
and U10410 (N_10410,N_7013,N_8037);
nand U10411 (N_10411,N_8812,N_7488);
nor U10412 (N_10412,N_6536,N_7243);
nand U10413 (N_10413,N_6192,N_8287);
nor U10414 (N_10414,N_8351,N_8501);
xnor U10415 (N_10415,N_8195,N_6936);
xnor U10416 (N_10416,N_7758,N_6712);
nor U10417 (N_10417,N_6488,N_7668);
nor U10418 (N_10418,N_8603,N_8622);
or U10419 (N_10419,N_7648,N_7328);
or U10420 (N_10420,N_7980,N_7045);
xor U10421 (N_10421,N_6552,N_7101);
or U10422 (N_10422,N_6831,N_7287);
nor U10423 (N_10423,N_6208,N_8897);
nor U10424 (N_10424,N_8519,N_6204);
or U10425 (N_10425,N_6122,N_7605);
and U10426 (N_10426,N_6529,N_7525);
and U10427 (N_10427,N_7239,N_7944);
and U10428 (N_10428,N_6064,N_7115);
and U10429 (N_10429,N_8148,N_8170);
and U10430 (N_10430,N_6956,N_8574);
and U10431 (N_10431,N_8822,N_6492);
and U10432 (N_10432,N_8261,N_7383);
and U10433 (N_10433,N_8012,N_8296);
nor U10434 (N_10434,N_6582,N_6863);
nor U10435 (N_10435,N_8707,N_8397);
nor U10436 (N_10436,N_6871,N_8769);
nand U10437 (N_10437,N_7029,N_7597);
nor U10438 (N_10438,N_7764,N_8998);
or U10439 (N_10439,N_7363,N_6779);
or U10440 (N_10440,N_8247,N_8221);
xor U10441 (N_10441,N_7193,N_6616);
and U10442 (N_10442,N_8007,N_8973);
nand U10443 (N_10443,N_7166,N_8766);
and U10444 (N_10444,N_7765,N_7207);
nor U10445 (N_10445,N_6199,N_6327);
and U10446 (N_10446,N_8087,N_7670);
nand U10447 (N_10447,N_6471,N_6890);
xor U10448 (N_10448,N_8517,N_7498);
nor U10449 (N_10449,N_7868,N_7354);
nor U10450 (N_10450,N_6374,N_8907);
nand U10451 (N_10451,N_7370,N_7049);
nor U10452 (N_10452,N_8417,N_8641);
nor U10453 (N_10453,N_6606,N_6953);
or U10454 (N_10454,N_8206,N_7697);
nor U10455 (N_10455,N_8733,N_6200);
and U10456 (N_10456,N_6977,N_6559);
nor U10457 (N_10457,N_6646,N_6669);
xor U10458 (N_10458,N_8301,N_7206);
or U10459 (N_10459,N_8088,N_7753);
nor U10460 (N_10460,N_6598,N_7728);
nand U10461 (N_10461,N_8107,N_8807);
nand U10462 (N_10462,N_7499,N_7673);
and U10463 (N_10463,N_7023,N_7796);
or U10464 (N_10464,N_7677,N_7707);
or U10465 (N_10465,N_6087,N_7491);
and U10466 (N_10466,N_6241,N_8473);
or U10467 (N_10467,N_8659,N_6878);
nand U10468 (N_10468,N_6091,N_7323);
xor U10469 (N_10469,N_8853,N_8665);
xnor U10470 (N_10470,N_6500,N_8911);
or U10471 (N_10471,N_8819,N_8789);
or U10472 (N_10472,N_6100,N_7312);
and U10473 (N_10473,N_6123,N_8871);
nor U10474 (N_10474,N_7971,N_6260);
and U10475 (N_10475,N_8459,N_6810);
nor U10476 (N_10476,N_7382,N_6840);
nor U10477 (N_10477,N_8082,N_6647);
nand U10478 (N_10478,N_6306,N_6618);
nor U10479 (N_10479,N_6042,N_8434);
or U10480 (N_10480,N_6867,N_7530);
nor U10481 (N_10481,N_6107,N_8157);
nor U10482 (N_10482,N_8566,N_8451);
or U10483 (N_10483,N_6537,N_6336);
or U10484 (N_10484,N_8755,N_8024);
or U10485 (N_10485,N_6392,N_8922);
or U10486 (N_10486,N_7831,N_7194);
nor U10487 (N_10487,N_7151,N_6273);
or U10488 (N_10488,N_8471,N_8530);
nand U10489 (N_10489,N_8474,N_6103);
or U10490 (N_10490,N_7923,N_7050);
or U10491 (N_10491,N_7235,N_8991);
and U10492 (N_10492,N_8627,N_8413);
nand U10493 (N_10493,N_6800,N_8878);
nand U10494 (N_10494,N_6243,N_6418);
nor U10495 (N_10495,N_6566,N_8116);
and U10496 (N_10496,N_7175,N_6038);
and U10497 (N_10497,N_8383,N_6900);
or U10498 (N_10498,N_8371,N_8536);
nor U10499 (N_10499,N_6416,N_7776);
and U10500 (N_10500,N_7674,N_7373);
nand U10501 (N_10501,N_6377,N_7080);
and U10502 (N_10502,N_8861,N_8161);
nor U10503 (N_10503,N_8850,N_7193);
xor U10504 (N_10504,N_7140,N_6027);
nand U10505 (N_10505,N_8661,N_7684);
or U10506 (N_10506,N_7823,N_6315);
xnor U10507 (N_10507,N_7948,N_7787);
nor U10508 (N_10508,N_7273,N_6038);
nand U10509 (N_10509,N_7222,N_6568);
nand U10510 (N_10510,N_7953,N_6776);
or U10511 (N_10511,N_7633,N_8682);
or U10512 (N_10512,N_6176,N_7783);
or U10513 (N_10513,N_7842,N_6329);
nor U10514 (N_10514,N_6568,N_6317);
nor U10515 (N_10515,N_7174,N_7363);
or U10516 (N_10516,N_7083,N_6534);
nand U10517 (N_10517,N_8601,N_6043);
nor U10518 (N_10518,N_7060,N_6689);
nand U10519 (N_10519,N_8098,N_6897);
xnor U10520 (N_10520,N_6207,N_7575);
nor U10521 (N_10521,N_6879,N_7806);
nor U10522 (N_10522,N_6419,N_6926);
and U10523 (N_10523,N_7420,N_7899);
nand U10524 (N_10524,N_7891,N_6046);
or U10525 (N_10525,N_7772,N_8936);
nand U10526 (N_10526,N_8008,N_6910);
nand U10527 (N_10527,N_6136,N_8542);
xor U10528 (N_10528,N_6218,N_7864);
xnor U10529 (N_10529,N_7171,N_6498);
nand U10530 (N_10530,N_6337,N_6282);
nor U10531 (N_10531,N_7323,N_8196);
or U10532 (N_10532,N_7167,N_6574);
xor U10533 (N_10533,N_7784,N_6391);
and U10534 (N_10534,N_8541,N_6022);
or U10535 (N_10535,N_7484,N_6548);
nand U10536 (N_10536,N_7281,N_7885);
nand U10537 (N_10537,N_6892,N_6890);
xnor U10538 (N_10538,N_6245,N_6991);
nand U10539 (N_10539,N_8567,N_8635);
nor U10540 (N_10540,N_6774,N_6586);
or U10541 (N_10541,N_6308,N_6765);
nor U10542 (N_10542,N_7908,N_6051);
or U10543 (N_10543,N_6689,N_6512);
and U10544 (N_10544,N_7808,N_7765);
nand U10545 (N_10545,N_7105,N_7793);
nor U10546 (N_10546,N_6133,N_7727);
xor U10547 (N_10547,N_7690,N_6697);
or U10548 (N_10548,N_6880,N_6295);
and U10549 (N_10549,N_7708,N_6281);
or U10550 (N_10550,N_7452,N_7625);
and U10551 (N_10551,N_8840,N_7341);
or U10552 (N_10552,N_8819,N_6924);
nor U10553 (N_10553,N_7522,N_8566);
nor U10554 (N_10554,N_8851,N_7954);
or U10555 (N_10555,N_8080,N_6888);
and U10556 (N_10556,N_8252,N_6888);
nand U10557 (N_10557,N_8313,N_6738);
and U10558 (N_10558,N_8441,N_8856);
xor U10559 (N_10559,N_6770,N_7733);
nor U10560 (N_10560,N_6451,N_8546);
or U10561 (N_10561,N_7219,N_7951);
and U10562 (N_10562,N_6466,N_6623);
or U10563 (N_10563,N_8488,N_7747);
or U10564 (N_10564,N_7163,N_8416);
and U10565 (N_10565,N_6415,N_8295);
and U10566 (N_10566,N_6253,N_6615);
and U10567 (N_10567,N_8056,N_8033);
nand U10568 (N_10568,N_6259,N_6304);
and U10569 (N_10569,N_8332,N_6719);
or U10570 (N_10570,N_8102,N_6260);
nor U10571 (N_10571,N_6755,N_8360);
or U10572 (N_10572,N_8360,N_7579);
or U10573 (N_10573,N_7286,N_8960);
and U10574 (N_10574,N_8718,N_8692);
nand U10575 (N_10575,N_8291,N_8696);
nor U10576 (N_10576,N_8577,N_8478);
and U10577 (N_10577,N_7827,N_8392);
or U10578 (N_10578,N_6300,N_8065);
nand U10579 (N_10579,N_6078,N_7911);
and U10580 (N_10580,N_7522,N_8965);
nand U10581 (N_10581,N_7734,N_7195);
or U10582 (N_10582,N_6405,N_6705);
and U10583 (N_10583,N_8968,N_6033);
nor U10584 (N_10584,N_6925,N_6131);
nand U10585 (N_10585,N_8921,N_8923);
nor U10586 (N_10586,N_8513,N_6584);
and U10587 (N_10587,N_8234,N_6447);
nor U10588 (N_10588,N_8046,N_8423);
xor U10589 (N_10589,N_7597,N_8542);
nand U10590 (N_10590,N_7537,N_8285);
and U10591 (N_10591,N_7374,N_6662);
nand U10592 (N_10592,N_8782,N_7683);
or U10593 (N_10593,N_8023,N_8463);
xor U10594 (N_10594,N_7000,N_8634);
nand U10595 (N_10595,N_6039,N_7174);
or U10596 (N_10596,N_6762,N_7875);
or U10597 (N_10597,N_7549,N_6991);
nor U10598 (N_10598,N_8820,N_8682);
nand U10599 (N_10599,N_7675,N_6788);
nand U10600 (N_10600,N_8843,N_8672);
nor U10601 (N_10601,N_8126,N_7415);
nand U10602 (N_10602,N_8316,N_7971);
nand U10603 (N_10603,N_7840,N_7796);
and U10604 (N_10604,N_7247,N_6244);
nor U10605 (N_10605,N_6811,N_6689);
or U10606 (N_10606,N_8920,N_8820);
nor U10607 (N_10607,N_6674,N_8379);
and U10608 (N_10608,N_6350,N_6080);
or U10609 (N_10609,N_8069,N_7925);
and U10610 (N_10610,N_7824,N_8140);
or U10611 (N_10611,N_8346,N_6359);
or U10612 (N_10612,N_6895,N_8492);
nor U10613 (N_10613,N_6569,N_6895);
and U10614 (N_10614,N_8204,N_8475);
nor U10615 (N_10615,N_7646,N_6211);
nor U10616 (N_10616,N_7786,N_8224);
or U10617 (N_10617,N_6791,N_8045);
nand U10618 (N_10618,N_6931,N_6305);
or U10619 (N_10619,N_6112,N_7531);
or U10620 (N_10620,N_8819,N_7286);
nand U10621 (N_10621,N_7107,N_8401);
xnor U10622 (N_10622,N_7021,N_7848);
and U10623 (N_10623,N_6438,N_7306);
or U10624 (N_10624,N_6291,N_8300);
xor U10625 (N_10625,N_7351,N_8965);
and U10626 (N_10626,N_7561,N_7170);
nand U10627 (N_10627,N_6647,N_8733);
nor U10628 (N_10628,N_8081,N_7335);
nand U10629 (N_10629,N_7234,N_8534);
nand U10630 (N_10630,N_7039,N_8253);
or U10631 (N_10631,N_8929,N_6780);
nor U10632 (N_10632,N_7461,N_6470);
nor U10633 (N_10633,N_7131,N_6742);
and U10634 (N_10634,N_6963,N_7516);
nand U10635 (N_10635,N_8103,N_6321);
nor U10636 (N_10636,N_7036,N_8403);
nor U10637 (N_10637,N_6218,N_8768);
nand U10638 (N_10638,N_6396,N_7584);
nand U10639 (N_10639,N_7022,N_8708);
nor U10640 (N_10640,N_7672,N_6200);
or U10641 (N_10641,N_6125,N_6076);
nand U10642 (N_10642,N_7745,N_7830);
nand U10643 (N_10643,N_8099,N_7157);
or U10644 (N_10644,N_8025,N_6581);
nor U10645 (N_10645,N_8810,N_7882);
and U10646 (N_10646,N_8081,N_7937);
nor U10647 (N_10647,N_7306,N_8440);
nand U10648 (N_10648,N_8357,N_8206);
nand U10649 (N_10649,N_6489,N_7353);
nor U10650 (N_10650,N_6421,N_6219);
nor U10651 (N_10651,N_6812,N_8233);
nor U10652 (N_10652,N_8350,N_6852);
or U10653 (N_10653,N_6463,N_8566);
nor U10654 (N_10654,N_6430,N_8793);
or U10655 (N_10655,N_7635,N_8810);
nand U10656 (N_10656,N_8958,N_8884);
nor U10657 (N_10657,N_8762,N_8233);
and U10658 (N_10658,N_8254,N_7032);
or U10659 (N_10659,N_8146,N_7191);
nand U10660 (N_10660,N_8830,N_6099);
nand U10661 (N_10661,N_7418,N_8484);
nor U10662 (N_10662,N_7212,N_8844);
and U10663 (N_10663,N_6693,N_8268);
nor U10664 (N_10664,N_8630,N_6770);
and U10665 (N_10665,N_8960,N_8243);
and U10666 (N_10666,N_8141,N_8689);
or U10667 (N_10667,N_7023,N_7269);
nand U10668 (N_10668,N_7609,N_6158);
and U10669 (N_10669,N_7741,N_8158);
or U10670 (N_10670,N_6753,N_6980);
nand U10671 (N_10671,N_6185,N_7749);
or U10672 (N_10672,N_7066,N_7368);
nand U10673 (N_10673,N_8838,N_6073);
or U10674 (N_10674,N_8868,N_6527);
or U10675 (N_10675,N_6448,N_8902);
nor U10676 (N_10676,N_8196,N_6819);
nor U10677 (N_10677,N_6773,N_7241);
xnor U10678 (N_10678,N_8799,N_7293);
nor U10679 (N_10679,N_7411,N_8521);
nand U10680 (N_10680,N_8750,N_6293);
and U10681 (N_10681,N_6800,N_6467);
or U10682 (N_10682,N_6064,N_8464);
and U10683 (N_10683,N_7007,N_6242);
and U10684 (N_10684,N_6188,N_8574);
xnor U10685 (N_10685,N_8983,N_8742);
and U10686 (N_10686,N_7052,N_7665);
or U10687 (N_10687,N_6557,N_7752);
nor U10688 (N_10688,N_6732,N_8224);
xnor U10689 (N_10689,N_8203,N_6367);
and U10690 (N_10690,N_7543,N_8387);
or U10691 (N_10691,N_7998,N_6815);
nand U10692 (N_10692,N_7541,N_6470);
nor U10693 (N_10693,N_7308,N_6390);
or U10694 (N_10694,N_6714,N_6026);
xor U10695 (N_10695,N_7007,N_7650);
nor U10696 (N_10696,N_6368,N_7500);
nand U10697 (N_10697,N_8309,N_7762);
nand U10698 (N_10698,N_8397,N_7274);
xnor U10699 (N_10699,N_7782,N_7123);
and U10700 (N_10700,N_8654,N_8807);
nor U10701 (N_10701,N_7054,N_7690);
xnor U10702 (N_10702,N_7325,N_7355);
nand U10703 (N_10703,N_7456,N_6766);
nand U10704 (N_10704,N_6386,N_7232);
and U10705 (N_10705,N_8310,N_7066);
and U10706 (N_10706,N_7627,N_7750);
and U10707 (N_10707,N_6970,N_7150);
nor U10708 (N_10708,N_7122,N_8365);
or U10709 (N_10709,N_8233,N_6003);
or U10710 (N_10710,N_7258,N_6893);
nand U10711 (N_10711,N_8098,N_6016);
and U10712 (N_10712,N_7071,N_8899);
nor U10713 (N_10713,N_6495,N_6007);
nor U10714 (N_10714,N_6087,N_7410);
and U10715 (N_10715,N_6186,N_7843);
nor U10716 (N_10716,N_8140,N_8604);
and U10717 (N_10717,N_6713,N_8658);
and U10718 (N_10718,N_7135,N_8738);
nor U10719 (N_10719,N_8204,N_8666);
nor U10720 (N_10720,N_8718,N_7277);
xnor U10721 (N_10721,N_8864,N_8359);
or U10722 (N_10722,N_7942,N_8368);
nor U10723 (N_10723,N_8717,N_8412);
nand U10724 (N_10724,N_6669,N_8651);
xor U10725 (N_10725,N_6534,N_7226);
xor U10726 (N_10726,N_6087,N_6760);
or U10727 (N_10727,N_6133,N_6156);
xor U10728 (N_10728,N_6629,N_8303);
nor U10729 (N_10729,N_6698,N_8797);
nand U10730 (N_10730,N_7341,N_6074);
nor U10731 (N_10731,N_8518,N_8798);
and U10732 (N_10732,N_7289,N_7087);
or U10733 (N_10733,N_6278,N_7158);
nand U10734 (N_10734,N_7185,N_6625);
or U10735 (N_10735,N_7133,N_7704);
nor U10736 (N_10736,N_7243,N_8754);
or U10737 (N_10737,N_7492,N_8781);
and U10738 (N_10738,N_8925,N_7914);
nor U10739 (N_10739,N_7010,N_8628);
nor U10740 (N_10740,N_6210,N_6574);
or U10741 (N_10741,N_8076,N_6858);
nand U10742 (N_10742,N_7466,N_7346);
nor U10743 (N_10743,N_6839,N_8638);
nand U10744 (N_10744,N_6300,N_7609);
and U10745 (N_10745,N_8142,N_8278);
nor U10746 (N_10746,N_6783,N_6325);
or U10747 (N_10747,N_6435,N_6112);
or U10748 (N_10748,N_8339,N_6577);
or U10749 (N_10749,N_6891,N_7279);
xor U10750 (N_10750,N_7497,N_7064);
and U10751 (N_10751,N_6415,N_6777);
nor U10752 (N_10752,N_7347,N_7452);
nand U10753 (N_10753,N_8695,N_6188);
nor U10754 (N_10754,N_7847,N_6741);
nor U10755 (N_10755,N_6604,N_8977);
nand U10756 (N_10756,N_6660,N_8611);
xnor U10757 (N_10757,N_8738,N_8519);
or U10758 (N_10758,N_8644,N_6484);
nand U10759 (N_10759,N_7886,N_8957);
and U10760 (N_10760,N_8255,N_6731);
nor U10761 (N_10761,N_6070,N_6267);
and U10762 (N_10762,N_8086,N_6354);
or U10763 (N_10763,N_6624,N_7385);
and U10764 (N_10764,N_6089,N_6211);
nand U10765 (N_10765,N_7892,N_7682);
or U10766 (N_10766,N_8491,N_7344);
or U10767 (N_10767,N_7179,N_7977);
xor U10768 (N_10768,N_8936,N_8308);
nor U10769 (N_10769,N_8691,N_6498);
or U10770 (N_10770,N_8448,N_6564);
xor U10771 (N_10771,N_8996,N_8670);
or U10772 (N_10772,N_7150,N_6391);
nor U10773 (N_10773,N_6991,N_8265);
and U10774 (N_10774,N_6679,N_7836);
or U10775 (N_10775,N_7702,N_8992);
nand U10776 (N_10776,N_6420,N_8160);
xor U10777 (N_10777,N_6083,N_6711);
and U10778 (N_10778,N_7756,N_6420);
nor U10779 (N_10779,N_6635,N_6492);
nor U10780 (N_10780,N_7810,N_7258);
or U10781 (N_10781,N_7297,N_8729);
and U10782 (N_10782,N_7617,N_8763);
nand U10783 (N_10783,N_7617,N_6828);
or U10784 (N_10784,N_6352,N_7139);
and U10785 (N_10785,N_7647,N_7183);
or U10786 (N_10786,N_6007,N_8091);
or U10787 (N_10787,N_6567,N_7999);
and U10788 (N_10788,N_6715,N_8282);
and U10789 (N_10789,N_6942,N_8795);
nor U10790 (N_10790,N_6301,N_7802);
or U10791 (N_10791,N_8786,N_6074);
or U10792 (N_10792,N_8013,N_8235);
nor U10793 (N_10793,N_6062,N_7731);
nand U10794 (N_10794,N_8252,N_8012);
nand U10795 (N_10795,N_8232,N_8389);
nand U10796 (N_10796,N_7703,N_6933);
nand U10797 (N_10797,N_6939,N_7933);
nand U10798 (N_10798,N_6829,N_6412);
and U10799 (N_10799,N_8192,N_6569);
nor U10800 (N_10800,N_8347,N_7770);
xnor U10801 (N_10801,N_7269,N_8131);
and U10802 (N_10802,N_8657,N_8156);
and U10803 (N_10803,N_6040,N_7857);
or U10804 (N_10804,N_8153,N_7743);
nor U10805 (N_10805,N_7343,N_6497);
and U10806 (N_10806,N_7529,N_6869);
nor U10807 (N_10807,N_7489,N_8151);
nor U10808 (N_10808,N_6312,N_8530);
nand U10809 (N_10809,N_7946,N_6218);
nand U10810 (N_10810,N_8216,N_8555);
and U10811 (N_10811,N_8681,N_7486);
nand U10812 (N_10812,N_6370,N_7158);
and U10813 (N_10813,N_6364,N_6836);
and U10814 (N_10814,N_6194,N_7012);
or U10815 (N_10815,N_7407,N_8223);
nor U10816 (N_10816,N_6136,N_7941);
nand U10817 (N_10817,N_8538,N_6535);
and U10818 (N_10818,N_8600,N_6318);
nand U10819 (N_10819,N_7108,N_6335);
xnor U10820 (N_10820,N_7082,N_8910);
nor U10821 (N_10821,N_6596,N_7646);
or U10822 (N_10822,N_8559,N_8086);
xor U10823 (N_10823,N_8733,N_7380);
nor U10824 (N_10824,N_8995,N_7598);
and U10825 (N_10825,N_7366,N_7210);
and U10826 (N_10826,N_8473,N_6124);
and U10827 (N_10827,N_8467,N_7470);
and U10828 (N_10828,N_7421,N_7164);
and U10829 (N_10829,N_7463,N_8399);
and U10830 (N_10830,N_8210,N_7286);
and U10831 (N_10831,N_7113,N_7340);
nand U10832 (N_10832,N_8762,N_8109);
nor U10833 (N_10833,N_8113,N_6469);
or U10834 (N_10834,N_7683,N_6933);
and U10835 (N_10835,N_8331,N_7980);
or U10836 (N_10836,N_8356,N_7098);
or U10837 (N_10837,N_7788,N_7450);
or U10838 (N_10838,N_8910,N_8731);
and U10839 (N_10839,N_7616,N_8356);
nor U10840 (N_10840,N_8873,N_8956);
or U10841 (N_10841,N_7472,N_6742);
or U10842 (N_10842,N_7670,N_6503);
or U10843 (N_10843,N_6451,N_8629);
or U10844 (N_10844,N_6454,N_6924);
or U10845 (N_10845,N_7670,N_7300);
or U10846 (N_10846,N_8624,N_6985);
xor U10847 (N_10847,N_7490,N_7055);
nor U10848 (N_10848,N_8473,N_6697);
or U10849 (N_10849,N_6876,N_8856);
or U10850 (N_10850,N_7711,N_7526);
and U10851 (N_10851,N_6384,N_6459);
or U10852 (N_10852,N_8063,N_6567);
or U10853 (N_10853,N_8084,N_6372);
or U10854 (N_10854,N_8628,N_6699);
nor U10855 (N_10855,N_8295,N_7465);
and U10856 (N_10856,N_6856,N_6173);
nor U10857 (N_10857,N_6466,N_7881);
or U10858 (N_10858,N_7783,N_8837);
or U10859 (N_10859,N_6990,N_7577);
nor U10860 (N_10860,N_6113,N_8211);
and U10861 (N_10861,N_6858,N_7397);
or U10862 (N_10862,N_7975,N_7176);
nor U10863 (N_10863,N_6728,N_6002);
nor U10864 (N_10864,N_7364,N_8497);
nand U10865 (N_10865,N_6129,N_8842);
and U10866 (N_10866,N_8988,N_7638);
nor U10867 (N_10867,N_8219,N_7385);
xnor U10868 (N_10868,N_7390,N_7710);
nor U10869 (N_10869,N_7008,N_6709);
xor U10870 (N_10870,N_8067,N_8521);
nor U10871 (N_10871,N_8656,N_7864);
nor U10872 (N_10872,N_6819,N_7065);
nor U10873 (N_10873,N_7588,N_8162);
nor U10874 (N_10874,N_7688,N_7781);
or U10875 (N_10875,N_8379,N_6428);
nor U10876 (N_10876,N_6654,N_7343);
nor U10877 (N_10877,N_6706,N_7621);
nand U10878 (N_10878,N_6781,N_8415);
and U10879 (N_10879,N_7751,N_8711);
or U10880 (N_10880,N_8001,N_7703);
nand U10881 (N_10881,N_7639,N_7621);
xnor U10882 (N_10882,N_6870,N_6695);
or U10883 (N_10883,N_7293,N_8280);
or U10884 (N_10884,N_8362,N_8947);
nor U10885 (N_10885,N_7582,N_8321);
nand U10886 (N_10886,N_8501,N_7381);
nor U10887 (N_10887,N_8079,N_7072);
nand U10888 (N_10888,N_8640,N_7263);
nand U10889 (N_10889,N_6933,N_7685);
or U10890 (N_10890,N_8005,N_7386);
or U10891 (N_10891,N_6863,N_8615);
nand U10892 (N_10892,N_8187,N_6819);
nand U10893 (N_10893,N_8628,N_7535);
and U10894 (N_10894,N_8284,N_6802);
xor U10895 (N_10895,N_6482,N_6931);
nor U10896 (N_10896,N_6243,N_7426);
nor U10897 (N_10897,N_7846,N_6152);
and U10898 (N_10898,N_6103,N_7148);
nand U10899 (N_10899,N_8227,N_6132);
and U10900 (N_10900,N_8080,N_7939);
and U10901 (N_10901,N_7546,N_6725);
nand U10902 (N_10902,N_8444,N_7265);
and U10903 (N_10903,N_6071,N_8145);
nand U10904 (N_10904,N_6458,N_6243);
or U10905 (N_10905,N_8804,N_8290);
and U10906 (N_10906,N_7226,N_7598);
or U10907 (N_10907,N_8135,N_8782);
and U10908 (N_10908,N_8386,N_7643);
and U10909 (N_10909,N_8162,N_7394);
nor U10910 (N_10910,N_8832,N_8453);
or U10911 (N_10911,N_7435,N_8931);
nand U10912 (N_10912,N_7451,N_7178);
nor U10913 (N_10913,N_6658,N_8431);
and U10914 (N_10914,N_7494,N_7181);
nand U10915 (N_10915,N_7792,N_8654);
and U10916 (N_10916,N_7609,N_6040);
or U10917 (N_10917,N_8112,N_6202);
nor U10918 (N_10918,N_8129,N_6467);
or U10919 (N_10919,N_8472,N_8775);
xor U10920 (N_10920,N_6122,N_6079);
and U10921 (N_10921,N_8469,N_8797);
nand U10922 (N_10922,N_7822,N_7565);
nor U10923 (N_10923,N_8963,N_7736);
nor U10924 (N_10924,N_8929,N_8468);
and U10925 (N_10925,N_7144,N_8713);
nor U10926 (N_10926,N_7420,N_8086);
nor U10927 (N_10927,N_6675,N_7980);
or U10928 (N_10928,N_7539,N_6025);
nand U10929 (N_10929,N_6365,N_7366);
nand U10930 (N_10930,N_6908,N_7084);
or U10931 (N_10931,N_8732,N_6800);
and U10932 (N_10932,N_6854,N_7025);
nand U10933 (N_10933,N_6195,N_8291);
and U10934 (N_10934,N_8806,N_7351);
nor U10935 (N_10935,N_6866,N_6663);
or U10936 (N_10936,N_8126,N_8454);
or U10937 (N_10937,N_8810,N_7140);
or U10938 (N_10938,N_6123,N_6002);
nand U10939 (N_10939,N_8659,N_6407);
nor U10940 (N_10940,N_8818,N_6532);
nor U10941 (N_10941,N_7987,N_6479);
and U10942 (N_10942,N_7244,N_8590);
or U10943 (N_10943,N_6631,N_6842);
and U10944 (N_10944,N_6335,N_6272);
nand U10945 (N_10945,N_7870,N_8600);
or U10946 (N_10946,N_8788,N_7395);
or U10947 (N_10947,N_7216,N_7055);
and U10948 (N_10948,N_8145,N_7829);
and U10949 (N_10949,N_6440,N_7210);
and U10950 (N_10950,N_6466,N_8387);
and U10951 (N_10951,N_7806,N_6712);
nand U10952 (N_10952,N_7624,N_7363);
or U10953 (N_10953,N_6720,N_6035);
nor U10954 (N_10954,N_8251,N_8837);
or U10955 (N_10955,N_6106,N_7690);
and U10956 (N_10956,N_8175,N_8145);
xnor U10957 (N_10957,N_6666,N_7276);
xor U10958 (N_10958,N_7755,N_7309);
and U10959 (N_10959,N_6898,N_7846);
nand U10960 (N_10960,N_6240,N_6928);
and U10961 (N_10961,N_6058,N_6517);
nand U10962 (N_10962,N_8251,N_6259);
and U10963 (N_10963,N_8752,N_7745);
and U10964 (N_10964,N_8187,N_7823);
xor U10965 (N_10965,N_7779,N_8094);
or U10966 (N_10966,N_8569,N_7016);
xnor U10967 (N_10967,N_8727,N_8940);
nand U10968 (N_10968,N_6213,N_8905);
nor U10969 (N_10969,N_6286,N_7651);
nor U10970 (N_10970,N_8202,N_6431);
or U10971 (N_10971,N_7545,N_7071);
or U10972 (N_10972,N_6018,N_7491);
or U10973 (N_10973,N_8992,N_7966);
xor U10974 (N_10974,N_7209,N_8436);
nand U10975 (N_10975,N_8994,N_7257);
and U10976 (N_10976,N_7743,N_7404);
nand U10977 (N_10977,N_6230,N_6874);
or U10978 (N_10978,N_6408,N_7640);
nor U10979 (N_10979,N_6743,N_6253);
nor U10980 (N_10980,N_8018,N_7898);
nand U10981 (N_10981,N_7022,N_7461);
or U10982 (N_10982,N_8456,N_6164);
and U10983 (N_10983,N_7177,N_7952);
and U10984 (N_10984,N_8409,N_8764);
and U10985 (N_10985,N_8363,N_6966);
nand U10986 (N_10986,N_8070,N_8536);
and U10987 (N_10987,N_7851,N_7593);
nand U10988 (N_10988,N_7252,N_6721);
and U10989 (N_10989,N_6140,N_7659);
nor U10990 (N_10990,N_8062,N_6641);
or U10991 (N_10991,N_6234,N_8140);
xnor U10992 (N_10992,N_7991,N_8941);
xor U10993 (N_10993,N_6326,N_7762);
nor U10994 (N_10994,N_6717,N_8299);
or U10995 (N_10995,N_7525,N_8570);
and U10996 (N_10996,N_6140,N_6364);
nand U10997 (N_10997,N_8148,N_7940);
nor U10998 (N_10998,N_8867,N_7985);
nor U10999 (N_10999,N_6151,N_8217);
xnor U11000 (N_11000,N_6684,N_7449);
or U11001 (N_11001,N_6597,N_6000);
and U11002 (N_11002,N_6379,N_6599);
nand U11003 (N_11003,N_7799,N_8512);
and U11004 (N_11004,N_6993,N_8956);
nand U11005 (N_11005,N_7758,N_6402);
or U11006 (N_11006,N_7160,N_8008);
nor U11007 (N_11007,N_6623,N_6545);
or U11008 (N_11008,N_6853,N_8628);
or U11009 (N_11009,N_8038,N_8586);
nand U11010 (N_11010,N_8491,N_8628);
or U11011 (N_11011,N_7313,N_8984);
xnor U11012 (N_11012,N_8819,N_7704);
or U11013 (N_11013,N_7431,N_6440);
and U11014 (N_11014,N_6939,N_6739);
and U11015 (N_11015,N_8104,N_6482);
and U11016 (N_11016,N_8832,N_6780);
or U11017 (N_11017,N_7879,N_8945);
nand U11018 (N_11018,N_7595,N_7920);
nor U11019 (N_11019,N_8171,N_6646);
nand U11020 (N_11020,N_8413,N_8073);
nand U11021 (N_11021,N_7893,N_8082);
and U11022 (N_11022,N_7177,N_6571);
nand U11023 (N_11023,N_7367,N_7578);
nor U11024 (N_11024,N_6269,N_7352);
and U11025 (N_11025,N_7665,N_8829);
and U11026 (N_11026,N_8283,N_6603);
nor U11027 (N_11027,N_7642,N_8362);
nand U11028 (N_11028,N_7489,N_7773);
or U11029 (N_11029,N_8347,N_8277);
nand U11030 (N_11030,N_7607,N_8360);
nand U11031 (N_11031,N_6743,N_7667);
nand U11032 (N_11032,N_6448,N_8883);
nand U11033 (N_11033,N_6035,N_6689);
nand U11034 (N_11034,N_6538,N_7405);
nor U11035 (N_11035,N_6977,N_8080);
nor U11036 (N_11036,N_6908,N_6626);
or U11037 (N_11037,N_8882,N_8596);
nand U11038 (N_11038,N_7237,N_7077);
and U11039 (N_11039,N_6190,N_8684);
nor U11040 (N_11040,N_7887,N_6853);
or U11041 (N_11041,N_7257,N_6462);
or U11042 (N_11042,N_7340,N_7382);
or U11043 (N_11043,N_8404,N_8169);
nand U11044 (N_11044,N_7131,N_7841);
xnor U11045 (N_11045,N_7849,N_8596);
or U11046 (N_11046,N_8062,N_7192);
nor U11047 (N_11047,N_8506,N_7644);
and U11048 (N_11048,N_7449,N_8956);
nor U11049 (N_11049,N_7240,N_8121);
and U11050 (N_11050,N_8833,N_7224);
xor U11051 (N_11051,N_6984,N_7231);
and U11052 (N_11052,N_8415,N_6605);
nand U11053 (N_11053,N_8034,N_8216);
or U11054 (N_11054,N_6463,N_7975);
and U11055 (N_11055,N_7241,N_8212);
and U11056 (N_11056,N_6716,N_8348);
and U11057 (N_11057,N_8567,N_6913);
and U11058 (N_11058,N_6408,N_8014);
nand U11059 (N_11059,N_7846,N_8409);
nor U11060 (N_11060,N_6486,N_7128);
nor U11061 (N_11061,N_6829,N_7092);
or U11062 (N_11062,N_6843,N_7546);
or U11063 (N_11063,N_8401,N_7376);
nor U11064 (N_11064,N_8500,N_7861);
or U11065 (N_11065,N_6311,N_7522);
xor U11066 (N_11066,N_6341,N_8421);
nor U11067 (N_11067,N_7227,N_6794);
nor U11068 (N_11068,N_8439,N_8884);
and U11069 (N_11069,N_6940,N_6246);
or U11070 (N_11070,N_7887,N_6576);
nor U11071 (N_11071,N_7169,N_6895);
nand U11072 (N_11072,N_8596,N_8738);
and U11073 (N_11073,N_6886,N_6057);
or U11074 (N_11074,N_7629,N_7146);
nand U11075 (N_11075,N_6015,N_8283);
nand U11076 (N_11076,N_7257,N_6256);
nor U11077 (N_11077,N_8552,N_8238);
or U11078 (N_11078,N_7256,N_7065);
nand U11079 (N_11079,N_8115,N_6169);
or U11080 (N_11080,N_6300,N_6133);
nor U11081 (N_11081,N_6623,N_6143);
or U11082 (N_11082,N_8008,N_6772);
nand U11083 (N_11083,N_8821,N_6110);
nor U11084 (N_11084,N_6679,N_8095);
and U11085 (N_11085,N_8562,N_8785);
and U11086 (N_11086,N_6714,N_8663);
nor U11087 (N_11087,N_7806,N_6800);
or U11088 (N_11088,N_6594,N_7880);
or U11089 (N_11089,N_7782,N_7430);
nand U11090 (N_11090,N_6698,N_6427);
nand U11091 (N_11091,N_6858,N_6695);
nor U11092 (N_11092,N_7527,N_8786);
nor U11093 (N_11093,N_7368,N_8559);
or U11094 (N_11094,N_7723,N_6069);
and U11095 (N_11095,N_8065,N_6761);
xor U11096 (N_11096,N_6228,N_6873);
or U11097 (N_11097,N_6122,N_7043);
nand U11098 (N_11098,N_6986,N_7474);
and U11099 (N_11099,N_6348,N_6344);
and U11100 (N_11100,N_7759,N_8832);
or U11101 (N_11101,N_8571,N_6305);
or U11102 (N_11102,N_8357,N_6864);
nor U11103 (N_11103,N_7288,N_6138);
nor U11104 (N_11104,N_6177,N_8070);
nand U11105 (N_11105,N_7948,N_8092);
or U11106 (N_11106,N_6206,N_8031);
and U11107 (N_11107,N_6259,N_7402);
and U11108 (N_11108,N_8895,N_6798);
or U11109 (N_11109,N_8476,N_7154);
nand U11110 (N_11110,N_7806,N_6384);
or U11111 (N_11111,N_8812,N_7703);
nand U11112 (N_11112,N_6403,N_7959);
or U11113 (N_11113,N_8814,N_8961);
nand U11114 (N_11114,N_8905,N_8623);
or U11115 (N_11115,N_6143,N_6448);
xor U11116 (N_11116,N_6764,N_6645);
nor U11117 (N_11117,N_8108,N_6668);
or U11118 (N_11118,N_6962,N_8997);
or U11119 (N_11119,N_6500,N_6789);
nor U11120 (N_11120,N_6306,N_6331);
nor U11121 (N_11121,N_6104,N_6017);
and U11122 (N_11122,N_6008,N_8041);
xor U11123 (N_11123,N_7820,N_8492);
nand U11124 (N_11124,N_6526,N_7963);
xor U11125 (N_11125,N_8003,N_7774);
and U11126 (N_11126,N_7341,N_8003);
or U11127 (N_11127,N_6678,N_8007);
and U11128 (N_11128,N_8946,N_6481);
or U11129 (N_11129,N_7441,N_8169);
nand U11130 (N_11130,N_7719,N_7570);
nor U11131 (N_11131,N_8695,N_6777);
nor U11132 (N_11132,N_8216,N_7002);
or U11133 (N_11133,N_7599,N_7032);
or U11134 (N_11134,N_6189,N_8694);
and U11135 (N_11135,N_7311,N_6569);
nor U11136 (N_11136,N_8973,N_6794);
and U11137 (N_11137,N_6899,N_7706);
or U11138 (N_11138,N_8446,N_6942);
and U11139 (N_11139,N_6242,N_7123);
nor U11140 (N_11140,N_6687,N_6662);
or U11141 (N_11141,N_6757,N_7521);
nand U11142 (N_11142,N_7198,N_6263);
and U11143 (N_11143,N_8506,N_8943);
or U11144 (N_11144,N_8624,N_6409);
and U11145 (N_11145,N_6593,N_8120);
and U11146 (N_11146,N_8839,N_6143);
xnor U11147 (N_11147,N_6459,N_7999);
nand U11148 (N_11148,N_8877,N_8018);
nor U11149 (N_11149,N_6175,N_7568);
nand U11150 (N_11150,N_6048,N_6973);
and U11151 (N_11151,N_6467,N_6398);
nor U11152 (N_11152,N_8680,N_6699);
and U11153 (N_11153,N_7246,N_8454);
and U11154 (N_11154,N_7797,N_6835);
nand U11155 (N_11155,N_7973,N_6669);
nor U11156 (N_11156,N_8757,N_6123);
nor U11157 (N_11157,N_6660,N_8076);
and U11158 (N_11158,N_8941,N_7367);
xor U11159 (N_11159,N_8755,N_8446);
nand U11160 (N_11160,N_8205,N_8356);
nand U11161 (N_11161,N_7291,N_7506);
xor U11162 (N_11162,N_7895,N_8667);
nand U11163 (N_11163,N_8569,N_8751);
nor U11164 (N_11164,N_7613,N_7604);
nor U11165 (N_11165,N_6443,N_8311);
and U11166 (N_11166,N_8889,N_8362);
and U11167 (N_11167,N_7985,N_8224);
and U11168 (N_11168,N_6668,N_8287);
nand U11169 (N_11169,N_6238,N_7574);
or U11170 (N_11170,N_8949,N_8530);
nor U11171 (N_11171,N_8602,N_8600);
nor U11172 (N_11172,N_6783,N_8510);
or U11173 (N_11173,N_6046,N_8244);
or U11174 (N_11174,N_6568,N_6076);
and U11175 (N_11175,N_8417,N_6025);
and U11176 (N_11176,N_7411,N_7287);
nor U11177 (N_11177,N_7027,N_8338);
nor U11178 (N_11178,N_7234,N_6919);
nor U11179 (N_11179,N_7229,N_7693);
and U11180 (N_11180,N_6996,N_7552);
and U11181 (N_11181,N_8161,N_8905);
nor U11182 (N_11182,N_7932,N_6165);
xor U11183 (N_11183,N_7341,N_6477);
or U11184 (N_11184,N_8444,N_7263);
nand U11185 (N_11185,N_6736,N_8083);
and U11186 (N_11186,N_8304,N_8514);
and U11187 (N_11187,N_6638,N_8177);
or U11188 (N_11188,N_8854,N_7556);
and U11189 (N_11189,N_6602,N_8066);
nor U11190 (N_11190,N_6361,N_8848);
or U11191 (N_11191,N_7298,N_7483);
or U11192 (N_11192,N_6391,N_7876);
nand U11193 (N_11193,N_6274,N_7505);
nor U11194 (N_11194,N_7776,N_8498);
nand U11195 (N_11195,N_6856,N_6636);
nor U11196 (N_11196,N_7542,N_8543);
and U11197 (N_11197,N_6444,N_8219);
and U11198 (N_11198,N_7600,N_8330);
or U11199 (N_11199,N_6312,N_8907);
and U11200 (N_11200,N_8350,N_7266);
nor U11201 (N_11201,N_8455,N_6471);
or U11202 (N_11202,N_6449,N_6463);
nand U11203 (N_11203,N_8421,N_8437);
nand U11204 (N_11204,N_6008,N_7605);
and U11205 (N_11205,N_7017,N_7076);
or U11206 (N_11206,N_7697,N_7853);
nand U11207 (N_11207,N_8723,N_8452);
nand U11208 (N_11208,N_7724,N_8551);
nand U11209 (N_11209,N_8111,N_6680);
and U11210 (N_11210,N_7355,N_7606);
nand U11211 (N_11211,N_8056,N_8817);
or U11212 (N_11212,N_8452,N_6961);
nand U11213 (N_11213,N_8771,N_7002);
and U11214 (N_11214,N_7467,N_8595);
and U11215 (N_11215,N_8352,N_8066);
or U11216 (N_11216,N_8272,N_7738);
nand U11217 (N_11217,N_8448,N_8557);
and U11218 (N_11218,N_8904,N_6666);
and U11219 (N_11219,N_7090,N_7870);
or U11220 (N_11220,N_7299,N_7752);
or U11221 (N_11221,N_6563,N_6330);
nand U11222 (N_11222,N_7785,N_8710);
nor U11223 (N_11223,N_6953,N_8503);
and U11224 (N_11224,N_6879,N_6501);
nor U11225 (N_11225,N_8862,N_6942);
nor U11226 (N_11226,N_6682,N_6768);
nand U11227 (N_11227,N_6538,N_6261);
nor U11228 (N_11228,N_7243,N_8099);
nor U11229 (N_11229,N_8111,N_8238);
or U11230 (N_11230,N_7985,N_7623);
and U11231 (N_11231,N_6047,N_7053);
nand U11232 (N_11232,N_6644,N_8961);
nor U11233 (N_11233,N_6900,N_7915);
nand U11234 (N_11234,N_7913,N_7370);
nor U11235 (N_11235,N_8219,N_8992);
nand U11236 (N_11236,N_6234,N_6957);
nor U11237 (N_11237,N_7690,N_8026);
and U11238 (N_11238,N_8087,N_7930);
and U11239 (N_11239,N_6739,N_7386);
or U11240 (N_11240,N_6926,N_7264);
or U11241 (N_11241,N_7539,N_6449);
nor U11242 (N_11242,N_6101,N_6894);
or U11243 (N_11243,N_7019,N_6418);
and U11244 (N_11244,N_6790,N_7935);
xor U11245 (N_11245,N_7850,N_6483);
and U11246 (N_11246,N_8029,N_8864);
nor U11247 (N_11247,N_6943,N_7799);
nor U11248 (N_11248,N_7474,N_8292);
xnor U11249 (N_11249,N_7381,N_7596);
nand U11250 (N_11250,N_7900,N_7625);
xnor U11251 (N_11251,N_7372,N_6891);
and U11252 (N_11252,N_7053,N_6616);
xnor U11253 (N_11253,N_6076,N_6722);
and U11254 (N_11254,N_6892,N_6207);
or U11255 (N_11255,N_8703,N_6519);
nor U11256 (N_11256,N_8966,N_6080);
or U11257 (N_11257,N_7561,N_6857);
nor U11258 (N_11258,N_7948,N_8558);
and U11259 (N_11259,N_6634,N_6793);
nand U11260 (N_11260,N_7517,N_7670);
nor U11261 (N_11261,N_7575,N_7747);
xnor U11262 (N_11262,N_7528,N_8371);
or U11263 (N_11263,N_8046,N_8385);
nor U11264 (N_11264,N_8304,N_6460);
and U11265 (N_11265,N_8784,N_6776);
or U11266 (N_11266,N_6675,N_7611);
and U11267 (N_11267,N_8800,N_7595);
or U11268 (N_11268,N_8265,N_8350);
nand U11269 (N_11269,N_8211,N_7539);
nand U11270 (N_11270,N_7761,N_6057);
nor U11271 (N_11271,N_8870,N_8760);
nor U11272 (N_11272,N_7122,N_6316);
or U11273 (N_11273,N_6658,N_6451);
or U11274 (N_11274,N_8800,N_8500);
or U11275 (N_11275,N_8222,N_7677);
nand U11276 (N_11276,N_7133,N_6262);
nand U11277 (N_11277,N_6243,N_7863);
nor U11278 (N_11278,N_8901,N_8397);
nor U11279 (N_11279,N_6190,N_7222);
or U11280 (N_11280,N_8845,N_6854);
xnor U11281 (N_11281,N_6934,N_8444);
or U11282 (N_11282,N_8828,N_8386);
nand U11283 (N_11283,N_6861,N_8155);
and U11284 (N_11284,N_8751,N_6923);
or U11285 (N_11285,N_8158,N_8149);
nand U11286 (N_11286,N_6895,N_8454);
xor U11287 (N_11287,N_8509,N_6328);
nor U11288 (N_11288,N_8611,N_7581);
nand U11289 (N_11289,N_6371,N_7347);
and U11290 (N_11290,N_6021,N_6000);
and U11291 (N_11291,N_6703,N_8758);
or U11292 (N_11292,N_7366,N_8178);
xnor U11293 (N_11293,N_6060,N_6327);
and U11294 (N_11294,N_7193,N_8188);
or U11295 (N_11295,N_7949,N_8758);
nand U11296 (N_11296,N_8512,N_8409);
and U11297 (N_11297,N_6289,N_6941);
and U11298 (N_11298,N_6827,N_6903);
nand U11299 (N_11299,N_8618,N_8342);
nand U11300 (N_11300,N_6716,N_8965);
xor U11301 (N_11301,N_6624,N_6400);
or U11302 (N_11302,N_6435,N_6545);
nand U11303 (N_11303,N_6736,N_6650);
or U11304 (N_11304,N_6731,N_6919);
nand U11305 (N_11305,N_7382,N_8835);
or U11306 (N_11306,N_7212,N_8059);
or U11307 (N_11307,N_7244,N_8387);
and U11308 (N_11308,N_6620,N_8482);
nand U11309 (N_11309,N_6470,N_7085);
and U11310 (N_11310,N_7674,N_6518);
nor U11311 (N_11311,N_8289,N_6642);
or U11312 (N_11312,N_6016,N_7968);
xor U11313 (N_11313,N_8983,N_7086);
or U11314 (N_11314,N_6657,N_6772);
and U11315 (N_11315,N_6735,N_6102);
and U11316 (N_11316,N_6370,N_7162);
or U11317 (N_11317,N_8474,N_6379);
or U11318 (N_11318,N_6845,N_8080);
nor U11319 (N_11319,N_8334,N_6678);
nand U11320 (N_11320,N_6479,N_7234);
or U11321 (N_11321,N_6965,N_6102);
nand U11322 (N_11322,N_6191,N_7727);
and U11323 (N_11323,N_7703,N_7285);
or U11324 (N_11324,N_7682,N_8958);
nand U11325 (N_11325,N_8657,N_6052);
and U11326 (N_11326,N_7042,N_8070);
and U11327 (N_11327,N_7623,N_7014);
nor U11328 (N_11328,N_7498,N_6285);
or U11329 (N_11329,N_6548,N_7424);
and U11330 (N_11330,N_6666,N_6372);
nor U11331 (N_11331,N_7109,N_6974);
nand U11332 (N_11332,N_8955,N_8041);
and U11333 (N_11333,N_7212,N_7611);
or U11334 (N_11334,N_6184,N_8372);
or U11335 (N_11335,N_8847,N_6944);
nand U11336 (N_11336,N_6071,N_8960);
xnor U11337 (N_11337,N_7288,N_6754);
or U11338 (N_11338,N_7902,N_8860);
nor U11339 (N_11339,N_7325,N_6977);
nor U11340 (N_11340,N_8135,N_6928);
and U11341 (N_11341,N_6287,N_6771);
or U11342 (N_11342,N_8415,N_7955);
and U11343 (N_11343,N_8480,N_7379);
nor U11344 (N_11344,N_8099,N_8512);
or U11345 (N_11345,N_7397,N_8681);
and U11346 (N_11346,N_6025,N_8526);
xor U11347 (N_11347,N_7660,N_8684);
and U11348 (N_11348,N_7431,N_8191);
and U11349 (N_11349,N_8833,N_7050);
or U11350 (N_11350,N_6073,N_7153);
nand U11351 (N_11351,N_7774,N_6710);
xor U11352 (N_11352,N_7955,N_6682);
or U11353 (N_11353,N_6298,N_8183);
and U11354 (N_11354,N_7214,N_7253);
xor U11355 (N_11355,N_7167,N_6901);
nor U11356 (N_11356,N_6585,N_8962);
and U11357 (N_11357,N_7863,N_8849);
or U11358 (N_11358,N_7798,N_8833);
nor U11359 (N_11359,N_6004,N_7960);
nor U11360 (N_11360,N_7608,N_7542);
nor U11361 (N_11361,N_7465,N_6270);
nand U11362 (N_11362,N_8799,N_6004);
nor U11363 (N_11363,N_7404,N_8517);
and U11364 (N_11364,N_6513,N_6534);
nor U11365 (N_11365,N_8635,N_7561);
nand U11366 (N_11366,N_7067,N_6476);
nor U11367 (N_11367,N_6477,N_7814);
and U11368 (N_11368,N_8932,N_7889);
or U11369 (N_11369,N_8800,N_8129);
and U11370 (N_11370,N_6960,N_6769);
or U11371 (N_11371,N_7376,N_6851);
xor U11372 (N_11372,N_8669,N_8278);
nand U11373 (N_11373,N_8258,N_8993);
and U11374 (N_11374,N_6988,N_7840);
nor U11375 (N_11375,N_6513,N_8014);
nor U11376 (N_11376,N_6854,N_7125);
nor U11377 (N_11377,N_6905,N_7522);
and U11378 (N_11378,N_7504,N_7144);
nor U11379 (N_11379,N_8367,N_7079);
nor U11380 (N_11380,N_8152,N_7165);
nor U11381 (N_11381,N_8505,N_6877);
and U11382 (N_11382,N_7833,N_7795);
nor U11383 (N_11383,N_8176,N_6823);
nor U11384 (N_11384,N_7146,N_8671);
xor U11385 (N_11385,N_8790,N_8415);
or U11386 (N_11386,N_7600,N_8636);
and U11387 (N_11387,N_7565,N_6619);
or U11388 (N_11388,N_8030,N_8813);
nand U11389 (N_11389,N_6798,N_6148);
or U11390 (N_11390,N_6167,N_6941);
or U11391 (N_11391,N_8311,N_7056);
or U11392 (N_11392,N_8714,N_6262);
or U11393 (N_11393,N_7595,N_7628);
nor U11394 (N_11394,N_7240,N_6687);
and U11395 (N_11395,N_7622,N_7489);
or U11396 (N_11396,N_8500,N_6086);
nor U11397 (N_11397,N_8901,N_7437);
xor U11398 (N_11398,N_7027,N_8983);
nor U11399 (N_11399,N_6132,N_6866);
and U11400 (N_11400,N_7063,N_6854);
or U11401 (N_11401,N_6446,N_8708);
or U11402 (N_11402,N_6662,N_7222);
nand U11403 (N_11403,N_6923,N_6302);
nor U11404 (N_11404,N_8153,N_7599);
xnor U11405 (N_11405,N_8676,N_8536);
or U11406 (N_11406,N_7949,N_7987);
and U11407 (N_11407,N_8138,N_7069);
xor U11408 (N_11408,N_7013,N_7432);
or U11409 (N_11409,N_6811,N_7712);
or U11410 (N_11410,N_7247,N_8038);
nand U11411 (N_11411,N_6449,N_7895);
and U11412 (N_11412,N_6755,N_8987);
and U11413 (N_11413,N_8674,N_8003);
nand U11414 (N_11414,N_6788,N_6582);
and U11415 (N_11415,N_8786,N_7208);
nor U11416 (N_11416,N_7786,N_6235);
nand U11417 (N_11417,N_7378,N_7320);
xor U11418 (N_11418,N_6926,N_7835);
nand U11419 (N_11419,N_7669,N_6840);
and U11420 (N_11420,N_7681,N_7226);
or U11421 (N_11421,N_7127,N_6533);
and U11422 (N_11422,N_8231,N_7920);
and U11423 (N_11423,N_7427,N_6440);
and U11424 (N_11424,N_6279,N_8628);
and U11425 (N_11425,N_7522,N_8828);
nor U11426 (N_11426,N_7595,N_8557);
nor U11427 (N_11427,N_7443,N_7340);
or U11428 (N_11428,N_6519,N_7573);
nand U11429 (N_11429,N_6120,N_7426);
or U11430 (N_11430,N_7299,N_6705);
nor U11431 (N_11431,N_8961,N_6408);
nor U11432 (N_11432,N_6771,N_7426);
or U11433 (N_11433,N_8801,N_8183);
or U11434 (N_11434,N_6191,N_6256);
or U11435 (N_11435,N_7513,N_7088);
nand U11436 (N_11436,N_6845,N_7523);
or U11437 (N_11437,N_8306,N_7032);
nor U11438 (N_11438,N_8036,N_8661);
or U11439 (N_11439,N_7521,N_7538);
and U11440 (N_11440,N_8261,N_8820);
nor U11441 (N_11441,N_7161,N_6140);
or U11442 (N_11442,N_7180,N_6059);
nor U11443 (N_11443,N_6709,N_6904);
xnor U11444 (N_11444,N_7749,N_8800);
or U11445 (N_11445,N_6461,N_7013);
or U11446 (N_11446,N_6834,N_7896);
or U11447 (N_11447,N_8814,N_6261);
and U11448 (N_11448,N_6633,N_6463);
nor U11449 (N_11449,N_6946,N_6439);
xor U11450 (N_11450,N_7721,N_7415);
nor U11451 (N_11451,N_7843,N_8814);
xnor U11452 (N_11452,N_6928,N_6645);
or U11453 (N_11453,N_7206,N_8609);
nand U11454 (N_11454,N_7186,N_6523);
nor U11455 (N_11455,N_7994,N_6329);
and U11456 (N_11456,N_6940,N_6467);
xnor U11457 (N_11457,N_6526,N_8382);
nand U11458 (N_11458,N_6881,N_6292);
nand U11459 (N_11459,N_7189,N_7778);
nor U11460 (N_11460,N_6934,N_7865);
xnor U11461 (N_11461,N_8225,N_8977);
or U11462 (N_11462,N_8853,N_6977);
nor U11463 (N_11463,N_7343,N_8894);
and U11464 (N_11464,N_6871,N_8758);
nor U11465 (N_11465,N_6989,N_8919);
and U11466 (N_11466,N_6117,N_6924);
or U11467 (N_11467,N_6266,N_6178);
and U11468 (N_11468,N_8325,N_8530);
or U11469 (N_11469,N_6844,N_7033);
xnor U11470 (N_11470,N_7353,N_7772);
nand U11471 (N_11471,N_6470,N_6602);
nand U11472 (N_11472,N_7184,N_7418);
or U11473 (N_11473,N_7312,N_6066);
and U11474 (N_11474,N_6277,N_6462);
nand U11475 (N_11475,N_6535,N_8971);
nand U11476 (N_11476,N_8907,N_7054);
xnor U11477 (N_11477,N_6623,N_6965);
nand U11478 (N_11478,N_7000,N_7307);
nor U11479 (N_11479,N_7517,N_7929);
and U11480 (N_11480,N_6295,N_8174);
and U11481 (N_11481,N_8172,N_6500);
and U11482 (N_11482,N_8668,N_8667);
nor U11483 (N_11483,N_7868,N_7884);
xor U11484 (N_11484,N_6851,N_8160);
nor U11485 (N_11485,N_8639,N_6975);
xnor U11486 (N_11486,N_7551,N_7618);
nand U11487 (N_11487,N_8112,N_6155);
and U11488 (N_11488,N_7092,N_6811);
nand U11489 (N_11489,N_7724,N_7616);
or U11490 (N_11490,N_7028,N_7806);
and U11491 (N_11491,N_8246,N_8517);
nand U11492 (N_11492,N_7042,N_6425);
or U11493 (N_11493,N_8202,N_8997);
nor U11494 (N_11494,N_8327,N_8241);
nand U11495 (N_11495,N_6378,N_6358);
nor U11496 (N_11496,N_6295,N_7230);
xnor U11497 (N_11497,N_8158,N_6980);
or U11498 (N_11498,N_8896,N_8795);
nor U11499 (N_11499,N_6528,N_7285);
or U11500 (N_11500,N_7546,N_8083);
or U11501 (N_11501,N_7308,N_8162);
nor U11502 (N_11502,N_8060,N_7073);
nand U11503 (N_11503,N_8547,N_7003);
nand U11504 (N_11504,N_7217,N_8212);
or U11505 (N_11505,N_6280,N_7957);
and U11506 (N_11506,N_8014,N_8547);
nor U11507 (N_11507,N_7886,N_6622);
and U11508 (N_11508,N_8289,N_6212);
or U11509 (N_11509,N_7267,N_6097);
nor U11510 (N_11510,N_6282,N_8168);
or U11511 (N_11511,N_7349,N_6122);
nor U11512 (N_11512,N_6020,N_8830);
or U11513 (N_11513,N_8211,N_6851);
or U11514 (N_11514,N_8743,N_7164);
nor U11515 (N_11515,N_8933,N_7036);
and U11516 (N_11516,N_6136,N_6380);
nor U11517 (N_11517,N_7180,N_7687);
nor U11518 (N_11518,N_6143,N_6398);
nor U11519 (N_11519,N_6450,N_7549);
and U11520 (N_11520,N_6688,N_8292);
and U11521 (N_11521,N_6337,N_7681);
and U11522 (N_11522,N_6489,N_7544);
nor U11523 (N_11523,N_7125,N_6219);
and U11524 (N_11524,N_8925,N_6206);
nor U11525 (N_11525,N_8857,N_8540);
or U11526 (N_11526,N_6115,N_8913);
and U11527 (N_11527,N_7560,N_7978);
or U11528 (N_11528,N_7742,N_7396);
xor U11529 (N_11529,N_6928,N_7594);
nand U11530 (N_11530,N_8057,N_8563);
nand U11531 (N_11531,N_8010,N_8387);
or U11532 (N_11532,N_6169,N_8095);
and U11533 (N_11533,N_7761,N_6076);
nor U11534 (N_11534,N_7718,N_8946);
and U11535 (N_11535,N_7784,N_8238);
nand U11536 (N_11536,N_6612,N_8324);
nand U11537 (N_11537,N_7974,N_6311);
and U11538 (N_11538,N_6139,N_6635);
nor U11539 (N_11539,N_8591,N_6355);
nor U11540 (N_11540,N_8364,N_7525);
and U11541 (N_11541,N_8873,N_8663);
nor U11542 (N_11542,N_6237,N_8522);
and U11543 (N_11543,N_6006,N_7423);
nand U11544 (N_11544,N_7956,N_8176);
and U11545 (N_11545,N_8269,N_7042);
and U11546 (N_11546,N_7634,N_6523);
nor U11547 (N_11547,N_7173,N_6892);
nor U11548 (N_11548,N_7256,N_8622);
or U11549 (N_11549,N_8687,N_7969);
nand U11550 (N_11550,N_6198,N_6136);
and U11551 (N_11551,N_7255,N_8514);
or U11552 (N_11552,N_7277,N_7297);
or U11553 (N_11553,N_6889,N_7859);
nand U11554 (N_11554,N_6844,N_8914);
or U11555 (N_11555,N_8377,N_6112);
nand U11556 (N_11556,N_7878,N_8993);
nor U11557 (N_11557,N_7917,N_8189);
xnor U11558 (N_11558,N_8595,N_6287);
and U11559 (N_11559,N_6229,N_8661);
xnor U11560 (N_11560,N_7128,N_6604);
nor U11561 (N_11561,N_7533,N_8928);
nand U11562 (N_11562,N_7275,N_8017);
and U11563 (N_11563,N_7944,N_7995);
and U11564 (N_11564,N_6808,N_7170);
nand U11565 (N_11565,N_7719,N_8440);
nor U11566 (N_11566,N_7805,N_7477);
or U11567 (N_11567,N_6257,N_6274);
xnor U11568 (N_11568,N_7426,N_6295);
and U11569 (N_11569,N_7041,N_6720);
or U11570 (N_11570,N_8401,N_6717);
and U11571 (N_11571,N_7744,N_7160);
xnor U11572 (N_11572,N_7320,N_7957);
and U11573 (N_11573,N_8686,N_6883);
and U11574 (N_11574,N_6211,N_6124);
nand U11575 (N_11575,N_8452,N_8281);
nand U11576 (N_11576,N_8462,N_6061);
xor U11577 (N_11577,N_7896,N_6548);
nand U11578 (N_11578,N_7332,N_6447);
nor U11579 (N_11579,N_8938,N_7094);
nand U11580 (N_11580,N_6651,N_6292);
nand U11581 (N_11581,N_7209,N_7447);
nor U11582 (N_11582,N_6356,N_6514);
or U11583 (N_11583,N_8868,N_7115);
xnor U11584 (N_11584,N_6237,N_8876);
and U11585 (N_11585,N_6700,N_6417);
nor U11586 (N_11586,N_6689,N_8357);
nand U11587 (N_11587,N_8130,N_7710);
or U11588 (N_11588,N_7566,N_7821);
and U11589 (N_11589,N_7519,N_6489);
nand U11590 (N_11590,N_7724,N_6911);
nor U11591 (N_11591,N_8100,N_8539);
nand U11592 (N_11592,N_8473,N_8318);
or U11593 (N_11593,N_7192,N_7513);
nor U11594 (N_11594,N_8024,N_6351);
xnor U11595 (N_11595,N_6088,N_8973);
nand U11596 (N_11596,N_6536,N_8671);
nor U11597 (N_11597,N_6112,N_8207);
xnor U11598 (N_11598,N_6297,N_7324);
or U11599 (N_11599,N_6397,N_8929);
and U11600 (N_11600,N_8962,N_6621);
nand U11601 (N_11601,N_6082,N_7106);
nor U11602 (N_11602,N_6448,N_6895);
or U11603 (N_11603,N_7006,N_8334);
nor U11604 (N_11604,N_6040,N_8458);
and U11605 (N_11605,N_7076,N_7667);
or U11606 (N_11606,N_7741,N_7099);
or U11607 (N_11607,N_8962,N_6652);
or U11608 (N_11608,N_6556,N_7385);
nand U11609 (N_11609,N_6179,N_8101);
nand U11610 (N_11610,N_7305,N_7270);
xnor U11611 (N_11611,N_7757,N_7693);
and U11612 (N_11612,N_7254,N_7718);
xor U11613 (N_11613,N_8227,N_8716);
nand U11614 (N_11614,N_7179,N_7999);
or U11615 (N_11615,N_7085,N_6149);
or U11616 (N_11616,N_8850,N_8937);
or U11617 (N_11617,N_7931,N_7860);
nor U11618 (N_11618,N_6425,N_6599);
nand U11619 (N_11619,N_6461,N_8877);
nand U11620 (N_11620,N_7403,N_6307);
nand U11621 (N_11621,N_6703,N_7518);
nor U11622 (N_11622,N_8270,N_6419);
nor U11623 (N_11623,N_8503,N_8108);
nor U11624 (N_11624,N_7749,N_8593);
xnor U11625 (N_11625,N_8548,N_8939);
and U11626 (N_11626,N_7994,N_6614);
nor U11627 (N_11627,N_6026,N_8742);
nand U11628 (N_11628,N_8511,N_7695);
nand U11629 (N_11629,N_6855,N_8621);
and U11630 (N_11630,N_7608,N_6502);
xor U11631 (N_11631,N_7493,N_6508);
nand U11632 (N_11632,N_6322,N_6161);
or U11633 (N_11633,N_7329,N_8071);
nor U11634 (N_11634,N_8837,N_6035);
nand U11635 (N_11635,N_8885,N_7916);
and U11636 (N_11636,N_8287,N_7701);
nand U11637 (N_11637,N_6399,N_6839);
nor U11638 (N_11638,N_8427,N_8541);
and U11639 (N_11639,N_8681,N_7965);
xnor U11640 (N_11640,N_7131,N_6713);
and U11641 (N_11641,N_8129,N_6714);
nand U11642 (N_11642,N_6304,N_6243);
nand U11643 (N_11643,N_6297,N_7523);
nor U11644 (N_11644,N_7107,N_8352);
nor U11645 (N_11645,N_7069,N_8810);
nand U11646 (N_11646,N_6972,N_8980);
nor U11647 (N_11647,N_6821,N_8644);
and U11648 (N_11648,N_7498,N_7581);
or U11649 (N_11649,N_7415,N_7929);
or U11650 (N_11650,N_7105,N_8799);
nor U11651 (N_11651,N_8756,N_7985);
or U11652 (N_11652,N_6184,N_8104);
xor U11653 (N_11653,N_7892,N_6300);
xnor U11654 (N_11654,N_8702,N_7262);
and U11655 (N_11655,N_8311,N_7678);
xor U11656 (N_11656,N_7793,N_6953);
nor U11657 (N_11657,N_8877,N_8636);
nor U11658 (N_11658,N_7314,N_7129);
nor U11659 (N_11659,N_8593,N_6709);
nand U11660 (N_11660,N_6913,N_7424);
and U11661 (N_11661,N_8523,N_6662);
or U11662 (N_11662,N_8096,N_8504);
xnor U11663 (N_11663,N_6844,N_7960);
nor U11664 (N_11664,N_6641,N_6803);
xor U11665 (N_11665,N_8719,N_7956);
and U11666 (N_11666,N_7406,N_7105);
or U11667 (N_11667,N_6343,N_6598);
nor U11668 (N_11668,N_7430,N_8429);
and U11669 (N_11669,N_7066,N_6421);
nand U11670 (N_11670,N_6978,N_6606);
or U11671 (N_11671,N_8766,N_8138);
or U11672 (N_11672,N_6327,N_7639);
nor U11673 (N_11673,N_8568,N_7480);
nor U11674 (N_11674,N_8792,N_7390);
xnor U11675 (N_11675,N_7305,N_7661);
xnor U11676 (N_11676,N_6678,N_6713);
and U11677 (N_11677,N_8131,N_6864);
and U11678 (N_11678,N_6894,N_6788);
nor U11679 (N_11679,N_7081,N_7536);
nor U11680 (N_11680,N_7467,N_7913);
or U11681 (N_11681,N_6307,N_8240);
nand U11682 (N_11682,N_7946,N_7504);
nand U11683 (N_11683,N_6624,N_8975);
or U11684 (N_11684,N_8595,N_8816);
nand U11685 (N_11685,N_6934,N_6335);
or U11686 (N_11686,N_7828,N_8453);
nand U11687 (N_11687,N_6117,N_7729);
and U11688 (N_11688,N_8104,N_6860);
or U11689 (N_11689,N_8007,N_6437);
and U11690 (N_11690,N_6203,N_8092);
and U11691 (N_11691,N_8036,N_6436);
nor U11692 (N_11692,N_7539,N_7995);
xnor U11693 (N_11693,N_7848,N_8984);
nor U11694 (N_11694,N_7485,N_6181);
xor U11695 (N_11695,N_8017,N_6561);
xor U11696 (N_11696,N_8879,N_6031);
xnor U11697 (N_11697,N_7113,N_6009);
xnor U11698 (N_11698,N_7895,N_6352);
nand U11699 (N_11699,N_6406,N_8375);
and U11700 (N_11700,N_8177,N_8661);
or U11701 (N_11701,N_7213,N_7733);
nor U11702 (N_11702,N_6383,N_6988);
or U11703 (N_11703,N_7988,N_8284);
or U11704 (N_11704,N_7316,N_6338);
nand U11705 (N_11705,N_6308,N_8946);
or U11706 (N_11706,N_7355,N_6838);
nand U11707 (N_11707,N_8522,N_8512);
or U11708 (N_11708,N_8740,N_8697);
nand U11709 (N_11709,N_8618,N_8884);
nor U11710 (N_11710,N_8043,N_8417);
nor U11711 (N_11711,N_7262,N_8654);
nand U11712 (N_11712,N_8740,N_8266);
and U11713 (N_11713,N_7019,N_6129);
and U11714 (N_11714,N_6963,N_8690);
nand U11715 (N_11715,N_7449,N_6818);
nor U11716 (N_11716,N_8033,N_6689);
xnor U11717 (N_11717,N_7311,N_6805);
nand U11718 (N_11718,N_6190,N_6967);
nand U11719 (N_11719,N_8906,N_7091);
nand U11720 (N_11720,N_8819,N_7662);
or U11721 (N_11721,N_8780,N_6890);
xor U11722 (N_11722,N_6972,N_7032);
nor U11723 (N_11723,N_6874,N_6355);
nand U11724 (N_11724,N_6306,N_8111);
nor U11725 (N_11725,N_8095,N_8881);
nand U11726 (N_11726,N_6948,N_7799);
or U11727 (N_11727,N_7445,N_8543);
xor U11728 (N_11728,N_7941,N_7625);
nand U11729 (N_11729,N_6296,N_7950);
and U11730 (N_11730,N_6015,N_7450);
nand U11731 (N_11731,N_6297,N_6400);
nor U11732 (N_11732,N_7438,N_6336);
nor U11733 (N_11733,N_7469,N_7003);
or U11734 (N_11734,N_8912,N_6269);
nand U11735 (N_11735,N_7706,N_8368);
nor U11736 (N_11736,N_8558,N_7972);
and U11737 (N_11737,N_8743,N_6996);
or U11738 (N_11738,N_8638,N_7911);
nor U11739 (N_11739,N_6268,N_6843);
or U11740 (N_11740,N_7057,N_8390);
nand U11741 (N_11741,N_8650,N_7489);
nand U11742 (N_11742,N_8192,N_7014);
and U11743 (N_11743,N_7087,N_7359);
and U11744 (N_11744,N_7627,N_8080);
and U11745 (N_11745,N_7060,N_6453);
or U11746 (N_11746,N_7280,N_7217);
or U11747 (N_11747,N_8310,N_8704);
nand U11748 (N_11748,N_6948,N_6822);
nor U11749 (N_11749,N_7329,N_8136);
or U11750 (N_11750,N_6849,N_6608);
nand U11751 (N_11751,N_6205,N_8315);
and U11752 (N_11752,N_6209,N_8557);
and U11753 (N_11753,N_7351,N_7988);
nand U11754 (N_11754,N_8812,N_6659);
and U11755 (N_11755,N_7971,N_8806);
nand U11756 (N_11756,N_6799,N_7030);
and U11757 (N_11757,N_6037,N_7024);
or U11758 (N_11758,N_6514,N_7416);
nand U11759 (N_11759,N_7426,N_8394);
and U11760 (N_11760,N_6030,N_8190);
or U11761 (N_11761,N_7922,N_8965);
nand U11762 (N_11762,N_7658,N_8221);
nand U11763 (N_11763,N_7385,N_6816);
or U11764 (N_11764,N_6937,N_8103);
nor U11765 (N_11765,N_7173,N_8811);
nor U11766 (N_11766,N_7765,N_8136);
nand U11767 (N_11767,N_7230,N_8757);
nand U11768 (N_11768,N_7565,N_7714);
nand U11769 (N_11769,N_8551,N_8848);
or U11770 (N_11770,N_8689,N_6715);
nor U11771 (N_11771,N_8764,N_6154);
nand U11772 (N_11772,N_7323,N_6992);
or U11773 (N_11773,N_8321,N_7438);
xor U11774 (N_11774,N_8887,N_7167);
and U11775 (N_11775,N_6719,N_7354);
and U11776 (N_11776,N_6038,N_7154);
or U11777 (N_11777,N_6652,N_8354);
nand U11778 (N_11778,N_7552,N_8198);
or U11779 (N_11779,N_8938,N_6514);
nor U11780 (N_11780,N_6845,N_8948);
or U11781 (N_11781,N_6213,N_7793);
and U11782 (N_11782,N_6545,N_6175);
or U11783 (N_11783,N_7028,N_6729);
or U11784 (N_11784,N_8966,N_7023);
nor U11785 (N_11785,N_7162,N_8625);
nor U11786 (N_11786,N_7107,N_7156);
and U11787 (N_11787,N_8365,N_7074);
nor U11788 (N_11788,N_6086,N_6292);
and U11789 (N_11789,N_6626,N_6091);
or U11790 (N_11790,N_6294,N_7315);
or U11791 (N_11791,N_7737,N_8124);
and U11792 (N_11792,N_7182,N_7624);
nor U11793 (N_11793,N_7104,N_8781);
nand U11794 (N_11794,N_7100,N_8960);
or U11795 (N_11795,N_8042,N_8866);
or U11796 (N_11796,N_6200,N_7468);
and U11797 (N_11797,N_8536,N_6877);
or U11798 (N_11798,N_8333,N_6554);
xor U11799 (N_11799,N_7664,N_8247);
xnor U11800 (N_11800,N_6748,N_8055);
or U11801 (N_11801,N_6698,N_8281);
nand U11802 (N_11802,N_6097,N_8533);
nor U11803 (N_11803,N_7551,N_7766);
or U11804 (N_11804,N_7198,N_7700);
or U11805 (N_11805,N_7230,N_8466);
and U11806 (N_11806,N_8185,N_8017);
xnor U11807 (N_11807,N_8475,N_8281);
or U11808 (N_11808,N_7873,N_6391);
nor U11809 (N_11809,N_7923,N_7137);
or U11810 (N_11810,N_8482,N_8383);
and U11811 (N_11811,N_6988,N_8440);
or U11812 (N_11812,N_7523,N_6106);
nor U11813 (N_11813,N_6656,N_6002);
nand U11814 (N_11814,N_7519,N_7804);
xnor U11815 (N_11815,N_7590,N_6654);
nand U11816 (N_11816,N_7642,N_7576);
nand U11817 (N_11817,N_7980,N_8947);
nand U11818 (N_11818,N_6424,N_6978);
and U11819 (N_11819,N_8976,N_7417);
and U11820 (N_11820,N_6358,N_7146);
and U11821 (N_11821,N_6281,N_8147);
nand U11822 (N_11822,N_8635,N_8686);
nand U11823 (N_11823,N_6804,N_6271);
xnor U11824 (N_11824,N_8706,N_6806);
and U11825 (N_11825,N_8194,N_7375);
nor U11826 (N_11826,N_8392,N_7223);
and U11827 (N_11827,N_8019,N_6437);
nor U11828 (N_11828,N_6727,N_6496);
or U11829 (N_11829,N_7158,N_7001);
or U11830 (N_11830,N_7283,N_6590);
and U11831 (N_11831,N_6438,N_7577);
nor U11832 (N_11832,N_6609,N_6965);
nand U11833 (N_11833,N_8825,N_7772);
xor U11834 (N_11834,N_6672,N_6289);
or U11835 (N_11835,N_6043,N_7323);
nand U11836 (N_11836,N_8871,N_8422);
nand U11837 (N_11837,N_8485,N_7457);
nor U11838 (N_11838,N_7470,N_8192);
nand U11839 (N_11839,N_6826,N_7332);
nand U11840 (N_11840,N_8301,N_7471);
or U11841 (N_11841,N_6773,N_7141);
and U11842 (N_11842,N_6407,N_7644);
nand U11843 (N_11843,N_7597,N_6709);
xor U11844 (N_11844,N_8048,N_8116);
nand U11845 (N_11845,N_8655,N_6715);
nor U11846 (N_11846,N_7895,N_8588);
or U11847 (N_11847,N_7578,N_8445);
xnor U11848 (N_11848,N_8953,N_7189);
nor U11849 (N_11849,N_7605,N_6377);
nor U11850 (N_11850,N_8862,N_8369);
nand U11851 (N_11851,N_6849,N_8621);
nand U11852 (N_11852,N_7069,N_7978);
nor U11853 (N_11853,N_6975,N_7857);
nand U11854 (N_11854,N_7077,N_7793);
and U11855 (N_11855,N_8373,N_7220);
nand U11856 (N_11856,N_8654,N_6234);
nor U11857 (N_11857,N_6581,N_7703);
and U11858 (N_11858,N_6829,N_7438);
or U11859 (N_11859,N_6442,N_8398);
nor U11860 (N_11860,N_7311,N_8559);
xnor U11861 (N_11861,N_8091,N_7562);
xor U11862 (N_11862,N_7631,N_7876);
nand U11863 (N_11863,N_6686,N_6993);
nor U11864 (N_11864,N_7056,N_7251);
or U11865 (N_11865,N_7128,N_8084);
and U11866 (N_11866,N_7002,N_8312);
nand U11867 (N_11867,N_6700,N_7133);
and U11868 (N_11868,N_7241,N_8293);
and U11869 (N_11869,N_6286,N_8830);
xnor U11870 (N_11870,N_6353,N_7564);
and U11871 (N_11871,N_7274,N_7238);
or U11872 (N_11872,N_6337,N_7058);
nand U11873 (N_11873,N_6441,N_8193);
nand U11874 (N_11874,N_7265,N_8197);
or U11875 (N_11875,N_7836,N_7147);
or U11876 (N_11876,N_7090,N_8557);
or U11877 (N_11877,N_7916,N_6462);
nand U11878 (N_11878,N_7733,N_8195);
nand U11879 (N_11879,N_6949,N_7965);
and U11880 (N_11880,N_6581,N_8755);
nand U11881 (N_11881,N_8127,N_6880);
nor U11882 (N_11882,N_6199,N_6197);
nor U11883 (N_11883,N_7960,N_8591);
nand U11884 (N_11884,N_8574,N_8512);
and U11885 (N_11885,N_6154,N_8585);
and U11886 (N_11886,N_7137,N_7861);
nand U11887 (N_11887,N_6395,N_7139);
nand U11888 (N_11888,N_6984,N_8851);
nand U11889 (N_11889,N_8823,N_8092);
nor U11890 (N_11890,N_7921,N_7438);
and U11891 (N_11891,N_8277,N_6616);
or U11892 (N_11892,N_6463,N_6024);
or U11893 (N_11893,N_6279,N_6595);
or U11894 (N_11894,N_7216,N_8162);
or U11895 (N_11895,N_8227,N_7261);
or U11896 (N_11896,N_8753,N_7771);
nor U11897 (N_11897,N_8392,N_6257);
nor U11898 (N_11898,N_7651,N_8762);
nand U11899 (N_11899,N_8446,N_7289);
nor U11900 (N_11900,N_8295,N_8977);
nand U11901 (N_11901,N_8803,N_8738);
or U11902 (N_11902,N_6631,N_6989);
and U11903 (N_11903,N_6940,N_8746);
xor U11904 (N_11904,N_7237,N_8674);
or U11905 (N_11905,N_6762,N_6679);
and U11906 (N_11906,N_6223,N_7293);
nand U11907 (N_11907,N_8288,N_7331);
and U11908 (N_11908,N_8856,N_7266);
xor U11909 (N_11909,N_7042,N_6152);
nor U11910 (N_11910,N_8597,N_6351);
and U11911 (N_11911,N_7750,N_7293);
xor U11912 (N_11912,N_8367,N_6560);
nand U11913 (N_11913,N_6024,N_8226);
xor U11914 (N_11914,N_8895,N_7066);
nand U11915 (N_11915,N_7027,N_6071);
and U11916 (N_11916,N_6243,N_6779);
and U11917 (N_11917,N_8697,N_7310);
nor U11918 (N_11918,N_8803,N_6226);
and U11919 (N_11919,N_7768,N_7196);
xor U11920 (N_11920,N_7946,N_8023);
nor U11921 (N_11921,N_7943,N_8847);
nor U11922 (N_11922,N_7179,N_8253);
nor U11923 (N_11923,N_7378,N_6170);
or U11924 (N_11924,N_8716,N_6284);
nor U11925 (N_11925,N_6080,N_7426);
nand U11926 (N_11926,N_6372,N_7362);
nor U11927 (N_11927,N_6820,N_7469);
or U11928 (N_11928,N_8989,N_6527);
or U11929 (N_11929,N_7941,N_6664);
nor U11930 (N_11930,N_6169,N_6743);
nor U11931 (N_11931,N_6761,N_8580);
xnor U11932 (N_11932,N_8793,N_6426);
nor U11933 (N_11933,N_7546,N_6630);
nand U11934 (N_11934,N_6815,N_6521);
xnor U11935 (N_11935,N_7612,N_8241);
and U11936 (N_11936,N_7716,N_7638);
nor U11937 (N_11937,N_7943,N_7551);
nand U11938 (N_11938,N_6249,N_7979);
nor U11939 (N_11939,N_8672,N_8637);
and U11940 (N_11940,N_6659,N_7442);
or U11941 (N_11941,N_8038,N_6820);
nand U11942 (N_11942,N_6326,N_7719);
nor U11943 (N_11943,N_6516,N_7716);
nor U11944 (N_11944,N_8904,N_7635);
or U11945 (N_11945,N_8582,N_8954);
and U11946 (N_11946,N_8754,N_6232);
nand U11947 (N_11947,N_8644,N_7971);
or U11948 (N_11948,N_7228,N_6961);
and U11949 (N_11949,N_6727,N_7668);
nand U11950 (N_11950,N_6551,N_8158);
nor U11951 (N_11951,N_6454,N_7124);
and U11952 (N_11952,N_7604,N_8622);
nand U11953 (N_11953,N_7842,N_8542);
xnor U11954 (N_11954,N_6951,N_7279);
or U11955 (N_11955,N_6111,N_8946);
xnor U11956 (N_11956,N_6142,N_6368);
and U11957 (N_11957,N_7809,N_8429);
or U11958 (N_11958,N_7461,N_6474);
and U11959 (N_11959,N_8634,N_7190);
nand U11960 (N_11960,N_6800,N_8987);
xor U11961 (N_11961,N_7774,N_6846);
or U11962 (N_11962,N_6560,N_8021);
or U11963 (N_11963,N_7844,N_8732);
and U11964 (N_11964,N_8989,N_6992);
and U11965 (N_11965,N_6007,N_7725);
and U11966 (N_11966,N_7834,N_7888);
nand U11967 (N_11967,N_6357,N_7425);
nand U11968 (N_11968,N_8336,N_7450);
xnor U11969 (N_11969,N_6358,N_8682);
or U11970 (N_11970,N_8364,N_6858);
nand U11971 (N_11971,N_8067,N_8762);
or U11972 (N_11972,N_6300,N_6692);
xnor U11973 (N_11973,N_7834,N_8043);
xor U11974 (N_11974,N_6771,N_6269);
and U11975 (N_11975,N_6251,N_7553);
xor U11976 (N_11976,N_7841,N_8485);
or U11977 (N_11977,N_8803,N_7521);
nand U11978 (N_11978,N_7991,N_6049);
and U11979 (N_11979,N_7998,N_6503);
and U11980 (N_11980,N_6134,N_7044);
or U11981 (N_11981,N_7672,N_6564);
and U11982 (N_11982,N_7110,N_6701);
nor U11983 (N_11983,N_6545,N_8224);
nor U11984 (N_11984,N_6360,N_7592);
or U11985 (N_11985,N_7170,N_6706);
and U11986 (N_11986,N_7210,N_8208);
nor U11987 (N_11987,N_8912,N_7101);
or U11988 (N_11988,N_6399,N_8155);
nor U11989 (N_11989,N_6678,N_7094);
nor U11990 (N_11990,N_8041,N_6342);
xnor U11991 (N_11991,N_6076,N_8059);
or U11992 (N_11992,N_6832,N_6189);
nand U11993 (N_11993,N_6579,N_8621);
nor U11994 (N_11994,N_8139,N_6958);
xor U11995 (N_11995,N_7556,N_7199);
nand U11996 (N_11996,N_6388,N_7142);
nor U11997 (N_11997,N_6319,N_8698);
or U11998 (N_11998,N_8860,N_8757);
nor U11999 (N_11999,N_7732,N_6824);
and U12000 (N_12000,N_11222,N_11260);
nand U12001 (N_12001,N_11698,N_11475);
or U12002 (N_12002,N_10068,N_9178);
nand U12003 (N_12003,N_11280,N_11223);
nor U12004 (N_12004,N_9455,N_9460);
nand U12005 (N_12005,N_10364,N_11881);
and U12006 (N_12006,N_9132,N_9692);
nand U12007 (N_12007,N_10144,N_10275);
and U12008 (N_12008,N_10266,N_11840);
and U12009 (N_12009,N_9166,N_10050);
xnor U12010 (N_12010,N_11586,N_9246);
nand U12011 (N_12011,N_10365,N_10646);
or U12012 (N_12012,N_9298,N_10340);
nor U12013 (N_12013,N_9661,N_10138);
or U12014 (N_12014,N_11438,N_11392);
xor U12015 (N_12015,N_10710,N_11358);
nand U12016 (N_12016,N_9792,N_10557);
or U12017 (N_12017,N_10383,N_10752);
xor U12018 (N_12018,N_10343,N_11926);
and U12019 (N_12019,N_11110,N_11111);
and U12020 (N_12020,N_9119,N_11718);
and U12021 (N_12021,N_9960,N_9948);
xor U12022 (N_12022,N_9799,N_11080);
xor U12023 (N_12023,N_9289,N_11179);
and U12024 (N_12024,N_11776,N_11020);
nand U12025 (N_12025,N_10886,N_10893);
xor U12026 (N_12026,N_10405,N_9883);
nor U12027 (N_12027,N_10105,N_10185);
nand U12028 (N_12028,N_10963,N_11990);
xor U12029 (N_12029,N_10910,N_10552);
xnor U12030 (N_12030,N_10374,N_11780);
nor U12031 (N_12031,N_9498,N_11794);
or U12032 (N_12032,N_11285,N_11725);
or U12033 (N_12033,N_11919,N_11030);
nor U12034 (N_12034,N_10992,N_9276);
and U12035 (N_12035,N_11953,N_9439);
and U12036 (N_12036,N_10629,N_10877);
and U12037 (N_12037,N_10356,N_9686);
nand U12038 (N_12038,N_10490,N_10297);
or U12039 (N_12039,N_10638,N_11202);
and U12040 (N_12040,N_11243,N_10290);
nand U12041 (N_12041,N_9318,N_9575);
xor U12042 (N_12042,N_11534,N_9270);
nor U12043 (N_12043,N_9077,N_10442);
nand U12044 (N_12044,N_10334,N_9974);
or U12045 (N_12045,N_10999,N_9005);
nand U12046 (N_12046,N_11356,N_9446);
or U12047 (N_12047,N_9622,N_10687);
or U12048 (N_12048,N_11536,N_9581);
nand U12049 (N_12049,N_10837,N_9539);
and U12050 (N_12050,N_11558,N_11726);
xnor U12051 (N_12051,N_11148,N_10924);
and U12052 (N_12052,N_9422,N_11906);
and U12053 (N_12053,N_11665,N_10930);
xnor U12054 (N_12054,N_10262,N_11598);
xnor U12055 (N_12055,N_11710,N_9537);
or U12056 (N_12056,N_9781,N_9436);
or U12057 (N_12057,N_9763,N_11487);
nand U12058 (N_12058,N_10065,N_9306);
nor U12059 (N_12059,N_11390,N_10039);
and U12060 (N_12060,N_10414,N_10090);
xnor U12061 (N_12061,N_9604,N_11562);
and U12062 (N_12062,N_9494,N_11181);
and U12063 (N_12063,N_10159,N_11644);
nor U12064 (N_12064,N_10941,N_9797);
or U12065 (N_12065,N_10288,N_9476);
and U12066 (N_12066,N_9521,N_11941);
or U12067 (N_12067,N_11137,N_11403);
and U12068 (N_12068,N_11958,N_9607);
and U12069 (N_12069,N_10219,N_10178);
nand U12070 (N_12070,N_10287,N_9734);
nor U12071 (N_12071,N_11631,N_9979);
nor U12072 (N_12072,N_9678,N_9061);
and U12073 (N_12073,N_11332,N_10212);
nand U12074 (N_12074,N_11311,N_10857);
and U12075 (N_12075,N_9050,N_9423);
nor U12076 (N_12076,N_9441,N_9742);
and U12077 (N_12077,N_9041,N_11180);
nor U12078 (N_12078,N_10098,N_10717);
nand U12079 (N_12079,N_9044,N_10804);
nand U12080 (N_12080,N_11295,N_9156);
nor U12081 (N_12081,N_10747,N_9552);
or U12082 (N_12082,N_9807,N_11380);
nor U12083 (N_12083,N_9813,N_11040);
nand U12084 (N_12084,N_10911,N_11081);
or U12085 (N_12085,N_9377,N_9698);
nor U12086 (N_12086,N_10619,N_11360);
or U12087 (N_12087,N_10677,N_9143);
nor U12088 (N_12088,N_10567,N_10753);
or U12089 (N_12089,N_9348,N_9546);
or U12090 (N_12090,N_10165,N_9594);
nand U12091 (N_12091,N_10095,N_10540);
nand U12092 (N_12092,N_10021,N_9310);
nand U12093 (N_12093,N_9060,N_11105);
or U12094 (N_12094,N_10038,N_9736);
nor U12095 (N_12095,N_10451,N_9032);
nor U12096 (N_12096,N_9187,N_11911);
nand U12097 (N_12097,N_10236,N_9589);
or U12098 (N_12098,N_11842,N_11150);
or U12099 (N_12099,N_9043,N_10816);
nor U12100 (N_12100,N_11834,N_9850);
nor U12101 (N_12101,N_10410,N_10495);
or U12102 (N_12102,N_10871,N_11581);
nand U12103 (N_12103,N_11944,N_10652);
and U12104 (N_12104,N_10951,N_11089);
or U12105 (N_12105,N_10624,N_11946);
nand U12106 (N_12106,N_11267,N_9179);
nor U12107 (N_12107,N_9654,N_9629);
nor U12108 (N_12108,N_10213,N_11957);
and U12109 (N_12109,N_10749,N_10461);
xor U12110 (N_12110,N_11277,N_9501);
nor U12111 (N_12111,N_10063,N_9645);
nand U12112 (N_12112,N_10264,N_9519);
or U12113 (N_12113,N_11022,N_11405);
nand U12114 (N_12114,N_11803,N_10000);
nand U12115 (N_12115,N_9320,N_9812);
and U12116 (N_12116,N_10788,N_11793);
nor U12117 (N_12117,N_11992,N_11658);
nor U12118 (N_12118,N_10667,N_10591);
nand U12119 (N_12119,N_9419,N_10062);
and U12120 (N_12120,N_10499,N_10534);
xnor U12121 (N_12121,N_11963,N_9258);
nand U12122 (N_12122,N_11977,N_9659);
nor U12123 (N_12123,N_10564,N_9479);
nor U12124 (N_12124,N_10579,N_9582);
and U12125 (N_12125,N_9769,N_11826);
and U12126 (N_12126,N_10504,N_11366);
or U12127 (N_12127,N_11373,N_9313);
nor U12128 (N_12128,N_10500,N_11686);
and U12129 (N_12129,N_9353,N_11535);
nor U12130 (N_12130,N_11668,N_9565);
and U12131 (N_12131,N_11350,N_11670);
xor U12132 (N_12132,N_10224,N_11024);
or U12133 (N_12133,N_11076,N_9252);
xnor U12134 (N_12134,N_11994,N_9725);
nand U12135 (N_12135,N_9766,N_11524);
nor U12136 (N_12136,N_10030,N_10437);
nor U12137 (N_12137,N_9121,N_9463);
or U12138 (N_12138,N_10277,N_9102);
nand U12139 (N_12139,N_9091,N_9819);
and U12140 (N_12140,N_11255,N_9155);
xnor U12141 (N_12141,N_11770,N_9100);
and U12142 (N_12142,N_9042,N_10370);
or U12143 (N_12143,N_9107,N_9406);
nand U12144 (N_12144,N_10813,N_9585);
and U12145 (N_12145,N_11003,N_9905);
and U12146 (N_12146,N_11531,N_10086);
or U12147 (N_12147,N_11626,N_9639);
nor U12148 (N_12148,N_10439,N_10465);
and U12149 (N_12149,N_10202,N_11979);
or U12150 (N_12150,N_10291,N_11584);
or U12151 (N_12151,N_11318,N_10382);
or U12152 (N_12152,N_10027,N_10254);
or U12153 (N_12153,N_11553,N_9198);
and U12154 (N_12154,N_9756,N_9347);
or U12155 (N_12155,N_10339,N_11334);
or U12156 (N_12156,N_11023,N_10338);
nor U12157 (N_12157,N_9677,N_10192);
or U12158 (N_12158,N_10328,N_11164);
or U12159 (N_12159,N_10840,N_10423);
or U12160 (N_12160,N_11763,N_11431);
and U12161 (N_12161,N_11655,N_10017);
nand U12162 (N_12162,N_10130,N_9976);
and U12163 (N_12163,N_11637,N_9990);
xnor U12164 (N_12164,N_10450,N_10831);
or U12165 (N_12165,N_9909,N_11322);
nor U12166 (N_12166,N_10389,N_10737);
and U12167 (N_12167,N_10241,N_10286);
or U12168 (N_12168,N_11005,N_9959);
xor U12169 (N_12169,N_10929,N_10161);
xor U12170 (N_12170,N_9307,N_11597);
or U12171 (N_12171,N_9130,N_11126);
and U12172 (N_12172,N_11094,N_10990);
xnor U12173 (N_12173,N_10913,N_10462);
nor U12174 (N_12174,N_9752,N_11661);
nand U12175 (N_12175,N_10974,N_10516);
nor U12176 (N_12176,N_10315,N_11629);
and U12177 (N_12177,N_11293,N_9690);
nand U12178 (N_12178,N_10734,N_10102);
and U12179 (N_12179,N_9437,N_9008);
nand U12180 (N_12180,N_11532,N_11479);
nand U12181 (N_12181,N_10836,N_9723);
xor U12182 (N_12182,N_11929,N_11666);
and U12183 (N_12183,N_10551,N_9177);
xnor U12184 (N_12184,N_11510,N_9997);
and U12185 (N_12185,N_11765,N_9169);
nor U12186 (N_12186,N_10467,N_11721);
nand U12187 (N_12187,N_10429,N_10659);
nor U12188 (N_12188,N_9346,N_11057);
nor U12189 (N_12189,N_10074,N_11874);
or U12190 (N_12190,N_9975,N_10613);
nand U12191 (N_12191,N_10509,N_9945);
and U12192 (N_12192,N_11732,N_10525);
or U12193 (N_12193,N_9058,N_10486);
or U12194 (N_12194,N_11972,N_9214);
or U12195 (N_12195,N_11846,N_11067);
and U12196 (N_12196,N_10321,N_11162);
or U12197 (N_12197,N_9683,N_11432);
xor U12198 (N_12198,N_11797,N_11653);
or U12199 (N_12199,N_10251,N_9830);
and U12200 (N_12200,N_10436,N_9737);
nor U12201 (N_12201,N_10255,N_11727);
nor U12202 (N_12202,N_10359,N_10520);
and U12203 (N_12203,N_10519,N_11887);
nand U12204 (N_12204,N_11901,N_11103);
xor U12205 (N_12205,N_11781,N_10890);
and U12206 (N_12206,N_11875,N_9915);
or U12207 (N_12207,N_9250,N_11753);
and U12208 (N_12208,N_10745,N_11000);
and U12209 (N_12209,N_10698,N_10563);
xnor U12210 (N_12210,N_10401,N_11805);
xnor U12211 (N_12211,N_9613,N_9577);
and U12212 (N_12212,N_11601,N_10764);
and U12213 (N_12213,N_9168,N_10846);
or U12214 (N_12214,N_9450,N_11983);
nor U12215 (N_12215,N_11169,N_10248);
nand U12216 (N_12216,N_11116,N_11577);
or U12217 (N_12217,N_10885,N_9136);
nand U12218 (N_12218,N_11493,N_9429);
nor U12219 (N_12219,N_10660,N_11809);
xor U12220 (N_12220,N_11075,N_9451);
nand U12221 (N_12221,N_9603,N_11595);
xnor U12222 (N_12222,N_11178,N_10744);
nor U12223 (N_12223,N_11592,N_11624);
nand U12224 (N_12224,N_9887,N_9308);
and U12225 (N_12225,N_11956,N_11888);
nor U12226 (N_12226,N_11071,N_10396);
and U12227 (N_12227,N_10601,N_10651);
or U12228 (N_12228,N_11298,N_10657);
nand U12229 (N_12229,N_11959,N_9006);
and U12230 (N_12230,N_10580,N_9878);
or U12231 (N_12231,N_11883,N_10977);
nand U12232 (N_12232,N_9610,N_11074);
or U12233 (N_12233,N_11968,N_11999);
xnor U12234 (N_12234,N_11671,N_9200);
or U12235 (N_12235,N_9785,N_10645);
nand U12236 (N_12236,N_10238,N_10766);
and U12237 (N_12237,N_9493,N_11530);
or U12238 (N_12238,N_10637,N_9188);
xor U12239 (N_12239,N_10526,N_11862);
or U12240 (N_12240,N_10748,N_10326);
xnor U12241 (N_12241,N_9069,N_10319);
or U12242 (N_12242,N_9359,N_9073);
nand U12243 (N_12243,N_10016,N_10197);
nand U12244 (N_12244,N_11918,N_10097);
or U12245 (N_12245,N_10539,N_11011);
nand U12246 (N_12246,N_9281,N_10047);
nand U12247 (N_12247,N_9949,N_9209);
nor U12248 (N_12248,N_10741,N_11242);
or U12249 (N_12249,N_11412,N_9832);
and U12250 (N_12250,N_11633,N_11903);
nand U12251 (N_12251,N_11033,N_10470);
and U12252 (N_12252,N_11096,N_11306);
nand U12253 (N_12253,N_10513,N_11750);
xnor U12254 (N_12254,N_9266,N_9162);
or U12255 (N_12255,N_10147,N_11095);
or U12256 (N_12256,N_9772,N_10609);
or U12257 (N_12257,N_10705,N_10997);
nand U12258 (N_12258,N_9167,N_10422);
nand U12259 (N_12259,N_9029,N_10289);
or U12260 (N_12260,N_9715,N_11772);
nand U12261 (N_12261,N_10092,N_9699);
and U12262 (N_12262,N_9477,N_11939);
nand U12263 (N_12263,N_11622,N_11467);
xnor U12264 (N_12264,N_9520,N_10426);
or U12265 (N_12265,N_10094,N_10046);
nor U12266 (N_12266,N_9146,N_10942);
and U12267 (N_12267,N_11490,N_10904);
nor U12268 (N_12268,N_9248,N_9025);
nor U12269 (N_12269,N_11927,N_10862);
or U12270 (N_12270,N_10909,N_11195);
or U12271 (N_12271,N_9074,N_11582);
or U12272 (N_12272,N_9696,N_11233);
xnor U12273 (N_12273,N_11864,N_11533);
nand U12274 (N_12274,N_10568,N_9732);
and U12275 (N_12275,N_10142,N_11786);
xor U12276 (N_12276,N_11821,N_11835);
or U12277 (N_12277,N_9040,N_10173);
or U12278 (N_12278,N_10103,N_11625);
nand U12279 (N_12279,N_11119,N_10154);
and U12280 (N_12280,N_11346,N_10253);
or U12281 (N_12281,N_10570,N_10785);
or U12282 (N_12282,N_11738,N_10765);
or U12283 (N_12283,N_9688,N_9910);
nor U12284 (N_12284,N_11440,N_11441);
nand U12285 (N_12285,N_11708,N_11287);
or U12286 (N_12286,N_10966,N_9083);
nor U12287 (N_12287,N_11494,N_11574);
nor U12288 (N_12288,N_10076,N_9516);
nor U12289 (N_12289,N_9870,N_11564);
nand U12290 (N_12290,N_9217,N_11509);
nor U12291 (N_12291,N_10633,N_9590);
nor U12292 (N_12292,N_11656,N_9784);
nand U12293 (N_12293,N_10919,N_9838);
or U12294 (N_12294,N_10282,N_11853);
nand U12295 (N_12295,N_11228,N_10618);
or U12296 (N_12296,N_11733,N_9658);
or U12297 (N_12297,N_9259,N_11792);
nor U12298 (N_12298,N_10614,N_10901);
nand U12299 (N_12299,N_9412,N_11021);
or U12300 (N_12300,N_9541,N_9300);
xnor U12301 (N_12301,N_10820,N_10949);
nand U12302 (N_12302,N_11799,N_11433);
or U12303 (N_12303,N_11612,N_9687);
and U12304 (N_12304,N_11940,N_9355);
nand U12305 (N_12305,N_11741,N_10456);
nor U12306 (N_12306,N_9434,N_11465);
nor U12307 (N_12307,N_11437,N_10441);
nor U12308 (N_12308,N_11385,N_11365);
nand U12309 (N_12309,N_9898,N_11871);
or U12310 (N_12310,N_9836,N_11302);
or U12311 (N_12311,N_10874,N_10345);
and U12312 (N_12312,N_9961,N_10398);
nor U12313 (N_12313,N_11652,N_9935);
and U12314 (N_12314,N_10166,N_10209);
or U12315 (N_12315,N_11965,N_9940);
nand U12316 (N_12316,N_9745,N_10043);
and U12317 (N_12317,N_11210,N_10797);
nor U12318 (N_12318,N_11908,N_11596);
or U12319 (N_12319,N_11559,N_10786);
xnor U12320 (N_12320,N_10313,N_11305);
or U12321 (N_12321,N_10243,N_9249);
nand U12322 (N_12322,N_9021,N_9183);
nand U12323 (N_12323,N_10767,N_9771);
and U12324 (N_12324,N_10543,N_10608);
or U12325 (N_12325,N_10453,N_9514);
and U12326 (N_12326,N_10109,N_9592);
nand U12327 (N_12327,N_9328,N_10220);
or U12328 (N_12328,N_11274,N_9007);
and U12329 (N_12329,N_11594,N_10952);
xnor U12330 (N_12330,N_10711,N_10029);
nand U12331 (N_12331,N_9694,N_11250);
nand U12332 (N_12332,N_11663,N_10231);
and U12333 (N_12333,N_11217,N_11639);
nor U12334 (N_12334,N_11042,N_11795);
nor U12335 (N_12335,N_11426,N_11702);
nand U12336 (N_12336,N_11331,N_11265);
or U12337 (N_12337,N_9731,N_11647);
nand U12338 (N_12338,N_9367,N_11225);
nor U12339 (N_12339,N_11616,N_9488);
nand U12340 (N_12340,N_10333,N_11697);
and U12341 (N_12341,N_10879,N_9420);
or U12342 (N_12342,N_11695,N_10079);
or U12343 (N_12343,N_9706,N_10239);
nand U12344 (N_12344,N_9216,N_9841);
and U12345 (N_12345,N_11141,N_11041);
nand U12346 (N_12346,N_9133,N_9324);
nor U12347 (N_12347,N_11495,N_9821);
nand U12348 (N_12348,N_11922,N_11989);
and U12349 (N_12349,N_11694,N_9504);
or U12350 (N_12350,N_10784,N_11514);
nor U12351 (N_12351,N_10245,N_10139);
nor U12352 (N_12352,N_10413,N_10800);
nor U12353 (N_12353,N_9265,N_11521);
and U12354 (N_12354,N_9657,N_11215);
xor U12355 (N_12355,N_10690,N_10607);
nand U12356 (N_12356,N_9794,N_10489);
and U12357 (N_12357,N_11900,N_9733);
and U12358 (N_12358,N_9978,N_9893);
and U12359 (N_12359,N_11478,N_11538);
xnor U12360 (N_12360,N_9971,N_9801);
or U12361 (N_12361,N_9424,N_9193);
nand U12362 (N_12362,N_10704,N_9457);
or U12363 (N_12363,N_11824,N_9055);
nand U12364 (N_12364,N_9633,N_11693);
or U12365 (N_12365,N_10894,N_11063);
nand U12366 (N_12366,N_11848,N_10632);
nand U12367 (N_12367,N_9376,N_9288);
nand U12368 (N_12368,N_9092,N_9160);
or U12369 (N_12369,N_10529,N_11272);
nor U12370 (N_12370,N_10428,N_10668);
xor U12371 (N_12371,N_10225,N_9815);
or U12372 (N_12372,N_9848,N_10216);
nor U12373 (N_12373,N_10179,N_9382);
xor U12374 (N_12374,N_9024,N_10556);
nor U12375 (N_12375,N_9888,N_9438);
nand U12376 (N_12376,N_10970,N_11610);
nand U12377 (N_12377,N_10042,N_11654);
and U12378 (N_12378,N_9793,N_11375);
nand U12379 (N_12379,N_9672,N_11086);
nor U12380 (N_12380,N_11312,N_11863);
and U12381 (N_12381,N_11251,N_11404);
nor U12382 (N_12382,N_10269,N_11966);
nor U12383 (N_12383,N_11731,N_9934);
or U12384 (N_12384,N_11383,N_11543);
nand U12385 (N_12385,N_9284,N_10560);
nor U12386 (N_12386,N_9663,N_11461);
and U12387 (N_12387,N_11909,N_11713);
nor U12388 (N_12388,N_11142,N_11129);
and U12389 (N_12389,N_9775,N_9876);
nand U12390 (N_12390,N_10627,N_10521);
nand U12391 (N_12391,N_11504,N_11314);
nor U12392 (N_12392,N_11491,N_11401);
nand U12393 (N_12393,N_9291,N_10073);
and U12394 (N_12394,N_11667,N_10488);
and U12395 (N_12395,N_9987,N_9808);
nor U12396 (N_12396,N_9621,N_10935);
nor U12397 (N_12397,N_11818,N_10869);
nor U12398 (N_12398,N_11008,N_10377);
and U12399 (N_12399,N_10380,N_10172);
or U12400 (N_12400,N_10409,N_11550);
nand U12401 (N_12401,N_10457,N_10517);
and U12402 (N_12402,N_11769,N_10841);
or U12403 (N_12403,N_9510,N_9523);
nor U12404 (N_12404,N_10325,N_10803);
and U12405 (N_12405,N_11266,N_9015);
nor U12406 (N_12406,N_11760,N_11097);
nand U12407 (N_12407,N_11851,N_10128);
nor U12408 (N_12408,N_10041,N_10246);
nand U12409 (N_12409,N_10561,N_11673);
or U12410 (N_12410,N_9037,N_11801);
or U12411 (N_12411,N_10850,N_10727);
nor U12412 (N_12412,N_9544,N_10975);
and U12413 (N_12413,N_11425,N_11035);
nor U12414 (N_12414,N_9835,N_9147);
nor U12415 (N_12415,N_9028,N_9947);
and U12416 (N_12416,N_9369,N_10485);
or U12417 (N_12417,N_10284,N_9472);
nand U12418 (N_12418,N_10308,N_9499);
and U12419 (N_12419,N_11855,N_9558);
or U12420 (N_12420,N_10505,N_11173);
and U12421 (N_12421,N_10615,N_11985);
nand U12422 (N_12422,N_9720,N_11269);
and U12423 (N_12423,N_9863,N_9803);
or U12424 (N_12424,N_11816,N_9986);
or U12425 (N_12425,N_11333,N_10671);
and U12426 (N_12426,N_10944,N_11893);
nand U12427 (N_12427,N_10684,N_9017);
and U12428 (N_12428,N_10124,N_9139);
or U12429 (N_12429,N_10536,N_9184);
nand U12430 (N_12430,N_10273,N_11349);
nand U12431 (N_12431,N_10839,N_10151);
nor U12432 (N_12432,N_9903,N_11472);
or U12433 (N_12433,N_9428,N_11613);
or U12434 (N_12434,N_11669,N_9128);
nor U12435 (N_12435,N_10337,N_9396);
and U12436 (N_12436,N_10912,N_11335);
nor U12437 (N_12437,N_11276,N_10385);
and U12438 (N_12438,N_11719,N_11800);
nor U12439 (N_12439,N_11471,N_10835);
or U12440 (N_12440,N_11297,N_10150);
nand U12441 (N_12441,N_9726,N_10427);
xor U12442 (N_12442,N_11028,N_9456);
and U12443 (N_12443,N_9398,N_11341);
or U12444 (N_12444,N_11205,N_10587);
nand U12445 (N_12445,N_11357,N_9220);
and U12446 (N_12446,N_10189,N_9236);
nand U12447 (N_12447,N_9082,N_9416);
or U12448 (N_12448,N_11705,N_9840);
or U12449 (N_12449,N_11323,N_11270);
nor U12450 (N_12450,N_10452,N_9665);
or U12451 (N_12451,N_9445,N_11427);
or U12452 (N_12452,N_11462,N_9115);
and U12453 (N_12453,N_9525,N_10025);
nand U12454 (N_12454,N_11006,N_10547);
xnor U12455 (N_12455,N_10654,N_10675);
nor U12456 (N_12456,N_10769,N_9616);
and U12457 (N_12457,N_9432,N_11703);
or U12458 (N_12458,N_11168,N_9556);
or U12459 (N_12459,N_11854,N_9648);
nor U12460 (N_12460,N_10542,N_10826);
or U12461 (N_12461,N_11976,N_10796);
xnor U12462 (N_12462,N_11359,N_11009);
nand U12463 (N_12463,N_11248,N_11604);
nand U12464 (N_12464,N_10293,N_10045);
and U12465 (N_12465,N_9517,N_11869);
xor U12466 (N_12466,N_9352,N_9913);
nor U12467 (N_12467,N_9485,N_11503);
xor U12468 (N_12468,N_9066,N_9929);
xor U12469 (N_12469,N_10257,N_11413);
and U12470 (N_12470,N_9591,N_11231);
or U12471 (N_12471,N_10593,N_9764);
nand U12472 (N_12472,N_10829,N_11327);
nand U12473 (N_12473,N_11811,N_10639);
xnor U12474 (N_12474,N_9453,N_11194);
and U12475 (N_12475,N_11676,N_9653);
nand U12476 (N_12476,N_10294,N_10887);
nand U12477 (N_12477,N_11832,N_9680);
or U12478 (N_12478,N_11961,N_11048);
and U12479 (N_12479,N_9148,N_9138);
nor U12480 (N_12480,N_9361,N_10384);
nand U12481 (N_12481,N_9194,N_9261);
nand U12482 (N_12482,N_9388,N_10415);
nand U12483 (N_12483,N_10058,N_9327);
nand U12484 (N_12484,N_9896,N_10362);
nand U12485 (N_12485,N_11515,N_9923);
nor U12486 (N_12486,N_10449,N_10342);
and U12487 (N_12487,N_9892,N_9461);
nor U12488 (N_12488,N_9708,N_10368);
nor U12489 (N_12489,N_11591,N_11570);
nor U12490 (N_12490,N_10702,N_9045);
nand U12491 (N_12491,N_10541,N_10795);
nor U12492 (N_12492,N_10152,N_10776);
nor U12493 (N_12493,N_10706,N_9031);
xor U12494 (N_12494,N_9564,N_11407);
nor U12495 (N_12495,N_11547,N_9914);
and U12496 (N_12496,N_10054,N_10920);
nand U12497 (N_12497,N_9334,N_9651);
nand U12498 (N_12498,N_11236,N_11207);
and U12499 (N_12499,N_11481,N_11696);
nor U12500 (N_12500,N_9968,N_11962);
and U12501 (N_12501,N_11500,N_10851);
and U12502 (N_12502,N_10242,N_9713);
or U12503 (N_12503,N_9917,N_10028);
nand U12504 (N_12504,N_10713,N_10487);
or U12505 (N_12505,N_10923,N_10898);
nand U12506 (N_12506,N_11160,N_10644);
nand U12507 (N_12507,N_9360,N_10164);
or U12508 (N_12508,N_11569,N_11756);
and U12509 (N_12509,N_9612,N_9695);
nor U12510 (N_12510,N_9538,N_9467);
or U12511 (N_12511,N_9027,N_11093);
and U12512 (N_12512,N_11975,N_9480);
nor U12513 (N_12513,N_10592,N_11127);
nor U12514 (N_12514,N_11072,N_11469);
and U12515 (N_12515,N_11920,N_9569);
nand U12516 (N_12516,N_11659,N_10739);
or U12517 (N_12517,N_9135,N_9458);
nor U12518 (N_12518,N_10096,N_10204);
nor U12519 (N_12519,N_9891,N_9491);
nor U12520 (N_12520,N_9164,N_9333);
nor U12521 (N_12521,N_10283,N_10181);
and U12522 (N_12522,N_9315,N_11599);
and U12523 (N_12523,N_10689,N_9440);
nor U12524 (N_12524,N_9608,N_11477);
and U12525 (N_12525,N_9003,N_11544);
nor U12526 (N_12526,N_9540,N_11970);
xor U12527 (N_12527,N_10718,N_9329);
nand U12528 (N_12528,N_11556,N_11294);
and U12529 (N_12529,N_9548,N_9536);
or U12530 (N_12530,N_11645,N_9191);
and U12531 (N_12531,N_10708,N_11566);
nand U12532 (N_12532,N_11018,N_11303);
or U12533 (N_12533,N_10678,N_10369);
nand U12534 (N_12534,N_9637,N_9972);
nor U12535 (N_12535,N_10686,N_9970);
or U12536 (N_12536,N_9111,N_10906);
nor U12537 (N_12537,N_9593,N_10817);
nand U12538 (N_12538,N_11384,N_11079);
and U12539 (N_12539,N_9056,N_10859);
nor U12540 (N_12540,N_9372,N_10824);
and U12541 (N_12541,N_11204,N_9402);
xnor U12542 (N_12542,N_11161,N_11059);
and U12543 (N_12543,N_10228,N_9567);
xnor U12544 (N_12544,N_10533,N_11641);
nor U12545 (N_12545,N_10845,N_10348);
nand U12546 (N_12546,N_11104,N_11165);
nand U12547 (N_12547,N_10674,N_11986);
and U12548 (N_12548,N_9760,N_10335);
or U12549 (N_12549,N_10169,N_11078);
and U12550 (N_12550,N_9062,N_10648);
or U12551 (N_12551,N_9255,N_11950);
or U12552 (N_12552,N_9068,N_9666);
nand U12553 (N_12553,N_11993,N_9381);
and U12554 (N_12554,N_11757,N_11775);
nor U12555 (N_12555,N_10562,N_10779);
nor U12556 (N_12556,N_11039,N_9798);
and U12557 (N_12557,N_11744,N_9795);
and U12558 (N_12558,N_9964,N_11034);
and U12559 (N_12559,N_10544,N_9175);
nor U12560 (N_12560,N_9181,N_11379);
nand U12561 (N_12561,N_9656,N_11418);
or U12562 (N_12562,N_9054,N_10976);
and U12563 (N_12563,N_10868,N_11381);
nor U12564 (N_12564,N_10656,N_9011);
and U12565 (N_12565,N_9993,N_10799);
nor U12566 (N_12566,N_9992,N_9205);
and U12567 (N_12567,N_9817,N_10565);
nand U12568 (N_12568,N_10832,N_11764);
and U12569 (N_12569,N_9816,N_10650);
nand U12570 (N_12570,N_11856,N_11117);
nand U12571 (N_12571,N_11395,N_10537);
and U12572 (N_12572,N_9150,N_11845);
nor U12573 (N_12573,N_11785,N_10066);
and U12574 (N_12574,N_10250,N_10889);
or U12575 (N_12575,N_10418,N_9251);
nor U12576 (N_12576,N_10088,N_11344);
nor U12577 (N_12577,N_9833,N_11729);
nor U12578 (N_12578,N_9356,N_9674);
and U12579 (N_12579,N_11084,N_9952);
and U12580 (N_12580,N_10936,N_10424);
or U12581 (N_12581,N_11038,N_10221);
nand U12582 (N_12582,N_11897,N_9967);
nor U12583 (N_12583,N_10407,N_10535);
and U12584 (N_12584,N_11788,N_10361);
nor U12585 (N_12585,N_9823,N_11674);
or U12586 (N_12586,N_10553,N_9197);
and U12587 (N_12587,N_11123,N_11371);
or U12588 (N_12588,N_9854,N_10602);
or U12589 (N_12589,N_9393,N_10945);
nand U12590 (N_12590,N_10483,N_9617);
nor U12591 (N_12591,N_10484,N_10760);
nor U12592 (N_12592,N_9026,N_9065);
xnor U12593 (N_12593,N_9554,N_9227);
nor U12594 (N_12594,N_10810,N_10372);
xor U12595 (N_12595,N_9553,N_9897);
nand U12596 (N_12596,N_11470,N_11054);
nand U12597 (N_12597,N_9998,N_11244);
or U12598 (N_12598,N_10214,N_10964);
or U12599 (N_12599,N_10137,N_11898);
xnor U12600 (N_12600,N_10494,N_11889);
nor U12601 (N_12601,N_10170,N_9285);
and U12602 (N_12602,N_9981,N_9820);
and U12603 (N_12603,N_11525,N_11640);
or U12604 (N_12604,N_11627,N_9627);
nand U12605 (N_12605,N_10672,N_10123);
nand U12606 (N_12606,N_10008,N_11787);
nor U12607 (N_12607,N_9882,N_10158);
nor U12608 (N_12608,N_10830,N_10538);
or U12609 (N_12609,N_11400,N_9405);
and U12610 (N_12610,N_9508,N_10307);
and U12611 (N_12611,N_11867,N_10444);
nand U12612 (N_12612,N_9740,N_11158);
nor U12613 (N_12613,N_10314,N_11108);
nand U12614 (N_12614,N_11421,N_10640);
or U12615 (N_12615,N_10420,N_10421);
xnor U12616 (N_12616,N_9322,N_9415);
or U12617 (N_12617,N_10261,N_10545);
or U12618 (N_12618,N_10881,N_9444);
or U12619 (N_12619,N_11839,N_9379);
xor U12620 (N_12620,N_9368,N_10458);
and U12621 (N_12621,N_9129,N_9606);
nor U12622 (N_12622,N_11124,N_9151);
or U12623 (N_12623,N_11010,N_10110);
nor U12624 (N_12624,N_11364,N_11709);
and U12625 (N_12625,N_11758,N_9743);
and U12626 (N_12626,N_10153,N_10233);
or U12627 (N_12627,N_10599,N_11203);
nand U12628 (N_12628,N_11125,N_11406);
and U12629 (N_12629,N_10798,N_10020);
or U12630 (N_12630,N_9459,N_11113);
nand U12631 (N_12631,N_9287,N_9547);
nor U12632 (N_12632,N_10709,N_10968);
nand U12633 (N_12633,N_11712,N_10448);
nand U12634 (N_12634,N_9944,N_9004);
nand U12635 (N_12635,N_11513,N_9649);
nand U12636 (N_12636,N_9773,N_9331);
xnor U12637 (N_12637,N_10510,N_11585);
nor U12638 (N_12638,N_10950,N_10106);
and U12639 (N_12639,N_9673,N_10834);
nor U12640 (N_12640,N_9623,N_10931);
xnor U12641 (N_12641,N_10358,N_10688);
nor U12642 (N_12642,N_10985,N_10603);
nand U12643 (N_12643,N_9710,N_11389);
or U12644 (N_12644,N_9067,N_10186);
or U12645 (N_12645,N_10725,N_10477);
and U12646 (N_12646,N_11955,N_10296);
or U12647 (N_12647,N_10168,N_10111);
or U12648 (N_12648,N_11254,N_9260);
nor U12649 (N_12649,N_10119,N_11838);
and U12650 (N_12650,N_9271,N_10378);
and U12651 (N_12651,N_11031,N_11062);
xnor U12652 (N_12652,N_11143,N_10203);
or U12653 (N_12653,N_9099,N_11352);
and U12654 (N_12654,N_11971,N_10928);
or U12655 (N_12655,N_11954,N_10967);
nand U12656 (N_12656,N_9345,N_9550);
nor U12657 (N_12657,N_10606,N_9371);
nor U12658 (N_12658,N_10497,N_10145);
and U12659 (N_12659,N_11420,N_11790);
nand U12660 (N_12660,N_11187,N_9362);
and U12661 (N_12661,N_11618,N_9526);
and U12662 (N_12662,N_10390,N_10127);
nand U12663 (N_12663,N_9304,N_10184);
or U12664 (N_12664,N_11445,N_11782);
nor U12665 (N_12665,N_9489,N_10626);
nand U12666 (N_12666,N_10699,N_11301);
and U12667 (N_12667,N_11147,N_9462);
nand U12668 (N_12668,N_9084,N_9875);
or U12669 (N_12669,N_10267,N_9806);
and U12670 (N_12670,N_11561,N_11759);
nand U12671 (N_12671,N_9165,N_9237);
xor U12672 (N_12672,N_10720,N_9305);
or U12673 (N_12673,N_9728,N_9118);
nand U12674 (N_12674,N_11910,N_11928);
or U12675 (N_12675,N_11414,N_9159);
or U12676 (N_12676,N_11565,N_10023);
xnor U12677 (N_12677,N_9988,N_11878);
nor U12678 (N_12678,N_9874,N_11523);
nand U12679 (N_12679,N_10381,N_11942);
and U12680 (N_12680,N_9410,N_10126);
xor U12681 (N_12681,N_10190,N_10515);
or U12682 (N_12682,N_11450,N_11263);
and U12683 (N_12683,N_11827,N_9879);
or U12684 (N_12684,N_11587,N_10682);
and U12685 (N_12685,N_9038,N_10195);
nand U12686 (N_12686,N_9262,N_9326);
or U12687 (N_12687,N_9966,N_11455);
xor U12688 (N_12688,N_9643,N_9779);
and U12689 (N_12689,N_10270,N_11716);
or U12690 (N_12690,N_10252,N_11932);
nand U12691 (N_12691,N_10496,N_11829);
nor U12692 (N_12692,N_10193,N_10347);
nand U12693 (N_12693,N_11498,N_10075);
and U12694 (N_12694,N_11519,N_11630);
or U12695 (N_12695,N_11367,N_10501);
or U12696 (N_12696,N_10351,N_9561);
and U12697 (N_12697,N_11091,N_11446);
nor U12698 (N_12698,N_11329,N_10061);
or U12699 (N_12699,N_10317,N_11088);
nor U12700 (N_12700,N_9886,N_10116);
nor U12701 (N_12701,N_9417,N_9400);
nand U12702 (N_12702,N_10812,N_10114);
nor U12703 (N_12703,N_9192,N_9991);
xnor U12704 (N_12704,N_9243,N_10726);
nand U12705 (N_12705,N_10162,N_9611);
and U12706 (N_12706,N_9586,N_9080);
nand U12707 (N_12707,N_11508,N_11984);
nor U12708 (N_12708,N_10980,N_10895);
or U12709 (N_12709,N_9994,N_11549);
nor U12710 (N_12710,N_11279,N_10693);
or U12711 (N_12711,N_9172,N_9873);
nor U12712 (N_12712,N_9847,N_9104);
or U12713 (N_12713,N_11229,N_9528);
nor U12714 (N_12714,N_9989,N_11988);
nor U12715 (N_12715,N_10336,N_11182);
nor U12716 (N_12716,N_9522,N_10956);
nand U12717 (N_12717,N_9861,N_9228);
nor U12718 (N_12718,N_10612,N_9578);
or U12719 (N_12719,N_11882,N_9053);
xor U12720 (N_12720,N_9566,N_9019);
nor U12721 (N_12721,N_11376,N_9524);
nand U12722 (N_12722,N_10777,N_11060);
or U12723 (N_12723,N_11372,N_11675);
and U12724 (N_12724,N_9842,N_10597);
or U12725 (N_12725,N_10454,N_11130);
and U12726 (N_12726,N_9238,N_10550);
nand U12727 (N_12727,N_10230,N_11745);
nand U12728 (N_12728,N_11967,N_9124);
and U12729 (N_12729,N_9933,N_9466);
nand U12730 (N_12730,N_10707,N_9682);
and U12731 (N_12731,N_11749,N_10084);
or U12732 (N_12732,N_10954,N_9557);
xnor U12733 (N_12733,N_9235,N_11083);
or U12734 (N_12734,N_10856,N_9922);
or U12735 (N_12735,N_11873,N_9885);
nand U12736 (N_12736,N_10438,N_10546);
and U12737 (N_12737,N_10780,N_10007);
nor U12738 (N_12738,N_9323,N_10012);
and U12739 (N_12739,N_11578,N_10425);
nand U12740 (N_12740,N_9230,N_9048);
xnor U12741 (N_12741,N_11434,N_10611);
nand U12742 (N_12742,N_9086,N_11345);
nor U12743 (N_12743,N_9512,N_11651);
and U12744 (N_12744,N_10735,N_10207);
and U12745 (N_12745,N_11628,N_10363);
nand U12746 (N_12746,N_10664,N_10666);
nor U12747 (N_12747,N_10987,N_10838);
nand U12748 (N_12748,N_11860,N_9219);
or U12749 (N_12749,N_10762,N_9101);
nand U12750 (N_12750,N_10392,N_11890);
or U12751 (N_12751,N_9685,N_9857);
and U12752 (N_12752,N_11227,N_10053);
or U12753 (N_12753,N_10048,N_9022);
or U12754 (N_12754,N_11843,N_11649);
xnor U12755 (N_12755,N_11737,N_11885);
nand U12756 (N_12756,N_9487,N_10117);
xor U12757 (N_12757,N_9717,N_10808);
xnor U12758 (N_12758,N_9675,N_11134);
and U12759 (N_12759,N_11691,N_10921);
nand U12760 (N_12760,N_9154,N_10443);
or U12761 (N_12761,N_11767,N_9096);
xnor U12762 (N_12762,N_9560,N_9384);
nand U12763 (N_12763,N_9085,N_9009);
nor U12764 (N_12764,N_10476,N_9856);
xnor U12765 (N_12765,N_10790,N_9822);
or U12766 (N_12766,N_9814,N_10625);
and U12767 (N_12767,N_11522,N_9263);
and U12768 (N_12768,N_9969,N_11796);
or U12769 (N_12769,N_10210,N_10249);
xnor U12770 (N_12770,N_10121,N_11982);
xor U12771 (N_12771,N_10433,N_9668);
and U12772 (N_12772,N_10044,N_11771);
nor U12773 (N_12773,N_9030,N_10300);
or U12774 (N_12774,N_11912,N_10171);
nor U12775 (N_12775,N_10115,N_11672);
xor U12776 (N_12776,N_10527,N_9454);
and U12777 (N_12777,N_11238,N_10412);
xor U12778 (N_12778,N_10996,N_10916);
and U12779 (N_12779,N_10040,N_11398);
nand U12780 (N_12780,N_10514,N_11936);
nand U12781 (N_12781,N_10814,N_11343);
xor U12782 (N_12782,N_9244,N_10771);
and U12783 (N_12783,N_11754,N_9701);
nor U12784 (N_12784,N_9709,N_10104);
nand U12785 (N_12785,N_9364,N_11393);
or U12786 (N_12786,N_10572,N_11783);
and U12787 (N_12787,N_10080,N_11145);
xnor U12788 (N_12788,N_9342,N_10825);
or U12789 (N_12789,N_10549,N_9290);
xor U12790 (N_12790,N_11964,N_9587);
and U12791 (N_12791,N_11361,N_11449);
and U12792 (N_12792,N_9254,N_10716);
nor U12793 (N_12793,N_9751,N_10235);
and U12794 (N_12794,N_9584,N_11736);
nand U12795 (N_12795,N_9302,N_11685);
nor U12796 (N_12796,N_11226,N_11723);
nor U12797 (N_12797,N_10595,N_11486);
xor U12798 (N_12798,N_9088,N_10331);
nand U12799 (N_12799,N_10994,N_11870);
nand U12800 (N_12800,N_10002,N_11099);
and U12801 (N_12801,N_9965,N_11100);
nor U12802 (N_12802,N_9864,N_9576);
nand U12803 (N_12803,N_9427,N_11580);
nand U12804 (N_12804,N_11224,N_11053);
and U12805 (N_12805,N_9618,N_9921);
or U12806 (N_12806,N_11257,N_9996);
nor U12807 (N_12807,N_11724,N_9225);
or U12808 (N_12808,N_10227,N_11002);
nor U12809 (N_12809,N_10959,N_9170);
and U12810 (N_12810,N_9932,N_9033);
and U12811 (N_12811,N_10683,N_10022);
or U12812 (N_12812,N_11635,N_9596);
or U12813 (N_12813,N_10460,N_10320);
and U12814 (N_12814,N_9010,N_11220);
nand U12815 (N_12815,N_11015,N_11157);
and U12816 (N_12816,N_11386,N_11552);
and U12817 (N_12817,N_10060,N_11810);
or U12818 (N_12818,N_10491,N_11489);
nand U12819 (N_12819,N_10344,N_9478);
nand U12820 (N_12820,N_9474,N_11830);
or U12821 (N_12821,N_10807,N_11717);
nand U12822 (N_12822,N_10805,N_10569);
or U12823 (N_12823,N_11463,N_11529);
nand U12824 (N_12824,N_9273,N_9714);
or U12825 (N_12825,N_10276,N_11139);
nand U12826 (N_12826,N_11234,N_11678);
and U12827 (N_12827,N_10217,N_9020);
nand U12828 (N_12828,N_11699,N_10847);
xnor U12829 (N_12829,N_10311,N_11948);
or U12830 (N_12830,N_11149,N_10631);
nor U12831 (N_12831,N_11052,N_11735);
xor U12832 (N_12832,N_11907,N_10112);
nand U12833 (N_12833,N_11027,N_11825);
xnor U12834 (N_12834,N_9113,N_10182);
nor U12835 (N_12835,N_9580,N_11505);
and U12836 (N_12836,N_10201,N_9319);
xnor U12837 (N_12837,N_10304,N_9064);
or U12838 (N_12838,N_11369,N_11634);
or U12839 (N_12839,N_11218,N_9796);
or U12840 (N_12840,N_10056,N_9224);
nand U12841 (N_12841,N_9365,N_10622);
or U12842 (N_12842,N_9647,N_9014);
or U12843 (N_12843,N_10724,N_11442);
or U12844 (N_12844,N_10663,N_9106);
nand U12845 (N_12845,N_9839,N_10258);
and U12846 (N_12846,N_11353,N_11714);
xnor U12847 (N_12847,N_9366,N_9518);
nand U12848 (N_12848,N_9335,N_11568);
nor U12849 (N_12849,N_11016,N_9747);
and U12850 (N_12850,N_10729,N_9641);
xnor U12851 (N_12851,N_9872,N_10107);
nor U12852 (N_12852,N_9486,N_11282);
or U12853 (N_12853,N_9503,N_11092);
xnor U12854 (N_12854,N_11391,N_9919);
or U12855 (N_12855,N_11252,N_9283);
or U12856 (N_12856,N_11328,N_10346);
nor U12857 (N_12857,N_11876,N_11156);
or U12858 (N_12858,N_10432,N_9693);
or U12859 (N_12859,N_10474,N_9780);
nand U12860 (N_12860,N_10176,N_10003);
or U12861 (N_12861,N_10167,N_10327);
and U12862 (N_12862,N_9317,N_11159);
or U12863 (N_12863,N_10554,N_10399);
nand U12864 (N_12864,N_11551,N_11278);
and U12865 (N_12865,N_9865,N_9631);
nor U12866 (N_12866,N_10581,N_11363);
nor U12867 (N_12867,N_9223,N_10240);
xnor U12868 (N_12868,N_9729,N_11087);
xor U12869 (N_12869,N_11309,N_10770);
nor U12870 (N_12870,N_9942,N_10867);
xnor U12871 (N_12871,N_9442,N_9013);
xor U12872 (N_12872,N_9280,N_10915);
nor U12873 (N_12873,N_11175,N_9430);
nand U12874 (N_12874,N_10818,N_10349);
nand U12875 (N_12875,N_11572,N_10087);
nand U12876 (N_12876,N_9811,N_11935);
or U12877 (N_12877,N_9846,N_10440);
or U12878 (N_12878,N_10466,N_11183);
nand U12879 (N_12879,N_10598,N_9605);
or U12880 (N_12880,N_9351,N_11777);
and U12881 (N_12881,N_11354,N_11043);
or U12882 (N_12882,N_9206,N_10531);
nor U12883 (N_12883,N_10828,N_9094);
nor U12884 (N_12884,N_9394,N_11424);
or U12885 (N_12885,N_11602,N_10278);
xnor U12886 (N_12886,N_10059,N_11485);
and U12887 (N_12887,N_11337,N_10089);
or U12888 (N_12888,N_9303,N_9039);
and U12889 (N_12889,N_10469,N_10940);
nor U12890 (N_12890,N_9983,N_11430);
or U12891 (N_12891,N_9471,N_11600);
and U12892 (N_12892,N_10594,N_10661);
nand U12893 (N_12893,N_10658,N_11290);
xnor U12894 (N_12894,N_9707,N_10018);
nor U12895 (N_12895,N_10670,N_10026);
nand U12896 (N_12896,N_10719,N_10984);
and U12897 (N_12897,N_10324,N_10833);
or U12898 (N_12898,N_10903,N_10965);
and U12899 (N_12899,N_11457,N_10108);
nor U12900 (N_12900,N_10013,N_9203);
nand U12901 (N_12901,N_10280,N_11483);
and U12902 (N_12902,N_10120,N_10113);
nand U12903 (N_12903,N_10610,N_10134);
xnor U12904 (N_12904,N_11497,N_11762);
xnor U12905 (N_12905,N_9447,N_9999);
and U12906 (N_12906,N_9925,N_9904);
and U12907 (N_12907,N_10600,N_9598);
or U12908 (N_12908,N_11214,N_11017);
nand U12909 (N_12909,N_11120,N_9232);
nand U12910 (N_12910,N_10681,N_11768);
or U12911 (N_12911,N_11240,N_9936);
and U12912 (N_12912,N_10035,N_9824);
or U12913 (N_12913,N_10256,N_10653);
nand U12914 (N_12914,N_9655,N_10353);
nand U12915 (N_12915,N_10306,N_11073);
or U12916 (N_12916,N_9818,N_11662);
xor U12917 (N_12917,N_9800,N_10532);
and U12918 (N_12918,N_11969,N_11815);
nand U12919 (N_12919,N_11296,N_11978);
nor U12920 (N_12920,N_11259,N_11448);
or U12921 (N_12921,N_11914,N_9931);
and U12922 (N_12922,N_10793,N_10417);
nand U12923 (N_12923,N_9375,N_11734);
nand U12924 (N_12924,N_10730,N_9390);
nand U12925 (N_12925,N_9035,N_11155);
nor U12926 (N_12926,N_9274,N_10360);
nand U12927 (N_12927,N_9385,N_9109);
nand U12928 (N_12928,N_10498,N_11114);
nand U12929 (N_12929,N_10001,N_10703);
and U12930 (N_12930,N_10875,N_11007);
or U12931 (N_12931,N_9063,N_11742);
nand U12932 (N_12932,N_11368,N_10691);
or U12933 (N_12933,N_11539,N_11981);
and U12934 (N_12934,N_9851,N_9153);
nor U12935 (N_12935,N_9515,N_11351);
xor U12936 (N_12936,N_9505,N_9047);
or U12937 (N_12937,N_9373,N_10732);
and U12938 (N_12938,N_9973,N_11032);
xor U12939 (N_12939,N_11219,N_9543);
nor U12940 (N_12940,N_10900,N_9902);
or U12941 (N_12941,N_11198,N_9609);
or U12942 (N_12942,N_11286,N_11995);
and U12943 (N_12943,N_10806,N_10843);
nor U12944 (N_12944,N_10435,N_11289);
nand U12945 (N_12945,N_11643,N_10628);
or U12946 (N_12946,N_11288,N_10100);
nor U12947 (N_12947,N_10459,N_11836);
nand U12948 (N_12948,N_9778,N_11447);
nand U12949 (N_12949,N_11444,N_11325);
or U12950 (N_12950,N_11915,N_10330);
or U12951 (N_12951,N_11814,N_10792);
or U12952 (N_12952,N_10072,N_11739);
or U12953 (N_12953,N_10863,N_11886);
nor U12954 (N_12954,N_11743,N_9906);
nand U12955 (N_12955,N_9826,N_9204);
nand U12956 (N_12956,N_9744,N_11239);
and U12957 (N_12957,N_10772,N_11338);
nor U12958 (N_12958,N_9679,N_10229);
and U12959 (N_12959,N_11892,N_11066);
or U12960 (N_12960,N_9549,N_9571);
nand U12961 (N_12961,N_10131,N_9739);
xnor U12962 (N_12962,N_10036,N_10281);
or U12963 (N_12963,N_9212,N_10902);
or U12964 (N_12964,N_10783,N_11304);
nand U12965 (N_12965,N_9977,N_9413);
nand U12966 (N_12966,N_11140,N_11453);
or U12967 (N_12967,N_9804,N_10375);
nor U12968 (N_12968,N_9511,N_11466);
or U12969 (N_12969,N_10391,N_10093);
and U12970 (N_12970,N_10218,N_9404);
nand U12971 (N_12971,N_10962,N_10758);
nor U12972 (N_12972,N_9233,N_11609);
or U12973 (N_12973,N_11423,N_11849);
or U12974 (N_12974,N_11520,N_11607);
and U12975 (N_12975,N_10298,N_11947);
nor U12976 (N_12976,N_10259,N_10917);
xnor U12977 (N_12977,N_9691,N_11684);
or U12978 (N_12978,N_11689,N_9776);
xnor U12979 (N_12979,N_10548,N_10492);
nor U12980 (N_12980,N_9619,N_10584);
or U12981 (N_12981,N_9635,N_10292);
nor U12982 (N_12982,N_11563,N_11933);
and U12983 (N_12983,N_9001,N_11949);
or U12984 (N_12984,N_9958,N_11324);
or U12985 (N_12985,N_11049,N_11593);
or U12986 (N_12986,N_9754,N_11952);
nand U12987 (N_12987,N_11546,N_10157);
or U12988 (N_12988,N_11879,N_10480);
nor U12989 (N_12989,N_10604,N_10789);
nand U12990 (N_12990,N_10854,N_9642);
and U12991 (N_12991,N_9809,N_10721);
or U12992 (N_12992,N_11813,N_11480);
or U12993 (N_12993,N_9357,N_11300);
nor U12994 (N_12994,N_9229,N_10665);
or U12995 (N_12995,N_10866,N_11991);
nor U12996 (N_12996,N_11025,N_10223);
or U12997 (N_12997,N_10187,N_9116);
nand U12998 (N_12998,N_9786,N_11082);
nand U12999 (N_12999,N_10888,N_11330);
xor U13000 (N_13000,N_9052,N_11388);
or U13001 (N_13001,N_11026,N_11464);
nor U13002 (N_13002,N_11050,N_11747);
nor U13003 (N_13003,N_11711,N_10332);
or U13004 (N_13004,N_9002,N_11492);
nand U13005 (N_13005,N_11571,N_10620);
or U13006 (N_13006,N_10135,N_11188);
nor U13007 (N_13007,N_11456,N_9496);
or U13008 (N_13008,N_10781,N_11623);
nor U13009 (N_13009,N_11896,N_10049);
or U13010 (N_13010,N_10998,N_9535);
nor U13011 (N_13011,N_9858,N_11488);
and U13012 (N_13012,N_9173,N_9127);
and U13013 (N_13013,N_11190,N_11683);
nand U13014 (N_13014,N_10010,N_10194);
and U13015 (N_13015,N_9341,N_11789);
and U13016 (N_13016,N_10873,N_9464);
or U13017 (N_13017,N_11237,N_10148);
nor U13018 (N_13018,N_10605,N_11784);
nand U13019 (N_13019,N_11291,N_9721);
nand U13020 (N_13020,N_9120,N_11077);
nor U13021 (N_13021,N_10132,N_9337);
nor U13022 (N_13022,N_10180,N_10673);
nor U13023 (N_13023,N_11567,N_9727);
nand U13024 (N_13024,N_10271,N_11590);
and U13025 (N_13025,N_9299,N_11321);
and U13026 (N_13026,N_11642,N_11807);
nand U13027 (N_13027,N_11315,N_10578);
nor U13028 (N_13028,N_9583,N_10695);
or U13029 (N_13029,N_9090,N_9401);
and U13030 (N_13030,N_9336,N_11131);
or U13031 (N_13031,N_10582,N_9788);
and U13032 (N_13032,N_9196,N_10005);
or U13033 (N_13033,N_10014,N_11545);
nor U13034 (N_13034,N_11603,N_9470);
or U13035 (N_13035,N_10588,N_9071);
and U13036 (N_13036,N_11191,N_9201);
nand U13037 (N_13037,N_9171,N_11185);
nand U13038 (N_13038,N_11037,N_9370);
and U13039 (N_13039,N_11923,N_9669);
nand U13040 (N_13040,N_9634,N_11013);
or U13041 (N_13041,N_11650,N_11452);
nand U13042 (N_13042,N_11755,N_10508);
nor U13043 (N_13043,N_10728,N_11362);
nor U13044 (N_13044,N_11812,N_10430);
xnor U13045 (N_13045,N_11715,N_11307);
and U13046 (N_13046,N_9628,N_11101);
and U13047 (N_13047,N_10479,N_10811);
nor U13048 (N_13048,N_10947,N_9414);
nand U13049 (N_13049,N_10925,N_11045);
and U13050 (N_13050,N_9142,N_10590);
or U13051 (N_13051,N_9805,N_11722);
xnor U13052 (N_13052,N_9908,N_11506);
xnor U13053 (N_13053,N_10263,N_10434);
nor U13054 (N_13054,N_11458,N_10309);
or U13055 (N_13055,N_9383,N_9036);
xor U13056 (N_13056,N_10692,N_11292);
nor U13057 (N_13057,N_9108,N_9810);
nor U13058 (N_13058,N_9757,N_10511);
nand U13059 (N_13059,N_10208,N_11436);
xor U13060 (N_13060,N_9295,N_11213);
nor U13061 (N_13061,N_9443,N_11540);
and U13062 (N_13062,N_10756,N_10024);
or U13063 (N_13063,N_9703,N_11937);
nor U13064 (N_13064,N_9343,N_9911);
nand U13065 (N_13065,N_11258,N_11443);
and U13066 (N_13066,N_10404,N_9078);
nor U13067 (N_13067,N_11336,N_10299);
nor U13068 (N_13068,N_11859,N_10616);
nand U13069 (N_13069,N_10696,N_10200);
nand U13070 (N_13070,N_11701,N_10848);
nand U13071 (N_13071,N_10322,N_9389);
and U13072 (N_13072,N_9330,N_11537);
nor U13073 (N_13073,N_10400,N_10183);
and U13074 (N_13074,N_11313,N_10402);
and U13075 (N_13075,N_9208,N_9684);
nand U13076 (N_13076,N_11894,N_11319);
nor U13077 (N_13077,N_10773,N_10493);
or U13078 (N_13078,N_9182,N_10891);
nand U13079 (N_13079,N_11271,N_9316);
nand U13080 (N_13080,N_9292,N_11107);
and U13081 (N_13081,N_10419,N_11679);
and U13082 (N_13082,N_10589,N_11858);
nand U13083 (N_13083,N_9765,N_9529);
nor U13084 (N_13084,N_9378,N_10234);
nor U13085 (N_13085,N_9755,N_9534);
and U13086 (N_13086,N_11283,N_10823);
and U13087 (N_13087,N_11707,N_9221);
nand U13088 (N_13088,N_9681,N_11144);
or U13089 (N_13089,N_9490,N_10763);
nor U13090 (N_13090,N_9123,N_10312);
and U13091 (N_13091,N_10472,N_10642);
nor U13092 (N_13092,N_11429,N_9871);
or U13093 (N_13093,N_10641,N_9241);
nand U13094 (N_13094,N_10722,N_10006);
and U13095 (N_13095,N_11261,N_10355);
nand U13096 (N_13096,N_9825,N_9293);
nand U13097 (N_13097,N_11512,N_10055);
and U13098 (N_13098,N_10155,N_10031);
or U13099 (N_13099,N_10892,N_11268);
nor U13100 (N_13100,N_10067,N_11284);
nor U13101 (N_13101,N_10226,N_10714);
nor U13102 (N_13102,N_11638,N_9664);
or U13103 (N_13103,N_10350,N_10196);
nor U13104 (N_13104,N_10101,N_9980);
nand U13105 (N_13105,N_10366,N_10815);
nand U13106 (N_13106,N_10723,N_9312);
nand U13107 (N_13107,N_9387,N_9358);
or U13108 (N_13108,N_11098,N_11435);
or U13109 (N_13109,N_10011,N_10746);
xnor U13110 (N_13110,N_10849,N_10731);
or U13111 (N_13111,N_11588,N_11808);
xor U13112 (N_13112,N_11192,N_9395);
nand U13113 (N_13113,N_9245,N_9239);
nor U13114 (N_13114,N_11047,N_10393);
and U13115 (N_13115,N_9105,N_10091);
nor U13116 (N_13116,N_10755,N_11473);
nand U13117 (N_13117,N_9777,N_9866);
and U13118 (N_13118,N_9636,N_9023);
nand U13119 (N_13119,N_9601,N_9652);
and U13120 (N_13120,N_9495,N_11193);
and U13121 (N_13121,N_10528,N_11516);
xor U13122 (N_13122,N_10884,N_9718);
nor U13123 (N_13123,N_9397,N_10634);
nand U13124 (N_13124,N_9533,N_9849);
or U13125 (N_13125,N_9845,N_11899);
nor U13126 (N_13126,N_11014,N_9555);
or U13127 (N_13127,N_10742,N_9761);
and U13128 (N_13128,N_11833,N_9667);
or U13129 (N_13129,N_10932,N_11904);
nand U13130 (N_13130,N_9630,N_10522);
or U13131 (N_13131,N_9513,N_9112);
and U13132 (N_13132,N_10323,N_9110);
nor U13133 (N_13133,N_9268,N_11692);
or U13134 (N_13134,N_10759,N_9632);
or U13135 (N_13135,N_10099,N_9889);
nand U13136 (N_13136,N_9380,N_11245);
xor U13137 (N_13137,N_9995,N_10305);
nand U13138 (N_13138,N_10934,N_9114);
nand U13139 (N_13139,N_11394,N_10395);
nand U13140 (N_13140,N_9711,N_11138);
xor U13141 (N_13141,N_10129,N_9530);
or U13142 (N_13142,N_10386,N_10222);
nand U13143 (N_13143,N_10078,N_9719);
nor U13144 (N_13144,N_11664,N_11945);
or U13145 (N_13145,N_9448,N_11135);
and U13146 (N_13146,N_11370,N_10174);
or U13147 (N_13147,N_10575,N_9894);
and U13148 (N_13148,N_10512,N_9075);
and U13149 (N_13149,N_11377,N_10523);
or U13150 (N_13150,N_10852,N_10318);
and U13151 (N_13151,N_10953,N_10743);
and U13152 (N_13152,N_10791,N_10635);
nand U13153 (N_13153,N_9660,N_11122);
nor U13154 (N_13154,N_9057,N_11857);
nand U13155 (N_13155,N_9912,N_11766);
and U13156 (N_13156,N_10478,N_10371);
nor U13157 (N_13157,N_11340,N_9145);
or U13158 (N_13158,N_11065,N_10978);
or U13159 (N_13159,N_9527,N_10530);
and U13160 (N_13160,N_11819,N_10948);
and U13161 (N_13161,N_11115,N_9240);
nand U13162 (N_13162,N_11614,N_10680);
nor U13163 (N_13163,N_11817,N_11249);
xnor U13164 (N_13164,N_10993,N_9507);
xor U13165 (N_13165,N_11044,N_9122);
or U13166 (N_13166,N_11058,N_11378);
nor U13167 (N_13167,N_10071,N_9614);
and U13168 (N_13168,N_11779,N_10070);
xor U13169 (N_13169,N_11275,N_11176);
or U13170 (N_13170,N_9483,N_11555);
and U13171 (N_13171,N_9532,N_9626);
nand U13172 (N_13172,N_10899,N_11166);
nor U13173 (N_13173,N_9750,N_10146);
nor U13174 (N_13174,N_10958,N_11230);
or U13175 (N_13175,N_9469,N_10357);
nor U13176 (N_13176,N_10118,N_11924);
nor U13177 (N_13177,N_10914,N_9829);
nand U13178 (N_13178,N_11617,N_10922);
nand U13179 (N_13179,N_11146,N_9880);
nor U13180 (N_13180,N_11677,N_10468);
nand U13181 (N_13181,N_9234,N_9768);
and U13182 (N_13182,N_9748,N_9218);
or U13183 (N_13183,N_10032,N_10503);
and U13184 (N_13184,N_9076,N_11374);
and U13185 (N_13185,N_9103,N_9789);
or U13186 (N_13186,N_10387,N_11055);
or U13187 (N_13187,N_10585,N_11527);
nand U13188 (N_13188,N_11451,N_11704);
xnor U13189 (N_13189,N_9753,N_9724);
nor U13190 (N_13190,N_10655,N_10274);
nor U13191 (N_13191,N_11730,N_10822);
nor U13192 (N_13192,N_11051,N_9275);
xor U13193 (N_13193,N_10870,N_11850);
and U13194 (N_13194,N_10373,N_11273);
or U13195 (N_13195,N_10937,N_9702);
and U13196 (N_13196,N_10761,N_11861);
xor U13197 (N_13197,N_9431,N_9853);
nand U13198 (N_13198,N_10285,N_9770);
or U13199 (N_13199,N_10938,N_9730);
and U13200 (N_13200,N_10265,N_9267);
nor U13201 (N_13201,N_11751,N_11606);
or U13202 (N_13202,N_9374,N_9783);
nor U13203 (N_13203,N_11902,N_9860);
nand U13204 (N_13204,N_10566,N_9141);
or U13205 (N_13205,N_10232,N_10768);
or U13206 (N_13206,N_9449,N_11209);
and U13207 (N_13207,N_9704,N_10617);
nor U13208 (N_13208,N_11660,N_9195);
nor U13209 (N_13209,N_11554,N_11128);
and U13210 (N_13210,N_11688,N_10821);
nor U13211 (N_13211,N_9481,N_11748);
nor U13212 (N_13212,N_11152,N_9468);
nor U13213 (N_13213,N_11980,N_10394);
nand U13214 (N_13214,N_9620,N_9862);
and U13215 (N_13215,N_11877,N_11526);
or U13216 (N_13216,N_9790,N_11012);
nor U13217 (N_13217,N_11706,N_9297);
or U13218 (N_13218,N_10676,N_11197);
nor U13219 (N_13219,N_10473,N_10211);
nor U13220 (N_13220,N_10447,N_9354);
or U13221 (N_13221,N_10464,N_11262);
nor U13222 (N_13222,N_10295,N_9542);
or U13223 (N_13223,N_11925,N_9098);
nand U13224 (N_13224,N_11186,N_10774);
nand U13225 (N_13225,N_9213,N_9562);
or U13226 (N_13226,N_9956,N_9256);
nand U13227 (N_13227,N_9963,N_9588);
nand U13228 (N_13228,N_11348,N_11264);
nand U13229 (N_13229,N_10329,N_10844);
nor U13230 (N_13230,N_9350,N_9937);
or U13231 (N_13231,N_9943,N_10083);
or U13232 (N_13232,N_9399,N_9403);
nand U13233 (N_13233,N_9081,N_10268);
xor U13234 (N_13234,N_11646,N_9900);
nand U13235 (N_13235,N_9962,N_9137);
or U13236 (N_13236,N_9072,N_11199);
nand U13237 (N_13237,N_10571,N_10802);
or U13238 (N_13238,N_10482,N_10897);
and U13239 (N_13239,N_9689,N_11880);
or U13240 (N_13240,N_9855,N_9916);
and U13241 (N_13241,N_9939,N_10787);
xnor U13242 (N_13242,N_11496,N_9152);
and U13243 (N_13243,N_10206,N_11905);
nor U13244 (N_13244,N_11998,N_9957);
or U13245 (N_13245,N_10260,N_11507);
nor U13246 (N_13246,N_9190,N_11528);
xnor U13247 (N_13247,N_9920,N_10019);
or U13248 (N_13248,N_10475,N_11090);
nand U13249 (N_13249,N_9638,N_10961);
xor U13250 (N_13250,N_11837,N_11036);
nor U13251 (N_13251,N_10876,N_10927);
or U13252 (N_13252,N_10406,N_11387);
or U13253 (N_13253,N_9435,N_10160);
or U13254 (N_13254,N_9492,N_11930);
xor U13255 (N_13255,N_9012,N_11872);
nor U13256 (N_13256,N_9722,N_9572);
xor U13257 (N_13257,N_10955,N_9573);
nand U13258 (N_13258,N_10643,N_9314);
nor U13259 (N_13259,N_10972,N_10446);
nand U13260 (N_13260,N_11560,N_10908);
or U13261 (N_13261,N_9834,N_9095);
nor U13262 (N_13262,N_10986,N_9231);
and U13263 (N_13263,N_11221,N_9749);
or U13264 (N_13264,N_9189,N_11133);
or U13265 (N_13265,N_9126,N_10596);
and U13266 (N_13266,N_10237,N_11281);
and U13267 (N_13267,N_10455,N_11987);
or U13268 (N_13268,N_11397,N_10272);
and U13269 (N_13269,N_11247,N_11605);
or U13270 (N_13270,N_10215,N_9202);
or U13271 (N_13271,N_11868,N_9409);
nor U13272 (N_13272,N_11476,N_11317);
and U13273 (N_13273,N_11844,N_11069);
nor U13274 (N_13274,N_9662,N_10883);
or U13275 (N_13275,N_9954,N_9500);
or U13276 (N_13276,N_10081,N_10191);
nand U13277 (N_13277,N_9895,N_11621);
nor U13278 (N_13278,N_11822,N_11206);
nand U13279 (N_13279,N_11153,N_9930);
or U13280 (N_13280,N_10577,N_11798);
and U13281 (N_13281,N_9046,N_9746);
and U13282 (N_13282,N_10057,N_11154);
nor U13283 (N_13283,N_10037,N_9735);
nand U13284 (N_13284,N_11163,N_9570);
nor U13285 (N_13285,N_10905,N_11070);
or U13286 (N_13286,N_11151,N_11382);
or U13287 (N_13287,N_9286,N_10700);
nor U13288 (N_13288,N_10507,N_9363);
nor U13289 (N_13289,N_10583,N_10649);
nor U13290 (N_13290,N_11973,N_9938);
nand U13291 (N_13291,N_10069,N_10809);
nand U13292 (N_13292,N_10983,N_11774);
nor U13293 (N_13293,N_9282,N_11761);
nand U13294 (N_13294,N_9670,N_10367);
xor U13295 (N_13295,N_9671,N_10751);
xnor U13296 (N_13296,N_9163,N_9296);
or U13297 (N_13297,N_11347,N_11974);
nand U13298 (N_13298,N_11619,N_9349);
or U13299 (N_13299,N_9161,N_9982);
nand U13300 (N_13300,N_9950,N_9000);
and U13301 (N_13301,N_10034,N_9433);
nor U13302 (N_13302,N_9391,N_9759);
nand U13303 (N_13303,N_10198,N_10969);
or U13304 (N_13304,N_10156,N_11773);
xor U13305 (N_13305,N_9199,N_10316);
or U13306 (N_13306,N_10697,N_9767);
nand U13307 (N_13307,N_9985,N_10801);
nand U13308 (N_13308,N_9852,N_10082);
and U13309 (N_13309,N_9421,N_11439);
and U13310 (N_13310,N_10205,N_9411);
nor U13311 (N_13311,N_11454,N_9144);
nor U13312 (N_13312,N_10085,N_10685);
xor U13313 (N_13313,N_9597,N_9738);
and U13314 (N_13314,N_10842,N_9386);
or U13315 (N_13315,N_10310,N_10064);
nand U13316 (N_13316,N_10341,N_10973);
and U13317 (N_13317,N_11831,N_10140);
and U13318 (N_13318,N_11611,N_11399);
or U13319 (N_13319,N_11934,N_9831);
and U13320 (N_13320,N_9140,N_11310);
or U13321 (N_13321,N_9877,N_9332);
and U13322 (N_13322,N_11019,N_9859);
or U13323 (N_13323,N_9185,N_11841);
nand U13324 (N_13324,N_11579,N_10524);
and U13325 (N_13325,N_11746,N_11200);
xnor U13326 (N_13326,N_10679,N_11482);
and U13327 (N_13327,N_10188,N_9301);
or U13328 (N_13328,N_11517,N_10506);
nor U13329 (N_13329,N_9311,N_10855);
and U13330 (N_13330,N_9955,N_9890);
and U13331 (N_13331,N_10009,N_9899);
or U13332 (N_13332,N_9774,N_11778);
nor U13333 (N_13333,N_9615,N_11419);
or U13334 (N_13334,N_9079,N_10960);
or U13335 (N_13335,N_9253,N_11246);
nor U13336 (N_13336,N_9712,N_11802);
nor U13337 (N_13337,N_10431,N_11001);
nand U13338 (N_13338,N_9568,N_9269);
or U13339 (N_13339,N_9644,N_9309);
xnor U13340 (N_13340,N_11943,N_11068);
and U13341 (N_13341,N_11396,N_11109);
nand U13342 (N_13342,N_9325,N_11996);
or U13343 (N_13343,N_10175,N_11687);
nor U13344 (N_13344,N_11170,N_9180);
nand U13345 (N_13345,N_9791,N_9506);
nand U13346 (N_13346,N_9222,N_11575);
nor U13347 (N_13347,N_11320,N_11326);
nor U13348 (N_13348,N_9131,N_10279);
nor U13349 (N_13349,N_9640,N_9884);
and U13350 (N_13350,N_11589,N_10558);
nor U13351 (N_13351,N_10051,N_10136);
and U13352 (N_13352,N_11913,N_9579);
and U13353 (N_13353,N_10865,N_9869);
or U13354 (N_13354,N_10244,N_9624);
xnor U13355 (N_13355,N_9563,N_9758);
or U13356 (N_13356,N_10995,N_11657);
and U13357 (N_13357,N_10882,N_10004);
xnor U13358 (N_13358,N_9953,N_10015);
or U13359 (N_13359,N_10853,N_11132);
nor U13360 (N_13360,N_10858,N_9828);
nand U13361 (N_13361,N_10199,N_9787);
nand U13362 (N_13362,N_10247,N_11459);
xor U13363 (N_13363,N_9827,N_11339);
xor U13364 (N_13364,N_9697,N_11997);
nand U13365 (N_13365,N_9016,N_10861);
and U13366 (N_13366,N_9157,N_10141);
nand U13367 (N_13367,N_10982,N_10177);
nand U13368 (N_13368,N_10991,N_9595);
or U13369 (N_13369,N_11501,N_11064);
and U13370 (N_13370,N_10750,N_10077);
nand U13371 (N_13371,N_11029,N_11061);
or U13372 (N_13372,N_10957,N_9802);
or U13373 (N_13373,N_10463,N_9125);
nor U13374 (N_13374,N_11791,N_9277);
nand U13375 (N_13375,N_10939,N_10586);
or U13376 (N_13376,N_9279,N_10989);
or U13377 (N_13377,N_11402,N_11583);
nand U13378 (N_13378,N_9928,N_11417);
xnor U13379 (N_13379,N_11342,N_9425);
and U13380 (N_13380,N_10445,N_9465);
and U13381 (N_13381,N_11256,N_11410);
or U13382 (N_13382,N_11960,N_10576);
and U13383 (N_13383,N_11866,N_11615);
or U13384 (N_13384,N_10481,N_10471);
nand U13385 (N_13385,N_11891,N_9901);
nand U13386 (N_13386,N_10778,N_11428);
or U13387 (N_13387,N_11184,N_9051);
nor U13388 (N_13388,N_11299,N_11499);
nor U13389 (N_13389,N_9545,N_9338);
xnor U13390 (N_13390,N_9340,N_11167);
and U13391 (N_13391,N_11408,N_9676);
nor U13392 (N_13392,N_10712,N_10647);
nor U13393 (N_13393,N_11004,N_11682);
and U13394 (N_13394,N_9867,N_11212);
nand U13395 (N_13395,N_9926,N_10408);
nor U13396 (N_13396,N_9093,N_10864);
nand U13397 (N_13397,N_10403,N_11232);
or U13398 (N_13398,N_9924,N_10918);
nor U13399 (N_13399,N_9497,N_10352);
or U13400 (N_13400,N_10979,N_11216);
and U13401 (N_13401,N_9186,N_10574);
or U13402 (N_13402,N_11241,N_9272);
nand U13403 (N_13403,N_9984,N_10933);
and U13404 (N_13404,N_11484,N_10878);
nand U13405 (N_13405,N_9149,N_10662);
xnor U13406 (N_13406,N_11518,N_11938);
nand U13407 (N_13407,N_9215,N_9907);
or U13408 (N_13408,N_9392,N_11355);
nor U13409 (N_13409,N_11576,N_9034);
and U13410 (N_13410,N_9344,N_9531);
or U13411 (N_13411,N_10518,N_11253);
or U13412 (N_13412,N_10926,N_9837);
and U13413 (N_13413,N_11172,N_11823);
nor U13414 (N_13414,N_11112,N_11415);
nor U13415 (N_13415,N_11852,N_10827);
or U13416 (N_13416,N_11820,N_11921);
nor U13417 (N_13417,N_9257,N_11409);
nand U13418 (N_13418,N_10794,N_9646);
nand U13419 (N_13419,N_9600,N_11917);
xnor U13420 (N_13420,N_10416,N_9158);
nand U13421 (N_13421,N_10819,N_11931);
and U13422 (N_13422,N_11740,N_11804);
nand U13423 (N_13423,N_11502,N_9087);
nor U13424 (N_13424,N_10757,N_11828);
nor U13425 (N_13425,N_11106,N_10740);
or U13426 (N_13426,N_9941,N_9407);
nor U13427 (N_13427,N_9484,N_10125);
nand U13428 (N_13428,N_11460,N_10133);
nor U13429 (N_13429,N_10860,N_11468);
nand U13430 (N_13430,N_9716,N_11847);
xnor U13431 (N_13431,N_9059,N_11895);
or U13432 (N_13432,N_9741,N_11085);
or U13433 (N_13433,N_9210,N_9602);
nand U13434 (N_13434,N_9018,N_9089);
nand U13435 (N_13435,N_11308,N_9599);
nor U13436 (N_13436,N_10033,N_10872);
or U13437 (N_13437,N_10701,N_11121);
and U13438 (N_13438,N_9176,N_9339);
or U13439 (N_13439,N_11951,N_9134);
and U13440 (N_13440,N_10630,N_10733);
nand U13441 (N_13441,N_10052,N_9625);
or U13442 (N_13442,N_9574,N_9705);
and U13443 (N_13443,N_9951,N_9408);
nor U13444 (N_13444,N_10775,N_10303);
or U13445 (N_13445,N_9551,N_10149);
or U13446 (N_13446,N_9844,N_11720);
nor U13447 (N_13447,N_10782,N_10981);
or U13448 (N_13448,N_9502,N_9070);
or U13449 (N_13449,N_9278,N_10354);
and U13450 (N_13450,N_9927,N_11700);
nor U13451 (N_13451,N_9482,N_11728);
nor U13452 (N_13452,N_10636,N_10573);
nor U13453 (N_13453,N_11177,N_10694);
and U13454 (N_13454,N_10880,N_9294);
nand U13455 (N_13455,N_10896,N_9247);
or U13456 (N_13456,N_11189,N_10738);
or U13457 (N_13457,N_10302,N_9211);
nor U13458 (N_13458,N_11174,N_9452);
nor U13459 (N_13459,N_11235,N_11548);
nand U13460 (N_13460,N_9843,N_10946);
nor U13461 (N_13461,N_9207,N_9473);
or U13462 (N_13462,N_11411,N_11865);
nor U13463 (N_13463,N_11916,N_9264);
nor U13464 (N_13464,N_9242,N_11316);
nor U13465 (N_13465,N_10143,N_9946);
nor U13466 (N_13466,N_11208,N_10907);
nand U13467 (N_13467,N_11196,N_9509);
and U13468 (N_13468,N_10988,N_11056);
nand U13469 (N_13469,N_9174,N_11201);
and U13470 (N_13470,N_9321,N_9881);
nand U13471 (N_13471,N_10971,N_10397);
nand U13472 (N_13472,N_9782,N_9650);
nor U13473 (N_13473,N_11680,N_11541);
or U13474 (N_13474,N_11884,N_10411);
nor U13475 (N_13475,N_11752,N_11118);
nor U13476 (N_13476,N_11211,N_10621);
xor U13477 (N_13477,N_9097,N_9918);
nand U13478 (N_13478,N_9475,N_9049);
nand U13479 (N_13479,N_9226,N_10623);
or U13480 (N_13480,N_11511,N_11416);
nor U13481 (N_13481,N_9762,N_10669);
nor U13482 (N_13482,N_9426,N_9700);
nand U13483 (N_13483,N_10163,N_11422);
and U13484 (N_13484,N_11573,N_10736);
and U13485 (N_13485,N_10122,N_10555);
nand U13486 (N_13486,N_10301,N_9868);
or U13487 (N_13487,N_11632,N_11690);
nor U13488 (N_13488,N_11136,N_11542);
and U13489 (N_13489,N_9418,N_11046);
nand U13490 (N_13490,N_9117,N_11648);
or U13491 (N_13491,N_10943,N_11608);
or U13492 (N_13492,N_11681,N_10559);
nor U13493 (N_13493,N_10715,N_11636);
and U13494 (N_13494,N_11102,N_10754);
nand U13495 (N_13495,N_10379,N_10502);
nor U13496 (N_13496,N_10376,N_11474);
nor U13497 (N_13497,N_11557,N_9559);
nor U13498 (N_13498,N_11620,N_11171);
and U13499 (N_13499,N_11806,N_10388);
nand U13500 (N_13500,N_11538,N_11000);
nor U13501 (N_13501,N_11375,N_11927);
or U13502 (N_13502,N_11514,N_11259);
xor U13503 (N_13503,N_11452,N_9062);
xnor U13504 (N_13504,N_11505,N_9337);
or U13505 (N_13505,N_9508,N_10843);
xnor U13506 (N_13506,N_10545,N_10933);
nand U13507 (N_13507,N_11836,N_10440);
xnor U13508 (N_13508,N_11122,N_11175);
nand U13509 (N_13509,N_11200,N_9888);
nand U13510 (N_13510,N_10904,N_11709);
nand U13511 (N_13511,N_10636,N_10537);
and U13512 (N_13512,N_9653,N_9936);
nand U13513 (N_13513,N_9554,N_10189);
nor U13514 (N_13514,N_10357,N_11946);
or U13515 (N_13515,N_10243,N_9837);
nor U13516 (N_13516,N_11675,N_10814);
or U13517 (N_13517,N_11682,N_10133);
nor U13518 (N_13518,N_10065,N_11796);
nand U13519 (N_13519,N_9035,N_9631);
nand U13520 (N_13520,N_9218,N_11580);
and U13521 (N_13521,N_9039,N_11672);
or U13522 (N_13522,N_10239,N_11697);
nand U13523 (N_13523,N_11988,N_11567);
xnor U13524 (N_13524,N_9362,N_11736);
or U13525 (N_13525,N_11387,N_9190);
nand U13526 (N_13526,N_11343,N_10825);
or U13527 (N_13527,N_10359,N_9306);
xor U13528 (N_13528,N_9224,N_9800);
and U13529 (N_13529,N_10714,N_11203);
nor U13530 (N_13530,N_11238,N_11133);
nor U13531 (N_13531,N_11687,N_10794);
nor U13532 (N_13532,N_9414,N_10309);
nand U13533 (N_13533,N_11721,N_9993);
and U13534 (N_13534,N_9959,N_11812);
or U13535 (N_13535,N_11075,N_11686);
or U13536 (N_13536,N_9117,N_11306);
and U13537 (N_13537,N_9402,N_11599);
nand U13538 (N_13538,N_11210,N_10855);
and U13539 (N_13539,N_11275,N_10072);
nand U13540 (N_13540,N_9852,N_9887);
or U13541 (N_13541,N_9512,N_9045);
or U13542 (N_13542,N_10222,N_10326);
xor U13543 (N_13543,N_9295,N_9330);
nand U13544 (N_13544,N_10437,N_10094);
nand U13545 (N_13545,N_11373,N_10668);
nand U13546 (N_13546,N_11685,N_10586);
nor U13547 (N_13547,N_9390,N_10653);
nand U13548 (N_13548,N_10075,N_9667);
nor U13549 (N_13549,N_10083,N_9504);
nor U13550 (N_13550,N_9202,N_11269);
nor U13551 (N_13551,N_9701,N_11865);
nand U13552 (N_13552,N_11526,N_11312);
nor U13553 (N_13553,N_11322,N_11558);
or U13554 (N_13554,N_11443,N_10090);
nor U13555 (N_13555,N_9891,N_10054);
and U13556 (N_13556,N_11740,N_11578);
nand U13557 (N_13557,N_10231,N_9975);
and U13558 (N_13558,N_11957,N_9964);
or U13559 (N_13559,N_9315,N_9368);
nand U13560 (N_13560,N_11621,N_11148);
or U13561 (N_13561,N_10766,N_10546);
nand U13562 (N_13562,N_9093,N_11816);
nand U13563 (N_13563,N_11977,N_11986);
and U13564 (N_13564,N_9051,N_10863);
nor U13565 (N_13565,N_11165,N_11044);
and U13566 (N_13566,N_10497,N_10643);
nor U13567 (N_13567,N_11743,N_9530);
nand U13568 (N_13568,N_10757,N_9329);
nor U13569 (N_13569,N_9807,N_9712);
or U13570 (N_13570,N_10954,N_9338);
or U13571 (N_13571,N_11435,N_9258);
nand U13572 (N_13572,N_9504,N_10338);
nand U13573 (N_13573,N_10713,N_9025);
nand U13574 (N_13574,N_10918,N_11395);
nor U13575 (N_13575,N_11461,N_11016);
nor U13576 (N_13576,N_9723,N_11442);
xnor U13577 (N_13577,N_9878,N_11729);
and U13578 (N_13578,N_10416,N_11360);
nor U13579 (N_13579,N_9360,N_9291);
xnor U13580 (N_13580,N_9262,N_9876);
nand U13581 (N_13581,N_10033,N_11533);
and U13582 (N_13582,N_9437,N_9060);
and U13583 (N_13583,N_11337,N_11978);
nor U13584 (N_13584,N_9619,N_11037);
nand U13585 (N_13585,N_11850,N_10121);
and U13586 (N_13586,N_9616,N_10920);
xnor U13587 (N_13587,N_9513,N_10370);
xnor U13588 (N_13588,N_10111,N_10828);
nor U13589 (N_13589,N_10165,N_10642);
and U13590 (N_13590,N_9004,N_9672);
nor U13591 (N_13591,N_11709,N_10431);
nand U13592 (N_13592,N_9879,N_9435);
or U13593 (N_13593,N_10536,N_9083);
and U13594 (N_13594,N_10306,N_11424);
nand U13595 (N_13595,N_9433,N_9102);
nand U13596 (N_13596,N_10948,N_9051);
nor U13597 (N_13597,N_11512,N_10121);
nand U13598 (N_13598,N_11284,N_9675);
nor U13599 (N_13599,N_9250,N_10242);
nand U13600 (N_13600,N_9466,N_11943);
xor U13601 (N_13601,N_11058,N_9332);
and U13602 (N_13602,N_9189,N_9166);
nor U13603 (N_13603,N_9667,N_11151);
or U13604 (N_13604,N_10477,N_9480);
nand U13605 (N_13605,N_10715,N_10950);
nand U13606 (N_13606,N_9493,N_11650);
xnor U13607 (N_13607,N_10176,N_11525);
nor U13608 (N_13608,N_11130,N_9991);
and U13609 (N_13609,N_9785,N_9638);
or U13610 (N_13610,N_9991,N_9755);
xor U13611 (N_13611,N_9103,N_11536);
xnor U13612 (N_13612,N_9352,N_11656);
and U13613 (N_13613,N_9458,N_11147);
or U13614 (N_13614,N_9328,N_11709);
nand U13615 (N_13615,N_9210,N_10192);
or U13616 (N_13616,N_11705,N_10004);
or U13617 (N_13617,N_11673,N_10178);
xor U13618 (N_13618,N_9474,N_11287);
or U13619 (N_13619,N_10412,N_11040);
or U13620 (N_13620,N_10370,N_10636);
or U13621 (N_13621,N_10485,N_9285);
nor U13622 (N_13622,N_11585,N_10175);
or U13623 (N_13623,N_10948,N_11684);
or U13624 (N_13624,N_10812,N_9806);
or U13625 (N_13625,N_10157,N_11467);
nor U13626 (N_13626,N_9788,N_10233);
or U13627 (N_13627,N_10509,N_10278);
or U13628 (N_13628,N_9968,N_11278);
or U13629 (N_13629,N_10102,N_10625);
or U13630 (N_13630,N_9121,N_9367);
or U13631 (N_13631,N_11432,N_11712);
or U13632 (N_13632,N_11708,N_11227);
and U13633 (N_13633,N_11076,N_9959);
xor U13634 (N_13634,N_10181,N_10974);
nor U13635 (N_13635,N_10392,N_11707);
nand U13636 (N_13636,N_9081,N_10258);
nand U13637 (N_13637,N_9066,N_10157);
nand U13638 (N_13638,N_9447,N_9132);
and U13639 (N_13639,N_11984,N_10664);
and U13640 (N_13640,N_9144,N_9913);
or U13641 (N_13641,N_9155,N_11880);
xor U13642 (N_13642,N_11924,N_10892);
and U13643 (N_13643,N_9410,N_10438);
and U13644 (N_13644,N_11627,N_10596);
nand U13645 (N_13645,N_9836,N_11135);
and U13646 (N_13646,N_10875,N_11472);
xor U13647 (N_13647,N_10309,N_11609);
nand U13648 (N_13648,N_11116,N_9415);
and U13649 (N_13649,N_9582,N_9007);
or U13650 (N_13650,N_9947,N_9479);
nand U13651 (N_13651,N_10502,N_10566);
or U13652 (N_13652,N_11652,N_10979);
and U13653 (N_13653,N_10604,N_10717);
nand U13654 (N_13654,N_11199,N_10067);
nor U13655 (N_13655,N_10891,N_9802);
nor U13656 (N_13656,N_10386,N_11378);
nor U13657 (N_13657,N_11655,N_9074);
or U13658 (N_13658,N_10902,N_10851);
nor U13659 (N_13659,N_10252,N_10723);
or U13660 (N_13660,N_9480,N_9378);
and U13661 (N_13661,N_11327,N_10260);
nor U13662 (N_13662,N_11705,N_9647);
nor U13663 (N_13663,N_10876,N_9085);
nand U13664 (N_13664,N_11545,N_11205);
or U13665 (N_13665,N_9249,N_10413);
and U13666 (N_13666,N_9735,N_10576);
nor U13667 (N_13667,N_9691,N_10269);
or U13668 (N_13668,N_9640,N_9492);
nor U13669 (N_13669,N_10453,N_10441);
and U13670 (N_13670,N_10028,N_10384);
and U13671 (N_13671,N_11299,N_11111);
nor U13672 (N_13672,N_10124,N_10110);
nor U13673 (N_13673,N_11252,N_9656);
and U13674 (N_13674,N_11533,N_10211);
or U13675 (N_13675,N_11711,N_10047);
nor U13676 (N_13676,N_11346,N_10451);
nor U13677 (N_13677,N_9787,N_11840);
or U13678 (N_13678,N_11337,N_9111);
and U13679 (N_13679,N_11046,N_10537);
xnor U13680 (N_13680,N_11052,N_9443);
nand U13681 (N_13681,N_11585,N_10377);
or U13682 (N_13682,N_11262,N_9581);
xor U13683 (N_13683,N_10778,N_11504);
and U13684 (N_13684,N_10798,N_9379);
nand U13685 (N_13685,N_9935,N_9652);
nor U13686 (N_13686,N_9219,N_11667);
and U13687 (N_13687,N_11048,N_9676);
nor U13688 (N_13688,N_10816,N_9329);
and U13689 (N_13689,N_11660,N_11806);
or U13690 (N_13690,N_9683,N_9744);
nand U13691 (N_13691,N_11676,N_9681);
nor U13692 (N_13692,N_9140,N_10178);
or U13693 (N_13693,N_10688,N_10793);
nand U13694 (N_13694,N_10757,N_9647);
nand U13695 (N_13695,N_9609,N_11104);
or U13696 (N_13696,N_10889,N_11575);
nor U13697 (N_13697,N_10824,N_9751);
or U13698 (N_13698,N_9434,N_10882);
or U13699 (N_13699,N_10245,N_11687);
nand U13700 (N_13700,N_9547,N_11682);
or U13701 (N_13701,N_10474,N_11079);
and U13702 (N_13702,N_9302,N_10738);
and U13703 (N_13703,N_10910,N_11369);
nand U13704 (N_13704,N_11872,N_10357);
or U13705 (N_13705,N_10229,N_9513);
nor U13706 (N_13706,N_9533,N_9247);
nor U13707 (N_13707,N_10225,N_9486);
xnor U13708 (N_13708,N_9129,N_10664);
nor U13709 (N_13709,N_11666,N_9827);
or U13710 (N_13710,N_10393,N_11446);
or U13711 (N_13711,N_11041,N_9496);
and U13712 (N_13712,N_11931,N_11024);
and U13713 (N_13713,N_11301,N_9106);
or U13714 (N_13714,N_11832,N_11934);
and U13715 (N_13715,N_9805,N_11843);
nand U13716 (N_13716,N_9921,N_11897);
and U13717 (N_13717,N_11627,N_9970);
nor U13718 (N_13718,N_11509,N_11169);
nor U13719 (N_13719,N_9933,N_11159);
xnor U13720 (N_13720,N_11064,N_10787);
and U13721 (N_13721,N_9592,N_11797);
nand U13722 (N_13722,N_11123,N_9688);
or U13723 (N_13723,N_9787,N_10863);
nor U13724 (N_13724,N_10018,N_10966);
nor U13725 (N_13725,N_10299,N_11649);
and U13726 (N_13726,N_9081,N_10662);
or U13727 (N_13727,N_11244,N_9980);
or U13728 (N_13728,N_10193,N_10586);
nor U13729 (N_13729,N_9722,N_10336);
or U13730 (N_13730,N_11010,N_10623);
or U13731 (N_13731,N_11880,N_9013);
nand U13732 (N_13732,N_11728,N_9637);
nor U13733 (N_13733,N_10404,N_10933);
xor U13734 (N_13734,N_11215,N_9099);
nor U13735 (N_13735,N_11818,N_9955);
or U13736 (N_13736,N_11123,N_11979);
nor U13737 (N_13737,N_9674,N_11563);
nand U13738 (N_13738,N_11147,N_9282);
nor U13739 (N_13739,N_11859,N_10291);
xor U13740 (N_13740,N_11598,N_11080);
and U13741 (N_13741,N_11545,N_10403);
and U13742 (N_13742,N_11910,N_9991);
nand U13743 (N_13743,N_9995,N_9117);
nand U13744 (N_13744,N_11119,N_11488);
nor U13745 (N_13745,N_10304,N_9129);
nand U13746 (N_13746,N_10529,N_11391);
xor U13747 (N_13747,N_9446,N_10418);
nand U13748 (N_13748,N_10230,N_11265);
nand U13749 (N_13749,N_11981,N_9254);
nand U13750 (N_13750,N_10640,N_11967);
nor U13751 (N_13751,N_10760,N_10883);
or U13752 (N_13752,N_11834,N_10685);
xnor U13753 (N_13753,N_9756,N_9974);
nand U13754 (N_13754,N_10894,N_11165);
nand U13755 (N_13755,N_10144,N_10908);
and U13756 (N_13756,N_10811,N_11760);
or U13757 (N_13757,N_11001,N_11118);
nand U13758 (N_13758,N_9901,N_10223);
and U13759 (N_13759,N_10361,N_11850);
nand U13760 (N_13760,N_11550,N_10222);
xor U13761 (N_13761,N_11566,N_11840);
and U13762 (N_13762,N_11752,N_9889);
nand U13763 (N_13763,N_10626,N_10086);
nand U13764 (N_13764,N_11198,N_10942);
or U13765 (N_13765,N_11973,N_10563);
nand U13766 (N_13766,N_11123,N_11750);
or U13767 (N_13767,N_9168,N_10031);
xor U13768 (N_13768,N_10201,N_9371);
and U13769 (N_13769,N_11845,N_9811);
or U13770 (N_13770,N_10909,N_10284);
nand U13771 (N_13771,N_10188,N_11751);
and U13772 (N_13772,N_10729,N_9878);
nand U13773 (N_13773,N_9091,N_11540);
nor U13774 (N_13774,N_9158,N_10373);
or U13775 (N_13775,N_11163,N_11898);
nand U13776 (N_13776,N_10324,N_10095);
or U13777 (N_13777,N_10912,N_10624);
nand U13778 (N_13778,N_9086,N_10337);
and U13779 (N_13779,N_10371,N_9809);
nor U13780 (N_13780,N_10343,N_10638);
or U13781 (N_13781,N_11165,N_9551);
nor U13782 (N_13782,N_10789,N_9439);
or U13783 (N_13783,N_9860,N_11787);
nand U13784 (N_13784,N_10311,N_10462);
or U13785 (N_13785,N_9390,N_9067);
nand U13786 (N_13786,N_10644,N_10825);
or U13787 (N_13787,N_9479,N_11985);
and U13788 (N_13788,N_9119,N_11563);
nand U13789 (N_13789,N_9138,N_11258);
and U13790 (N_13790,N_9576,N_10571);
nor U13791 (N_13791,N_9757,N_9038);
or U13792 (N_13792,N_10289,N_11357);
or U13793 (N_13793,N_10695,N_9592);
nor U13794 (N_13794,N_11102,N_10207);
nor U13795 (N_13795,N_11140,N_9316);
nand U13796 (N_13796,N_11964,N_11111);
and U13797 (N_13797,N_10077,N_10179);
xor U13798 (N_13798,N_9232,N_11868);
nor U13799 (N_13799,N_9802,N_11169);
or U13800 (N_13800,N_10132,N_11306);
nor U13801 (N_13801,N_11485,N_10984);
nor U13802 (N_13802,N_11413,N_9542);
or U13803 (N_13803,N_9379,N_10822);
or U13804 (N_13804,N_10046,N_10431);
and U13805 (N_13805,N_9449,N_10869);
xor U13806 (N_13806,N_11721,N_9309);
and U13807 (N_13807,N_11052,N_11497);
nor U13808 (N_13808,N_10356,N_9711);
or U13809 (N_13809,N_11228,N_9750);
and U13810 (N_13810,N_11026,N_10351);
nor U13811 (N_13811,N_11194,N_9654);
nor U13812 (N_13812,N_10601,N_9916);
and U13813 (N_13813,N_9751,N_11909);
nand U13814 (N_13814,N_9635,N_10228);
nand U13815 (N_13815,N_11299,N_9058);
and U13816 (N_13816,N_9188,N_11748);
and U13817 (N_13817,N_10316,N_11268);
and U13818 (N_13818,N_11446,N_9395);
or U13819 (N_13819,N_9189,N_11304);
nand U13820 (N_13820,N_11581,N_10898);
nor U13821 (N_13821,N_9415,N_9790);
and U13822 (N_13822,N_9847,N_9705);
nand U13823 (N_13823,N_10685,N_10275);
and U13824 (N_13824,N_9912,N_9979);
or U13825 (N_13825,N_9319,N_11396);
nand U13826 (N_13826,N_11931,N_9947);
and U13827 (N_13827,N_10275,N_11441);
nor U13828 (N_13828,N_9851,N_11650);
nand U13829 (N_13829,N_11684,N_10902);
nor U13830 (N_13830,N_9316,N_11189);
nor U13831 (N_13831,N_9977,N_11171);
nand U13832 (N_13832,N_10430,N_10680);
nor U13833 (N_13833,N_9717,N_10992);
xor U13834 (N_13834,N_9736,N_9410);
and U13835 (N_13835,N_11937,N_9037);
nor U13836 (N_13836,N_9695,N_9546);
nand U13837 (N_13837,N_9074,N_11307);
nand U13838 (N_13838,N_9096,N_10655);
nand U13839 (N_13839,N_11198,N_9883);
or U13840 (N_13840,N_10773,N_11585);
nor U13841 (N_13841,N_11600,N_9085);
nand U13842 (N_13842,N_9810,N_9196);
or U13843 (N_13843,N_9745,N_10710);
or U13844 (N_13844,N_9443,N_10891);
or U13845 (N_13845,N_9341,N_9593);
nand U13846 (N_13846,N_11247,N_9283);
nand U13847 (N_13847,N_11924,N_11385);
and U13848 (N_13848,N_11373,N_11209);
or U13849 (N_13849,N_11013,N_10533);
and U13850 (N_13850,N_9148,N_10804);
xnor U13851 (N_13851,N_11642,N_9026);
nor U13852 (N_13852,N_10945,N_11203);
or U13853 (N_13853,N_10561,N_9348);
nor U13854 (N_13854,N_9460,N_10201);
or U13855 (N_13855,N_9758,N_9025);
nand U13856 (N_13856,N_11956,N_10295);
and U13857 (N_13857,N_11379,N_10351);
or U13858 (N_13858,N_9512,N_10552);
or U13859 (N_13859,N_11592,N_11296);
nor U13860 (N_13860,N_10323,N_11676);
nor U13861 (N_13861,N_9475,N_10829);
and U13862 (N_13862,N_11169,N_11499);
nor U13863 (N_13863,N_9246,N_9119);
or U13864 (N_13864,N_9394,N_10960);
or U13865 (N_13865,N_10892,N_10642);
nor U13866 (N_13866,N_9879,N_10103);
and U13867 (N_13867,N_9243,N_9820);
or U13868 (N_13868,N_11056,N_9985);
xnor U13869 (N_13869,N_9994,N_10321);
nor U13870 (N_13870,N_10651,N_11401);
xnor U13871 (N_13871,N_10169,N_10318);
and U13872 (N_13872,N_9576,N_11627);
or U13873 (N_13873,N_11083,N_9077);
or U13874 (N_13874,N_10193,N_11965);
xnor U13875 (N_13875,N_11611,N_9379);
or U13876 (N_13876,N_10099,N_10027);
nor U13877 (N_13877,N_11040,N_9331);
and U13878 (N_13878,N_11837,N_9139);
nand U13879 (N_13879,N_10903,N_11048);
and U13880 (N_13880,N_10368,N_9639);
nand U13881 (N_13881,N_10398,N_10311);
nor U13882 (N_13882,N_9289,N_11657);
nor U13883 (N_13883,N_11659,N_11117);
xnor U13884 (N_13884,N_11115,N_10041);
nor U13885 (N_13885,N_9991,N_10745);
xor U13886 (N_13886,N_9979,N_11996);
xnor U13887 (N_13887,N_11214,N_10642);
nor U13888 (N_13888,N_9812,N_9305);
nand U13889 (N_13889,N_10811,N_9289);
and U13890 (N_13890,N_11723,N_11456);
nand U13891 (N_13891,N_10031,N_9128);
and U13892 (N_13892,N_11769,N_10269);
nand U13893 (N_13893,N_10982,N_11110);
nand U13894 (N_13894,N_10160,N_11050);
nor U13895 (N_13895,N_9210,N_10116);
or U13896 (N_13896,N_11249,N_9018);
nand U13897 (N_13897,N_10525,N_9333);
nor U13898 (N_13898,N_9357,N_9522);
or U13899 (N_13899,N_11441,N_9222);
nand U13900 (N_13900,N_11371,N_9728);
or U13901 (N_13901,N_10956,N_11725);
xor U13902 (N_13902,N_10714,N_10558);
nor U13903 (N_13903,N_10779,N_11905);
and U13904 (N_13904,N_11288,N_11399);
xor U13905 (N_13905,N_11666,N_9848);
and U13906 (N_13906,N_9591,N_10320);
xnor U13907 (N_13907,N_11353,N_11762);
nor U13908 (N_13908,N_11584,N_10055);
or U13909 (N_13909,N_11451,N_10576);
nor U13910 (N_13910,N_11881,N_10446);
or U13911 (N_13911,N_9067,N_10966);
or U13912 (N_13912,N_10631,N_10380);
and U13913 (N_13913,N_10716,N_9837);
and U13914 (N_13914,N_9257,N_10495);
or U13915 (N_13915,N_9043,N_10992);
or U13916 (N_13916,N_11299,N_11059);
nor U13917 (N_13917,N_11854,N_9588);
or U13918 (N_13918,N_11102,N_9749);
and U13919 (N_13919,N_11864,N_11669);
or U13920 (N_13920,N_9419,N_11297);
nand U13921 (N_13921,N_10054,N_10304);
nor U13922 (N_13922,N_10858,N_10044);
and U13923 (N_13923,N_10346,N_9409);
nor U13924 (N_13924,N_9136,N_10140);
xnor U13925 (N_13925,N_10813,N_10917);
and U13926 (N_13926,N_9502,N_11803);
xnor U13927 (N_13927,N_11488,N_10804);
and U13928 (N_13928,N_11406,N_11335);
or U13929 (N_13929,N_11329,N_11505);
and U13930 (N_13930,N_10671,N_9505);
or U13931 (N_13931,N_9726,N_11896);
and U13932 (N_13932,N_9245,N_9112);
or U13933 (N_13933,N_9209,N_9715);
nor U13934 (N_13934,N_10473,N_10391);
or U13935 (N_13935,N_9476,N_10283);
nor U13936 (N_13936,N_9775,N_10192);
nor U13937 (N_13937,N_11425,N_9577);
and U13938 (N_13938,N_10731,N_11337);
nor U13939 (N_13939,N_11701,N_9734);
or U13940 (N_13940,N_10001,N_11388);
or U13941 (N_13941,N_11358,N_9954);
nand U13942 (N_13942,N_10552,N_9552);
nor U13943 (N_13943,N_11128,N_9871);
nand U13944 (N_13944,N_9976,N_11767);
nand U13945 (N_13945,N_9456,N_11312);
nand U13946 (N_13946,N_9556,N_9798);
or U13947 (N_13947,N_10275,N_10653);
xnor U13948 (N_13948,N_11287,N_10589);
xor U13949 (N_13949,N_11530,N_9725);
or U13950 (N_13950,N_10126,N_9462);
xnor U13951 (N_13951,N_11650,N_10533);
nand U13952 (N_13952,N_9379,N_11433);
or U13953 (N_13953,N_11454,N_11399);
xor U13954 (N_13954,N_10795,N_9937);
nand U13955 (N_13955,N_11405,N_10585);
and U13956 (N_13956,N_9174,N_10819);
and U13957 (N_13957,N_9124,N_11592);
or U13958 (N_13958,N_9922,N_10764);
xor U13959 (N_13959,N_9236,N_11670);
or U13960 (N_13960,N_9629,N_9661);
and U13961 (N_13961,N_9958,N_9980);
and U13962 (N_13962,N_10432,N_10637);
xnor U13963 (N_13963,N_11077,N_9162);
or U13964 (N_13964,N_11300,N_9441);
and U13965 (N_13965,N_11310,N_11247);
nor U13966 (N_13966,N_10518,N_10954);
or U13967 (N_13967,N_10627,N_9549);
or U13968 (N_13968,N_10697,N_11569);
and U13969 (N_13969,N_11667,N_10721);
nor U13970 (N_13970,N_9572,N_10735);
and U13971 (N_13971,N_10453,N_11844);
or U13972 (N_13972,N_11366,N_9211);
nand U13973 (N_13973,N_10274,N_9400);
nor U13974 (N_13974,N_11310,N_11723);
xnor U13975 (N_13975,N_9715,N_10059);
nor U13976 (N_13976,N_9065,N_11997);
nor U13977 (N_13977,N_9090,N_9870);
nand U13978 (N_13978,N_10849,N_11843);
or U13979 (N_13979,N_11331,N_10340);
and U13980 (N_13980,N_11469,N_9443);
xor U13981 (N_13981,N_11302,N_10502);
nand U13982 (N_13982,N_11396,N_11965);
or U13983 (N_13983,N_9156,N_11235);
xor U13984 (N_13984,N_11901,N_11980);
nor U13985 (N_13985,N_10092,N_9220);
or U13986 (N_13986,N_9565,N_9923);
nor U13987 (N_13987,N_9532,N_11969);
or U13988 (N_13988,N_10645,N_9355);
nor U13989 (N_13989,N_9271,N_9099);
or U13990 (N_13990,N_10759,N_11128);
and U13991 (N_13991,N_9406,N_10632);
or U13992 (N_13992,N_10616,N_11054);
nand U13993 (N_13993,N_9707,N_11115);
xnor U13994 (N_13994,N_11895,N_11380);
or U13995 (N_13995,N_9904,N_9980);
and U13996 (N_13996,N_9001,N_9838);
nor U13997 (N_13997,N_10550,N_11639);
and U13998 (N_13998,N_11281,N_11185);
and U13999 (N_13999,N_9564,N_9335);
nand U14000 (N_14000,N_11233,N_9079);
and U14001 (N_14001,N_10184,N_11401);
or U14002 (N_14002,N_9110,N_10963);
or U14003 (N_14003,N_10813,N_10894);
nor U14004 (N_14004,N_9569,N_10562);
and U14005 (N_14005,N_11592,N_10588);
nand U14006 (N_14006,N_10568,N_9189);
nand U14007 (N_14007,N_10157,N_11299);
xor U14008 (N_14008,N_11733,N_10464);
nand U14009 (N_14009,N_10751,N_9993);
nand U14010 (N_14010,N_9767,N_9967);
or U14011 (N_14011,N_9071,N_11445);
xor U14012 (N_14012,N_11213,N_9535);
nor U14013 (N_14013,N_11042,N_11583);
nand U14014 (N_14014,N_11027,N_9467);
nand U14015 (N_14015,N_10271,N_9173);
nor U14016 (N_14016,N_11854,N_11396);
nand U14017 (N_14017,N_10602,N_10448);
and U14018 (N_14018,N_10116,N_9919);
nor U14019 (N_14019,N_10262,N_10849);
and U14020 (N_14020,N_9942,N_11858);
or U14021 (N_14021,N_9631,N_10001);
nand U14022 (N_14022,N_10430,N_10875);
nor U14023 (N_14023,N_10620,N_10611);
or U14024 (N_14024,N_11616,N_10717);
nor U14025 (N_14025,N_10526,N_10410);
nor U14026 (N_14026,N_11190,N_10197);
xnor U14027 (N_14027,N_10118,N_10860);
and U14028 (N_14028,N_10933,N_11516);
and U14029 (N_14029,N_10446,N_11508);
and U14030 (N_14030,N_10059,N_9537);
and U14031 (N_14031,N_9141,N_11414);
and U14032 (N_14032,N_11117,N_11430);
xnor U14033 (N_14033,N_10320,N_11030);
or U14034 (N_14034,N_10148,N_9456);
nor U14035 (N_14035,N_10108,N_10507);
nor U14036 (N_14036,N_10483,N_11968);
or U14037 (N_14037,N_9119,N_10920);
xor U14038 (N_14038,N_11725,N_11013);
nand U14039 (N_14039,N_9734,N_10160);
nor U14040 (N_14040,N_11186,N_9200);
and U14041 (N_14041,N_10499,N_11710);
or U14042 (N_14042,N_9769,N_10389);
and U14043 (N_14043,N_11396,N_9637);
or U14044 (N_14044,N_11506,N_11777);
nor U14045 (N_14045,N_10171,N_10196);
and U14046 (N_14046,N_10366,N_10022);
nor U14047 (N_14047,N_9055,N_11491);
and U14048 (N_14048,N_9120,N_11534);
xor U14049 (N_14049,N_10071,N_10443);
nand U14050 (N_14050,N_11513,N_9637);
nor U14051 (N_14051,N_9863,N_9320);
or U14052 (N_14052,N_10745,N_11851);
or U14053 (N_14053,N_10752,N_10405);
nand U14054 (N_14054,N_11591,N_11748);
or U14055 (N_14055,N_10283,N_11292);
and U14056 (N_14056,N_11138,N_9042);
and U14057 (N_14057,N_10130,N_11521);
nand U14058 (N_14058,N_11485,N_10573);
nor U14059 (N_14059,N_10912,N_10276);
and U14060 (N_14060,N_11134,N_10867);
xnor U14061 (N_14061,N_11624,N_11240);
xor U14062 (N_14062,N_11303,N_10249);
xor U14063 (N_14063,N_10908,N_11881);
nand U14064 (N_14064,N_10232,N_11562);
and U14065 (N_14065,N_10078,N_9589);
or U14066 (N_14066,N_9009,N_11100);
xor U14067 (N_14067,N_9713,N_11688);
nand U14068 (N_14068,N_10417,N_10794);
nand U14069 (N_14069,N_11209,N_10487);
nand U14070 (N_14070,N_10715,N_9041);
and U14071 (N_14071,N_11299,N_11537);
or U14072 (N_14072,N_11531,N_10897);
xnor U14073 (N_14073,N_11687,N_9198);
nand U14074 (N_14074,N_9870,N_10106);
or U14075 (N_14075,N_9858,N_9101);
and U14076 (N_14076,N_11771,N_11429);
or U14077 (N_14077,N_11690,N_9021);
or U14078 (N_14078,N_9291,N_10920);
xnor U14079 (N_14079,N_9960,N_11573);
or U14080 (N_14080,N_10749,N_9631);
nor U14081 (N_14081,N_11213,N_10562);
nor U14082 (N_14082,N_11721,N_9159);
and U14083 (N_14083,N_10398,N_11612);
or U14084 (N_14084,N_10147,N_9039);
and U14085 (N_14085,N_11570,N_11287);
and U14086 (N_14086,N_9586,N_11300);
nor U14087 (N_14087,N_10283,N_11938);
and U14088 (N_14088,N_10650,N_10179);
and U14089 (N_14089,N_9479,N_9062);
and U14090 (N_14090,N_10732,N_11850);
and U14091 (N_14091,N_10170,N_10555);
nor U14092 (N_14092,N_10304,N_9452);
xor U14093 (N_14093,N_10787,N_11032);
nor U14094 (N_14094,N_9315,N_9118);
nand U14095 (N_14095,N_11313,N_10193);
nor U14096 (N_14096,N_10768,N_10275);
nand U14097 (N_14097,N_11918,N_9558);
or U14098 (N_14098,N_10472,N_9969);
and U14099 (N_14099,N_11104,N_11642);
nor U14100 (N_14100,N_11447,N_10348);
nand U14101 (N_14101,N_9496,N_11008);
and U14102 (N_14102,N_9821,N_11422);
nand U14103 (N_14103,N_9222,N_9556);
xnor U14104 (N_14104,N_9920,N_11024);
and U14105 (N_14105,N_9794,N_9601);
nand U14106 (N_14106,N_11501,N_10735);
or U14107 (N_14107,N_9376,N_9800);
nand U14108 (N_14108,N_11152,N_9977);
nor U14109 (N_14109,N_10060,N_10263);
nand U14110 (N_14110,N_11296,N_9243);
and U14111 (N_14111,N_10766,N_10449);
nand U14112 (N_14112,N_9432,N_11633);
xnor U14113 (N_14113,N_9530,N_11327);
xnor U14114 (N_14114,N_11967,N_11326);
or U14115 (N_14115,N_11966,N_9524);
xor U14116 (N_14116,N_11582,N_10902);
nor U14117 (N_14117,N_11743,N_11167);
nand U14118 (N_14118,N_10776,N_10446);
and U14119 (N_14119,N_10317,N_9745);
nand U14120 (N_14120,N_10010,N_11822);
or U14121 (N_14121,N_11152,N_10717);
xor U14122 (N_14122,N_10336,N_9535);
nor U14123 (N_14123,N_11801,N_11222);
and U14124 (N_14124,N_11472,N_9481);
or U14125 (N_14125,N_11901,N_10743);
and U14126 (N_14126,N_9241,N_11033);
nand U14127 (N_14127,N_11532,N_9835);
nand U14128 (N_14128,N_10478,N_9530);
nand U14129 (N_14129,N_11943,N_10038);
and U14130 (N_14130,N_10774,N_11662);
and U14131 (N_14131,N_9824,N_9964);
nand U14132 (N_14132,N_9914,N_9436);
nand U14133 (N_14133,N_9321,N_9083);
and U14134 (N_14134,N_10875,N_9181);
and U14135 (N_14135,N_9862,N_10105);
and U14136 (N_14136,N_10775,N_11194);
or U14137 (N_14137,N_9238,N_9842);
or U14138 (N_14138,N_11516,N_9699);
nor U14139 (N_14139,N_11695,N_10931);
or U14140 (N_14140,N_9881,N_11282);
nand U14141 (N_14141,N_9013,N_11044);
xor U14142 (N_14142,N_10843,N_11526);
and U14143 (N_14143,N_11470,N_9340);
nor U14144 (N_14144,N_11610,N_11430);
xnor U14145 (N_14145,N_9134,N_11045);
or U14146 (N_14146,N_10225,N_9883);
and U14147 (N_14147,N_9246,N_11565);
nor U14148 (N_14148,N_10226,N_9249);
and U14149 (N_14149,N_11546,N_9189);
nor U14150 (N_14150,N_9276,N_9974);
and U14151 (N_14151,N_10065,N_9894);
or U14152 (N_14152,N_9899,N_11715);
nor U14153 (N_14153,N_9216,N_9044);
nor U14154 (N_14154,N_11667,N_9241);
or U14155 (N_14155,N_11153,N_9409);
and U14156 (N_14156,N_9047,N_11335);
nor U14157 (N_14157,N_10262,N_10083);
and U14158 (N_14158,N_11839,N_11987);
and U14159 (N_14159,N_9496,N_11251);
or U14160 (N_14160,N_9388,N_9342);
and U14161 (N_14161,N_11875,N_11714);
xnor U14162 (N_14162,N_10324,N_9443);
or U14163 (N_14163,N_11251,N_9015);
or U14164 (N_14164,N_11878,N_9527);
or U14165 (N_14165,N_10483,N_9644);
nor U14166 (N_14166,N_10759,N_11530);
nor U14167 (N_14167,N_9732,N_9301);
nand U14168 (N_14168,N_9968,N_9990);
or U14169 (N_14169,N_9447,N_10662);
nor U14170 (N_14170,N_11358,N_10010);
or U14171 (N_14171,N_9975,N_9545);
nor U14172 (N_14172,N_9681,N_9201);
nand U14173 (N_14173,N_10327,N_9927);
nand U14174 (N_14174,N_11003,N_10991);
nor U14175 (N_14175,N_9486,N_11736);
and U14176 (N_14176,N_10663,N_9325);
or U14177 (N_14177,N_9264,N_9016);
nor U14178 (N_14178,N_11009,N_9849);
and U14179 (N_14179,N_10464,N_10766);
xor U14180 (N_14180,N_9136,N_9153);
nand U14181 (N_14181,N_9282,N_10696);
nor U14182 (N_14182,N_11034,N_10097);
nor U14183 (N_14183,N_11299,N_9792);
nand U14184 (N_14184,N_9212,N_11263);
or U14185 (N_14185,N_9141,N_9839);
or U14186 (N_14186,N_9223,N_11879);
and U14187 (N_14187,N_11390,N_9731);
xnor U14188 (N_14188,N_9582,N_11431);
and U14189 (N_14189,N_11162,N_10884);
and U14190 (N_14190,N_9415,N_9535);
nand U14191 (N_14191,N_9510,N_9382);
or U14192 (N_14192,N_10097,N_10336);
and U14193 (N_14193,N_11720,N_10300);
nand U14194 (N_14194,N_9409,N_9078);
nor U14195 (N_14195,N_11597,N_10703);
xnor U14196 (N_14196,N_9044,N_10103);
and U14197 (N_14197,N_9728,N_11913);
and U14198 (N_14198,N_9410,N_10838);
nand U14199 (N_14199,N_10833,N_11272);
or U14200 (N_14200,N_9515,N_9929);
and U14201 (N_14201,N_10816,N_9364);
or U14202 (N_14202,N_9048,N_10046);
or U14203 (N_14203,N_10682,N_11326);
and U14204 (N_14204,N_11032,N_9677);
and U14205 (N_14205,N_11489,N_11161);
or U14206 (N_14206,N_10415,N_10177);
nand U14207 (N_14207,N_11131,N_10061);
nor U14208 (N_14208,N_9973,N_11754);
or U14209 (N_14209,N_11513,N_11431);
or U14210 (N_14210,N_9958,N_11459);
or U14211 (N_14211,N_11967,N_10327);
nor U14212 (N_14212,N_10112,N_10352);
nand U14213 (N_14213,N_10574,N_11767);
nor U14214 (N_14214,N_10042,N_11029);
xnor U14215 (N_14215,N_9693,N_9750);
or U14216 (N_14216,N_9740,N_9639);
xnor U14217 (N_14217,N_11363,N_11659);
nand U14218 (N_14218,N_11708,N_11895);
nand U14219 (N_14219,N_10981,N_9385);
nand U14220 (N_14220,N_11524,N_9144);
nand U14221 (N_14221,N_10188,N_10275);
or U14222 (N_14222,N_11471,N_11371);
and U14223 (N_14223,N_10190,N_9650);
or U14224 (N_14224,N_10636,N_9133);
nand U14225 (N_14225,N_9865,N_11797);
xor U14226 (N_14226,N_10118,N_10978);
xor U14227 (N_14227,N_9866,N_9116);
or U14228 (N_14228,N_9340,N_11669);
nand U14229 (N_14229,N_9679,N_10674);
xnor U14230 (N_14230,N_10306,N_10507);
xnor U14231 (N_14231,N_10037,N_9833);
and U14232 (N_14232,N_10626,N_9479);
and U14233 (N_14233,N_10700,N_9170);
xnor U14234 (N_14234,N_10714,N_10631);
or U14235 (N_14235,N_11839,N_11217);
xor U14236 (N_14236,N_11995,N_10450);
or U14237 (N_14237,N_10387,N_11256);
xor U14238 (N_14238,N_10918,N_10405);
and U14239 (N_14239,N_9876,N_11697);
nand U14240 (N_14240,N_9895,N_9894);
nor U14241 (N_14241,N_10617,N_11104);
and U14242 (N_14242,N_9760,N_11904);
or U14243 (N_14243,N_11722,N_9743);
nor U14244 (N_14244,N_11874,N_10018);
or U14245 (N_14245,N_11740,N_9522);
nor U14246 (N_14246,N_10173,N_10338);
or U14247 (N_14247,N_10273,N_10102);
and U14248 (N_14248,N_9784,N_11173);
nor U14249 (N_14249,N_11201,N_9971);
xor U14250 (N_14250,N_10416,N_10630);
and U14251 (N_14251,N_9309,N_10161);
nor U14252 (N_14252,N_10685,N_11874);
nor U14253 (N_14253,N_10199,N_9826);
nor U14254 (N_14254,N_9262,N_9578);
nor U14255 (N_14255,N_11116,N_11139);
nor U14256 (N_14256,N_10472,N_9625);
xnor U14257 (N_14257,N_9510,N_9927);
nand U14258 (N_14258,N_11412,N_11916);
or U14259 (N_14259,N_9062,N_9433);
nand U14260 (N_14260,N_10385,N_10455);
and U14261 (N_14261,N_9412,N_10870);
or U14262 (N_14262,N_10114,N_11166);
nand U14263 (N_14263,N_9699,N_11525);
nand U14264 (N_14264,N_11586,N_11038);
or U14265 (N_14265,N_11402,N_11870);
nand U14266 (N_14266,N_9088,N_9199);
nand U14267 (N_14267,N_11424,N_9803);
nand U14268 (N_14268,N_10810,N_11091);
nand U14269 (N_14269,N_10140,N_11660);
and U14270 (N_14270,N_11167,N_9266);
and U14271 (N_14271,N_10886,N_9742);
or U14272 (N_14272,N_9325,N_9651);
and U14273 (N_14273,N_10144,N_9848);
nor U14274 (N_14274,N_10475,N_11826);
or U14275 (N_14275,N_9695,N_11228);
or U14276 (N_14276,N_10729,N_11580);
or U14277 (N_14277,N_10021,N_9283);
xor U14278 (N_14278,N_9739,N_10102);
or U14279 (N_14279,N_9298,N_10367);
or U14280 (N_14280,N_9696,N_10658);
and U14281 (N_14281,N_9266,N_9137);
or U14282 (N_14282,N_10415,N_9183);
and U14283 (N_14283,N_11371,N_9902);
xor U14284 (N_14284,N_9982,N_11284);
or U14285 (N_14285,N_9697,N_9809);
or U14286 (N_14286,N_9736,N_10820);
and U14287 (N_14287,N_11337,N_9356);
xnor U14288 (N_14288,N_11097,N_11639);
and U14289 (N_14289,N_11156,N_10229);
xor U14290 (N_14290,N_10087,N_10073);
nor U14291 (N_14291,N_9241,N_9259);
and U14292 (N_14292,N_9765,N_11016);
or U14293 (N_14293,N_9989,N_10289);
or U14294 (N_14294,N_9307,N_11126);
and U14295 (N_14295,N_9958,N_11964);
nor U14296 (N_14296,N_10345,N_11483);
or U14297 (N_14297,N_10832,N_11100);
nand U14298 (N_14298,N_11488,N_10763);
and U14299 (N_14299,N_11623,N_10810);
nor U14300 (N_14300,N_10133,N_10490);
nand U14301 (N_14301,N_10705,N_9544);
xor U14302 (N_14302,N_9660,N_11511);
nor U14303 (N_14303,N_11447,N_10529);
nand U14304 (N_14304,N_11686,N_9257);
and U14305 (N_14305,N_10663,N_9726);
xnor U14306 (N_14306,N_9407,N_11274);
or U14307 (N_14307,N_9223,N_9348);
nand U14308 (N_14308,N_10403,N_10578);
nand U14309 (N_14309,N_11034,N_11498);
or U14310 (N_14310,N_10297,N_9746);
and U14311 (N_14311,N_9255,N_9458);
or U14312 (N_14312,N_10915,N_10643);
nor U14313 (N_14313,N_9034,N_10598);
xor U14314 (N_14314,N_11786,N_10639);
or U14315 (N_14315,N_10749,N_11618);
and U14316 (N_14316,N_9371,N_11558);
nor U14317 (N_14317,N_9452,N_9835);
nand U14318 (N_14318,N_11264,N_9707);
or U14319 (N_14319,N_10619,N_9635);
nor U14320 (N_14320,N_9193,N_9215);
and U14321 (N_14321,N_10977,N_10677);
xnor U14322 (N_14322,N_9234,N_9414);
xnor U14323 (N_14323,N_11849,N_9003);
and U14324 (N_14324,N_9156,N_10811);
or U14325 (N_14325,N_9211,N_11473);
and U14326 (N_14326,N_11420,N_9298);
xor U14327 (N_14327,N_10355,N_9100);
or U14328 (N_14328,N_11481,N_11333);
nor U14329 (N_14329,N_10724,N_9520);
or U14330 (N_14330,N_11135,N_9347);
nor U14331 (N_14331,N_9792,N_11051);
xnor U14332 (N_14332,N_10710,N_9591);
and U14333 (N_14333,N_9462,N_9524);
xnor U14334 (N_14334,N_9237,N_10510);
nand U14335 (N_14335,N_11505,N_10154);
or U14336 (N_14336,N_9505,N_11013);
and U14337 (N_14337,N_9462,N_10086);
nor U14338 (N_14338,N_11285,N_10387);
nand U14339 (N_14339,N_11230,N_11187);
and U14340 (N_14340,N_10121,N_11389);
or U14341 (N_14341,N_10054,N_10479);
or U14342 (N_14342,N_11385,N_9148);
nor U14343 (N_14343,N_11912,N_11655);
nand U14344 (N_14344,N_9507,N_11740);
nand U14345 (N_14345,N_9195,N_10268);
or U14346 (N_14346,N_9144,N_10156);
nor U14347 (N_14347,N_9747,N_10563);
and U14348 (N_14348,N_11859,N_11655);
nand U14349 (N_14349,N_10422,N_11989);
and U14350 (N_14350,N_11568,N_9923);
nor U14351 (N_14351,N_9159,N_10172);
or U14352 (N_14352,N_9958,N_10703);
and U14353 (N_14353,N_9269,N_11687);
nand U14354 (N_14354,N_10666,N_10557);
nand U14355 (N_14355,N_11050,N_9102);
or U14356 (N_14356,N_10734,N_10751);
and U14357 (N_14357,N_11066,N_11462);
and U14358 (N_14358,N_9070,N_10015);
nand U14359 (N_14359,N_10903,N_9850);
and U14360 (N_14360,N_11262,N_9671);
and U14361 (N_14361,N_10031,N_9022);
or U14362 (N_14362,N_9675,N_11919);
nor U14363 (N_14363,N_11888,N_11927);
nand U14364 (N_14364,N_10323,N_9647);
nand U14365 (N_14365,N_11312,N_11351);
nand U14366 (N_14366,N_11357,N_11972);
or U14367 (N_14367,N_10785,N_9261);
or U14368 (N_14368,N_9250,N_9097);
nor U14369 (N_14369,N_11303,N_9884);
and U14370 (N_14370,N_10321,N_10235);
or U14371 (N_14371,N_9878,N_11980);
and U14372 (N_14372,N_11663,N_10360);
nor U14373 (N_14373,N_11147,N_11733);
nand U14374 (N_14374,N_9836,N_9503);
nor U14375 (N_14375,N_10589,N_11255);
nor U14376 (N_14376,N_11247,N_11855);
or U14377 (N_14377,N_9272,N_9561);
or U14378 (N_14378,N_10226,N_9302);
nor U14379 (N_14379,N_10142,N_10690);
xnor U14380 (N_14380,N_10282,N_11745);
nor U14381 (N_14381,N_10818,N_11392);
nor U14382 (N_14382,N_10232,N_9356);
or U14383 (N_14383,N_10051,N_9137);
nor U14384 (N_14384,N_10322,N_11685);
or U14385 (N_14385,N_9014,N_11012);
and U14386 (N_14386,N_10431,N_10271);
or U14387 (N_14387,N_10892,N_9857);
nor U14388 (N_14388,N_10734,N_11749);
and U14389 (N_14389,N_9295,N_10504);
and U14390 (N_14390,N_9906,N_11265);
nand U14391 (N_14391,N_9156,N_10423);
or U14392 (N_14392,N_10111,N_11318);
xnor U14393 (N_14393,N_9080,N_11602);
and U14394 (N_14394,N_9014,N_9825);
nand U14395 (N_14395,N_11207,N_11179);
nand U14396 (N_14396,N_9713,N_11268);
or U14397 (N_14397,N_10538,N_11305);
and U14398 (N_14398,N_10017,N_9015);
nand U14399 (N_14399,N_11431,N_11259);
nand U14400 (N_14400,N_10661,N_9505);
or U14401 (N_14401,N_9863,N_10478);
or U14402 (N_14402,N_9732,N_10823);
or U14403 (N_14403,N_9338,N_9454);
and U14404 (N_14404,N_9273,N_9010);
nand U14405 (N_14405,N_10490,N_9666);
nand U14406 (N_14406,N_11528,N_9287);
and U14407 (N_14407,N_9163,N_9603);
nor U14408 (N_14408,N_10860,N_9256);
nor U14409 (N_14409,N_9109,N_11176);
nor U14410 (N_14410,N_11786,N_11976);
nand U14411 (N_14411,N_10201,N_9800);
nand U14412 (N_14412,N_9413,N_9722);
or U14413 (N_14413,N_11601,N_10867);
nand U14414 (N_14414,N_11857,N_9235);
and U14415 (N_14415,N_9569,N_9295);
or U14416 (N_14416,N_11036,N_10941);
and U14417 (N_14417,N_10923,N_10029);
nand U14418 (N_14418,N_11976,N_11571);
and U14419 (N_14419,N_11465,N_11844);
nor U14420 (N_14420,N_11870,N_9750);
nor U14421 (N_14421,N_11896,N_10551);
and U14422 (N_14422,N_9066,N_9573);
nor U14423 (N_14423,N_9355,N_11322);
nor U14424 (N_14424,N_9573,N_10485);
xnor U14425 (N_14425,N_11751,N_9748);
and U14426 (N_14426,N_9462,N_11330);
and U14427 (N_14427,N_11372,N_9686);
nand U14428 (N_14428,N_10263,N_10173);
or U14429 (N_14429,N_9701,N_10583);
nor U14430 (N_14430,N_10524,N_10401);
and U14431 (N_14431,N_9077,N_11440);
and U14432 (N_14432,N_11849,N_11592);
and U14433 (N_14433,N_10675,N_9191);
and U14434 (N_14434,N_11435,N_10864);
xnor U14435 (N_14435,N_9335,N_11971);
nor U14436 (N_14436,N_9348,N_10496);
nor U14437 (N_14437,N_9750,N_9986);
xnor U14438 (N_14438,N_11997,N_9061);
or U14439 (N_14439,N_9709,N_10215);
xnor U14440 (N_14440,N_9629,N_9252);
nand U14441 (N_14441,N_11348,N_9249);
or U14442 (N_14442,N_10313,N_9305);
nor U14443 (N_14443,N_10984,N_10483);
xor U14444 (N_14444,N_11241,N_9946);
xor U14445 (N_14445,N_11387,N_11551);
or U14446 (N_14446,N_10300,N_10220);
and U14447 (N_14447,N_11950,N_11552);
nand U14448 (N_14448,N_11978,N_9702);
xnor U14449 (N_14449,N_9128,N_10529);
and U14450 (N_14450,N_9573,N_9879);
nand U14451 (N_14451,N_11719,N_10493);
nor U14452 (N_14452,N_9553,N_11273);
nor U14453 (N_14453,N_10941,N_9344);
nor U14454 (N_14454,N_11662,N_9249);
nand U14455 (N_14455,N_11789,N_9603);
or U14456 (N_14456,N_9170,N_11334);
nor U14457 (N_14457,N_10573,N_9160);
and U14458 (N_14458,N_9689,N_11504);
xnor U14459 (N_14459,N_10346,N_10435);
xnor U14460 (N_14460,N_10619,N_11858);
nor U14461 (N_14461,N_10170,N_11475);
nand U14462 (N_14462,N_10833,N_10254);
nand U14463 (N_14463,N_10995,N_10777);
nand U14464 (N_14464,N_10596,N_9985);
nor U14465 (N_14465,N_10250,N_9996);
nand U14466 (N_14466,N_11590,N_10593);
nor U14467 (N_14467,N_9525,N_9317);
and U14468 (N_14468,N_10687,N_9429);
nor U14469 (N_14469,N_11886,N_11904);
and U14470 (N_14470,N_11084,N_10699);
or U14471 (N_14471,N_11199,N_9947);
nand U14472 (N_14472,N_10131,N_9521);
and U14473 (N_14473,N_9434,N_9810);
and U14474 (N_14474,N_11719,N_9509);
nor U14475 (N_14475,N_10354,N_11548);
and U14476 (N_14476,N_11351,N_9040);
or U14477 (N_14477,N_11691,N_11893);
or U14478 (N_14478,N_10456,N_9556);
or U14479 (N_14479,N_9740,N_9658);
nor U14480 (N_14480,N_11668,N_11136);
and U14481 (N_14481,N_9211,N_10978);
xor U14482 (N_14482,N_11013,N_10542);
nand U14483 (N_14483,N_9544,N_10087);
and U14484 (N_14484,N_10547,N_11336);
nor U14485 (N_14485,N_11403,N_10022);
or U14486 (N_14486,N_10708,N_11928);
nand U14487 (N_14487,N_10693,N_9187);
nand U14488 (N_14488,N_10470,N_10956);
or U14489 (N_14489,N_9132,N_11332);
nand U14490 (N_14490,N_11558,N_9537);
or U14491 (N_14491,N_10413,N_9507);
xnor U14492 (N_14492,N_10075,N_9346);
or U14493 (N_14493,N_9002,N_9994);
nor U14494 (N_14494,N_11235,N_9827);
nand U14495 (N_14495,N_10647,N_10590);
nand U14496 (N_14496,N_9146,N_10175);
or U14497 (N_14497,N_10348,N_9946);
xor U14498 (N_14498,N_10493,N_11781);
or U14499 (N_14499,N_10303,N_9746);
nand U14500 (N_14500,N_9181,N_9816);
or U14501 (N_14501,N_9835,N_11316);
and U14502 (N_14502,N_9577,N_10761);
nand U14503 (N_14503,N_9818,N_10618);
or U14504 (N_14504,N_10917,N_9323);
nand U14505 (N_14505,N_11113,N_9961);
or U14506 (N_14506,N_9148,N_10943);
or U14507 (N_14507,N_9970,N_10872);
and U14508 (N_14508,N_9547,N_9132);
and U14509 (N_14509,N_11159,N_10817);
nor U14510 (N_14510,N_10899,N_10140);
and U14511 (N_14511,N_9162,N_10315);
nor U14512 (N_14512,N_10482,N_11199);
xnor U14513 (N_14513,N_9801,N_9772);
and U14514 (N_14514,N_10806,N_10230);
nand U14515 (N_14515,N_11593,N_11943);
nor U14516 (N_14516,N_11766,N_9496);
and U14517 (N_14517,N_9906,N_11806);
and U14518 (N_14518,N_11450,N_9612);
xor U14519 (N_14519,N_9534,N_9581);
or U14520 (N_14520,N_11458,N_11189);
nor U14521 (N_14521,N_9511,N_9143);
nand U14522 (N_14522,N_10524,N_10933);
or U14523 (N_14523,N_11215,N_10875);
nand U14524 (N_14524,N_9351,N_10215);
and U14525 (N_14525,N_9062,N_10676);
or U14526 (N_14526,N_10214,N_10691);
nand U14527 (N_14527,N_9304,N_9024);
and U14528 (N_14528,N_9627,N_11205);
and U14529 (N_14529,N_10792,N_11009);
nand U14530 (N_14530,N_11683,N_9950);
or U14531 (N_14531,N_9443,N_11749);
and U14532 (N_14532,N_11976,N_10571);
xor U14533 (N_14533,N_10078,N_9004);
and U14534 (N_14534,N_10910,N_10774);
or U14535 (N_14535,N_10187,N_11461);
nand U14536 (N_14536,N_10179,N_9370);
nand U14537 (N_14537,N_10721,N_10218);
or U14538 (N_14538,N_10981,N_9572);
nand U14539 (N_14539,N_10154,N_9139);
and U14540 (N_14540,N_10569,N_10240);
nor U14541 (N_14541,N_10285,N_10016);
nand U14542 (N_14542,N_9437,N_9605);
nor U14543 (N_14543,N_10545,N_10051);
nand U14544 (N_14544,N_10614,N_11696);
nand U14545 (N_14545,N_9825,N_11664);
or U14546 (N_14546,N_11726,N_10457);
or U14547 (N_14547,N_9701,N_10254);
and U14548 (N_14548,N_11843,N_11775);
nand U14549 (N_14549,N_10916,N_11737);
and U14550 (N_14550,N_11692,N_9141);
xnor U14551 (N_14551,N_9351,N_10055);
or U14552 (N_14552,N_9352,N_9347);
nand U14553 (N_14553,N_11396,N_9479);
nand U14554 (N_14554,N_10360,N_11628);
xor U14555 (N_14555,N_10506,N_10479);
nand U14556 (N_14556,N_10176,N_9069);
nor U14557 (N_14557,N_10851,N_10873);
nor U14558 (N_14558,N_9392,N_10477);
and U14559 (N_14559,N_9760,N_11166);
nor U14560 (N_14560,N_11568,N_11036);
or U14561 (N_14561,N_9640,N_10765);
and U14562 (N_14562,N_11814,N_10653);
or U14563 (N_14563,N_10300,N_10586);
xnor U14564 (N_14564,N_10362,N_9311);
xor U14565 (N_14565,N_9615,N_10611);
or U14566 (N_14566,N_11919,N_9288);
nor U14567 (N_14567,N_9264,N_9493);
and U14568 (N_14568,N_10558,N_11741);
or U14569 (N_14569,N_10910,N_9635);
and U14570 (N_14570,N_11173,N_10400);
nand U14571 (N_14571,N_9336,N_11597);
nand U14572 (N_14572,N_11500,N_9709);
nor U14573 (N_14573,N_10525,N_10801);
and U14574 (N_14574,N_10145,N_11825);
nor U14575 (N_14575,N_10673,N_11865);
and U14576 (N_14576,N_11913,N_11707);
or U14577 (N_14577,N_11795,N_9201);
nand U14578 (N_14578,N_10739,N_11202);
or U14579 (N_14579,N_10812,N_10466);
or U14580 (N_14580,N_10916,N_11475);
nor U14581 (N_14581,N_9271,N_10578);
or U14582 (N_14582,N_10487,N_10905);
and U14583 (N_14583,N_10743,N_11818);
or U14584 (N_14584,N_10113,N_11446);
and U14585 (N_14585,N_11692,N_10216);
nor U14586 (N_14586,N_10363,N_10774);
nor U14587 (N_14587,N_10038,N_10519);
xor U14588 (N_14588,N_11700,N_9964);
and U14589 (N_14589,N_11467,N_9040);
and U14590 (N_14590,N_9755,N_11467);
nand U14591 (N_14591,N_11707,N_11168);
nand U14592 (N_14592,N_9767,N_9984);
or U14593 (N_14593,N_9662,N_10166);
nand U14594 (N_14594,N_10610,N_9702);
and U14595 (N_14595,N_9563,N_9020);
and U14596 (N_14596,N_10450,N_10542);
xor U14597 (N_14597,N_10057,N_9803);
nand U14598 (N_14598,N_9986,N_11183);
nand U14599 (N_14599,N_10592,N_11039);
nor U14600 (N_14600,N_11232,N_9316);
and U14601 (N_14601,N_11075,N_9423);
or U14602 (N_14602,N_11290,N_10258);
xnor U14603 (N_14603,N_9089,N_11541);
or U14604 (N_14604,N_9739,N_11303);
nor U14605 (N_14605,N_11770,N_11702);
and U14606 (N_14606,N_10620,N_10413);
and U14607 (N_14607,N_11456,N_10888);
nor U14608 (N_14608,N_10237,N_10398);
nand U14609 (N_14609,N_9019,N_11096);
nand U14610 (N_14610,N_9076,N_10288);
nor U14611 (N_14611,N_10294,N_9309);
and U14612 (N_14612,N_11983,N_10922);
and U14613 (N_14613,N_10152,N_9357);
or U14614 (N_14614,N_9641,N_9192);
nand U14615 (N_14615,N_9105,N_10500);
and U14616 (N_14616,N_10303,N_11950);
nor U14617 (N_14617,N_11546,N_9899);
or U14618 (N_14618,N_10304,N_11942);
nand U14619 (N_14619,N_9547,N_10557);
or U14620 (N_14620,N_10165,N_9218);
xor U14621 (N_14621,N_11383,N_10790);
nor U14622 (N_14622,N_11358,N_9445);
nor U14623 (N_14623,N_11576,N_10279);
nor U14624 (N_14624,N_10686,N_10329);
nand U14625 (N_14625,N_9202,N_10855);
xnor U14626 (N_14626,N_11968,N_10522);
nand U14627 (N_14627,N_10079,N_9829);
and U14628 (N_14628,N_11802,N_9057);
and U14629 (N_14629,N_9851,N_9699);
nor U14630 (N_14630,N_11654,N_10927);
nand U14631 (N_14631,N_10139,N_11446);
and U14632 (N_14632,N_9231,N_10713);
nand U14633 (N_14633,N_11564,N_11607);
and U14634 (N_14634,N_10116,N_11944);
or U14635 (N_14635,N_10719,N_9039);
or U14636 (N_14636,N_9418,N_11798);
nand U14637 (N_14637,N_9740,N_9319);
nand U14638 (N_14638,N_11701,N_11122);
nor U14639 (N_14639,N_9028,N_10244);
nand U14640 (N_14640,N_11540,N_11895);
nor U14641 (N_14641,N_11640,N_10100);
or U14642 (N_14642,N_9357,N_10701);
nand U14643 (N_14643,N_10050,N_11689);
and U14644 (N_14644,N_10823,N_10181);
nor U14645 (N_14645,N_10306,N_9177);
nor U14646 (N_14646,N_10739,N_9608);
nand U14647 (N_14647,N_10038,N_9831);
and U14648 (N_14648,N_10878,N_9583);
xnor U14649 (N_14649,N_10896,N_9305);
and U14650 (N_14650,N_10489,N_9598);
or U14651 (N_14651,N_9256,N_10096);
and U14652 (N_14652,N_9193,N_9385);
nand U14653 (N_14653,N_11021,N_10765);
xnor U14654 (N_14654,N_11340,N_10484);
or U14655 (N_14655,N_9386,N_11373);
nor U14656 (N_14656,N_10995,N_11617);
nor U14657 (N_14657,N_9319,N_11534);
or U14658 (N_14658,N_10810,N_9315);
nand U14659 (N_14659,N_9056,N_10404);
xor U14660 (N_14660,N_10440,N_10408);
and U14661 (N_14661,N_10175,N_11529);
nor U14662 (N_14662,N_11707,N_9653);
and U14663 (N_14663,N_10094,N_11256);
or U14664 (N_14664,N_9117,N_10745);
and U14665 (N_14665,N_11604,N_9387);
nand U14666 (N_14666,N_9818,N_10052);
nor U14667 (N_14667,N_10731,N_11346);
or U14668 (N_14668,N_10620,N_11539);
or U14669 (N_14669,N_9315,N_10937);
nand U14670 (N_14670,N_11005,N_11038);
nor U14671 (N_14671,N_11089,N_10481);
nor U14672 (N_14672,N_10287,N_10779);
nor U14673 (N_14673,N_9469,N_10413);
and U14674 (N_14674,N_9842,N_10529);
and U14675 (N_14675,N_9895,N_11754);
nand U14676 (N_14676,N_9657,N_10962);
nand U14677 (N_14677,N_11209,N_9776);
nor U14678 (N_14678,N_10559,N_10930);
nand U14679 (N_14679,N_11214,N_11543);
and U14680 (N_14680,N_10775,N_9704);
nor U14681 (N_14681,N_10258,N_11094);
or U14682 (N_14682,N_11360,N_9385);
and U14683 (N_14683,N_10757,N_10775);
nand U14684 (N_14684,N_11207,N_10782);
nand U14685 (N_14685,N_10972,N_10691);
and U14686 (N_14686,N_10403,N_9312);
and U14687 (N_14687,N_10508,N_11234);
and U14688 (N_14688,N_10604,N_9380);
nor U14689 (N_14689,N_9603,N_9279);
nand U14690 (N_14690,N_10985,N_10592);
or U14691 (N_14691,N_11911,N_11824);
nand U14692 (N_14692,N_11412,N_11971);
and U14693 (N_14693,N_10195,N_9083);
nor U14694 (N_14694,N_11733,N_9808);
and U14695 (N_14695,N_9094,N_11139);
nand U14696 (N_14696,N_11839,N_9828);
nand U14697 (N_14697,N_9786,N_10495);
nor U14698 (N_14698,N_10143,N_11417);
xnor U14699 (N_14699,N_9622,N_11855);
xor U14700 (N_14700,N_11088,N_9619);
nor U14701 (N_14701,N_10707,N_11148);
nand U14702 (N_14702,N_10438,N_10107);
or U14703 (N_14703,N_11193,N_10371);
and U14704 (N_14704,N_11065,N_9977);
nor U14705 (N_14705,N_11582,N_11620);
nor U14706 (N_14706,N_11676,N_9663);
nor U14707 (N_14707,N_9389,N_10545);
nand U14708 (N_14708,N_11260,N_10100);
and U14709 (N_14709,N_9100,N_11569);
nor U14710 (N_14710,N_11527,N_10967);
and U14711 (N_14711,N_9320,N_9539);
nor U14712 (N_14712,N_11578,N_9804);
nor U14713 (N_14713,N_10579,N_9505);
xnor U14714 (N_14714,N_10184,N_9355);
or U14715 (N_14715,N_11458,N_9420);
nor U14716 (N_14716,N_9347,N_9080);
nor U14717 (N_14717,N_9135,N_10899);
nor U14718 (N_14718,N_11891,N_10708);
or U14719 (N_14719,N_10641,N_11815);
and U14720 (N_14720,N_9562,N_9115);
nor U14721 (N_14721,N_11825,N_11609);
nor U14722 (N_14722,N_9723,N_10459);
or U14723 (N_14723,N_9827,N_10095);
and U14724 (N_14724,N_11056,N_9106);
or U14725 (N_14725,N_9085,N_11842);
or U14726 (N_14726,N_10083,N_9258);
or U14727 (N_14727,N_9861,N_11619);
or U14728 (N_14728,N_9332,N_9895);
and U14729 (N_14729,N_9843,N_10732);
nand U14730 (N_14730,N_10843,N_9194);
nor U14731 (N_14731,N_11916,N_10922);
nor U14732 (N_14732,N_10484,N_10640);
nand U14733 (N_14733,N_11644,N_10503);
or U14734 (N_14734,N_10218,N_11475);
or U14735 (N_14735,N_10645,N_11291);
or U14736 (N_14736,N_11233,N_10346);
and U14737 (N_14737,N_11006,N_11772);
or U14738 (N_14738,N_9541,N_11918);
and U14739 (N_14739,N_9290,N_9428);
and U14740 (N_14740,N_9132,N_9015);
or U14741 (N_14741,N_10071,N_9436);
and U14742 (N_14742,N_9929,N_9703);
or U14743 (N_14743,N_11899,N_11430);
nand U14744 (N_14744,N_9999,N_9808);
xnor U14745 (N_14745,N_9419,N_9326);
or U14746 (N_14746,N_10809,N_11724);
nor U14747 (N_14747,N_9963,N_9605);
and U14748 (N_14748,N_10375,N_11450);
nand U14749 (N_14749,N_10700,N_9820);
nand U14750 (N_14750,N_9690,N_11889);
and U14751 (N_14751,N_11282,N_11080);
or U14752 (N_14752,N_9032,N_11458);
nor U14753 (N_14753,N_11729,N_9533);
xor U14754 (N_14754,N_11387,N_9460);
or U14755 (N_14755,N_11917,N_11644);
and U14756 (N_14756,N_9197,N_10525);
or U14757 (N_14757,N_10704,N_11859);
nand U14758 (N_14758,N_9629,N_9282);
and U14759 (N_14759,N_10027,N_10564);
and U14760 (N_14760,N_11398,N_10043);
nand U14761 (N_14761,N_11866,N_11030);
or U14762 (N_14762,N_9600,N_10655);
or U14763 (N_14763,N_9069,N_11332);
or U14764 (N_14764,N_10091,N_11571);
nand U14765 (N_14765,N_10155,N_11011);
or U14766 (N_14766,N_11314,N_10125);
and U14767 (N_14767,N_10561,N_9531);
or U14768 (N_14768,N_9677,N_9024);
nand U14769 (N_14769,N_10885,N_11251);
or U14770 (N_14770,N_9902,N_11618);
and U14771 (N_14771,N_11979,N_9021);
xor U14772 (N_14772,N_9285,N_10282);
nand U14773 (N_14773,N_11779,N_10690);
and U14774 (N_14774,N_10009,N_10629);
and U14775 (N_14775,N_11850,N_11116);
and U14776 (N_14776,N_11703,N_9781);
nand U14777 (N_14777,N_9016,N_9100);
and U14778 (N_14778,N_11429,N_10203);
nor U14779 (N_14779,N_10762,N_11545);
nor U14780 (N_14780,N_10513,N_10972);
nand U14781 (N_14781,N_9793,N_9312);
nor U14782 (N_14782,N_11285,N_10538);
or U14783 (N_14783,N_11597,N_9067);
xnor U14784 (N_14784,N_9542,N_10299);
and U14785 (N_14785,N_11527,N_9388);
or U14786 (N_14786,N_9840,N_11752);
nand U14787 (N_14787,N_10191,N_11021);
nor U14788 (N_14788,N_9527,N_9188);
nor U14789 (N_14789,N_10302,N_9652);
or U14790 (N_14790,N_10456,N_11951);
nand U14791 (N_14791,N_11644,N_11367);
nand U14792 (N_14792,N_9878,N_11467);
nand U14793 (N_14793,N_9924,N_10342);
nand U14794 (N_14794,N_11521,N_10409);
nand U14795 (N_14795,N_11203,N_11934);
and U14796 (N_14796,N_9543,N_10859);
or U14797 (N_14797,N_9525,N_10559);
xnor U14798 (N_14798,N_9340,N_10855);
nor U14799 (N_14799,N_10588,N_11705);
nand U14800 (N_14800,N_9321,N_9950);
and U14801 (N_14801,N_11361,N_10922);
xor U14802 (N_14802,N_10505,N_10440);
or U14803 (N_14803,N_11377,N_9126);
nand U14804 (N_14804,N_10105,N_11211);
and U14805 (N_14805,N_9270,N_11897);
or U14806 (N_14806,N_9052,N_9595);
or U14807 (N_14807,N_10506,N_10117);
nor U14808 (N_14808,N_11016,N_10760);
nand U14809 (N_14809,N_11427,N_9145);
xnor U14810 (N_14810,N_9258,N_11971);
or U14811 (N_14811,N_9815,N_9732);
nor U14812 (N_14812,N_10431,N_11862);
xnor U14813 (N_14813,N_11207,N_11173);
and U14814 (N_14814,N_9359,N_11003);
or U14815 (N_14815,N_11422,N_11988);
nand U14816 (N_14816,N_10366,N_11149);
and U14817 (N_14817,N_11385,N_11113);
nor U14818 (N_14818,N_9657,N_11116);
xor U14819 (N_14819,N_9717,N_11256);
xnor U14820 (N_14820,N_10058,N_11099);
and U14821 (N_14821,N_11371,N_9929);
and U14822 (N_14822,N_10850,N_10074);
nor U14823 (N_14823,N_10857,N_11080);
nand U14824 (N_14824,N_10725,N_11837);
nor U14825 (N_14825,N_9286,N_9063);
nor U14826 (N_14826,N_9128,N_9497);
nor U14827 (N_14827,N_11872,N_10204);
or U14828 (N_14828,N_10845,N_9268);
nand U14829 (N_14829,N_10516,N_10194);
and U14830 (N_14830,N_9574,N_10908);
nand U14831 (N_14831,N_11544,N_10915);
or U14832 (N_14832,N_10511,N_11456);
and U14833 (N_14833,N_10754,N_10310);
nor U14834 (N_14834,N_10384,N_11882);
or U14835 (N_14835,N_11218,N_11785);
nor U14836 (N_14836,N_9114,N_9004);
xor U14837 (N_14837,N_11884,N_11406);
nand U14838 (N_14838,N_10312,N_10761);
nand U14839 (N_14839,N_11738,N_10833);
and U14840 (N_14840,N_10873,N_9927);
nand U14841 (N_14841,N_9512,N_11113);
or U14842 (N_14842,N_11276,N_10644);
or U14843 (N_14843,N_10524,N_9596);
nand U14844 (N_14844,N_11089,N_9742);
nand U14845 (N_14845,N_11354,N_11325);
or U14846 (N_14846,N_11597,N_9063);
nand U14847 (N_14847,N_9209,N_9233);
and U14848 (N_14848,N_9131,N_11259);
or U14849 (N_14849,N_11002,N_11655);
nand U14850 (N_14850,N_10387,N_9602);
or U14851 (N_14851,N_11540,N_10229);
nor U14852 (N_14852,N_9584,N_9094);
or U14853 (N_14853,N_9978,N_11053);
and U14854 (N_14854,N_11278,N_9480);
and U14855 (N_14855,N_9342,N_10309);
xnor U14856 (N_14856,N_11126,N_10733);
xnor U14857 (N_14857,N_11249,N_9896);
nand U14858 (N_14858,N_11037,N_11019);
and U14859 (N_14859,N_10841,N_9823);
and U14860 (N_14860,N_9130,N_10137);
nor U14861 (N_14861,N_9579,N_11357);
nor U14862 (N_14862,N_9293,N_10428);
xor U14863 (N_14863,N_11643,N_11374);
nand U14864 (N_14864,N_9023,N_10118);
or U14865 (N_14865,N_10278,N_10953);
nor U14866 (N_14866,N_9750,N_9540);
xor U14867 (N_14867,N_11225,N_11571);
nand U14868 (N_14868,N_11730,N_11017);
nor U14869 (N_14869,N_10819,N_11453);
nand U14870 (N_14870,N_11841,N_9105);
nor U14871 (N_14871,N_9912,N_10336);
nor U14872 (N_14872,N_9624,N_10224);
nor U14873 (N_14873,N_10250,N_10018);
or U14874 (N_14874,N_11556,N_11170);
nor U14875 (N_14875,N_9088,N_9222);
xor U14876 (N_14876,N_11809,N_10388);
or U14877 (N_14877,N_11476,N_10978);
or U14878 (N_14878,N_9507,N_9169);
and U14879 (N_14879,N_9615,N_9105);
and U14880 (N_14880,N_11432,N_11185);
xnor U14881 (N_14881,N_10546,N_11318);
nor U14882 (N_14882,N_11372,N_9869);
or U14883 (N_14883,N_9392,N_9274);
and U14884 (N_14884,N_10260,N_10968);
nor U14885 (N_14885,N_10208,N_10921);
nor U14886 (N_14886,N_10380,N_10183);
and U14887 (N_14887,N_9474,N_9469);
nor U14888 (N_14888,N_10755,N_9407);
nor U14889 (N_14889,N_9013,N_11692);
xnor U14890 (N_14890,N_9211,N_11226);
and U14891 (N_14891,N_10383,N_9577);
nand U14892 (N_14892,N_11302,N_11890);
nor U14893 (N_14893,N_10620,N_9297);
and U14894 (N_14894,N_9640,N_11343);
nor U14895 (N_14895,N_9982,N_10219);
or U14896 (N_14896,N_9793,N_9168);
and U14897 (N_14897,N_10198,N_11106);
and U14898 (N_14898,N_9078,N_9669);
and U14899 (N_14899,N_10603,N_9423);
nor U14900 (N_14900,N_11495,N_10089);
or U14901 (N_14901,N_11329,N_9672);
nand U14902 (N_14902,N_9359,N_11199);
or U14903 (N_14903,N_10650,N_11211);
and U14904 (N_14904,N_11333,N_9956);
or U14905 (N_14905,N_10113,N_11997);
and U14906 (N_14906,N_9619,N_11958);
nand U14907 (N_14907,N_9272,N_9247);
nand U14908 (N_14908,N_9854,N_9551);
and U14909 (N_14909,N_10403,N_11322);
nor U14910 (N_14910,N_10003,N_10659);
nor U14911 (N_14911,N_9187,N_9142);
nor U14912 (N_14912,N_9992,N_10349);
xnor U14913 (N_14913,N_9614,N_9647);
nor U14914 (N_14914,N_10061,N_9771);
and U14915 (N_14915,N_11766,N_11305);
and U14916 (N_14916,N_11094,N_10368);
and U14917 (N_14917,N_9929,N_10426);
or U14918 (N_14918,N_11277,N_9611);
or U14919 (N_14919,N_10670,N_11318);
xnor U14920 (N_14920,N_10743,N_11710);
nor U14921 (N_14921,N_11904,N_10844);
or U14922 (N_14922,N_9953,N_9765);
or U14923 (N_14923,N_10502,N_9094);
nor U14924 (N_14924,N_11018,N_10952);
nor U14925 (N_14925,N_10230,N_11708);
nor U14926 (N_14926,N_9817,N_10857);
xnor U14927 (N_14927,N_11714,N_9971);
or U14928 (N_14928,N_11426,N_11956);
xnor U14929 (N_14929,N_10100,N_10777);
or U14930 (N_14930,N_9583,N_11710);
or U14931 (N_14931,N_11743,N_9795);
nor U14932 (N_14932,N_11881,N_11586);
or U14933 (N_14933,N_9639,N_11610);
xor U14934 (N_14934,N_10853,N_11732);
and U14935 (N_14935,N_11450,N_9102);
nor U14936 (N_14936,N_9681,N_10346);
nand U14937 (N_14937,N_10253,N_11747);
and U14938 (N_14938,N_9635,N_11269);
nor U14939 (N_14939,N_11468,N_10539);
or U14940 (N_14940,N_10438,N_10830);
nand U14941 (N_14941,N_11986,N_9578);
and U14942 (N_14942,N_9740,N_11323);
xor U14943 (N_14943,N_10486,N_9262);
or U14944 (N_14944,N_9882,N_11918);
and U14945 (N_14945,N_11050,N_11828);
or U14946 (N_14946,N_9744,N_9176);
xnor U14947 (N_14947,N_9012,N_11438);
nand U14948 (N_14948,N_10504,N_11550);
or U14949 (N_14949,N_11332,N_9524);
nand U14950 (N_14950,N_9714,N_10116);
or U14951 (N_14951,N_11643,N_9830);
and U14952 (N_14952,N_11682,N_10878);
or U14953 (N_14953,N_11527,N_9902);
and U14954 (N_14954,N_11264,N_10273);
or U14955 (N_14955,N_11333,N_11329);
xnor U14956 (N_14956,N_11465,N_11293);
nand U14957 (N_14957,N_9924,N_10465);
xor U14958 (N_14958,N_11795,N_9915);
and U14959 (N_14959,N_11339,N_10936);
nor U14960 (N_14960,N_9868,N_9691);
nand U14961 (N_14961,N_10960,N_9133);
and U14962 (N_14962,N_9169,N_10037);
or U14963 (N_14963,N_9518,N_9295);
and U14964 (N_14964,N_10160,N_9287);
nand U14965 (N_14965,N_11651,N_9976);
and U14966 (N_14966,N_10067,N_10402);
and U14967 (N_14967,N_9482,N_9415);
nor U14968 (N_14968,N_10046,N_11192);
nand U14969 (N_14969,N_10487,N_11003);
or U14970 (N_14970,N_9382,N_9799);
nand U14971 (N_14971,N_9079,N_9559);
or U14972 (N_14972,N_10042,N_10513);
nor U14973 (N_14973,N_9500,N_9828);
xnor U14974 (N_14974,N_9981,N_10243);
nand U14975 (N_14975,N_10401,N_11272);
nand U14976 (N_14976,N_10643,N_9635);
or U14977 (N_14977,N_10266,N_10431);
nand U14978 (N_14978,N_9552,N_10216);
nor U14979 (N_14979,N_10480,N_11242);
nand U14980 (N_14980,N_9982,N_11622);
and U14981 (N_14981,N_11459,N_10419);
nand U14982 (N_14982,N_10712,N_9949);
or U14983 (N_14983,N_9962,N_10444);
xnor U14984 (N_14984,N_11352,N_11064);
nand U14985 (N_14985,N_9125,N_11765);
xnor U14986 (N_14986,N_9315,N_10750);
nand U14987 (N_14987,N_11441,N_11429);
nand U14988 (N_14988,N_10992,N_11523);
and U14989 (N_14989,N_11752,N_11490);
xor U14990 (N_14990,N_9976,N_11880);
xor U14991 (N_14991,N_11583,N_9930);
xor U14992 (N_14992,N_11960,N_11081);
nand U14993 (N_14993,N_9700,N_11122);
and U14994 (N_14994,N_10204,N_10645);
nand U14995 (N_14995,N_10804,N_10236);
xnor U14996 (N_14996,N_9512,N_9869);
nor U14997 (N_14997,N_10791,N_11614);
xor U14998 (N_14998,N_9759,N_9141);
or U14999 (N_14999,N_11055,N_10396);
and UO_0 (O_0,N_14383,N_12875);
nor UO_1 (O_1,N_12155,N_12646);
or UO_2 (O_2,N_14122,N_12200);
and UO_3 (O_3,N_12435,N_14505);
and UO_4 (O_4,N_12041,N_14341);
or UO_5 (O_5,N_12710,N_12375);
nand UO_6 (O_6,N_14470,N_13754);
or UO_7 (O_7,N_13508,N_13771);
xnor UO_8 (O_8,N_12832,N_14321);
xor UO_9 (O_9,N_13221,N_12417);
nand UO_10 (O_10,N_12960,N_13320);
or UO_11 (O_11,N_14213,N_12240);
nand UO_12 (O_12,N_14354,N_13365);
and UO_13 (O_13,N_13848,N_12172);
and UO_14 (O_14,N_13056,N_12608);
or UO_15 (O_15,N_14103,N_12777);
or UO_16 (O_16,N_14432,N_12458);
nand UO_17 (O_17,N_12560,N_12889);
xnor UO_18 (O_18,N_14583,N_14855);
nand UO_19 (O_19,N_14082,N_12291);
or UO_20 (O_20,N_14899,N_12070);
or UO_21 (O_21,N_14154,N_13307);
and UO_22 (O_22,N_14486,N_14148);
xnor UO_23 (O_23,N_12830,N_14004);
nor UO_24 (O_24,N_13305,N_12851);
and UO_25 (O_25,N_14933,N_12000);
nand UO_26 (O_26,N_12446,N_13660);
nand UO_27 (O_27,N_13512,N_12266);
or UO_28 (O_28,N_12311,N_14145);
nand UO_29 (O_29,N_13162,N_12469);
and UO_30 (O_30,N_12885,N_14248);
nor UO_31 (O_31,N_14089,N_12700);
xor UO_32 (O_32,N_14329,N_12938);
nand UO_33 (O_33,N_12053,N_12756);
nand UO_34 (O_34,N_13861,N_13743);
nand UO_35 (O_35,N_14740,N_14619);
nor UO_36 (O_36,N_12223,N_13270);
and UO_37 (O_37,N_13435,N_14837);
and UO_38 (O_38,N_14072,N_13643);
and UO_39 (O_39,N_13337,N_14070);
nor UO_40 (O_40,N_12628,N_12871);
nor UO_41 (O_41,N_13967,N_13783);
or UO_42 (O_42,N_12891,N_13709);
xnor UO_43 (O_43,N_12774,N_14053);
or UO_44 (O_44,N_12737,N_12917);
nor UO_45 (O_45,N_13716,N_12619);
and UO_46 (O_46,N_14522,N_14935);
and UO_47 (O_47,N_14296,N_14284);
and UO_48 (O_48,N_12002,N_14345);
and UO_49 (O_49,N_12431,N_12129);
or UO_50 (O_50,N_12984,N_13577);
xnor UO_51 (O_51,N_14726,N_14652);
or UO_52 (O_52,N_14706,N_14628);
xnor UO_53 (O_53,N_14451,N_14625);
or UO_54 (O_54,N_14724,N_12703);
and UO_55 (O_55,N_12970,N_14775);
xnor UO_56 (O_56,N_13515,N_14768);
or UO_57 (O_57,N_13010,N_12482);
nor UO_58 (O_58,N_14143,N_12072);
xnor UO_59 (O_59,N_14428,N_12990);
and UO_60 (O_60,N_14924,N_13186);
and UO_61 (O_61,N_14830,N_12668);
and UO_62 (O_62,N_13628,N_13913);
nor UO_63 (O_63,N_14362,N_14828);
xor UO_64 (O_64,N_12135,N_13686);
nor UO_65 (O_65,N_13419,N_13616);
and UO_66 (O_66,N_14887,N_12963);
and UO_67 (O_67,N_13853,N_13016);
and UO_68 (O_68,N_12733,N_14635);
or UO_69 (O_69,N_13361,N_13450);
nor UO_70 (O_70,N_14964,N_12570);
nor UO_71 (O_71,N_12078,N_12670);
or UO_72 (O_72,N_14340,N_13411);
and UO_73 (O_73,N_14208,N_12962);
or UO_74 (O_74,N_13585,N_13864);
or UO_75 (O_75,N_14790,N_13963);
or UO_76 (O_76,N_12232,N_14506);
or UO_77 (O_77,N_13812,N_12309);
nor UO_78 (O_78,N_13103,N_13413);
xnor UO_79 (O_79,N_14204,N_13784);
or UO_80 (O_80,N_13164,N_12250);
and UO_81 (O_81,N_14422,N_12828);
and UO_82 (O_82,N_13373,N_14045);
and UO_83 (O_83,N_12447,N_12075);
or UO_84 (O_84,N_13766,N_13761);
and UO_85 (O_85,N_13328,N_14403);
or UO_86 (O_86,N_14821,N_14377);
and UO_87 (O_87,N_13637,N_13332);
nand UO_88 (O_88,N_13844,N_14541);
or UO_89 (O_89,N_14744,N_14269);
nand UO_90 (O_90,N_14916,N_12429);
nand UO_91 (O_91,N_12811,N_12182);
and UO_92 (O_92,N_14511,N_12669);
and UO_93 (O_93,N_12799,N_12350);
nor UO_94 (O_94,N_13691,N_13827);
nor UO_95 (O_95,N_13318,N_14299);
xor UO_96 (O_96,N_13323,N_12788);
nand UO_97 (O_97,N_14934,N_12790);
nand UO_98 (O_98,N_13146,N_14315);
xor UO_99 (O_99,N_12996,N_13917);
nor UO_100 (O_100,N_14127,N_13541);
nand UO_101 (O_101,N_12982,N_13813);
and UO_102 (O_102,N_14263,N_13656);
nor UO_103 (O_103,N_13747,N_14474);
or UO_104 (O_104,N_12983,N_13206);
and UO_105 (O_105,N_13204,N_13817);
or UO_106 (O_106,N_12198,N_14244);
nor UO_107 (O_107,N_12042,N_13354);
and UO_108 (O_108,N_12210,N_14512);
nand UO_109 (O_109,N_13017,N_13054);
nand UO_110 (O_110,N_14438,N_13926);
or UO_111 (O_111,N_13145,N_13887);
nor UO_112 (O_112,N_14287,N_13339);
nand UO_113 (O_113,N_14491,N_12927);
nor UO_114 (O_114,N_12787,N_13382);
nor UO_115 (O_115,N_14712,N_13961);
xnor UO_116 (O_116,N_12762,N_12679);
nand UO_117 (O_117,N_13936,N_14226);
nor UO_118 (O_118,N_14551,N_13989);
or UO_119 (O_119,N_13938,N_13454);
nand UO_120 (O_120,N_13797,N_13654);
nor UO_121 (O_121,N_14995,N_14503);
or UO_122 (O_122,N_14693,N_12086);
and UO_123 (O_123,N_14499,N_12015);
nand UO_124 (O_124,N_12113,N_13526);
and UO_125 (O_125,N_12330,N_13424);
nor UO_126 (O_126,N_13004,N_12823);
or UO_127 (O_127,N_14202,N_14741);
or UO_128 (O_128,N_12284,N_14643);
or UO_129 (O_129,N_13529,N_13977);
or UO_130 (O_130,N_12360,N_12865);
nand UO_131 (O_131,N_13978,N_14447);
and UO_132 (O_132,N_13184,N_14391);
or UO_133 (O_133,N_12562,N_13499);
nand UO_134 (O_134,N_13561,N_12079);
or UO_135 (O_135,N_14002,N_14854);
nand UO_136 (O_136,N_13914,N_14465);
nor UO_137 (O_137,N_13059,N_14424);
nand UO_138 (O_138,N_13476,N_12986);
nand UO_139 (O_139,N_13724,N_13493);
nand UO_140 (O_140,N_12459,N_12196);
xor UO_141 (O_141,N_14752,N_12486);
xnor UO_142 (O_142,N_14832,N_12021);
nand UO_143 (O_143,N_12886,N_14835);
nand UO_144 (O_144,N_13680,N_13708);
and UO_145 (O_145,N_12207,N_13890);
nor UO_146 (O_146,N_14717,N_12862);
or UO_147 (O_147,N_13288,N_14142);
nor UO_148 (O_148,N_13255,N_13975);
and UO_149 (O_149,N_12226,N_14336);
nor UO_150 (O_150,N_12112,N_14399);
nor UO_151 (O_151,N_14586,N_14765);
nand UO_152 (O_152,N_14071,N_13471);
nand UO_153 (O_153,N_12726,N_14613);
nand UO_154 (O_154,N_13799,N_14650);
or UO_155 (O_155,N_13289,N_14124);
nor UO_156 (O_156,N_13316,N_14910);
and UO_157 (O_157,N_13400,N_13895);
or UO_158 (O_158,N_12414,N_12090);
and UO_159 (O_159,N_12228,N_12299);
nor UO_160 (O_160,N_14543,N_12222);
and UO_161 (O_161,N_14792,N_12060);
or UO_162 (O_162,N_14324,N_13891);
nand UO_163 (O_163,N_12876,N_14896);
nor UO_164 (O_164,N_14048,N_14530);
and UO_165 (O_165,N_13360,N_13552);
or UO_166 (O_166,N_13941,N_13213);
xnor UO_167 (O_167,N_13688,N_14889);
nand UO_168 (O_168,N_12229,N_14032);
nand UO_169 (O_169,N_13500,N_13148);
or UO_170 (O_170,N_12418,N_12943);
nand UO_171 (O_171,N_12369,N_14331);
nand UO_172 (O_172,N_14086,N_14773);
and UO_173 (O_173,N_12348,N_13317);
and UO_174 (O_174,N_13315,N_13062);
and UO_175 (O_175,N_14814,N_14257);
and UO_176 (O_176,N_12604,N_12084);
xnor UO_177 (O_177,N_12390,N_12321);
and UO_178 (O_178,N_14747,N_12211);
and UO_179 (O_179,N_14128,N_13612);
and UO_180 (O_180,N_13960,N_12270);
nand UO_181 (O_181,N_12366,N_12528);
and UO_182 (O_182,N_13292,N_13242);
nand UO_183 (O_183,N_13809,N_13939);
nand UO_184 (O_184,N_13933,N_12100);
nor UO_185 (O_185,N_12826,N_14681);
xnor UO_186 (O_186,N_13085,N_13753);
xnor UO_187 (O_187,N_13501,N_13112);
or UO_188 (O_188,N_14801,N_12387);
xnor UO_189 (O_189,N_13284,N_14390);
xor UO_190 (O_190,N_13083,N_12630);
and UO_191 (O_191,N_14357,N_14267);
or UO_192 (O_192,N_12205,N_14076);
or UO_193 (O_193,N_12306,N_14621);
or UO_194 (O_194,N_12197,N_14963);
and UO_195 (O_195,N_12747,N_12289);
or UO_196 (O_196,N_13847,N_13582);
nand UO_197 (O_197,N_12224,N_12835);
and UO_198 (O_198,N_14947,N_14904);
and UO_199 (O_199,N_12263,N_14567);
and UO_200 (O_200,N_13586,N_13014);
and UO_201 (O_201,N_14359,N_13590);
nand UO_202 (O_202,N_14888,N_14540);
nor UO_203 (O_203,N_13735,N_13009);
xor UO_204 (O_204,N_14157,N_12692);
nand UO_205 (O_205,N_12098,N_13675);
xor UO_206 (O_206,N_14015,N_13828);
and UO_207 (O_207,N_14245,N_12576);
or UO_208 (O_208,N_12355,N_12452);
and UO_209 (O_209,N_13983,N_12616);
nand UO_210 (O_210,N_14075,N_13097);
and UO_211 (O_211,N_12731,N_14679);
or UO_212 (O_212,N_14605,N_13734);
nand UO_213 (O_213,N_14212,N_13326);
or UO_214 (O_214,N_14985,N_14193);
nor UO_215 (O_215,N_12336,N_12281);
nor UO_216 (O_216,N_13094,N_14364);
or UO_217 (O_217,N_12852,N_12613);
or UO_218 (O_218,N_14787,N_12230);
xor UO_219 (O_219,N_14365,N_12433);
or UO_220 (O_220,N_14303,N_13196);
or UO_221 (O_221,N_13915,N_14783);
nand UO_222 (O_222,N_12988,N_14492);
or UO_223 (O_223,N_14538,N_12667);
and UO_224 (O_224,N_14845,N_14028);
nand UO_225 (O_225,N_14882,N_12994);
or UO_226 (O_226,N_13905,N_14493);
nor UO_227 (O_227,N_12904,N_14982);
or UO_228 (O_228,N_14966,N_14817);
xor UO_229 (O_229,N_13102,N_13235);
or UO_230 (O_230,N_13952,N_14640);
and UO_231 (O_231,N_13523,N_14636);
xor UO_232 (O_232,N_14062,N_14903);
nor UO_233 (O_233,N_13543,N_12916);
or UO_234 (O_234,N_13547,N_12978);
or UO_235 (O_235,N_14848,N_13077);
and UO_236 (O_236,N_12940,N_13495);
nand UO_237 (O_237,N_14862,N_14126);
nor UO_238 (O_238,N_13984,N_12382);
nand UO_239 (O_239,N_12145,N_12279);
nor UO_240 (O_240,N_12579,N_13446);
nor UO_241 (O_241,N_13521,N_12082);
nor UO_242 (O_242,N_14800,N_13567);
or UO_243 (O_243,N_12900,N_13385);
nor UO_244 (O_244,N_14729,N_13445);
and UO_245 (O_245,N_14979,N_14769);
nand UO_246 (O_246,N_14667,N_12288);
xnor UO_247 (O_247,N_14130,N_13718);
or UO_248 (O_248,N_14956,N_13756);
nand UO_249 (O_249,N_12688,N_12467);
or UO_250 (O_250,N_13272,N_13862);
nor UO_251 (O_251,N_13796,N_13825);
and UO_252 (O_252,N_14881,N_13222);
nor UO_253 (O_253,N_14444,N_13957);
or UO_254 (O_254,N_14430,N_13979);
nor UO_255 (O_255,N_13490,N_12523);
nor UO_256 (O_256,N_13554,N_12739);
nor UO_257 (O_257,N_13275,N_13849);
nor UO_258 (O_258,N_12683,N_12219);
or UO_259 (O_259,N_14151,N_12440);
or UO_260 (O_260,N_12157,N_14440);
nand UO_261 (O_261,N_12640,N_12519);
nor UO_262 (O_262,N_12815,N_12913);
nor UO_263 (O_263,N_12052,N_12543);
nor UO_264 (O_264,N_12738,N_14866);
or UO_265 (O_265,N_13626,N_12681);
xor UO_266 (O_266,N_14579,N_14961);
or UO_267 (O_267,N_12349,N_13180);
and UO_268 (O_268,N_14252,N_13532);
nand UO_269 (O_269,N_13069,N_13909);
or UO_270 (O_270,N_12147,N_14595);
and UO_271 (O_271,N_12705,N_12095);
or UO_272 (O_272,N_12019,N_13576);
nand UO_273 (O_273,N_14016,N_13719);
nor UO_274 (O_274,N_12478,N_13945);
or UO_275 (O_275,N_12445,N_14408);
nand UO_276 (O_276,N_14131,N_14313);
and UO_277 (O_277,N_13026,N_12723);
and UO_278 (O_278,N_14095,N_12529);
nor UO_279 (O_279,N_14040,N_12092);
nor UO_280 (O_280,N_14475,N_13035);
nand UO_281 (O_281,N_12255,N_12393);
and UO_282 (O_282,N_12868,N_14268);
and UO_283 (O_283,N_14155,N_14826);
nor UO_284 (O_284,N_12819,N_14820);
nand UO_285 (O_285,N_14107,N_12806);
and UO_286 (O_286,N_12972,N_14373);
nand UO_287 (O_287,N_12989,N_12183);
and UO_288 (O_288,N_12173,N_13821);
nand UO_289 (O_289,N_12073,N_13555);
nor UO_290 (O_290,N_13782,N_13140);
nand UO_291 (O_291,N_12293,N_14137);
and UO_292 (O_292,N_14558,N_13473);
and UO_293 (O_293,N_12138,N_13283);
nand UO_294 (O_294,N_13605,N_14634);
nor UO_295 (O_295,N_13133,N_14784);
nor UO_296 (O_296,N_14818,N_14429);
nor UO_297 (O_297,N_13299,N_12967);
and UO_298 (O_298,N_13095,N_12014);
and UO_299 (O_299,N_14958,N_12323);
nor UO_300 (O_300,N_12062,N_13048);
nand UO_301 (O_301,N_14182,N_13568);
nor UO_302 (O_302,N_14527,N_14000);
and UO_303 (O_303,N_12834,N_12001);
xor UO_304 (O_304,N_13138,N_13301);
or UO_305 (O_305,N_13349,N_14066);
nand UO_306 (O_306,N_14805,N_12404);
and UO_307 (O_307,N_14811,N_12637);
or UO_308 (O_308,N_13182,N_14423);
and UO_309 (O_309,N_12471,N_13396);
nand UO_310 (O_310,N_13233,N_12845);
nor UO_311 (O_311,N_12328,N_14501);
nand UO_312 (O_312,N_12671,N_13266);
nand UO_313 (O_313,N_12857,N_14316);
nand UO_314 (O_314,N_14623,N_12782);
nor UO_315 (O_315,N_13306,N_13453);
and UO_316 (O_316,N_14225,N_12099);
and UO_317 (O_317,N_12812,N_13815);
or UO_318 (O_318,N_14946,N_12559);
nand UO_319 (O_319,N_13243,N_12011);
nand UO_320 (O_320,N_14535,N_12934);
or UO_321 (O_321,N_13099,N_13658);
nor UO_322 (O_322,N_14594,N_13550);
nor UO_323 (O_323,N_12653,N_14654);
nor UO_324 (O_324,N_13179,N_12143);
nand UO_325 (O_325,N_14203,N_13229);
nand UO_326 (O_326,N_13748,N_12480);
nor UO_327 (O_327,N_14645,N_12758);
nand UO_328 (O_328,N_14519,N_14046);
nor UO_329 (O_329,N_13417,N_14270);
nor UO_330 (O_330,N_14980,N_14256);
nand UO_331 (O_331,N_13540,N_14701);
xnor UO_332 (O_332,N_12606,N_14617);
nand UO_333 (O_333,N_13937,N_14144);
or UO_334 (O_334,N_13623,N_13236);
nand UO_335 (O_335,N_13281,N_12676);
or UO_336 (O_336,N_12745,N_13902);
nor UO_337 (O_337,N_12612,N_14894);
and UO_338 (O_338,N_13431,N_14153);
xnor UO_339 (O_339,N_14192,N_12055);
nor UO_340 (O_340,N_12434,N_13614);
xor UO_341 (O_341,N_12159,N_13487);
and UO_342 (O_342,N_13898,N_14973);
or UO_343 (O_343,N_13496,N_13882);
and UO_344 (O_344,N_13502,N_13723);
or UO_345 (O_345,N_13313,N_13434);
or UO_346 (O_346,N_12779,N_14473);
nand UO_347 (O_347,N_12632,N_14042);
nor UO_348 (O_348,N_14996,N_14426);
nor UO_349 (O_349,N_12995,N_14080);
nor UO_350 (O_350,N_13667,N_12939);
and UO_351 (O_351,N_14368,N_14547);
or UO_352 (O_352,N_13234,N_14104);
nand UO_353 (O_353,N_12206,N_12253);
or UO_354 (O_354,N_13263,N_14561);
or UO_355 (O_355,N_12771,N_12622);
or UO_356 (O_356,N_14656,N_12221);
nand UO_357 (O_357,N_14249,N_12016);
or UO_358 (O_358,N_14839,N_14581);
nor UO_359 (O_359,N_14965,N_14109);
or UO_360 (O_360,N_13956,N_12831);
nor UO_361 (O_361,N_13990,N_14034);
or UO_362 (O_362,N_13881,N_13468);
xnor UO_363 (O_363,N_13930,N_14689);
nor UO_364 (O_364,N_12557,N_13449);
nor UO_365 (O_365,N_13795,N_14385);
xnor UO_366 (O_366,N_14745,N_12937);
or UO_367 (O_367,N_12381,N_12957);
nand UO_368 (O_368,N_14384,N_13273);
nand UO_369 (O_369,N_14049,N_14960);
and UO_370 (O_370,N_14648,N_13203);
xor UO_371 (O_371,N_13447,N_12907);
nand UO_372 (O_372,N_12331,N_13443);
or UO_373 (O_373,N_14106,N_12575);
and UO_374 (O_374,N_14056,N_13730);
and UO_375 (O_375,N_14928,N_13985);
nor UO_376 (O_376,N_12423,N_14708);
xnor UO_377 (O_377,N_12912,N_14785);
and UO_378 (O_378,N_12372,N_12880);
nor UO_379 (O_379,N_12450,N_13402);
nand UO_380 (O_380,N_14850,N_14720);
or UO_381 (O_381,N_14394,N_13603);
nor UO_382 (O_382,N_12502,N_12897);
and UO_383 (O_383,N_14258,N_12441);
and UO_384 (O_384,N_13710,N_14565);
nor UO_385 (O_385,N_12477,N_12531);
nor UO_386 (O_386,N_14190,N_12649);
nor UO_387 (O_387,N_13149,N_13820);
nand UO_388 (O_388,N_12798,N_12615);
xor UO_389 (O_389,N_14698,N_12740);
and UO_390 (O_390,N_13257,N_13268);
and UO_391 (O_391,N_12827,N_12689);
nor UO_392 (O_392,N_14929,N_13157);
or UO_393 (O_393,N_14917,N_14378);
nand UO_394 (O_394,N_13207,N_14201);
nand UO_395 (O_395,N_14907,N_13001);
nand UO_396 (O_396,N_13042,N_14813);
nor UO_397 (O_397,N_12898,N_14312);
xnor UO_398 (O_398,N_14678,N_14140);
or UO_399 (O_399,N_13033,N_14932);
or UO_400 (O_400,N_13696,N_13465);
xor UO_401 (O_401,N_14999,N_14749);
xor UO_402 (O_402,N_14508,N_14367);
or UO_403 (O_403,N_14663,N_12357);
nor UO_404 (O_404,N_13625,N_13214);
nor UO_405 (O_405,N_13463,N_12454);
nor UO_406 (O_406,N_12672,N_12032);
or UO_407 (O_407,N_14990,N_14181);
nor UO_408 (O_408,N_14366,N_13995);
nor UO_409 (O_409,N_13093,N_14178);
xnor UO_410 (O_410,N_13139,N_12734);
and UO_411 (O_411,N_14962,N_13608);
or UO_412 (O_412,N_12924,N_14702);
nor UO_413 (O_413,N_13073,N_12192);
nor UO_414 (O_414,N_12796,N_13197);
or UO_415 (O_415,N_13110,N_12861);
nor UO_416 (O_416,N_14149,N_13976);
or UO_417 (O_417,N_14184,N_12151);
nand UO_418 (O_418,N_13972,N_14794);
or UO_419 (O_419,N_12058,N_12430);
and UO_420 (O_420,N_12461,N_12856);
xor UO_421 (O_421,N_12903,N_12674);
xor UO_422 (O_422,N_12189,N_14893);
and UO_423 (O_423,N_13712,N_13535);
and UO_424 (O_424,N_13019,N_14959);
nor UO_425 (O_425,N_14191,N_14931);
and UO_426 (O_426,N_13269,N_14224);
and UO_427 (O_427,N_12872,N_12936);
and UO_428 (O_428,N_13169,N_13556);
nor UO_429 (O_429,N_14230,N_13362);
and UO_430 (O_430,N_14529,N_13666);
nand UO_431 (O_431,N_13202,N_12706);
nor UO_432 (O_432,N_12506,N_13383);
nand UO_433 (O_433,N_12470,N_14975);
xnor UO_434 (O_434,N_12773,N_12314);
nor UO_435 (O_435,N_14864,N_12840);
xnor UO_436 (O_436,N_14734,N_12961);
and UO_437 (O_437,N_13030,N_14065);
nor UO_438 (O_438,N_13951,N_13505);
nand UO_439 (O_439,N_12757,N_12633);
and UO_440 (O_440,N_13147,N_12475);
nand UO_441 (O_441,N_13872,N_14139);
xor UO_442 (O_442,N_12376,N_14305);
nand UO_443 (O_443,N_12245,N_14349);
nor UO_444 (O_444,N_12029,N_13353);
nor UO_445 (O_445,N_13919,N_14500);
and UO_446 (O_446,N_12048,N_12325);
and UO_447 (O_447,N_12666,N_13657);
or UO_448 (O_448,N_13615,N_14326);
and UO_449 (O_449,N_13791,N_14715);
or UO_450 (O_450,N_13226,N_14057);
or UO_451 (O_451,N_13790,N_12074);
and UO_452 (O_452,N_13650,N_14951);
xor UO_453 (O_453,N_14480,N_12005);
or UO_454 (O_454,N_12617,N_13684);
and UO_455 (O_455,N_14274,N_14327);
nor UO_456 (O_456,N_14719,N_14463);
and UO_457 (O_457,N_13805,N_12030);
nor UO_458 (O_458,N_12709,N_14232);
or UO_459 (O_459,N_14302,N_13829);
nand UO_460 (O_460,N_14084,N_14993);
and UO_461 (O_461,N_12103,N_12783);
nor UO_462 (O_462,N_12356,N_12769);
nand UO_463 (O_463,N_14168,N_14496);
nand UO_464 (O_464,N_12169,N_13553);
xor UO_465 (O_465,N_13211,N_14926);
nand UO_466 (O_466,N_13282,N_14163);
xnor UO_467 (O_467,N_14670,N_14912);
nor UO_468 (O_468,N_13928,N_14936);
xor UO_469 (O_469,N_13144,N_13948);
and UO_470 (O_470,N_12123,N_12332);
nor UO_471 (O_471,N_14402,N_14819);
nand UO_472 (O_472,N_13717,N_14686);
nor UO_473 (O_473,N_14264,N_13906);
nor UO_474 (O_474,N_12054,N_12026);
nor UO_475 (O_475,N_12379,N_14945);
or UO_476 (O_476,N_14020,N_14639);
nor UO_477 (O_477,N_14011,N_13868);
xor UO_478 (O_478,N_12193,N_13368);
or UO_479 (O_479,N_12691,N_14886);
nor UO_480 (O_480,N_12577,N_13770);
nor UO_481 (O_481,N_13092,N_14593);
nor UO_482 (O_482,N_14050,N_12879);
or UO_483 (O_483,N_14770,N_14471);
xnor UO_484 (O_484,N_13163,N_14031);
nor UO_485 (O_485,N_14054,N_14531);
nor UO_486 (O_486,N_13918,N_13441);
nand UO_487 (O_487,N_13810,N_13806);
nand UO_488 (O_488,N_13607,N_13604);
nor UO_489 (O_489,N_12941,N_12539);
nand UO_490 (O_490,N_13044,N_12027);
or UO_491 (O_491,N_13037,N_13751);
or UO_492 (O_492,N_12954,N_12023);
nand UO_493 (O_493,N_12385,N_13061);
nand UO_494 (O_494,N_13433,N_13973);
or UO_495 (O_495,N_14575,N_12453);
nor UO_496 (O_496,N_14118,N_14214);
and UO_497 (O_497,N_13692,N_13715);
nand UO_498 (O_498,N_14343,N_13397);
or UO_499 (O_499,N_13423,N_13785);
nand UO_500 (O_500,N_13794,N_12620);
and UO_501 (O_501,N_13321,N_13889);
or UO_502 (O_502,N_12171,N_13296);
or UO_503 (O_503,N_13894,N_12490);
and UO_504 (O_504,N_14766,N_13338);
nor UO_505 (O_505,N_12918,N_12322);
and UO_506 (O_506,N_13006,N_14897);
nand UO_507 (O_507,N_12968,N_12252);
nor UO_508 (O_508,N_13798,N_13994);
and UO_509 (O_509,N_13811,N_14525);
nand UO_510 (O_510,N_12665,N_13792);
nand UO_511 (O_511,N_13072,N_14664);
nor UO_512 (O_512,N_14607,N_13057);
or UO_513 (O_513,N_13104,N_12128);
nand UO_514 (O_514,N_14620,N_13551);
and UO_515 (O_515,N_12344,N_13240);
and UO_516 (O_516,N_12069,N_13293);
nor UO_517 (O_517,N_12362,N_14294);
and UO_518 (O_518,N_13822,N_12346);
and UO_519 (O_519,N_12582,N_14563);
and UO_520 (O_520,N_14913,N_12491);
and UO_521 (O_521,N_14025,N_14700);
nor UO_522 (O_522,N_13218,N_14406);
nand UO_523 (O_523,N_12775,N_12951);
nor UO_524 (O_524,N_13549,N_12034);
nand UO_525 (O_525,N_13879,N_12776);
and UO_526 (O_526,N_13008,N_14393);
nor UO_527 (O_527,N_14604,N_13673);
or UO_528 (O_528,N_12096,N_13329);
and UO_529 (O_529,N_12334,N_14035);
or UO_530 (O_530,N_14560,N_13854);
or UO_531 (O_531,N_14351,N_13036);
and UO_532 (O_532,N_14166,N_14552);
nand UO_533 (O_533,N_12584,N_12500);
nand UO_534 (O_534,N_13377,N_14578);
and UO_535 (O_535,N_14370,N_12377);
or UO_536 (O_536,N_12424,N_12300);
and UO_537 (O_537,N_12618,N_12693);
and UO_538 (O_538,N_12624,N_13132);
nor UO_539 (O_539,N_12165,N_12824);
nand UO_540 (O_540,N_13412,N_12167);
or UO_541 (O_541,N_14314,N_12077);
nand UO_542 (O_542,N_12839,N_13425);
xor UO_543 (O_543,N_13461,N_13166);
nand UO_544 (O_544,N_12191,N_13781);
or UO_545 (O_545,N_12438,N_14459);
or UO_546 (O_546,N_14952,N_13314);
or UO_547 (O_547,N_12690,N_13507);
and UO_548 (O_548,N_14233,N_12553);
nand UO_549 (O_549,N_12154,N_14983);
nand UO_550 (O_550,N_12651,N_14713);
nand UO_551 (O_551,N_13841,N_13219);
nand UO_552 (O_552,N_14310,N_13969);
or UO_553 (O_553,N_12911,N_13787);
and UO_554 (O_554,N_14710,N_14793);
xnor UO_555 (O_555,N_12466,N_13459);
and UO_556 (O_556,N_13665,N_13005);
and UO_557 (O_557,N_13651,N_13228);
nand UO_558 (O_558,N_12524,N_12025);
nor UO_559 (O_559,N_14646,N_13034);
xor UO_560 (O_560,N_12287,N_12849);
and UO_561 (O_561,N_12698,N_12378);
nor UO_562 (O_562,N_13713,N_14063);
nand UO_563 (O_563,N_14461,N_12102);
or UO_564 (O_564,N_13720,N_14984);
and UO_565 (O_565,N_13826,N_12801);
or UO_566 (O_566,N_13359,N_12901);
or UO_567 (O_567,N_13738,N_12186);
nand UO_568 (O_568,N_13183,N_12662);
xnor UO_569 (O_569,N_14467,N_13729);
and UO_570 (O_570,N_13509,N_12124);
xor UO_571 (O_571,N_13047,N_14725);
nor UO_572 (O_572,N_14441,N_12233);
nor UO_573 (O_573,N_14344,N_13776);
and UO_574 (O_574,N_13388,N_13150);
or UO_575 (O_575,N_14748,N_14568);
and UO_576 (O_576,N_12597,N_14259);
nand UO_577 (O_577,N_13528,N_12574);
or UO_578 (O_578,N_13498,N_13803);
nor UO_579 (O_579,N_13420,N_12437);
nor UO_580 (O_580,N_14220,N_12109);
nand UO_581 (O_581,N_13901,N_13171);
and UO_582 (O_582,N_12699,N_13391);
nand UO_583 (O_583,N_13893,N_14774);
and UO_584 (O_584,N_13676,N_12512);
nand UO_585 (O_585,N_12347,N_12784);
nor UO_586 (O_586,N_13655,N_12902);
nor UO_587 (O_587,N_12541,N_13105);
nor UO_588 (O_588,N_12141,N_13611);
and UO_589 (O_589,N_14753,N_12772);
nand UO_590 (O_590,N_12735,N_12083);
nand UO_591 (O_591,N_13265,N_13950);
or UO_592 (O_592,N_12800,N_12131);
and UO_593 (O_593,N_14711,N_13662);
or UO_594 (O_594,N_12719,N_14788);
or UO_595 (O_595,N_14986,N_14867);
and UO_596 (O_596,N_14870,N_13745);
nand UO_597 (O_597,N_12647,N_13910);
and UO_598 (O_598,N_14275,N_12384);
or UO_599 (O_599,N_13253,N_14211);
nand UO_600 (O_600,N_12678,N_12022);
nand UO_601 (O_601,N_13697,N_12492);
and UO_602 (O_602,N_14549,N_14834);
and UO_603 (O_603,N_14798,N_14597);
nor UO_604 (O_604,N_12484,N_14925);
nor UO_605 (O_605,N_13290,N_13352);
and UO_606 (O_606,N_14342,N_13760);
xnor UO_607 (O_607,N_12590,N_14443);
nor UO_608 (O_608,N_14240,N_14550);
nor UO_609 (O_609,N_13965,N_12530);
or UO_610 (O_610,N_14685,N_12324);
xnor UO_611 (O_611,N_13303,N_14074);
or UO_612 (O_612,N_13871,N_12687);
and UO_613 (O_613,N_13661,N_13224);
and UO_614 (O_614,N_14436,N_14949);
xor UO_615 (O_615,N_14347,N_14055);
xor UO_616 (O_616,N_12271,N_12877);
xor UO_617 (O_617,N_14282,N_13920);
or UO_618 (O_618,N_14954,N_13970);
and UO_619 (O_619,N_12317,N_13393);
nand UO_620 (O_620,N_14013,N_13845);
nand UO_621 (O_621,N_13514,N_14059);
nor UO_622 (O_622,N_14466,N_13562);
xor UO_623 (O_623,N_12354,N_13833);
or UO_624 (O_624,N_14930,N_12724);
nor UO_625 (O_625,N_12449,N_14997);
or UO_626 (O_626,N_12754,N_14205);
nand UO_627 (O_627,N_14714,N_13262);
and UO_628 (O_628,N_12542,N_12750);
nand UO_629 (O_629,N_13244,N_13897);
or UO_630 (O_630,N_13426,N_14513);
nor UO_631 (O_631,N_13621,N_13379);
nor UO_632 (O_632,N_12926,N_13295);
nand UO_633 (O_633,N_14180,N_13935);
nand UO_634 (O_634,N_13421,N_14759);
nor UO_635 (O_635,N_12101,N_12514);
and UO_636 (O_636,N_13310,N_12144);
and UO_637 (O_637,N_14455,N_12659);
nand UO_638 (O_638,N_12535,N_13800);
and UO_639 (O_639,N_13633,N_12554);
or UO_640 (O_640,N_13700,N_12256);
and UO_641 (O_641,N_14566,N_13837);
nor UO_642 (O_642,N_12190,N_12673);
nand UO_643 (O_643,N_14577,N_13635);
or UO_644 (O_644,N_12974,N_14323);
and UO_645 (O_645,N_14877,N_14602);
and UO_646 (O_646,N_12752,N_12566);
nand UO_647 (O_647,N_12040,N_12540);
and UO_648 (O_648,N_12370,N_13107);
nor UO_649 (O_649,N_12339,N_12714);
xnor UO_650 (O_650,N_12254,N_12340);
and UO_651 (O_651,N_12125,N_13479);
or UO_652 (O_652,N_13230,N_13609);
and UO_653 (O_653,N_12277,N_14043);
nand UO_654 (O_654,N_14102,N_14521);
and UO_655 (O_655,N_14695,N_12307);
nor UO_656 (O_656,N_12993,N_14977);
nand UO_657 (O_657,N_14632,N_12234);
and UO_658 (O_658,N_13599,N_14914);
and UO_659 (O_659,N_12361,N_14570);
nor UO_660 (O_660,N_14998,N_14942);
or UO_661 (O_661,N_14721,N_14757);
and UO_662 (O_662,N_14994,N_12807);
nand UO_663 (O_663,N_12593,N_14038);
and UO_664 (O_664,N_14019,N_14281);
or UO_665 (O_665,N_14414,N_12854);
nand UO_666 (O_666,N_14703,N_12150);
xor UO_667 (O_667,N_14659,N_14842);
or UO_668 (O_668,N_12786,N_14456);
and UO_669 (O_669,N_14520,N_12627);
or UO_670 (O_670,N_12368,N_12405);
and UO_671 (O_671,N_14051,N_14401);
nand UO_672 (O_672,N_14271,N_13742);
nand UO_673 (O_673,N_14534,N_12712);
nand UO_674 (O_674,N_12805,N_14776);
nor UO_675 (O_675,N_12236,N_14216);
and UO_676 (O_676,N_13513,N_14442);
nand UO_677 (O_677,N_13530,N_14039);
nor UO_678 (O_678,N_13167,N_12586);
and UO_679 (O_679,N_14592,N_14450);
nand UO_680 (O_680,N_13689,N_14386);
or UO_681 (O_681,N_13118,N_12202);
nor UO_682 (O_682,N_14407,N_14810);
or UO_683 (O_683,N_12093,N_13869);
nor UO_684 (O_684,N_14601,N_12364);
and UO_685 (O_685,N_13726,N_12704);
nor UO_686 (O_686,N_14472,N_13068);
and UO_687 (O_687,N_14671,N_14388);
and UO_688 (O_688,N_14627,N_12187);
nand UO_689 (O_689,N_12581,N_13988);
or UO_690 (O_690,N_14021,N_14337);
and UO_691 (O_691,N_13823,N_13981);
xnor UO_692 (O_692,N_14298,N_13602);
xnor UO_693 (O_693,N_13405,N_14857);
nor UO_694 (O_694,N_13544,N_13594);
and UO_695 (O_695,N_12338,N_14981);
or UO_696 (O_696,N_12407,N_12718);
nand UO_697 (O_697,N_13653,N_13571);
nor UO_698 (O_698,N_12081,N_14510);
nor UO_699 (O_699,N_12890,N_13309);
nand UO_700 (O_700,N_13123,N_13707);
and UO_701 (O_701,N_12971,N_13108);
or UO_702 (O_702,N_13750,N_13032);
nor UO_703 (O_703,N_14006,N_13063);
xnor UO_704 (O_704,N_12213,N_13198);
or UO_705 (O_705,N_13237,N_13160);
and UO_706 (O_706,N_12049,N_12607);
and UO_707 (O_707,N_13830,N_13191);
nand UO_708 (O_708,N_13762,N_12711);
or UO_709 (O_709,N_14243,N_13758);
and UO_710 (O_710,N_13261,N_14791);
nor UO_711 (O_711,N_13460,N_12516);
and UO_712 (O_712,N_13636,N_14528);
and UO_713 (O_713,N_14416,N_12132);
or UO_714 (O_714,N_13966,N_14718);
or UO_715 (O_715,N_12297,N_12327);
or UO_716 (O_716,N_12122,N_14871);
nand UO_717 (O_717,N_12071,N_13474);
nor UO_718 (O_718,N_13856,N_12652);
nor UO_719 (O_719,N_12785,N_12351);
and UO_720 (O_720,N_12987,N_13081);
nand UO_721 (O_721,N_12031,N_14108);
nand UO_722 (O_722,N_14262,N_13020);
xor UO_723 (O_723,N_14113,N_12498);
nor UO_724 (O_724,N_14772,N_13596);
or UO_725 (O_725,N_14199,N_13041);
nor UO_726 (O_726,N_13174,N_12802);
and UO_727 (O_727,N_14033,N_12406);
nand UO_728 (O_728,N_14539,N_12950);
or UO_729 (O_729,N_14389,N_13201);
or UO_730 (O_730,N_12257,N_13217);
nand UO_731 (O_731,N_14273,N_14751);
and UO_732 (O_732,N_13126,N_14007);
nand UO_733 (O_733,N_14058,N_12549);
or UO_734 (O_734,N_12545,N_14895);
nand UO_735 (O_735,N_14900,N_14290);
nand UO_736 (O_736,N_13722,N_12425);
xnor UO_737 (O_737,N_14615,N_13477);
nand UO_738 (O_738,N_12345,N_12946);
nor UO_739 (O_739,N_14380,N_13071);
nand UO_740 (O_740,N_12696,N_12547);
or UO_741 (O_741,N_12959,N_14379);
or UO_742 (O_742,N_14352,N_13135);
nand UO_743 (O_743,N_14068,N_13374);
or UO_744 (O_744,N_12285,N_12392);
or UO_745 (O_745,N_13251,N_14827);
nand UO_746 (O_746,N_13892,N_13406);
nor UO_747 (O_747,N_14940,N_14484);
nor UO_748 (O_748,N_14196,N_13524);
nor UO_749 (O_749,N_13324,N_13511);
or UO_750 (O_750,N_12399,N_14194);
nor UO_751 (O_751,N_12463,N_14489);
and UO_752 (O_752,N_12464,N_14185);
xor UO_753 (O_753,N_14161,N_14545);
and UO_754 (O_754,N_13859,N_12007);
or UO_755 (O_755,N_12766,N_12133);
and UO_756 (O_756,N_14666,N_12208);
nand UO_757 (O_757,N_13591,N_14024);
or UO_758 (O_758,N_12743,N_12497);
and UO_759 (O_759,N_12059,N_13899);
and UO_760 (O_760,N_13807,N_13117);
or UO_761 (O_761,N_14957,N_13409);
nor UO_762 (O_762,N_12881,N_14129);
nor UO_763 (O_763,N_13319,N_13190);
nor UO_764 (O_764,N_14374,N_14723);
nor UO_765 (O_765,N_13154,N_12427);
or UO_766 (O_766,N_14120,N_13437);
or UO_767 (O_767,N_14164,N_14387);
or UO_768 (O_768,N_14919,N_14657);
and UO_769 (O_769,N_14200,N_12869);
nor UO_770 (O_770,N_14815,N_14927);
nor UO_771 (O_771,N_12018,N_14419);
nor UO_772 (O_772,N_13022,N_12403);
nor UO_773 (O_773,N_12227,N_13245);
xor UO_774 (O_774,N_12174,N_12629);
and UO_775 (O_775,N_13838,N_12822);
nand UO_776 (O_776,N_13404,N_13418);
nand UO_777 (O_777,N_13464,N_12534);
nor UO_778 (O_778,N_13091,N_14589);
xnor UO_779 (O_779,N_14988,N_13451);
nand UO_780 (O_780,N_14876,N_12874);
nor UO_781 (O_781,N_13390,N_14400);
nand UO_782 (O_782,N_13298,N_12009);
and UO_783 (O_783,N_13699,N_12468);
nor UO_784 (O_784,N_13286,N_14482);
nor UO_785 (O_785,N_12749,N_12755);
or UO_786 (O_786,N_13051,N_14093);
xor UO_787 (O_787,N_13536,N_13223);
and UO_788 (O_788,N_14227,N_13331);
xor UO_789 (O_789,N_13232,N_12225);
nor UO_790 (O_790,N_12451,N_13348);
nor UO_791 (O_791,N_13765,N_14223);
nand UO_792 (O_792,N_12568,N_13089);
or UO_793 (O_793,N_13834,N_12111);
and UO_794 (O_794,N_13581,N_12057);
or UO_795 (O_795,N_12684,N_12115);
or UO_796 (O_796,N_12682,N_13986);
or UO_797 (O_797,N_12546,N_14733);
xnor UO_798 (O_798,N_13786,N_12472);
nor UO_799 (O_799,N_12091,N_12761);
nand UO_800 (O_800,N_13870,N_14761);
nor UO_801 (O_801,N_13639,N_13070);
nand UO_802 (O_802,N_13386,N_13086);
and UO_803 (O_803,N_12292,N_14622);
nand UO_804 (O_804,N_12412,N_14026);
and UO_805 (O_805,N_12408,N_13137);
or UO_806 (O_806,N_14060,N_13569);
nand UO_807 (O_807,N_12804,N_14454);
nor UO_808 (O_808,N_14439,N_14653);
xor UO_809 (O_809,N_13278,N_13560);
and UO_810 (O_810,N_13074,N_13682);
nor UO_811 (O_811,N_14238,N_14699);
or UO_812 (O_812,N_12969,N_12024);
nand UO_813 (O_813,N_12817,N_12623);
nor UO_814 (O_814,N_13200,N_12922);
nor UO_815 (O_815,N_13208,N_14099);
xor UO_816 (O_816,N_14921,N_14458);
xor UO_817 (O_817,N_14684,N_13227);
or UO_818 (O_818,N_14255,N_13249);
and UO_819 (O_819,N_14110,N_12080);
nand UO_820 (O_820,N_12896,N_12038);
nor UO_821 (O_821,N_14825,N_14844);
nand UO_822 (O_822,N_14135,N_13067);
nor UO_823 (O_823,N_12268,N_14333);
or UO_824 (O_824,N_13589,N_14722);
xor UO_825 (O_825,N_13038,N_12481);
or UO_826 (O_826,N_13701,N_13597);
nor UO_827 (O_827,N_13472,N_13046);
nor UO_828 (O_828,N_13127,N_12126);
and UO_829 (O_829,N_13279,N_13155);
nand UO_830 (O_830,N_12850,N_14584);
nand UO_831 (O_831,N_12146,N_14582);
nand UO_832 (O_832,N_13982,N_12396);
nor UO_833 (O_833,N_13679,N_12895);
nand UO_834 (O_834,N_14278,N_12333);
or UO_835 (O_835,N_13737,N_14564);
or UO_836 (O_836,N_13343,N_12148);
and UO_837 (O_837,N_12595,N_14782);
and UO_838 (O_838,N_13857,N_12789);
or UO_839 (O_839,N_12727,N_13971);
nor UO_840 (O_840,N_14802,N_13294);
nor UO_841 (O_841,N_12686,N_13640);
xor UO_842 (O_842,N_13695,N_14300);
nor UO_843 (O_843,N_14600,N_13334);
or UO_844 (O_844,N_13271,N_14266);
or UO_845 (O_845,N_13176,N_14250);
nor UO_846 (O_846,N_13151,N_12130);
and UO_847 (O_847,N_13744,N_12517);
and UO_848 (O_848,N_14174,N_14001);
nor UO_849 (O_849,N_12415,N_13350);
nor UO_850 (O_850,N_12503,N_13055);
nand UO_851 (O_851,N_12127,N_14160);
xnor UO_852 (O_852,N_12702,N_14803);
nor UO_853 (O_853,N_14651,N_13013);
or UO_854 (O_854,N_14437,N_14234);
and UO_855 (O_855,N_13789,N_14969);
nor UO_856 (O_856,N_14739,N_13565);
or UO_857 (O_857,N_14081,N_12258);
nand UO_858 (O_858,N_14972,N_12864);
or UO_859 (O_859,N_12899,N_13486);
nor UO_860 (O_860,N_13678,N_12076);
or UO_861 (O_861,N_13613,N_13846);
and UO_862 (O_862,N_12394,N_12863);
and UO_863 (O_863,N_12400,N_14392);
or UO_864 (O_864,N_13389,N_12220);
xor UO_865 (O_865,N_13415,N_14410);
nor UO_866 (O_866,N_14304,N_14941);
or UO_867 (O_867,N_12722,N_12641);
nor UO_868 (O_868,N_14799,N_12035);
nand UO_869 (O_869,N_13333,N_13668);
nand UO_870 (O_870,N_12932,N_12286);
and UO_871 (O_871,N_13188,N_12045);
nand UO_872 (O_872,N_12283,N_13646);
or UO_873 (O_873,N_13403,N_12953);
nor UO_874 (O_874,N_12087,N_12302);
or UO_875 (O_875,N_12846,N_12310);
xnor UO_876 (O_876,N_14696,N_12658);
nand UO_877 (O_877,N_13000,N_12118);
nor UO_878 (O_878,N_14320,N_12457);
nor UO_879 (O_879,N_12611,N_12888);
nor UO_880 (O_880,N_14229,N_13900);
nor UO_881 (O_881,N_12563,N_13860);
nand UO_882 (O_882,N_13357,N_14008);
or UO_883 (O_883,N_14683,N_12697);
xnor UO_884 (O_884,N_13545,N_14334);
and UO_885 (O_885,N_14858,N_14328);
and UO_886 (O_886,N_14141,N_14674);
nand UO_887 (O_887,N_13302,N_14265);
nand UO_888 (O_888,N_12797,N_13356);
nor UO_889 (O_889,N_12028,N_13078);
nor UO_890 (O_890,N_12603,N_13579);
or UO_891 (O_891,N_14865,N_12908);
and UO_892 (O_892,N_13084,N_13997);
or UO_893 (O_893,N_12820,N_14176);
and UO_894 (O_894,N_13082,N_12767);
nor UO_895 (O_895,N_14533,N_14779);
nand UO_896 (O_896,N_13024,N_14730);
or UO_897 (O_897,N_12448,N_14923);
and UO_898 (O_898,N_12260,N_14911);
xor UO_899 (O_899,N_14829,N_12108);
xor UO_900 (O_900,N_14187,N_14875);
and UO_901 (O_901,N_13482,N_14272);
nor UO_902 (O_902,N_14123,N_13921);
and UO_903 (O_903,N_12335,N_13134);
and UO_904 (O_904,N_12716,N_13492);
or UO_905 (O_905,N_14955,N_13767);
nor UO_906 (O_906,N_14251,N_12583);
nand UO_907 (O_907,N_13181,N_12780);
or UO_908 (O_908,N_13076,N_12981);
and UO_909 (O_909,N_12556,N_12510);
and UO_910 (O_910,N_13638,N_14381);
nor UO_911 (O_911,N_12443,N_14434);
xor UO_912 (O_912,N_12239,N_14395);
nand UO_913 (O_913,N_14198,N_14138);
or UO_914 (O_914,N_14523,N_14286);
and UO_915 (O_915,N_14404,N_14569);
or UO_916 (O_916,N_12537,N_13079);
or UO_917 (O_917,N_13711,N_12139);
nor UO_918 (O_918,N_13346,N_12914);
or UO_919 (O_919,N_13764,N_13671);
nand UO_920 (O_920,N_14780,N_14609);
nand UO_921 (O_921,N_14005,N_12262);
nor UO_922 (O_922,N_14427,N_12532);
nand UO_923 (O_923,N_12956,N_14778);
xnor UO_924 (O_924,N_13131,N_12178);
xor UO_925 (O_925,N_14536,N_12621);
nor UO_926 (O_926,N_14415,N_14083);
or UO_927 (O_927,N_13618,N_14052);
and UO_928 (O_928,N_14449,N_12695);
or UO_929 (O_929,N_13987,N_12214);
and UO_930 (O_930,N_13398,N_12567);
or UO_931 (O_931,N_14322,N_12920);
and UO_932 (O_932,N_12097,N_14078);
and UO_933 (O_933,N_13100,N_13949);
or UO_934 (O_934,N_13878,N_13335);
and UO_935 (O_935,N_13998,N_13136);
nor UO_936 (O_936,N_14092,N_13080);
nor UO_937 (O_937,N_14348,N_13814);
and UO_938 (O_938,N_13021,N_14167);
xor UO_939 (O_939,N_13775,N_13757);
nand UO_940 (O_940,N_14874,N_13246);
xnor UO_941 (O_941,N_14795,N_14494);
nor UO_942 (O_942,N_14162,N_14908);
and UO_943 (O_943,N_14125,N_14165);
and UO_944 (O_944,N_13470,N_12701);
and UO_945 (O_945,N_14177,N_14731);
nor UO_946 (O_946,N_14611,N_14027);
or UO_947 (O_947,N_13755,N_13165);
nand UO_948 (O_948,N_14079,N_13239);
and UO_949 (O_949,N_13908,N_14353);
or UO_950 (O_950,N_13842,N_14464);
nand UO_951 (O_951,N_13548,N_13534);
xor UO_952 (O_952,N_12352,N_12386);
nand UO_953 (O_953,N_14544,N_13311);
or UO_954 (O_954,N_13158,N_12487);
and UO_955 (O_955,N_13225,N_13539);
and UO_956 (O_956,N_13336,N_13168);
nor UO_957 (O_957,N_13370,N_14396);
nor UO_958 (O_958,N_14146,N_13448);
nor UO_959 (O_959,N_12039,N_12215);
nor UO_960 (O_960,N_14433,N_14460);
and UO_961 (O_961,N_13351,N_12044);
or UO_962 (O_962,N_13885,N_14219);
nand UO_963 (O_963,N_12507,N_13300);
nand UO_964 (O_964,N_12436,N_12442);
nand UO_965 (O_965,N_13488,N_12813);
nor UO_966 (O_966,N_13210,N_14105);
or UO_967 (O_967,N_14808,N_13574);
and UO_968 (O_968,N_14879,N_14360);
nor UO_969 (O_969,N_14490,N_14497);
xor UO_970 (O_970,N_14728,N_12495);
and UO_971 (O_971,N_13531,N_14301);
and UO_972 (O_972,N_12713,N_14487);
xor UO_973 (O_973,N_12626,N_14405);
xor UO_974 (O_974,N_14989,N_12803);
nand UO_975 (O_975,N_12421,N_12342);
and UO_976 (O_976,N_12318,N_14295);
and UO_977 (O_977,N_13015,N_14939);
or UO_978 (O_978,N_13216,N_14210);
nor UO_979 (O_979,N_13436,N_12909);
nor UO_980 (O_980,N_13677,N_14716);
nor UO_981 (O_981,N_13252,N_12645);
nand UO_982 (O_982,N_14309,N_14970);
nand UO_983 (O_983,N_13876,N_12708);
nor UO_984 (O_984,N_13944,N_12844);
nor UO_985 (O_985,N_13706,N_12276);
nand UO_986 (O_986,N_12374,N_12929);
and UO_987 (O_987,N_14156,N_12244);
nand UO_988 (O_988,N_13649,N_13371);
or UO_989 (O_989,N_13772,N_13573);
or UO_990 (O_990,N_12163,N_12661);
and UO_991 (O_991,N_12110,N_13570);
nand UO_992 (O_992,N_12625,N_13510);
or UO_993 (O_993,N_14096,N_13355);
xor UO_994 (O_994,N_12536,N_13205);
xnor UO_995 (O_995,N_12591,N_13291);
or UO_996 (O_996,N_12675,N_13267);
and UO_997 (O_997,N_14237,N_12952);
nand UO_998 (O_998,N_13380,N_12156);
nand UO_999 (O_999,N_12664,N_12114);
and UO_1000 (O_1000,N_14987,N_12838);
or UO_1001 (O_1001,N_14175,N_12760);
or UO_1002 (O_1002,N_13416,N_14100);
nor UO_1003 (O_1003,N_13494,N_14338);
and UO_1004 (O_1004,N_14481,N_14922);
nand UO_1005 (O_1005,N_14572,N_13025);
nand UO_1006 (O_1006,N_13129,N_12273);
nor UO_1007 (O_1007,N_14242,N_13414);
nor UO_1008 (O_1008,N_12729,N_13992);
nand UO_1009 (O_1009,N_12509,N_14868);
nor UO_1010 (O_1010,N_13358,N_13903);
nor UO_1011 (O_1011,N_14548,N_14762);
nor UO_1012 (O_1012,N_13557,N_12859);
nand UO_1013 (O_1013,N_14809,N_14629);
xnor UO_1014 (O_1014,N_13922,N_14346);
and UO_1015 (O_1015,N_13912,N_13832);
nand UO_1016 (O_1016,N_12842,N_14088);
and UO_1017 (O_1017,N_12882,N_13739);
and UO_1018 (O_1018,N_13090,N_13247);
nor UO_1019 (O_1019,N_12161,N_14691);
xor UO_1020 (O_1020,N_12373,N_12884);
or UO_1021 (O_1021,N_12966,N_12106);
nand UO_1022 (O_1022,N_13664,N_13342);
or UO_1023 (O_1023,N_12493,N_14483);
nor UO_1024 (O_1024,N_13159,N_12976);
nor UO_1025 (O_1025,N_14291,N_12180);
and UO_1026 (O_1026,N_14277,N_12367);
or UO_1027 (O_1027,N_13325,N_14111);
or UO_1028 (O_1028,N_13693,N_12068);
xnor UO_1029 (O_1029,N_12275,N_12462);
or UO_1030 (O_1030,N_14682,N_12598);
and UO_1031 (O_1031,N_13002,N_12274);
nor UO_1032 (O_1032,N_12003,N_12496);
nand UO_1033 (O_1033,N_12791,N_13974);
nand UO_1034 (O_1034,N_12238,N_13520);
nand UO_1035 (O_1035,N_14041,N_13111);
nor UO_1036 (O_1036,N_13843,N_14116);
or UO_1037 (O_1037,N_12588,N_13522);
nand UO_1038 (O_1038,N_13410,N_13106);
and UO_1039 (O_1039,N_13363,N_14279);
or UO_1040 (O_1040,N_12685,N_12736);
xor UO_1041 (O_1041,N_12814,N_14195);
nor UO_1042 (O_1042,N_14292,N_12958);
and UO_1043 (O_1043,N_12089,N_13156);
or UO_1044 (O_1044,N_14445,N_14293);
nor UO_1045 (O_1045,N_12061,N_12316);
xnor UO_1046 (O_1046,N_13672,N_12237);
xor UO_1047 (O_1047,N_13430,N_14849);
or UO_1048 (O_1048,N_12513,N_12358);
nor UO_1049 (O_1049,N_14308,N_13587);
or UO_1050 (O_1050,N_13277,N_14836);
and UO_1051 (O_1051,N_12548,N_14902);
nor UO_1052 (O_1052,N_12176,N_12764);
or UO_1053 (O_1053,N_13194,N_14953);
nand UO_1054 (O_1054,N_12928,N_14261);
or UO_1055 (O_1055,N_13780,N_13801);
nor UO_1056 (O_1056,N_13875,N_14976);
or UO_1057 (O_1057,N_14159,N_12181);
nand UO_1058 (O_1058,N_13489,N_13087);
nand UO_1059 (O_1059,N_13874,N_13773);
xnor UO_1060 (O_1060,N_13546,N_13345);
nor UO_1061 (O_1061,N_12520,N_13804);
and UO_1062 (O_1062,N_12251,N_14526);
or UO_1063 (O_1063,N_14169,N_14446);
and UO_1064 (O_1064,N_12088,N_12636);
or UO_1065 (O_1065,N_13703,N_14115);
xor UO_1066 (O_1066,N_13779,N_12184);
or UO_1067 (O_1067,N_13125,N_13934);
and UO_1068 (O_1068,N_14588,N_12551);
or UO_1069 (O_1069,N_12010,N_12298);
and UO_1070 (O_1070,N_14767,N_14288);
and UO_1071 (O_1071,N_14974,N_13011);
or UO_1072 (O_1072,N_12383,N_12601);
nor UO_1073 (O_1073,N_12067,N_13049);
and UO_1074 (O_1074,N_12892,N_14786);
and UO_1075 (O_1075,N_12343,N_12858);
and UO_1076 (O_1076,N_13212,N_14197);
nand UO_1077 (O_1077,N_14114,N_12413);
xnor UO_1078 (O_1078,N_13517,N_13456);
nor UO_1079 (O_1079,N_13119,N_12533);
xnor UO_1080 (O_1080,N_13043,N_12763);
nand UO_1081 (O_1081,N_14892,N_12992);
and UO_1082 (O_1082,N_12999,N_14476);
nor UO_1083 (O_1083,N_13731,N_14694);
or UO_1084 (O_1084,N_14880,N_14756);
and UO_1085 (O_1085,N_13066,N_13999);
nor UO_1086 (O_1086,N_13045,N_14003);
or UO_1087 (O_1087,N_12587,N_14777);
or UO_1088 (O_1088,N_14909,N_14094);
xnor UO_1089 (O_1089,N_14992,N_13968);
or UO_1090 (O_1090,N_12295,N_14576);
and UO_1091 (O_1091,N_13485,N_14542);
nand UO_1092 (O_1092,N_12063,N_12930);
xnor UO_1093 (O_1093,N_13863,N_13260);
or UO_1094 (O_1094,N_13583,N_14147);
nand UO_1095 (O_1095,N_14372,N_13768);
nor UO_1096 (O_1096,N_13769,N_14283);
nand UO_1097 (O_1097,N_12923,N_13469);
and UO_1098 (O_1098,N_13619,N_12218);
nor UO_1099 (O_1099,N_13475,N_12409);
and UO_1100 (O_1100,N_13942,N_12149);
or UO_1101 (O_1101,N_13542,N_13122);
nand UO_1102 (O_1102,N_13774,N_14260);
nor UO_1103 (O_1103,N_13192,N_12732);
or UO_1104 (O_1104,N_12809,N_12479);
and UO_1105 (O_1105,N_14633,N_13384);
xor UO_1106 (O_1106,N_14179,N_12085);
or UO_1107 (O_1107,N_13442,N_13883);
nor UO_1108 (O_1108,N_13185,N_12066);
and UO_1109 (O_1109,N_13504,N_13564);
nor UO_1110 (O_1110,N_14630,N_14209);
and UO_1111 (O_1111,N_14218,N_12465);
nand UO_1112 (O_1112,N_13818,N_14840);
nor UO_1113 (O_1113,N_13601,N_12639);
xnor UO_1114 (O_1114,N_14873,N_12428);
and UO_1115 (O_1115,N_13378,N_13483);
or UO_1116 (O_1116,N_12305,N_12065);
and UO_1117 (O_1117,N_13088,N_14610);
nor UO_1118 (O_1118,N_14585,N_13178);
or UO_1119 (O_1119,N_12781,N_14603);
and UO_1120 (O_1120,N_12246,N_12499);
and UO_1121 (O_1121,N_12663,N_13652);
and UO_1122 (O_1122,N_14557,N_14517);
or UO_1123 (O_1123,N_13575,N_12494);
and UO_1124 (O_1124,N_14358,N_13209);
nand UO_1125 (O_1125,N_13778,N_14488);
nor UO_1126 (O_1126,N_12525,N_14841);
nor UO_1127 (O_1127,N_13369,N_13698);
xor UO_1128 (O_1128,N_12140,N_14010);
or UO_1129 (O_1129,N_14853,N_14417);
nand UO_1130 (O_1130,N_13752,N_14618);
or UO_1131 (O_1131,N_12474,N_12439);
and UO_1132 (O_1132,N_12915,N_13480);
nand UO_1133 (O_1133,N_12301,N_13259);
and UO_1134 (O_1134,N_12759,N_14246);
and UO_1135 (O_1135,N_14647,N_13702);
and UO_1136 (O_1136,N_14938,N_13040);
and UO_1137 (O_1137,N_12249,N_14971);
or UO_1138 (O_1138,N_12175,N_14514);
nand UO_1139 (O_1139,N_12280,N_12998);
nand UO_1140 (O_1140,N_12572,N_12216);
or UO_1141 (O_1141,N_13120,N_14217);
and UO_1142 (O_1142,N_14891,N_14732);
nand UO_1143 (O_1143,N_14658,N_12319);
nand UO_1144 (O_1144,N_13629,N_13641);
xnor UO_1145 (O_1145,N_12363,N_13375);
or UO_1146 (O_1146,N_13991,N_13907);
nor UO_1147 (O_1147,N_13690,N_12195);
nor UO_1148 (O_1148,N_12680,N_12580);
and UO_1149 (O_1149,N_12555,N_14967);
nand UO_1150 (O_1150,N_13929,N_14241);
xor UO_1151 (O_1151,N_12947,N_14047);
and UO_1152 (O_1152,N_12209,N_14950);
or UO_1153 (O_1153,N_14421,N_14044);
nand UO_1154 (O_1154,N_13193,N_13851);
xor UO_1155 (O_1155,N_14524,N_14742);
nor UO_1156 (O_1156,N_12720,N_13142);
and UO_1157 (O_1157,N_13852,N_14590);
or UO_1158 (O_1158,N_12422,N_12836);
or UO_1159 (O_1159,N_12980,N_12770);
nand UO_1160 (O_1160,N_12137,N_13598);
and UO_1161 (O_1161,N_12473,N_12655);
or UO_1162 (O_1162,N_12303,N_12511);
or UO_1163 (O_1163,N_13736,N_13627);
and UO_1164 (O_1164,N_13427,N_13759);
or UO_1165 (O_1165,N_14171,N_13518);
nor UO_1166 (O_1166,N_13258,N_13669);
and UO_1167 (O_1167,N_14823,N_12518);
or UO_1168 (O_1168,N_14097,N_13931);
nor UO_1169 (O_1169,N_13462,N_12168);
xnor UO_1170 (O_1170,N_14098,N_14136);
nor UO_1171 (O_1171,N_14215,N_12848);
and UO_1172 (O_1172,N_13075,N_12359);
nor UO_1173 (O_1173,N_13631,N_14690);
or UO_1174 (O_1174,N_13128,N_12558);
nor UO_1175 (O_1175,N_14649,N_14479);
and UO_1176 (O_1176,N_14418,N_13927);
or UO_1177 (O_1177,N_12841,N_14369);
nand UO_1178 (O_1178,N_12326,N_12117);
nor UO_1179 (O_1179,N_12643,N_12860);
or UO_1180 (O_1180,N_12185,N_14608);
nand UO_1181 (O_1181,N_13058,N_13466);
and UO_1182 (O_1182,N_14134,N_12573);
or UO_1183 (O_1183,N_12282,N_14755);
nand UO_1184 (O_1184,N_12294,N_12248);
and UO_1185 (O_1185,N_14188,N_13888);
or UO_1186 (O_1186,N_14030,N_13663);
nor UO_1187 (O_1187,N_13422,N_13141);
xnor UO_1188 (O_1188,N_13130,N_12715);
or UO_1189 (O_1189,N_13831,N_13161);
and UO_1190 (O_1190,N_12610,N_13364);
and UO_1191 (O_1191,N_13606,N_14420);
and UO_1192 (O_1192,N_12105,N_12008);
nand UO_1193 (O_1193,N_14319,N_13962);
or UO_1194 (O_1194,N_12419,N_14206);
or UO_1195 (O_1195,N_13124,N_12847);
or UO_1196 (O_1196,N_14553,N_14280);
nor UO_1197 (O_1197,N_12158,N_13685);
and UO_1198 (O_1198,N_12043,N_13714);
or UO_1199 (O_1199,N_12485,N_13238);
and UO_1200 (O_1200,N_14743,N_14641);
nor UO_1201 (O_1201,N_12121,N_14598);
nand UO_1202 (O_1202,N_12721,N_12505);
and UO_1203 (O_1203,N_12046,N_13537);
or UO_1204 (O_1204,N_12657,N_14596);
and UO_1205 (O_1205,N_14727,N_13634);
nor UO_1206 (O_1206,N_14642,N_12867);
nand UO_1207 (O_1207,N_13274,N_12201);
nand UO_1208 (O_1208,N_14361,N_13458);
and UO_1209 (O_1209,N_13394,N_12935);
nor UO_1210 (O_1210,N_12265,N_12707);
nor UO_1211 (O_1211,N_13993,N_13381);
and UO_1212 (O_1212,N_12164,N_14061);
or UO_1213 (O_1213,N_13659,N_13578);
nor UO_1214 (O_1214,N_14991,N_12793);
nand UO_1215 (O_1215,N_13280,N_13438);
nand UO_1216 (O_1216,N_14254,N_13955);
xnor UO_1217 (O_1217,N_14860,N_13855);
nor UO_1218 (O_1218,N_12837,N_12521);
nor UO_1219 (O_1219,N_12594,N_14468);
nand UO_1220 (O_1220,N_14754,N_13432);
nor UO_1221 (O_1221,N_14189,N_14705);
xnor UO_1222 (O_1222,N_13516,N_12119);
xor UO_1223 (O_1223,N_12037,N_12402);
or UO_1224 (O_1224,N_14843,N_12460);
xnor UO_1225 (O_1225,N_14655,N_13399);
or UO_1226 (O_1226,N_13559,N_14872);
and UO_1227 (O_1227,N_13254,N_13028);
nor UO_1228 (O_1228,N_13367,N_14509);
or UO_1229 (O_1229,N_14978,N_12391);
or UO_1230 (O_1230,N_13452,N_12944);
and UO_1231 (O_1231,N_13617,N_13387);
nand UO_1232 (O_1232,N_12544,N_13746);
nor UO_1233 (O_1233,N_14943,N_12398);
nor UO_1234 (O_1234,N_13187,N_12614);
nand UO_1235 (O_1235,N_13728,N_12247);
xnor UO_1236 (O_1236,N_14847,N_13098);
xor UO_1237 (O_1237,N_13428,N_14023);
nand UO_1238 (O_1238,N_13648,N_13808);
and UO_1239 (O_1239,N_14885,N_14186);
or UO_1240 (O_1240,N_13642,N_14121);
or UO_1241 (O_1241,N_13344,N_13964);
nor UO_1242 (O_1242,N_12188,N_13566);
nand UO_1243 (O_1243,N_13839,N_12051);
nor UO_1244 (O_1244,N_12020,N_13491);
nor UO_1245 (O_1245,N_14101,N_14571);
nand UO_1246 (O_1246,N_14562,N_12810);
xnor UO_1247 (O_1247,N_14285,N_12056);
nor UO_1248 (O_1248,N_13304,N_14644);
nor UO_1249 (O_1249,N_12561,N_12337);
xnor UO_1250 (O_1250,N_13533,N_14626);
or UO_1251 (O_1251,N_14350,N_14411);
or UO_1252 (O_1252,N_13816,N_14307);
nor UO_1253 (O_1253,N_12748,N_12033);
nor UO_1254 (O_1254,N_14587,N_14807);
nor UO_1255 (O_1255,N_14453,N_13484);
nand UO_1256 (O_1256,N_12550,N_13376);
and UO_1257 (O_1257,N_13681,N_12341);
xnor UO_1258 (O_1258,N_13340,N_12526);
nand UO_1259 (O_1259,N_12816,N_14133);
nor UO_1260 (O_1260,N_14631,N_13115);
nor UO_1261 (O_1261,N_13395,N_12329);
nor UO_1262 (O_1262,N_12893,N_14375);
xnor UO_1263 (O_1263,N_14736,N_12050);
nor UO_1264 (O_1264,N_13896,N_13959);
and UO_1265 (O_1265,N_12585,N_13439);
xor UO_1266 (O_1266,N_13858,N_14863);
xnor UO_1267 (O_1267,N_14660,N_12179);
nand UO_1268 (O_1268,N_14915,N_13592);
and UO_1269 (O_1269,N_12600,N_13256);
or UO_1270 (O_1270,N_12241,N_12677);
and UO_1271 (O_1271,N_14036,N_14797);
xnor UO_1272 (O_1272,N_14838,N_12742);
nand UO_1273 (O_1273,N_14709,N_14675);
nor UO_1274 (O_1274,N_14462,N_12694);
nand UO_1275 (O_1275,N_14037,N_13610);
nor UO_1276 (O_1276,N_12571,N_12975);
or UO_1277 (O_1277,N_14637,N_12906);
or UO_1278 (O_1278,N_12064,N_13401);
or UO_1279 (O_1279,N_14425,N_14737);
nand UO_1280 (O_1280,N_12308,N_12808);
and UO_1281 (O_1281,N_12501,N_13114);
xor UO_1282 (O_1282,N_12931,N_14325);
or UO_1283 (O_1283,N_14824,N_14771);
xor UO_1284 (O_1284,N_13113,N_13285);
xor UO_1285 (O_1285,N_13632,N_13250);
and UO_1286 (O_1286,N_14228,N_12476);
or UO_1287 (O_1287,N_12231,N_13865);
nor UO_1288 (O_1288,N_13153,N_14546);
nor UO_1289 (O_1289,N_13064,N_13873);
nand UO_1290 (O_1290,N_13620,N_12631);
and UO_1291 (O_1291,N_12426,N_14398);
or UO_1292 (O_1292,N_14231,N_12380);
nand UO_1293 (O_1293,N_12948,N_14859);
nand UO_1294 (O_1294,N_12235,N_12753);
and UO_1295 (O_1295,N_14363,N_12596);
and UO_1296 (O_1296,N_14009,N_13109);
nor UO_1297 (O_1297,N_12410,N_14017);
xnor UO_1298 (O_1298,N_12654,N_12609);
and UO_1299 (O_1299,N_12455,N_14332);
or UO_1300 (O_1300,N_14477,N_13173);
nand UO_1301 (O_1301,N_13012,N_13050);
or UO_1302 (O_1302,N_12921,N_13911);
xnor UO_1303 (O_1303,N_14469,N_13904);
nor UO_1304 (O_1304,N_14172,N_14306);
and UO_1305 (O_1305,N_13347,N_13705);
xnor UO_1306 (O_1306,N_13172,N_13940);
xor UO_1307 (O_1307,N_14668,N_13003);
nor UO_1308 (O_1308,N_13152,N_13264);
nand UO_1309 (O_1309,N_12866,N_13916);
and UO_1310 (O_1310,N_13563,N_12203);
nor UO_1311 (O_1311,N_13497,N_12264);
and UO_1312 (O_1312,N_14317,N_13175);
nor UO_1313 (O_1313,N_12883,N_13199);
or UO_1314 (O_1314,N_12635,N_14119);
nand UO_1315 (O_1315,N_14064,N_13372);
nor UO_1316 (O_1316,N_14673,N_13503);
nor UO_1317 (O_1317,N_12411,N_12818);
nand UO_1318 (O_1318,N_13877,N_13867);
or UO_1319 (O_1319,N_14382,N_12242);
xnor UO_1320 (O_1320,N_12395,N_12508);
and UO_1321 (O_1321,N_12504,N_13341);
nand UO_1322 (O_1322,N_13248,N_14069);
nand UO_1323 (O_1323,N_12006,N_12116);
and UO_1324 (O_1324,N_14158,N_14944);
or UO_1325 (O_1325,N_12004,N_12152);
nand UO_1326 (O_1326,N_12104,N_12765);
nand UO_1327 (O_1327,N_13429,N_14516);
or UO_1328 (O_1328,N_12744,N_14207);
nor UO_1329 (O_1329,N_12134,N_13725);
and UO_1330 (O_1330,N_14554,N_12036);
and UO_1331 (O_1331,N_12538,N_13886);
and UO_1332 (O_1332,N_13732,N_14591);
nor UO_1333 (O_1333,N_14090,N_12047);
xor UO_1334 (O_1334,N_14085,N_13170);
xnor UO_1335 (O_1335,N_12778,N_14431);
nand UO_1336 (O_1336,N_13980,N_12527);
nor UO_1337 (O_1337,N_13440,N_14672);
nor UO_1338 (O_1338,N_14559,N_14661);
nor UO_1339 (O_1339,N_14764,N_14532);
and UO_1340 (O_1340,N_13953,N_12243);
nor UO_1341 (O_1341,N_14758,N_14937);
nor UO_1342 (O_1342,N_13645,N_14884);
or UO_1343 (O_1343,N_13802,N_13053);
nand UO_1344 (O_1344,N_14435,N_12979);
xnor UO_1345 (O_1345,N_14573,N_13819);
nand UO_1346 (O_1346,N_12843,N_13408);
nand UO_1347 (O_1347,N_14556,N_14898);
nor UO_1348 (O_1348,N_14452,N_13478);
and UO_1349 (O_1349,N_14781,N_14515);
nor UO_1350 (O_1350,N_12634,N_13231);
or UO_1351 (O_1351,N_12432,N_12873);
or UO_1352 (O_1352,N_14498,N_12153);
nor UO_1353 (O_1353,N_14852,N_12094);
xnor UO_1354 (O_1354,N_12855,N_12656);
nand UO_1355 (O_1355,N_14330,N_12365);
nor UO_1356 (O_1356,N_13836,N_14018);
or UO_1357 (O_1357,N_12853,N_14856);
nand UO_1358 (O_1358,N_13793,N_14253);
xor UO_1359 (O_1359,N_13683,N_12569);
and UO_1360 (O_1360,N_14833,N_14339);
nand UO_1361 (O_1361,N_13763,N_12973);
and UO_1362 (O_1362,N_14485,N_12304);
xnor UO_1363 (O_1363,N_14746,N_12829);
or UO_1364 (O_1364,N_14239,N_14356);
and UO_1365 (O_1365,N_12388,N_13023);
nand UO_1366 (O_1366,N_12792,N_14495);
and UO_1367 (O_1367,N_14851,N_12870);
nand UO_1368 (O_1368,N_12489,N_13039);
nor UO_1369 (O_1369,N_13506,N_13946);
or UO_1370 (O_1370,N_14409,N_13444);
nor UO_1371 (O_1371,N_12942,N_12794);
nand UO_1372 (O_1372,N_12012,N_14890);
and UO_1373 (O_1373,N_13687,N_12017);
nor UO_1374 (O_1374,N_14518,N_13007);
or UO_1375 (O_1375,N_12389,N_12170);
xnor UO_1376 (O_1376,N_13143,N_14247);
nand UO_1377 (O_1377,N_13327,N_13880);
xor UO_1378 (O_1378,N_13600,N_13932);
nand UO_1379 (O_1379,N_13052,N_12945);
xor UO_1380 (O_1380,N_14173,N_13297);
and UO_1381 (O_1381,N_13096,N_14861);
xnor UO_1382 (O_1382,N_12313,N_13525);
nor UO_1383 (O_1383,N_14376,N_14235);
or UO_1384 (O_1384,N_12833,N_14612);
or UO_1385 (O_1385,N_14087,N_14638);
or UO_1386 (O_1386,N_14412,N_12267);
nor UO_1387 (O_1387,N_13694,N_13924);
nand UO_1388 (O_1388,N_13029,N_14112);
or UO_1389 (O_1389,N_14665,N_13670);
or UO_1390 (O_1390,N_12564,N_14738);
nor UO_1391 (O_1391,N_14707,N_13741);
and UO_1392 (O_1392,N_13558,N_14236);
or UO_1393 (O_1393,N_12910,N_13588);
nor UO_1394 (O_1394,N_13455,N_14555);
or UO_1395 (O_1395,N_13366,N_14806);
and UO_1396 (O_1396,N_13519,N_14297);
nor UO_1397 (O_1397,N_13189,N_13840);
or UO_1398 (O_1398,N_13177,N_13947);
or UO_1399 (O_1399,N_13060,N_14831);
nand UO_1400 (O_1400,N_14677,N_14676);
and UO_1401 (O_1401,N_12977,N_13287);
and UO_1402 (O_1402,N_12644,N_14918);
and UO_1403 (O_1403,N_14796,N_14457);
nand UO_1404 (O_1404,N_12204,N_14335);
or UO_1405 (O_1405,N_12768,N_14804);
or UO_1406 (O_1406,N_13195,N_13630);
nor UO_1407 (O_1407,N_12964,N_13407);
or UO_1408 (O_1408,N_12589,N_14760);
nor UO_1409 (O_1409,N_12578,N_14448);
nand UO_1410 (O_1410,N_14692,N_12985);
or UO_1411 (O_1411,N_12592,N_13580);
nand UO_1412 (O_1412,N_13943,N_12107);
and UO_1413 (O_1413,N_12991,N_12320);
nand UO_1414 (O_1414,N_13884,N_12728);
nand UO_1415 (O_1415,N_14704,N_14222);
nor UO_1416 (O_1416,N_14697,N_13740);
or UO_1417 (O_1417,N_13467,N_13527);
and UO_1418 (O_1418,N_14968,N_12261);
or UO_1419 (O_1419,N_12933,N_12194);
nor UO_1420 (O_1420,N_14680,N_13215);
nand UO_1421 (O_1421,N_12162,N_12160);
and UO_1422 (O_1422,N_12290,N_14221);
nand UO_1423 (O_1423,N_13027,N_13777);
and UO_1424 (O_1424,N_12949,N_14662);
xor UO_1425 (O_1425,N_12565,N_14789);
nor UO_1426 (O_1426,N_14580,N_14906);
and UO_1427 (O_1427,N_14883,N_14022);
nand UO_1428 (O_1428,N_12730,N_13850);
nor UO_1429 (O_1429,N_12136,N_12142);
nor UO_1430 (O_1430,N_12997,N_12212);
and UO_1431 (O_1431,N_13457,N_14478);
nor UO_1432 (O_1432,N_12965,N_12552);
and UO_1433 (O_1433,N_13593,N_14150);
nand UO_1434 (O_1434,N_14012,N_13624);
nand UO_1435 (O_1435,N_14606,N_12741);
nand UO_1436 (O_1436,N_14067,N_13572);
or UO_1437 (O_1437,N_13308,N_12456);
xnor UO_1438 (O_1438,N_14152,N_12642);
nor UO_1439 (O_1439,N_12488,N_12717);
nor UO_1440 (O_1440,N_14355,N_14616);
and UO_1441 (O_1441,N_13958,N_12515);
and UO_1442 (O_1442,N_14507,N_12894);
or UO_1443 (O_1443,N_12272,N_12353);
nor UO_1444 (O_1444,N_12650,N_13031);
nand UO_1445 (O_1445,N_13749,N_14077);
and UO_1446 (O_1446,N_13923,N_14822);
nor UO_1447 (O_1447,N_13721,N_12483);
nor UO_1448 (O_1448,N_14276,N_12955);
xor UO_1449 (O_1449,N_12269,N_13312);
and UO_1450 (O_1450,N_14073,N_12660);
nor UO_1451 (O_1451,N_13622,N_14183);
and UO_1452 (O_1452,N_12259,N_14905);
or UO_1453 (O_1453,N_13595,N_13322);
nor UO_1454 (O_1454,N_12120,N_13538);
nand UO_1455 (O_1455,N_12397,N_13674);
xor UO_1456 (O_1456,N_14920,N_14311);
nor UO_1457 (O_1457,N_13065,N_13866);
xor UO_1458 (O_1458,N_12217,N_14289);
or UO_1459 (O_1459,N_12919,N_14816);
and UO_1460 (O_1460,N_13954,N_12371);
xor UO_1461 (O_1461,N_13925,N_12746);
or UO_1462 (O_1462,N_12905,N_13788);
nor UO_1463 (O_1463,N_12602,N_12401);
or UO_1464 (O_1464,N_12648,N_14687);
nor UO_1465 (O_1465,N_14574,N_13276);
or UO_1466 (O_1466,N_12420,N_12638);
nand UO_1467 (O_1467,N_12416,N_14614);
and UO_1468 (O_1468,N_12166,N_13727);
nor UO_1469 (O_1469,N_14878,N_14624);
or UO_1470 (O_1470,N_14750,N_12199);
nor UO_1471 (O_1471,N_14599,N_12751);
nand UO_1472 (O_1472,N_14091,N_13996);
nand UO_1473 (O_1473,N_12522,N_14846);
nand UO_1474 (O_1474,N_12599,N_14735);
xor UO_1475 (O_1475,N_14371,N_13018);
nor UO_1476 (O_1476,N_14132,N_14812);
xor UO_1477 (O_1477,N_13704,N_12725);
nand UO_1478 (O_1478,N_14901,N_12312);
or UO_1479 (O_1479,N_12315,N_12278);
or UO_1480 (O_1480,N_14504,N_12177);
and UO_1481 (O_1481,N_12925,N_12795);
and UO_1482 (O_1482,N_14763,N_13481);
and UO_1483 (O_1483,N_14170,N_13644);
or UO_1484 (O_1484,N_13392,N_12821);
or UO_1485 (O_1485,N_14537,N_13647);
xor UO_1486 (O_1486,N_12887,N_14688);
xor UO_1487 (O_1487,N_14014,N_14397);
nand UO_1488 (O_1488,N_12296,N_14948);
or UO_1489 (O_1489,N_13733,N_13241);
and UO_1490 (O_1490,N_14413,N_12444);
nand UO_1491 (O_1491,N_13824,N_12013);
nor UO_1492 (O_1492,N_13116,N_13835);
or UO_1493 (O_1493,N_14669,N_13330);
or UO_1494 (O_1494,N_14869,N_14318);
nand UO_1495 (O_1495,N_12825,N_14117);
xor UO_1496 (O_1496,N_13220,N_13584);
nand UO_1497 (O_1497,N_14029,N_12878);
and UO_1498 (O_1498,N_14502,N_13101);
nor UO_1499 (O_1499,N_12605,N_13121);
nor UO_1500 (O_1500,N_12077,N_12794);
or UO_1501 (O_1501,N_12215,N_13415);
xnor UO_1502 (O_1502,N_12475,N_12941);
xor UO_1503 (O_1503,N_13635,N_13620);
nor UO_1504 (O_1504,N_12339,N_13394);
nor UO_1505 (O_1505,N_12948,N_12995);
nor UO_1506 (O_1506,N_12844,N_12265);
and UO_1507 (O_1507,N_12925,N_13250);
xor UO_1508 (O_1508,N_14472,N_12559);
and UO_1509 (O_1509,N_14393,N_12631);
xnor UO_1510 (O_1510,N_13234,N_12617);
nor UO_1511 (O_1511,N_12132,N_12323);
nor UO_1512 (O_1512,N_14253,N_12171);
xnor UO_1513 (O_1513,N_13261,N_12624);
and UO_1514 (O_1514,N_14067,N_13196);
and UO_1515 (O_1515,N_13200,N_12979);
or UO_1516 (O_1516,N_12980,N_12457);
nor UO_1517 (O_1517,N_13924,N_14404);
nor UO_1518 (O_1518,N_13489,N_14649);
nand UO_1519 (O_1519,N_13505,N_13961);
or UO_1520 (O_1520,N_14994,N_12945);
and UO_1521 (O_1521,N_13844,N_13459);
nor UO_1522 (O_1522,N_14660,N_14983);
nand UO_1523 (O_1523,N_12453,N_13739);
nand UO_1524 (O_1524,N_14068,N_12373);
nand UO_1525 (O_1525,N_12808,N_12533);
nor UO_1526 (O_1526,N_14437,N_12272);
nor UO_1527 (O_1527,N_14399,N_12549);
nand UO_1528 (O_1528,N_12100,N_12161);
nand UO_1529 (O_1529,N_12415,N_14567);
nor UO_1530 (O_1530,N_12925,N_12086);
nand UO_1531 (O_1531,N_12930,N_14507);
nand UO_1532 (O_1532,N_13687,N_12101);
or UO_1533 (O_1533,N_13296,N_14175);
nor UO_1534 (O_1534,N_13920,N_12916);
nand UO_1535 (O_1535,N_13648,N_12362);
nor UO_1536 (O_1536,N_12491,N_14091);
nand UO_1537 (O_1537,N_14777,N_13136);
and UO_1538 (O_1538,N_13879,N_14783);
or UO_1539 (O_1539,N_13307,N_13805);
nor UO_1540 (O_1540,N_14019,N_12464);
or UO_1541 (O_1541,N_14901,N_13817);
and UO_1542 (O_1542,N_13104,N_12255);
nand UO_1543 (O_1543,N_14728,N_12548);
nand UO_1544 (O_1544,N_14585,N_14734);
xnor UO_1545 (O_1545,N_13395,N_13079);
or UO_1546 (O_1546,N_13432,N_14557);
nand UO_1547 (O_1547,N_12225,N_13518);
and UO_1548 (O_1548,N_14692,N_14163);
xor UO_1549 (O_1549,N_13737,N_12530);
nand UO_1550 (O_1550,N_13631,N_14605);
or UO_1551 (O_1551,N_12648,N_14543);
nand UO_1552 (O_1552,N_14179,N_12594);
or UO_1553 (O_1553,N_14187,N_12759);
nor UO_1554 (O_1554,N_12848,N_13058);
nor UO_1555 (O_1555,N_14429,N_14458);
xor UO_1556 (O_1556,N_14756,N_14901);
and UO_1557 (O_1557,N_13426,N_13048);
nand UO_1558 (O_1558,N_12131,N_12335);
nand UO_1559 (O_1559,N_14594,N_14839);
nand UO_1560 (O_1560,N_12039,N_14076);
or UO_1561 (O_1561,N_14138,N_14968);
and UO_1562 (O_1562,N_12042,N_12402);
nor UO_1563 (O_1563,N_14089,N_12223);
and UO_1564 (O_1564,N_13546,N_12670);
nand UO_1565 (O_1565,N_14677,N_14516);
nand UO_1566 (O_1566,N_13074,N_14942);
nand UO_1567 (O_1567,N_12105,N_14575);
and UO_1568 (O_1568,N_13712,N_12874);
xnor UO_1569 (O_1569,N_14367,N_14331);
nand UO_1570 (O_1570,N_14491,N_13697);
or UO_1571 (O_1571,N_13042,N_13487);
or UO_1572 (O_1572,N_13780,N_13891);
nand UO_1573 (O_1573,N_14485,N_12094);
nand UO_1574 (O_1574,N_12007,N_14728);
nor UO_1575 (O_1575,N_12265,N_14957);
or UO_1576 (O_1576,N_14633,N_13316);
or UO_1577 (O_1577,N_13532,N_12093);
xor UO_1578 (O_1578,N_13442,N_14986);
and UO_1579 (O_1579,N_14999,N_14276);
and UO_1580 (O_1580,N_12976,N_14649);
or UO_1581 (O_1581,N_14671,N_14309);
or UO_1582 (O_1582,N_13954,N_14779);
nand UO_1583 (O_1583,N_13882,N_12099);
and UO_1584 (O_1584,N_12954,N_13540);
or UO_1585 (O_1585,N_13726,N_14291);
or UO_1586 (O_1586,N_12868,N_12811);
nor UO_1587 (O_1587,N_14757,N_14194);
xor UO_1588 (O_1588,N_14612,N_12712);
and UO_1589 (O_1589,N_12882,N_14363);
nand UO_1590 (O_1590,N_13181,N_13437);
nor UO_1591 (O_1591,N_12502,N_14565);
and UO_1592 (O_1592,N_13178,N_14533);
nand UO_1593 (O_1593,N_14034,N_14450);
and UO_1594 (O_1594,N_13645,N_14846);
or UO_1595 (O_1595,N_14229,N_13046);
and UO_1596 (O_1596,N_14023,N_13111);
nor UO_1597 (O_1597,N_14211,N_14041);
nor UO_1598 (O_1598,N_12099,N_12098);
and UO_1599 (O_1599,N_13407,N_14006);
and UO_1600 (O_1600,N_14278,N_13460);
nor UO_1601 (O_1601,N_14251,N_12248);
or UO_1602 (O_1602,N_14813,N_14345);
or UO_1603 (O_1603,N_13083,N_12257);
and UO_1604 (O_1604,N_12713,N_13060);
nor UO_1605 (O_1605,N_12927,N_13259);
xnor UO_1606 (O_1606,N_13819,N_14776);
nor UO_1607 (O_1607,N_14438,N_14738);
xnor UO_1608 (O_1608,N_14027,N_14247);
and UO_1609 (O_1609,N_14127,N_12532);
nand UO_1610 (O_1610,N_14295,N_12119);
nor UO_1611 (O_1611,N_13816,N_13533);
nor UO_1612 (O_1612,N_13189,N_13435);
xnor UO_1613 (O_1613,N_14347,N_13113);
and UO_1614 (O_1614,N_14447,N_13464);
nand UO_1615 (O_1615,N_14541,N_13731);
nor UO_1616 (O_1616,N_14468,N_14526);
nand UO_1617 (O_1617,N_12426,N_12102);
or UO_1618 (O_1618,N_12442,N_12502);
and UO_1619 (O_1619,N_14347,N_12811);
or UO_1620 (O_1620,N_13780,N_13048);
nor UO_1621 (O_1621,N_14596,N_13697);
nand UO_1622 (O_1622,N_12627,N_12030);
nand UO_1623 (O_1623,N_12344,N_13542);
and UO_1624 (O_1624,N_12623,N_14924);
xnor UO_1625 (O_1625,N_13799,N_12749);
nand UO_1626 (O_1626,N_12011,N_12839);
or UO_1627 (O_1627,N_14448,N_13040);
nor UO_1628 (O_1628,N_14309,N_14890);
nor UO_1629 (O_1629,N_12467,N_12881);
nand UO_1630 (O_1630,N_13862,N_13596);
nor UO_1631 (O_1631,N_13569,N_13563);
nand UO_1632 (O_1632,N_14139,N_13278);
nand UO_1633 (O_1633,N_12161,N_13449);
and UO_1634 (O_1634,N_14219,N_13459);
or UO_1635 (O_1635,N_14178,N_12464);
or UO_1636 (O_1636,N_14012,N_14680);
xnor UO_1637 (O_1637,N_12358,N_14829);
and UO_1638 (O_1638,N_14318,N_12326);
or UO_1639 (O_1639,N_13392,N_13710);
xor UO_1640 (O_1640,N_12743,N_12391);
xnor UO_1641 (O_1641,N_14965,N_12273);
and UO_1642 (O_1642,N_12097,N_14580);
or UO_1643 (O_1643,N_13456,N_13009);
nand UO_1644 (O_1644,N_12550,N_13630);
and UO_1645 (O_1645,N_13282,N_14383);
and UO_1646 (O_1646,N_13099,N_14260);
or UO_1647 (O_1647,N_13446,N_12885);
nand UO_1648 (O_1648,N_12012,N_14325);
or UO_1649 (O_1649,N_13990,N_13476);
or UO_1650 (O_1650,N_12238,N_14855);
nor UO_1651 (O_1651,N_13462,N_13656);
and UO_1652 (O_1652,N_12176,N_13423);
nand UO_1653 (O_1653,N_14270,N_12635);
nor UO_1654 (O_1654,N_12105,N_12748);
and UO_1655 (O_1655,N_13460,N_13012);
xor UO_1656 (O_1656,N_13022,N_13486);
nor UO_1657 (O_1657,N_13951,N_12461);
nor UO_1658 (O_1658,N_14129,N_14119);
and UO_1659 (O_1659,N_14478,N_14621);
or UO_1660 (O_1660,N_12148,N_12456);
nand UO_1661 (O_1661,N_14015,N_12401);
nor UO_1662 (O_1662,N_12003,N_14039);
nand UO_1663 (O_1663,N_13328,N_13403);
nor UO_1664 (O_1664,N_14926,N_12512);
nand UO_1665 (O_1665,N_13952,N_14848);
xnor UO_1666 (O_1666,N_12251,N_13096);
nand UO_1667 (O_1667,N_12905,N_13383);
nand UO_1668 (O_1668,N_13069,N_14548);
xor UO_1669 (O_1669,N_14453,N_14594);
or UO_1670 (O_1670,N_14820,N_12820);
nor UO_1671 (O_1671,N_12549,N_12457);
nand UO_1672 (O_1672,N_14528,N_14836);
or UO_1673 (O_1673,N_13236,N_14886);
nand UO_1674 (O_1674,N_13910,N_13159);
nor UO_1675 (O_1675,N_12563,N_12737);
xor UO_1676 (O_1676,N_14198,N_14371);
nand UO_1677 (O_1677,N_14503,N_12671);
or UO_1678 (O_1678,N_14139,N_12603);
and UO_1679 (O_1679,N_13608,N_13927);
and UO_1680 (O_1680,N_13499,N_14357);
and UO_1681 (O_1681,N_14442,N_14621);
nor UO_1682 (O_1682,N_12266,N_13984);
and UO_1683 (O_1683,N_14966,N_14371);
xor UO_1684 (O_1684,N_12690,N_13331);
nor UO_1685 (O_1685,N_14824,N_12642);
nand UO_1686 (O_1686,N_14962,N_13017);
and UO_1687 (O_1687,N_12853,N_13484);
nor UO_1688 (O_1688,N_12325,N_13000);
and UO_1689 (O_1689,N_12128,N_14467);
and UO_1690 (O_1690,N_13370,N_14062);
nor UO_1691 (O_1691,N_14518,N_12698);
or UO_1692 (O_1692,N_12236,N_14203);
nand UO_1693 (O_1693,N_14452,N_12940);
or UO_1694 (O_1694,N_14503,N_12734);
or UO_1695 (O_1695,N_13064,N_14102);
xor UO_1696 (O_1696,N_12179,N_13430);
and UO_1697 (O_1697,N_14542,N_14196);
xnor UO_1698 (O_1698,N_14919,N_12137);
or UO_1699 (O_1699,N_14265,N_13412);
or UO_1700 (O_1700,N_12323,N_12733);
nor UO_1701 (O_1701,N_14644,N_14741);
and UO_1702 (O_1702,N_13451,N_14429);
xor UO_1703 (O_1703,N_14665,N_12333);
and UO_1704 (O_1704,N_14548,N_12806);
and UO_1705 (O_1705,N_14820,N_12344);
or UO_1706 (O_1706,N_13128,N_14795);
nand UO_1707 (O_1707,N_13335,N_12399);
and UO_1708 (O_1708,N_12563,N_13337);
nand UO_1709 (O_1709,N_14406,N_13896);
nor UO_1710 (O_1710,N_14707,N_12752);
nor UO_1711 (O_1711,N_12441,N_12222);
or UO_1712 (O_1712,N_13021,N_13735);
and UO_1713 (O_1713,N_14533,N_13438);
nor UO_1714 (O_1714,N_14379,N_12255);
and UO_1715 (O_1715,N_12756,N_14554);
nor UO_1716 (O_1716,N_14699,N_12992);
or UO_1717 (O_1717,N_12672,N_12532);
xor UO_1718 (O_1718,N_12335,N_14401);
or UO_1719 (O_1719,N_13586,N_12570);
and UO_1720 (O_1720,N_12984,N_14803);
and UO_1721 (O_1721,N_14502,N_12543);
or UO_1722 (O_1722,N_12990,N_12833);
or UO_1723 (O_1723,N_13754,N_14115);
nand UO_1724 (O_1724,N_13484,N_12528);
nand UO_1725 (O_1725,N_13086,N_13207);
and UO_1726 (O_1726,N_13632,N_13618);
or UO_1727 (O_1727,N_12399,N_12592);
nand UO_1728 (O_1728,N_14397,N_13077);
or UO_1729 (O_1729,N_12657,N_14907);
nor UO_1730 (O_1730,N_12493,N_12469);
or UO_1731 (O_1731,N_14720,N_13814);
nor UO_1732 (O_1732,N_14982,N_13688);
nand UO_1733 (O_1733,N_12100,N_14593);
nand UO_1734 (O_1734,N_12415,N_14928);
nand UO_1735 (O_1735,N_14423,N_13801);
xnor UO_1736 (O_1736,N_14168,N_14033);
xnor UO_1737 (O_1737,N_12189,N_12165);
and UO_1738 (O_1738,N_14167,N_13836);
or UO_1739 (O_1739,N_13552,N_13668);
xnor UO_1740 (O_1740,N_14456,N_13959);
or UO_1741 (O_1741,N_12854,N_12537);
and UO_1742 (O_1742,N_12099,N_14510);
nor UO_1743 (O_1743,N_13513,N_12205);
nor UO_1744 (O_1744,N_12593,N_14780);
or UO_1745 (O_1745,N_13834,N_13151);
nor UO_1746 (O_1746,N_12307,N_14032);
nand UO_1747 (O_1747,N_14956,N_13005);
nor UO_1748 (O_1748,N_12337,N_12522);
or UO_1749 (O_1749,N_13427,N_13965);
or UO_1750 (O_1750,N_14134,N_14369);
and UO_1751 (O_1751,N_12143,N_14479);
and UO_1752 (O_1752,N_13947,N_13753);
and UO_1753 (O_1753,N_14270,N_12413);
xor UO_1754 (O_1754,N_14112,N_14909);
nand UO_1755 (O_1755,N_14122,N_14331);
and UO_1756 (O_1756,N_13771,N_14536);
or UO_1757 (O_1757,N_13479,N_14028);
or UO_1758 (O_1758,N_14490,N_13458);
nand UO_1759 (O_1759,N_13365,N_12075);
or UO_1760 (O_1760,N_13182,N_12844);
nand UO_1761 (O_1761,N_13726,N_13373);
nor UO_1762 (O_1762,N_12331,N_12188);
and UO_1763 (O_1763,N_12180,N_14083);
nand UO_1764 (O_1764,N_14433,N_14184);
and UO_1765 (O_1765,N_14234,N_13004);
nor UO_1766 (O_1766,N_13892,N_14961);
and UO_1767 (O_1767,N_12160,N_12338);
or UO_1768 (O_1768,N_13542,N_12034);
nor UO_1769 (O_1769,N_12876,N_12940);
and UO_1770 (O_1770,N_13400,N_14714);
nor UO_1771 (O_1771,N_13697,N_14135);
or UO_1772 (O_1772,N_14961,N_13801);
or UO_1773 (O_1773,N_12925,N_12916);
nor UO_1774 (O_1774,N_12853,N_12445);
xnor UO_1775 (O_1775,N_13667,N_13423);
nand UO_1776 (O_1776,N_13570,N_13706);
and UO_1777 (O_1777,N_14892,N_13501);
nand UO_1778 (O_1778,N_13159,N_14494);
or UO_1779 (O_1779,N_14526,N_13993);
nand UO_1780 (O_1780,N_13362,N_12058);
nor UO_1781 (O_1781,N_12698,N_12355);
and UO_1782 (O_1782,N_13449,N_13198);
nand UO_1783 (O_1783,N_12756,N_13655);
nor UO_1784 (O_1784,N_13819,N_14337);
and UO_1785 (O_1785,N_12963,N_13320);
or UO_1786 (O_1786,N_12231,N_14952);
nand UO_1787 (O_1787,N_13768,N_14394);
nand UO_1788 (O_1788,N_14131,N_14507);
nand UO_1789 (O_1789,N_13061,N_13677);
or UO_1790 (O_1790,N_14963,N_13363);
or UO_1791 (O_1791,N_13247,N_12002);
nand UO_1792 (O_1792,N_12194,N_14422);
or UO_1793 (O_1793,N_13822,N_14153);
nor UO_1794 (O_1794,N_12577,N_12251);
and UO_1795 (O_1795,N_13806,N_12593);
nor UO_1796 (O_1796,N_14917,N_14489);
xor UO_1797 (O_1797,N_13038,N_12541);
nand UO_1798 (O_1798,N_13276,N_12701);
and UO_1799 (O_1799,N_12231,N_14618);
and UO_1800 (O_1800,N_13625,N_13843);
xnor UO_1801 (O_1801,N_13607,N_14699);
and UO_1802 (O_1802,N_12730,N_13594);
and UO_1803 (O_1803,N_14823,N_14626);
xnor UO_1804 (O_1804,N_12663,N_14682);
xnor UO_1805 (O_1805,N_14647,N_13658);
or UO_1806 (O_1806,N_12710,N_12488);
xor UO_1807 (O_1807,N_12140,N_13341);
nor UO_1808 (O_1808,N_12573,N_13391);
nor UO_1809 (O_1809,N_14342,N_12721);
nand UO_1810 (O_1810,N_12901,N_14017);
nand UO_1811 (O_1811,N_13248,N_13921);
nor UO_1812 (O_1812,N_13513,N_13542);
xor UO_1813 (O_1813,N_12408,N_12910);
and UO_1814 (O_1814,N_12112,N_12542);
xor UO_1815 (O_1815,N_12191,N_14093);
nor UO_1816 (O_1816,N_14025,N_13400);
nand UO_1817 (O_1817,N_12672,N_12063);
or UO_1818 (O_1818,N_14311,N_12722);
and UO_1819 (O_1819,N_13208,N_13476);
nor UO_1820 (O_1820,N_14244,N_14785);
and UO_1821 (O_1821,N_13576,N_14581);
and UO_1822 (O_1822,N_12741,N_13308);
or UO_1823 (O_1823,N_12797,N_14211);
nor UO_1824 (O_1824,N_13500,N_14874);
nor UO_1825 (O_1825,N_13784,N_14614);
or UO_1826 (O_1826,N_14275,N_12620);
or UO_1827 (O_1827,N_12736,N_12937);
or UO_1828 (O_1828,N_12027,N_14309);
nand UO_1829 (O_1829,N_12850,N_12233);
nand UO_1830 (O_1830,N_13079,N_13518);
and UO_1831 (O_1831,N_14483,N_12488);
and UO_1832 (O_1832,N_14300,N_12117);
nand UO_1833 (O_1833,N_14257,N_14029);
or UO_1834 (O_1834,N_12562,N_12580);
nand UO_1835 (O_1835,N_13156,N_12689);
or UO_1836 (O_1836,N_13527,N_13920);
nor UO_1837 (O_1837,N_14119,N_12163);
nand UO_1838 (O_1838,N_14249,N_13170);
xnor UO_1839 (O_1839,N_13134,N_12780);
and UO_1840 (O_1840,N_12551,N_14567);
or UO_1841 (O_1841,N_14603,N_14187);
nor UO_1842 (O_1842,N_12404,N_14099);
or UO_1843 (O_1843,N_12581,N_12553);
nor UO_1844 (O_1844,N_12355,N_12125);
nand UO_1845 (O_1845,N_12775,N_13553);
xor UO_1846 (O_1846,N_13000,N_12644);
nor UO_1847 (O_1847,N_14003,N_14770);
nand UO_1848 (O_1848,N_14311,N_14754);
nor UO_1849 (O_1849,N_14933,N_14931);
nand UO_1850 (O_1850,N_13914,N_14386);
and UO_1851 (O_1851,N_12040,N_12988);
nand UO_1852 (O_1852,N_12107,N_13868);
nor UO_1853 (O_1853,N_13469,N_14789);
xor UO_1854 (O_1854,N_12355,N_13617);
nor UO_1855 (O_1855,N_13770,N_12426);
or UO_1856 (O_1856,N_12765,N_12768);
nand UO_1857 (O_1857,N_14131,N_14412);
and UO_1858 (O_1858,N_14035,N_14738);
or UO_1859 (O_1859,N_13065,N_12506);
and UO_1860 (O_1860,N_12276,N_14773);
xnor UO_1861 (O_1861,N_12330,N_14692);
nand UO_1862 (O_1862,N_13983,N_14655);
nor UO_1863 (O_1863,N_13903,N_13996);
nand UO_1864 (O_1864,N_13035,N_13050);
and UO_1865 (O_1865,N_14476,N_12119);
and UO_1866 (O_1866,N_12696,N_13455);
and UO_1867 (O_1867,N_14098,N_14698);
or UO_1868 (O_1868,N_14603,N_13045);
or UO_1869 (O_1869,N_13363,N_12119);
nor UO_1870 (O_1870,N_14098,N_12130);
nand UO_1871 (O_1871,N_13419,N_12766);
or UO_1872 (O_1872,N_13848,N_14857);
nand UO_1873 (O_1873,N_13853,N_13470);
or UO_1874 (O_1874,N_12266,N_13235);
or UO_1875 (O_1875,N_14558,N_13594);
nand UO_1876 (O_1876,N_12343,N_13120);
xor UO_1877 (O_1877,N_12706,N_14948);
or UO_1878 (O_1878,N_14842,N_13782);
nor UO_1879 (O_1879,N_14420,N_12318);
nand UO_1880 (O_1880,N_14176,N_12562);
and UO_1881 (O_1881,N_14612,N_13246);
and UO_1882 (O_1882,N_12237,N_14343);
and UO_1883 (O_1883,N_13340,N_13826);
nand UO_1884 (O_1884,N_12295,N_13804);
nand UO_1885 (O_1885,N_14908,N_12797);
or UO_1886 (O_1886,N_13015,N_12333);
or UO_1887 (O_1887,N_12597,N_14818);
nand UO_1888 (O_1888,N_14269,N_13044);
nor UO_1889 (O_1889,N_13809,N_13090);
nand UO_1890 (O_1890,N_14275,N_14113);
nand UO_1891 (O_1891,N_14715,N_12573);
and UO_1892 (O_1892,N_14541,N_12816);
nor UO_1893 (O_1893,N_12471,N_13057);
nand UO_1894 (O_1894,N_13120,N_14125);
nand UO_1895 (O_1895,N_13608,N_12027);
nor UO_1896 (O_1896,N_13253,N_14776);
or UO_1897 (O_1897,N_14319,N_14728);
and UO_1898 (O_1898,N_13942,N_13585);
nor UO_1899 (O_1899,N_13047,N_14076);
nand UO_1900 (O_1900,N_13820,N_13604);
and UO_1901 (O_1901,N_12358,N_14867);
nor UO_1902 (O_1902,N_13311,N_13284);
or UO_1903 (O_1903,N_13379,N_14068);
xnor UO_1904 (O_1904,N_13315,N_13685);
nand UO_1905 (O_1905,N_12434,N_13015);
or UO_1906 (O_1906,N_12316,N_14032);
xnor UO_1907 (O_1907,N_13678,N_14499);
or UO_1908 (O_1908,N_13785,N_13995);
xor UO_1909 (O_1909,N_13475,N_13371);
nor UO_1910 (O_1910,N_14663,N_12004);
nand UO_1911 (O_1911,N_12159,N_12144);
and UO_1912 (O_1912,N_13685,N_12644);
nor UO_1913 (O_1913,N_14550,N_14480);
nor UO_1914 (O_1914,N_13535,N_14795);
nor UO_1915 (O_1915,N_14661,N_13927);
xnor UO_1916 (O_1916,N_12966,N_13833);
nand UO_1917 (O_1917,N_13524,N_13662);
or UO_1918 (O_1918,N_14787,N_13505);
or UO_1919 (O_1919,N_13336,N_13026);
nor UO_1920 (O_1920,N_14646,N_12624);
xor UO_1921 (O_1921,N_13205,N_14896);
nand UO_1922 (O_1922,N_14438,N_12504);
or UO_1923 (O_1923,N_14066,N_12468);
xor UO_1924 (O_1924,N_12595,N_13980);
nand UO_1925 (O_1925,N_14207,N_13408);
nor UO_1926 (O_1926,N_12394,N_12530);
and UO_1927 (O_1927,N_12144,N_12129);
nand UO_1928 (O_1928,N_14880,N_14665);
or UO_1929 (O_1929,N_14719,N_12472);
nand UO_1930 (O_1930,N_13620,N_12842);
nand UO_1931 (O_1931,N_13631,N_12190);
or UO_1932 (O_1932,N_12149,N_13303);
or UO_1933 (O_1933,N_13935,N_13291);
or UO_1934 (O_1934,N_14138,N_13808);
nand UO_1935 (O_1935,N_14497,N_13434);
or UO_1936 (O_1936,N_14466,N_12514);
and UO_1937 (O_1937,N_14799,N_14536);
nor UO_1938 (O_1938,N_13745,N_12220);
or UO_1939 (O_1939,N_13882,N_13431);
nand UO_1940 (O_1940,N_13218,N_13773);
nand UO_1941 (O_1941,N_14173,N_13121);
nand UO_1942 (O_1942,N_13737,N_12600);
or UO_1943 (O_1943,N_13924,N_14178);
nor UO_1944 (O_1944,N_13943,N_14100);
or UO_1945 (O_1945,N_12292,N_14730);
and UO_1946 (O_1946,N_12598,N_13246);
and UO_1947 (O_1947,N_13100,N_13242);
or UO_1948 (O_1948,N_12452,N_13976);
xnor UO_1949 (O_1949,N_13424,N_12548);
xor UO_1950 (O_1950,N_13919,N_14292);
xnor UO_1951 (O_1951,N_14101,N_12504);
and UO_1952 (O_1952,N_14290,N_14179);
nand UO_1953 (O_1953,N_12880,N_12028);
and UO_1954 (O_1954,N_13986,N_13030);
nor UO_1955 (O_1955,N_13711,N_14285);
nand UO_1956 (O_1956,N_12635,N_12364);
nand UO_1957 (O_1957,N_12017,N_14517);
nor UO_1958 (O_1958,N_13723,N_14044);
and UO_1959 (O_1959,N_13953,N_12103);
nor UO_1960 (O_1960,N_14053,N_12992);
or UO_1961 (O_1961,N_13187,N_12774);
or UO_1962 (O_1962,N_13447,N_12601);
nand UO_1963 (O_1963,N_13112,N_12267);
or UO_1964 (O_1964,N_13823,N_12079);
and UO_1965 (O_1965,N_13278,N_13374);
or UO_1966 (O_1966,N_14587,N_12703);
and UO_1967 (O_1967,N_12784,N_13527);
nand UO_1968 (O_1968,N_14893,N_12855);
nor UO_1969 (O_1969,N_12100,N_12786);
xor UO_1970 (O_1970,N_13821,N_14590);
xnor UO_1971 (O_1971,N_14715,N_12668);
nor UO_1972 (O_1972,N_12484,N_13268);
nor UO_1973 (O_1973,N_13567,N_14273);
nor UO_1974 (O_1974,N_13544,N_13791);
nand UO_1975 (O_1975,N_13132,N_13830);
or UO_1976 (O_1976,N_12670,N_12096);
nand UO_1977 (O_1977,N_14258,N_12545);
or UO_1978 (O_1978,N_12445,N_13299);
and UO_1979 (O_1979,N_14558,N_13397);
nand UO_1980 (O_1980,N_14094,N_13523);
nor UO_1981 (O_1981,N_14843,N_13244);
and UO_1982 (O_1982,N_13404,N_14753);
nor UO_1983 (O_1983,N_13436,N_13659);
and UO_1984 (O_1984,N_13101,N_13509);
and UO_1985 (O_1985,N_13064,N_13801);
xor UO_1986 (O_1986,N_13935,N_13373);
or UO_1987 (O_1987,N_13617,N_13463);
or UO_1988 (O_1988,N_14851,N_12677);
and UO_1989 (O_1989,N_12563,N_13944);
nand UO_1990 (O_1990,N_12473,N_12246);
nand UO_1991 (O_1991,N_14391,N_14050);
or UO_1992 (O_1992,N_12804,N_12869);
nand UO_1993 (O_1993,N_14517,N_14935);
or UO_1994 (O_1994,N_14427,N_12303);
and UO_1995 (O_1995,N_14000,N_14778);
and UO_1996 (O_1996,N_14957,N_12736);
or UO_1997 (O_1997,N_13818,N_14701);
nand UO_1998 (O_1998,N_13235,N_14886);
and UO_1999 (O_1999,N_13400,N_12016);
endmodule