module basic_1000_10000_1500_10_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_194,In_435);
or U1 (N_1,In_350,In_181);
and U2 (N_2,In_385,In_580);
nand U3 (N_3,In_178,In_4);
or U4 (N_4,In_746,In_203);
nand U5 (N_5,In_268,In_843);
or U6 (N_6,In_893,In_852);
or U7 (N_7,In_67,In_359);
nor U8 (N_8,In_701,In_293);
and U9 (N_9,In_406,In_726);
and U10 (N_10,In_933,In_470);
nor U11 (N_11,In_180,In_379);
or U12 (N_12,In_763,In_753);
nand U13 (N_13,In_501,In_845);
or U14 (N_14,In_747,In_770);
nand U15 (N_15,In_986,In_801);
or U16 (N_16,In_642,In_785);
nand U17 (N_17,In_963,In_583);
or U18 (N_18,In_579,In_212);
nand U19 (N_19,In_946,In_516);
nand U20 (N_20,In_585,In_23);
or U21 (N_21,In_36,In_916);
nand U22 (N_22,In_388,In_721);
and U23 (N_23,In_771,In_650);
nand U24 (N_24,In_632,In_233);
or U25 (N_25,In_519,In_183);
and U26 (N_26,In_641,In_241);
or U27 (N_27,In_577,In_676);
and U28 (N_28,In_965,In_133);
nand U29 (N_29,In_720,In_330);
nand U30 (N_30,In_961,In_670);
nand U31 (N_31,In_790,In_578);
nor U32 (N_32,In_321,In_329);
nor U33 (N_33,In_510,In_56);
or U34 (N_34,In_266,In_745);
nor U35 (N_35,In_989,In_99);
and U36 (N_36,In_815,In_381);
nor U37 (N_37,In_227,In_731);
nor U38 (N_38,In_775,In_619);
nor U39 (N_39,In_975,In_484);
and U40 (N_40,In_325,In_467);
nand U41 (N_41,In_112,In_306);
nand U42 (N_42,In_283,In_299);
nand U43 (N_43,In_547,In_12);
or U44 (N_44,In_688,In_3);
and U45 (N_45,In_430,In_103);
nor U46 (N_46,In_750,In_201);
nand U47 (N_47,In_728,In_977);
xnor U48 (N_48,In_479,In_628);
nand U49 (N_49,In_533,In_654);
nand U50 (N_50,In_985,In_289);
nand U51 (N_51,In_554,In_104);
nor U52 (N_52,In_396,In_981);
or U53 (N_53,In_626,In_341);
nor U54 (N_54,In_923,In_93);
nor U55 (N_55,In_73,In_47);
nand U56 (N_56,In_0,In_395);
nand U57 (N_57,In_429,In_620);
or U58 (N_58,In_298,In_394);
xnor U59 (N_59,In_738,In_873);
or U60 (N_60,In_444,In_851);
nand U61 (N_61,In_348,In_187);
or U62 (N_62,In_779,In_618);
nor U63 (N_63,In_734,In_562);
nand U64 (N_64,In_869,In_652);
and U65 (N_65,In_326,In_380);
nor U66 (N_66,In_534,In_639);
nand U67 (N_67,In_725,In_54);
xor U68 (N_68,In_79,In_523);
nand U69 (N_69,In_612,In_634);
or U70 (N_70,In_145,In_62);
and U71 (N_71,In_453,In_482);
or U72 (N_72,In_709,In_862);
xnor U73 (N_73,In_20,In_796);
nand U74 (N_74,In_239,In_651);
or U75 (N_75,In_84,In_448);
nand U76 (N_76,In_89,In_949);
nor U77 (N_77,In_269,In_575);
nor U78 (N_78,In_777,In_378);
nand U79 (N_79,In_727,In_419);
and U80 (N_80,In_814,In_878);
and U81 (N_81,In_952,In_912);
and U82 (N_82,In_765,In_653);
nand U83 (N_83,In_433,In_190);
nor U84 (N_84,In_18,In_68);
and U85 (N_85,In_640,In_566);
or U86 (N_86,In_410,In_597);
and U87 (N_87,In_384,In_972);
or U88 (N_88,In_234,In_169);
nand U89 (N_89,In_897,In_80);
nand U90 (N_90,In_886,In_70);
nor U91 (N_91,In_673,In_892);
nand U92 (N_92,In_553,In_317);
or U93 (N_93,In_52,In_987);
nor U94 (N_94,In_625,In_557);
nor U95 (N_95,In_32,In_392);
nand U96 (N_96,In_476,In_64);
and U97 (N_97,In_969,In_459);
and U98 (N_98,In_764,In_28);
and U99 (N_99,In_156,In_899);
nand U100 (N_100,In_638,In_550);
and U101 (N_101,In_454,In_911);
or U102 (N_102,In_860,In_581);
nand U103 (N_103,In_131,In_623);
nor U104 (N_104,In_215,In_92);
and U105 (N_105,In_407,In_440);
nand U106 (N_106,In_698,In_914);
or U107 (N_107,In_16,In_805);
or U108 (N_108,In_937,In_449);
and U109 (N_109,In_402,In_858);
or U110 (N_110,In_695,In_188);
or U111 (N_111,In_465,In_11);
or U112 (N_112,In_106,In_702);
nand U113 (N_113,In_500,In_736);
and U114 (N_114,In_278,In_784);
or U115 (N_115,In_332,In_393);
nand U116 (N_116,In_364,In_30);
and U117 (N_117,In_879,In_61);
nor U118 (N_118,In_552,In_200);
and U119 (N_119,In_783,In_284);
nor U120 (N_120,In_22,In_950);
nand U121 (N_121,In_599,In_262);
nand U122 (N_122,In_960,In_520);
nand U123 (N_123,In_416,In_428);
and U124 (N_124,In_789,In_953);
or U125 (N_125,In_957,In_903);
or U126 (N_126,In_489,In_883);
nor U127 (N_127,In_399,In_565);
and U128 (N_128,In_872,In_646);
nor U129 (N_129,In_60,In_165);
nand U130 (N_130,In_424,In_542);
or U131 (N_131,In_441,In_39);
nand U132 (N_132,In_954,In_930);
nor U133 (N_133,In_870,In_466);
nor U134 (N_134,In_65,In_596);
nor U135 (N_135,In_759,In_132);
nor U136 (N_136,In_323,In_866);
or U137 (N_137,In_630,In_90);
nor U138 (N_138,In_902,In_423);
nor U139 (N_139,In_383,In_877);
or U140 (N_140,In_808,In_98);
or U141 (N_141,In_182,In_367);
nand U142 (N_142,In_584,In_842);
nor U143 (N_143,In_72,In_915);
or U144 (N_144,In_797,In_335);
nand U145 (N_145,In_817,In_778);
or U146 (N_146,In_158,In_199);
nand U147 (N_147,In_636,In_229);
nor U148 (N_148,In_781,In_270);
and U149 (N_149,In_569,In_195);
nand U150 (N_150,In_613,In_824);
and U151 (N_151,In_69,In_198);
nor U152 (N_152,In_264,In_622);
and U153 (N_153,In_174,In_443);
nor U154 (N_154,In_8,In_744);
or U155 (N_155,In_603,In_925);
or U156 (N_156,In_799,In_594);
or U157 (N_157,In_287,In_286);
nand U158 (N_158,In_776,In_807);
nand U159 (N_159,In_791,In_446);
and U160 (N_160,In_551,In_514);
or U161 (N_161,In_526,In_617);
or U162 (N_162,In_255,In_437);
and U163 (N_163,In_760,In_486);
nor U164 (N_164,In_927,In_389);
nor U165 (N_165,In_285,In_863);
or U166 (N_166,In_600,In_249);
nor U167 (N_167,In_179,In_58);
nand U168 (N_168,In_222,In_48);
nor U169 (N_169,In_855,In_978);
or U170 (N_170,In_942,In_463);
and U171 (N_171,In_715,In_460);
or U172 (N_172,In_485,In_59);
nand U173 (N_173,In_172,In_624);
nor U174 (N_174,In_273,In_492);
nand U175 (N_175,In_697,In_109);
or U176 (N_176,In_220,In_157);
nor U177 (N_177,In_811,In_888);
and U178 (N_178,In_177,In_49);
or U179 (N_179,In_762,In_794);
nand U180 (N_180,In_924,In_88);
nand U181 (N_181,In_757,In_480);
and U182 (N_182,In_368,In_397);
and U183 (N_183,In_196,In_205);
and U184 (N_184,In_15,In_120);
nor U185 (N_185,In_244,In_539);
and U186 (N_186,In_793,In_409);
and U187 (N_187,In_769,In_462);
nand U188 (N_188,In_962,In_202);
or U189 (N_189,In_366,In_162);
nand U190 (N_190,In_537,In_191);
and U191 (N_191,In_309,In_515);
nand U192 (N_192,In_959,In_828);
nor U193 (N_193,In_607,In_729);
or U194 (N_194,In_295,In_904);
nor U195 (N_195,In_216,In_78);
nand U196 (N_196,In_331,In_668);
nand U197 (N_197,In_261,In_371);
xor U198 (N_198,In_71,In_345);
nand U199 (N_199,In_792,In_358);
nand U200 (N_200,In_365,In_153);
and U201 (N_201,In_629,In_431);
and U202 (N_202,In_563,In_19);
nor U203 (N_203,In_710,In_742);
and U204 (N_204,In_766,In_475);
nand U205 (N_205,In_502,In_703);
and U206 (N_206,In_493,In_576);
and U207 (N_207,In_38,In_898);
and U208 (N_208,In_496,In_943);
nor U209 (N_209,In_895,In_722);
or U210 (N_210,In_528,In_517);
and U211 (N_211,In_490,In_823);
nor U212 (N_212,In_655,In_356);
or U213 (N_213,In_574,In_300);
and U214 (N_214,In_31,In_144);
or U215 (N_215,In_250,In_43);
and U216 (N_216,In_684,In_140);
nor U217 (N_217,In_102,In_881);
and U218 (N_218,In_693,In_818);
and U219 (N_219,In_118,In_730);
and U220 (N_220,In_451,In_798);
and U221 (N_221,In_82,In_901);
or U222 (N_222,In_175,In_737);
and U223 (N_223,In_267,In_931);
nand U224 (N_224,In_339,In_361);
nor U225 (N_225,In_457,In_593);
and U226 (N_226,In_235,In_46);
nor U227 (N_227,In_966,In_932);
nor U228 (N_228,In_839,In_614);
or U229 (N_229,In_998,In_859);
and U230 (N_230,In_561,In_686);
and U231 (N_231,In_377,In_748);
xor U232 (N_232,In_427,In_647);
nand U233 (N_233,In_846,In_982);
nand U234 (N_234,In_787,In_310);
and U235 (N_235,In_105,In_768);
or U236 (N_236,In_474,In_13);
nand U237 (N_237,In_974,In_675);
nand U238 (N_238,In_7,In_248);
or U239 (N_239,In_935,In_920);
or U240 (N_240,In_166,In_219);
or U241 (N_241,In_277,In_94);
or U242 (N_242,In_861,In_327);
and U243 (N_243,In_403,In_50);
nor U244 (N_244,In_307,In_1);
nand U245 (N_245,In_346,In_832);
or U246 (N_246,In_148,In_100);
and U247 (N_247,In_311,In_592);
nand U248 (N_248,In_591,In_292);
and U249 (N_249,In_601,In_360);
nor U250 (N_250,In_302,In_447);
nand U251 (N_251,In_155,In_136);
or U252 (N_252,In_404,In_25);
or U253 (N_253,In_204,In_874);
and U254 (N_254,In_279,In_679);
nand U255 (N_255,In_724,In_840);
and U256 (N_256,In_193,In_35);
nand U257 (N_257,In_473,In_51);
and U258 (N_258,In_735,In_138);
and U259 (N_259,In_649,In_9);
and U260 (N_260,In_328,In_885);
nor U261 (N_261,In_271,In_812);
or U262 (N_262,In_240,In_964);
and U263 (N_263,In_876,In_926);
nor U264 (N_264,In_442,In_340);
or U265 (N_265,In_308,In_938);
nand U266 (N_266,In_648,In_108);
nor U267 (N_267,In_756,In_522);
and U268 (N_268,In_405,In_555);
nor U269 (N_269,In_304,In_983);
xor U270 (N_270,In_141,In_86);
and U271 (N_271,In_582,In_53);
nor U272 (N_272,In_408,In_170);
or U273 (N_273,In_816,In_232);
or U274 (N_274,In_909,In_588);
or U275 (N_275,In_272,In_129);
nand U276 (N_276,In_838,In_417);
nor U277 (N_277,In_868,In_682);
nand U278 (N_278,In_320,In_806);
or U279 (N_279,In_259,In_472);
nand U280 (N_280,In_280,In_590);
nor U281 (N_281,In_251,In_546);
nor U282 (N_282,In_936,In_513);
and U283 (N_283,In_706,In_545);
and U284 (N_284,In_711,In_436);
and U285 (N_285,In_875,In_767);
nor U286 (N_286,In_246,In_586);
and U287 (N_287,In_506,In_864);
nor U288 (N_288,In_362,In_343);
and U289 (N_289,In_33,In_572);
nor U290 (N_290,In_570,In_921);
nor U291 (N_291,In_751,In_687);
nor U292 (N_292,In_303,In_413);
nor U293 (N_293,In_324,In_226);
or U294 (N_294,In_438,In_87);
or U295 (N_295,In_281,In_115);
or U296 (N_296,In_247,In_627);
and U297 (N_297,In_544,In_678);
nor U298 (N_298,In_802,In_319);
nor U299 (N_299,In_143,In_334);
nor U300 (N_300,In_230,In_835);
nor U301 (N_301,In_81,In_605);
and U302 (N_302,In_207,In_602);
nand U303 (N_303,In_713,In_994);
nor U304 (N_304,In_833,In_521);
nand U305 (N_305,In_970,In_819);
nor U306 (N_306,In_529,In_354);
nor U307 (N_307,In_956,In_130);
nor U308 (N_308,In_161,In_663);
and U309 (N_309,In_439,In_37);
or U310 (N_310,In_681,In_236);
or U311 (N_311,In_732,In_567);
nor U312 (N_312,In_524,In_150);
or U313 (N_313,In_610,In_316);
xnor U314 (N_314,In_40,In_666);
nand U315 (N_315,In_315,In_900);
or U316 (N_316,In_836,In_907);
nor U317 (N_317,In_253,In_504);
or U318 (N_318,In_211,In_225);
xnor U319 (N_319,In_976,In_615);
nor U320 (N_320,In_882,In_26);
nand U321 (N_321,In_674,In_314);
nor U322 (N_322,In_896,In_352);
nand U323 (N_323,In_887,In_24);
nand U324 (N_324,In_206,In_386);
and U325 (N_325,In_980,In_77);
nor U326 (N_326,In_997,In_616);
and U327 (N_327,In_29,In_871);
nor U328 (N_328,In_126,In_644);
nand U329 (N_329,In_186,In_471);
and U330 (N_330,In_786,In_689);
nand U331 (N_331,In_2,In_979);
nor U332 (N_332,In_418,In_214);
or U333 (N_333,In_996,In_305);
nor U334 (N_334,In_712,In_645);
nor U335 (N_335,In_739,In_256);
or U336 (N_336,In_841,In_740);
nor U337 (N_337,In_42,In_425);
or U338 (N_338,In_434,In_322);
and U339 (N_339,In_27,In_714);
nor U340 (N_340,In_609,In_124);
or U341 (N_341,In_774,In_825);
nor U342 (N_342,In_243,In_680);
nor U343 (N_343,In_421,In_867);
or U344 (N_344,In_173,In_559);
nor U345 (N_345,In_971,In_116);
or U346 (N_346,In_830,In_844);
or U347 (N_347,In_755,In_683);
and U348 (N_348,In_564,In_992);
nor U349 (N_349,In_662,In_258);
nand U350 (N_350,In_497,In_951);
or U351 (N_351,In_483,In_160);
or U352 (N_352,In_910,In_197);
or U353 (N_353,In_213,In_928);
or U354 (N_354,In_967,In_420);
and U355 (N_355,In_355,In_531);
nor U356 (N_356,In_121,In_856);
nor U357 (N_357,In_123,In_139);
and U358 (N_358,In_660,In_958);
nor U359 (N_359,In_664,In_469);
and U360 (N_360,In_210,In_587);
or U361 (N_361,In_97,In_149);
nor U362 (N_362,In_192,In_464);
nand U363 (N_363,In_918,In_826);
nor U364 (N_364,In_163,In_290);
and U365 (N_365,In_543,In_254);
or U366 (N_366,In_387,In_282);
nand U367 (N_367,In_458,In_414);
and U368 (N_368,In_91,In_41);
nand U369 (N_369,In_333,In_549);
or U370 (N_370,In_595,In_445);
nor U371 (N_371,In_669,In_690);
and U372 (N_372,In_518,In_375);
nand U373 (N_373,In_494,In_571);
and U374 (N_374,In_491,In_95);
or U375 (N_375,In_917,In_478);
nand U376 (N_376,In_127,In_849);
and U377 (N_377,In_973,In_880);
or U378 (N_378,In_890,In_891);
or U379 (N_379,In_821,In_391);
and U380 (N_380,In_66,In_656);
or U381 (N_381,In_257,In_6);
nor U382 (N_382,In_773,In_837);
nor U383 (N_383,In_906,In_780);
or U384 (N_384,In_372,In_677);
or U385 (N_385,In_934,In_694);
or U386 (N_386,In_57,In_337);
or U387 (N_387,In_318,In_382);
or U388 (N_388,In_540,In_294);
and U389 (N_389,In_168,In_661);
nor U390 (N_390,In_154,In_301);
nand U391 (N_391,In_374,In_415);
and U392 (N_392,In_993,In_733);
or U393 (N_393,In_535,In_568);
nand U394 (N_394,In_541,In_412);
nand U395 (N_395,In_370,In_850);
nor U396 (N_396,In_658,In_237);
nor U397 (N_397,In_185,In_498);
or U398 (N_398,In_122,In_275);
or U399 (N_399,In_530,In_176);
and U400 (N_400,In_558,In_525);
nor U401 (N_401,In_548,In_10);
or U402 (N_402,In_865,In_889);
nor U403 (N_403,In_813,In_344);
nor U404 (N_404,In_336,In_633);
nor U405 (N_405,In_263,In_608);
and U406 (N_406,In_782,In_621);
nand U407 (N_407,In_487,In_400);
nor U408 (N_408,In_357,In_948);
and U409 (N_409,In_164,In_589);
and U410 (N_410,In_699,In_884);
nor U411 (N_411,In_342,In_940);
nand U412 (N_412,In_991,In_822);
or U413 (N_413,In_184,In_265);
and U414 (N_414,In_17,In_96);
xor U415 (N_415,In_665,In_810);
nand U416 (N_416,In_376,In_338);
nand U417 (N_417,In_809,In_908);
and U418 (N_418,In_398,In_719);
or U419 (N_419,In_83,In_14);
nand U420 (N_420,In_125,In_44);
or U421 (N_421,In_988,In_159);
nand U422 (N_422,In_135,In_635);
nand U423 (N_423,In_455,In_45);
xnor U424 (N_424,In_146,In_119);
and U425 (N_425,In_167,In_718);
or U426 (N_426,In_507,In_426);
or U427 (N_427,In_831,In_503);
or U428 (N_428,In_401,In_76);
nand U429 (N_429,In_228,In_853);
nand U430 (N_430,In_829,In_231);
nand U431 (N_431,In_134,In_291);
nor U432 (N_432,In_913,In_827);
nor U433 (N_433,In_351,In_717);
or U434 (N_434,In_795,In_527);
nand U435 (N_435,In_260,In_353);
nand U436 (N_436,In_509,In_708);
and U437 (N_437,In_854,In_101);
and U438 (N_438,In_631,In_857);
or U439 (N_439,In_481,In_152);
and U440 (N_440,In_208,In_984);
nor U441 (N_441,In_499,In_276);
and U442 (N_442,In_508,In_968);
and U443 (N_443,In_707,In_758);
or U444 (N_444,In_114,In_606);
nor U445 (N_445,In_313,In_598);
and U446 (N_446,In_894,In_692);
and U447 (N_447,In_788,In_848);
nand U448 (N_448,In_117,In_369);
and U449 (N_449,In_238,In_604);
and U450 (N_450,In_667,In_752);
or U451 (N_451,In_941,In_671);
nand U452 (N_452,In_512,In_560);
and U453 (N_453,In_700,In_245);
nor U454 (N_454,In_171,In_34);
nor U455 (N_455,In_704,In_922);
or U456 (N_456,In_432,In_696);
and U457 (N_457,In_716,In_349);
and U458 (N_458,In_221,In_456);
and U459 (N_459,In_312,In_691);
xnor U460 (N_460,In_74,In_209);
or U461 (N_461,In_761,In_111);
nand U462 (N_462,In_800,In_637);
nand U463 (N_463,In_63,In_363);
nand U464 (N_464,In_55,In_743);
or U465 (N_465,In_511,In_274);
nand U466 (N_466,In_990,In_189);
and U467 (N_467,In_297,In_741);
nor U468 (N_468,In_411,In_296);
nor U469 (N_469,In_373,In_820);
and U470 (N_470,In_422,In_450);
nand U471 (N_471,In_75,In_939);
nor U472 (N_472,In_390,In_224);
nand U473 (N_473,In_944,In_488);
nand U474 (N_474,In_659,In_611);
or U475 (N_475,In_929,In_505);
and U476 (N_476,In_288,In_672);
nand U477 (N_477,In_999,In_919);
nor U478 (N_478,In_538,In_749);
nand U479 (N_479,In_477,In_573);
nor U480 (N_480,In_834,In_5);
or U481 (N_481,In_803,In_223);
or U482 (N_482,In_772,In_556);
and U483 (N_483,In_21,In_705);
or U484 (N_484,In_113,In_468);
and U485 (N_485,In_657,In_804);
or U486 (N_486,In_495,In_128);
nor U487 (N_487,In_685,In_142);
nand U488 (N_488,In_85,In_252);
nor U489 (N_489,In_147,In_532);
nor U490 (N_490,In_347,In_107);
or U491 (N_491,In_995,In_137);
nor U492 (N_492,In_955,In_452);
nor U493 (N_493,In_945,In_947);
nand U494 (N_494,In_151,In_723);
nor U495 (N_495,In_536,In_905);
or U496 (N_496,In_218,In_110);
and U497 (N_497,In_754,In_242);
or U498 (N_498,In_643,In_847);
or U499 (N_499,In_217,In_461);
nand U500 (N_500,In_743,In_2);
nand U501 (N_501,In_615,In_51);
or U502 (N_502,In_974,In_706);
and U503 (N_503,In_497,In_43);
nor U504 (N_504,In_350,In_567);
nand U505 (N_505,In_734,In_541);
or U506 (N_506,In_391,In_231);
nor U507 (N_507,In_951,In_478);
nor U508 (N_508,In_771,In_104);
or U509 (N_509,In_660,In_602);
nor U510 (N_510,In_344,In_489);
nor U511 (N_511,In_165,In_38);
nand U512 (N_512,In_737,In_107);
and U513 (N_513,In_19,In_700);
and U514 (N_514,In_707,In_775);
or U515 (N_515,In_389,In_826);
nor U516 (N_516,In_187,In_79);
nand U517 (N_517,In_654,In_863);
or U518 (N_518,In_690,In_803);
or U519 (N_519,In_31,In_864);
and U520 (N_520,In_833,In_109);
or U521 (N_521,In_312,In_705);
or U522 (N_522,In_117,In_63);
nand U523 (N_523,In_969,In_18);
nand U524 (N_524,In_837,In_370);
nor U525 (N_525,In_51,In_204);
or U526 (N_526,In_326,In_50);
nand U527 (N_527,In_418,In_727);
and U528 (N_528,In_144,In_298);
nor U529 (N_529,In_666,In_511);
and U530 (N_530,In_611,In_648);
xor U531 (N_531,In_410,In_782);
and U532 (N_532,In_901,In_144);
or U533 (N_533,In_306,In_678);
nand U534 (N_534,In_337,In_501);
or U535 (N_535,In_93,In_123);
nor U536 (N_536,In_781,In_660);
nor U537 (N_537,In_644,In_623);
xnor U538 (N_538,In_631,In_100);
and U539 (N_539,In_363,In_595);
and U540 (N_540,In_95,In_875);
and U541 (N_541,In_530,In_919);
or U542 (N_542,In_909,In_289);
nor U543 (N_543,In_516,In_716);
nand U544 (N_544,In_809,In_424);
and U545 (N_545,In_749,In_62);
nand U546 (N_546,In_901,In_745);
nand U547 (N_547,In_517,In_91);
nand U548 (N_548,In_134,In_462);
nand U549 (N_549,In_827,In_265);
nor U550 (N_550,In_432,In_726);
and U551 (N_551,In_962,In_592);
nor U552 (N_552,In_678,In_496);
nand U553 (N_553,In_801,In_642);
nor U554 (N_554,In_385,In_634);
nand U555 (N_555,In_834,In_636);
nand U556 (N_556,In_467,In_870);
nand U557 (N_557,In_152,In_124);
or U558 (N_558,In_125,In_134);
and U559 (N_559,In_617,In_727);
or U560 (N_560,In_952,In_782);
nand U561 (N_561,In_220,In_47);
nor U562 (N_562,In_137,In_673);
or U563 (N_563,In_571,In_26);
or U564 (N_564,In_442,In_969);
nand U565 (N_565,In_193,In_275);
nand U566 (N_566,In_338,In_275);
or U567 (N_567,In_927,In_961);
nor U568 (N_568,In_230,In_957);
or U569 (N_569,In_933,In_109);
or U570 (N_570,In_740,In_748);
nor U571 (N_571,In_344,In_697);
nor U572 (N_572,In_516,In_315);
nor U573 (N_573,In_455,In_423);
and U574 (N_574,In_907,In_793);
and U575 (N_575,In_904,In_828);
or U576 (N_576,In_500,In_323);
nand U577 (N_577,In_795,In_87);
nand U578 (N_578,In_74,In_298);
nor U579 (N_579,In_735,In_205);
nand U580 (N_580,In_894,In_19);
nand U581 (N_581,In_143,In_319);
and U582 (N_582,In_282,In_193);
and U583 (N_583,In_965,In_437);
or U584 (N_584,In_58,In_782);
nor U585 (N_585,In_124,In_471);
nand U586 (N_586,In_48,In_341);
nand U587 (N_587,In_144,In_400);
nor U588 (N_588,In_918,In_792);
or U589 (N_589,In_982,In_871);
nor U590 (N_590,In_380,In_1);
or U591 (N_591,In_200,In_570);
nand U592 (N_592,In_253,In_139);
nor U593 (N_593,In_339,In_210);
nand U594 (N_594,In_102,In_321);
nand U595 (N_595,In_535,In_845);
nor U596 (N_596,In_904,In_625);
and U597 (N_597,In_311,In_831);
nand U598 (N_598,In_219,In_820);
and U599 (N_599,In_5,In_278);
nand U600 (N_600,In_768,In_142);
nor U601 (N_601,In_787,In_356);
and U602 (N_602,In_56,In_11);
nand U603 (N_603,In_30,In_611);
and U604 (N_604,In_102,In_997);
nand U605 (N_605,In_625,In_681);
and U606 (N_606,In_397,In_469);
nand U607 (N_607,In_840,In_228);
nand U608 (N_608,In_919,In_282);
nand U609 (N_609,In_883,In_543);
nand U610 (N_610,In_810,In_700);
nand U611 (N_611,In_885,In_627);
nand U612 (N_612,In_270,In_523);
nand U613 (N_613,In_655,In_603);
or U614 (N_614,In_158,In_714);
nand U615 (N_615,In_449,In_158);
nand U616 (N_616,In_93,In_346);
and U617 (N_617,In_204,In_95);
and U618 (N_618,In_306,In_793);
and U619 (N_619,In_615,In_423);
and U620 (N_620,In_383,In_614);
nor U621 (N_621,In_957,In_40);
nor U622 (N_622,In_742,In_404);
nand U623 (N_623,In_379,In_873);
nand U624 (N_624,In_875,In_922);
and U625 (N_625,In_774,In_369);
nand U626 (N_626,In_498,In_779);
nor U627 (N_627,In_409,In_231);
or U628 (N_628,In_879,In_533);
nor U629 (N_629,In_689,In_852);
or U630 (N_630,In_142,In_510);
nor U631 (N_631,In_873,In_825);
nand U632 (N_632,In_446,In_387);
nand U633 (N_633,In_445,In_919);
xor U634 (N_634,In_284,In_505);
nor U635 (N_635,In_188,In_448);
or U636 (N_636,In_955,In_110);
nand U637 (N_637,In_378,In_416);
nor U638 (N_638,In_508,In_100);
nand U639 (N_639,In_662,In_873);
or U640 (N_640,In_11,In_580);
nor U641 (N_641,In_791,In_669);
nor U642 (N_642,In_225,In_899);
and U643 (N_643,In_305,In_412);
nor U644 (N_644,In_587,In_737);
or U645 (N_645,In_915,In_196);
or U646 (N_646,In_808,In_921);
nand U647 (N_647,In_839,In_785);
and U648 (N_648,In_551,In_678);
and U649 (N_649,In_203,In_313);
nor U650 (N_650,In_465,In_741);
and U651 (N_651,In_856,In_279);
or U652 (N_652,In_501,In_383);
nand U653 (N_653,In_402,In_678);
nand U654 (N_654,In_708,In_914);
or U655 (N_655,In_484,In_50);
nor U656 (N_656,In_512,In_844);
nor U657 (N_657,In_66,In_919);
and U658 (N_658,In_180,In_999);
and U659 (N_659,In_522,In_292);
or U660 (N_660,In_691,In_592);
nor U661 (N_661,In_302,In_111);
and U662 (N_662,In_493,In_304);
and U663 (N_663,In_138,In_675);
nor U664 (N_664,In_585,In_997);
nand U665 (N_665,In_320,In_688);
or U666 (N_666,In_887,In_374);
nand U667 (N_667,In_907,In_380);
nand U668 (N_668,In_255,In_828);
or U669 (N_669,In_333,In_547);
nor U670 (N_670,In_153,In_327);
and U671 (N_671,In_110,In_660);
nand U672 (N_672,In_331,In_399);
and U673 (N_673,In_215,In_468);
nor U674 (N_674,In_782,In_871);
or U675 (N_675,In_437,In_742);
nor U676 (N_676,In_693,In_30);
nor U677 (N_677,In_218,In_666);
and U678 (N_678,In_816,In_742);
nor U679 (N_679,In_688,In_382);
nor U680 (N_680,In_868,In_468);
nor U681 (N_681,In_882,In_450);
nand U682 (N_682,In_476,In_74);
and U683 (N_683,In_372,In_272);
or U684 (N_684,In_700,In_678);
or U685 (N_685,In_657,In_558);
and U686 (N_686,In_998,In_616);
and U687 (N_687,In_222,In_999);
nand U688 (N_688,In_249,In_621);
or U689 (N_689,In_134,In_580);
or U690 (N_690,In_785,In_569);
or U691 (N_691,In_392,In_567);
nor U692 (N_692,In_985,In_687);
xnor U693 (N_693,In_208,In_343);
nand U694 (N_694,In_405,In_530);
nor U695 (N_695,In_632,In_324);
or U696 (N_696,In_456,In_849);
and U697 (N_697,In_478,In_658);
or U698 (N_698,In_938,In_375);
or U699 (N_699,In_365,In_745);
and U700 (N_700,In_536,In_383);
and U701 (N_701,In_379,In_496);
or U702 (N_702,In_752,In_623);
nand U703 (N_703,In_37,In_278);
nand U704 (N_704,In_802,In_377);
and U705 (N_705,In_334,In_151);
nor U706 (N_706,In_656,In_144);
nor U707 (N_707,In_917,In_20);
nor U708 (N_708,In_273,In_252);
and U709 (N_709,In_394,In_823);
nand U710 (N_710,In_618,In_546);
and U711 (N_711,In_26,In_21);
and U712 (N_712,In_757,In_473);
or U713 (N_713,In_122,In_329);
nor U714 (N_714,In_359,In_143);
or U715 (N_715,In_783,In_381);
xnor U716 (N_716,In_407,In_49);
nor U717 (N_717,In_360,In_699);
nor U718 (N_718,In_482,In_435);
nor U719 (N_719,In_961,In_910);
nand U720 (N_720,In_673,In_868);
nand U721 (N_721,In_750,In_841);
or U722 (N_722,In_466,In_939);
nor U723 (N_723,In_550,In_989);
or U724 (N_724,In_810,In_151);
or U725 (N_725,In_219,In_991);
nand U726 (N_726,In_966,In_779);
and U727 (N_727,In_255,In_294);
nor U728 (N_728,In_189,In_735);
nand U729 (N_729,In_823,In_766);
or U730 (N_730,In_287,In_614);
and U731 (N_731,In_614,In_806);
nor U732 (N_732,In_196,In_202);
nand U733 (N_733,In_818,In_500);
and U734 (N_734,In_148,In_592);
nand U735 (N_735,In_605,In_556);
nand U736 (N_736,In_894,In_50);
and U737 (N_737,In_844,In_658);
nor U738 (N_738,In_169,In_55);
or U739 (N_739,In_943,In_461);
or U740 (N_740,In_805,In_65);
nand U741 (N_741,In_504,In_375);
nor U742 (N_742,In_217,In_403);
and U743 (N_743,In_465,In_178);
and U744 (N_744,In_417,In_681);
or U745 (N_745,In_411,In_266);
xor U746 (N_746,In_19,In_675);
nand U747 (N_747,In_884,In_33);
xnor U748 (N_748,In_305,In_14);
nor U749 (N_749,In_192,In_528);
and U750 (N_750,In_918,In_588);
and U751 (N_751,In_20,In_914);
nand U752 (N_752,In_116,In_400);
or U753 (N_753,In_427,In_757);
and U754 (N_754,In_896,In_506);
xor U755 (N_755,In_367,In_207);
and U756 (N_756,In_599,In_743);
nand U757 (N_757,In_834,In_11);
and U758 (N_758,In_537,In_883);
or U759 (N_759,In_6,In_337);
or U760 (N_760,In_3,In_445);
nand U761 (N_761,In_926,In_643);
xor U762 (N_762,In_311,In_579);
and U763 (N_763,In_26,In_460);
or U764 (N_764,In_788,In_25);
and U765 (N_765,In_698,In_737);
or U766 (N_766,In_7,In_860);
and U767 (N_767,In_469,In_993);
nand U768 (N_768,In_833,In_693);
or U769 (N_769,In_335,In_713);
or U770 (N_770,In_54,In_560);
or U771 (N_771,In_784,In_782);
nand U772 (N_772,In_609,In_416);
nand U773 (N_773,In_663,In_107);
nand U774 (N_774,In_477,In_562);
or U775 (N_775,In_841,In_382);
and U776 (N_776,In_204,In_133);
and U777 (N_777,In_688,In_531);
and U778 (N_778,In_427,In_860);
and U779 (N_779,In_158,In_373);
nor U780 (N_780,In_708,In_464);
and U781 (N_781,In_431,In_31);
and U782 (N_782,In_405,In_422);
or U783 (N_783,In_814,In_612);
nor U784 (N_784,In_569,In_638);
and U785 (N_785,In_558,In_207);
or U786 (N_786,In_640,In_570);
nor U787 (N_787,In_417,In_658);
or U788 (N_788,In_615,In_779);
or U789 (N_789,In_489,In_599);
or U790 (N_790,In_7,In_927);
xor U791 (N_791,In_217,In_970);
nand U792 (N_792,In_312,In_638);
and U793 (N_793,In_136,In_811);
nand U794 (N_794,In_462,In_655);
and U795 (N_795,In_256,In_855);
or U796 (N_796,In_147,In_392);
nor U797 (N_797,In_736,In_418);
nand U798 (N_798,In_391,In_547);
nor U799 (N_799,In_836,In_420);
and U800 (N_800,In_405,In_104);
or U801 (N_801,In_440,In_251);
nand U802 (N_802,In_281,In_785);
nor U803 (N_803,In_596,In_790);
or U804 (N_804,In_119,In_797);
and U805 (N_805,In_672,In_306);
nand U806 (N_806,In_503,In_174);
nand U807 (N_807,In_42,In_769);
nor U808 (N_808,In_431,In_753);
nor U809 (N_809,In_367,In_449);
and U810 (N_810,In_794,In_263);
or U811 (N_811,In_578,In_957);
xor U812 (N_812,In_540,In_633);
or U813 (N_813,In_738,In_510);
nor U814 (N_814,In_373,In_723);
or U815 (N_815,In_343,In_888);
or U816 (N_816,In_754,In_166);
nor U817 (N_817,In_921,In_615);
nand U818 (N_818,In_573,In_858);
nor U819 (N_819,In_18,In_236);
or U820 (N_820,In_347,In_401);
and U821 (N_821,In_992,In_322);
and U822 (N_822,In_17,In_982);
and U823 (N_823,In_197,In_997);
and U824 (N_824,In_646,In_4);
or U825 (N_825,In_730,In_354);
and U826 (N_826,In_562,In_539);
nand U827 (N_827,In_903,In_564);
or U828 (N_828,In_382,In_119);
or U829 (N_829,In_747,In_227);
nand U830 (N_830,In_133,In_363);
or U831 (N_831,In_391,In_746);
or U832 (N_832,In_539,In_267);
and U833 (N_833,In_341,In_163);
and U834 (N_834,In_402,In_901);
nor U835 (N_835,In_871,In_516);
or U836 (N_836,In_5,In_860);
nor U837 (N_837,In_479,In_95);
nor U838 (N_838,In_913,In_625);
nand U839 (N_839,In_549,In_411);
or U840 (N_840,In_552,In_276);
nand U841 (N_841,In_395,In_549);
or U842 (N_842,In_737,In_717);
nor U843 (N_843,In_858,In_691);
and U844 (N_844,In_488,In_160);
nor U845 (N_845,In_608,In_293);
nand U846 (N_846,In_311,In_361);
nand U847 (N_847,In_667,In_823);
or U848 (N_848,In_516,In_373);
nand U849 (N_849,In_914,In_595);
nor U850 (N_850,In_431,In_406);
xor U851 (N_851,In_626,In_538);
nor U852 (N_852,In_662,In_158);
nor U853 (N_853,In_943,In_777);
and U854 (N_854,In_417,In_541);
nor U855 (N_855,In_789,In_147);
nor U856 (N_856,In_452,In_382);
nor U857 (N_857,In_490,In_151);
nand U858 (N_858,In_613,In_330);
or U859 (N_859,In_792,In_278);
xor U860 (N_860,In_516,In_675);
nor U861 (N_861,In_318,In_500);
and U862 (N_862,In_754,In_857);
xor U863 (N_863,In_937,In_877);
and U864 (N_864,In_857,In_826);
or U865 (N_865,In_363,In_577);
and U866 (N_866,In_997,In_712);
and U867 (N_867,In_663,In_177);
and U868 (N_868,In_765,In_244);
or U869 (N_869,In_962,In_708);
xor U870 (N_870,In_570,In_239);
or U871 (N_871,In_350,In_429);
nand U872 (N_872,In_680,In_772);
nand U873 (N_873,In_560,In_399);
nand U874 (N_874,In_905,In_890);
nand U875 (N_875,In_691,In_582);
or U876 (N_876,In_332,In_241);
and U877 (N_877,In_114,In_278);
and U878 (N_878,In_792,In_144);
nand U879 (N_879,In_661,In_146);
or U880 (N_880,In_31,In_915);
and U881 (N_881,In_637,In_124);
nand U882 (N_882,In_297,In_595);
and U883 (N_883,In_399,In_364);
or U884 (N_884,In_423,In_957);
or U885 (N_885,In_796,In_278);
nand U886 (N_886,In_505,In_115);
xnor U887 (N_887,In_705,In_56);
nor U888 (N_888,In_79,In_939);
nor U889 (N_889,In_513,In_360);
or U890 (N_890,In_693,In_744);
and U891 (N_891,In_120,In_201);
nor U892 (N_892,In_157,In_341);
or U893 (N_893,In_792,In_63);
and U894 (N_894,In_770,In_121);
or U895 (N_895,In_671,In_685);
or U896 (N_896,In_10,In_373);
nor U897 (N_897,In_468,In_825);
or U898 (N_898,In_848,In_349);
and U899 (N_899,In_92,In_216);
and U900 (N_900,In_381,In_467);
and U901 (N_901,In_750,In_457);
and U902 (N_902,In_509,In_59);
nand U903 (N_903,In_477,In_306);
nor U904 (N_904,In_155,In_29);
nor U905 (N_905,In_477,In_889);
nor U906 (N_906,In_740,In_695);
or U907 (N_907,In_17,In_359);
or U908 (N_908,In_917,In_726);
and U909 (N_909,In_271,In_858);
nor U910 (N_910,In_706,In_670);
nand U911 (N_911,In_430,In_963);
and U912 (N_912,In_647,In_395);
or U913 (N_913,In_82,In_719);
and U914 (N_914,In_921,In_359);
or U915 (N_915,In_968,In_476);
nor U916 (N_916,In_855,In_22);
and U917 (N_917,In_106,In_856);
xor U918 (N_918,In_48,In_180);
nor U919 (N_919,In_310,In_308);
nor U920 (N_920,In_760,In_136);
nand U921 (N_921,In_774,In_633);
nor U922 (N_922,In_605,In_234);
and U923 (N_923,In_488,In_196);
and U924 (N_924,In_577,In_413);
and U925 (N_925,In_211,In_710);
and U926 (N_926,In_68,In_586);
and U927 (N_927,In_617,In_72);
nor U928 (N_928,In_279,In_839);
nor U929 (N_929,In_434,In_340);
or U930 (N_930,In_481,In_967);
and U931 (N_931,In_206,In_768);
or U932 (N_932,In_764,In_396);
or U933 (N_933,In_587,In_824);
and U934 (N_934,In_942,In_881);
nor U935 (N_935,In_954,In_918);
and U936 (N_936,In_695,In_372);
nand U937 (N_937,In_835,In_696);
nor U938 (N_938,In_854,In_94);
and U939 (N_939,In_72,In_433);
nor U940 (N_940,In_436,In_392);
and U941 (N_941,In_678,In_973);
nand U942 (N_942,In_359,In_530);
nand U943 (N_943,In_92,In_340);
nand U944 (N_944,In_819,In_781);
or U945 (N_945,In_664,In_189);
and U946 (N_946,In_611,In_567);
and U947 (N_947,In_207,In_561);
or U948 (N_948,In_325,In_326);
and U949 (N_949,In_187,In_536);
or U950 (N_950,In_779,In_163);
or U951 (N_951,In_20,In_967);
or U952 (N_952,In_932,In_174);
and U953 (N_953,In_869,In_364);
nor U954 (N_954,In_28,In_435);
and U955 (N_955,In_277,In_65);
xnor U956 (N_956,In_145,In_732);
or U957 (N_957,In_792,In_609);
nand U958 (N_958,In_185,In_219);
nor U959 (N_959,In_91,In_12);
xor U960 (N_960,In_95,In_354);
nor U961 (N_961,In_121,In_167);
or U962 (N_962,In_148,In_733);
nand U963 (N_963,In_473,In_107);
nor U964 (N_964,In_614,In_195);
or U965 (N_965,In_85,In_289);
nand U966 (N_966,In_565,In_175);
or U967 (N_967,In_716,In_358);
xnor U968 (N_968,In_453,In_86);
and U969 (N_969,In_696,In_839);
xnor U970 (N_970,In_67,In_624);
or U971 (N_971,In_155,In_418);
or U972 (N_972,In_569,In_965);
or U973 (N_973,In_161,In_341);
and U974 (N_974,In_749,In_665);
and U975 (N_975,In_73,In_530);
or U976 (N_976,In_852,In_693);
nand U977 (N_977,In_769,In_666);
nand U978 (N_978,In_821,In_321);
nor U979 (N_979,In_926,In_708);
nor U980 (N_980,In_94,In_250);
and U981 (N_981,In_509,In_601);
and U982 (N_982,In_996,In_69);
nor U983 (N_983,In_389,In_306);
nand U984 (N_984,In_553,In_948);
and U985 (N_985,In_249,In_268);
nor U986 (N_986,In_328,In_315);
and U987 (N_987,In_387,In_547);
nor U988 (N_988,In_473,In_836);
or U989 (N_989,In_55,In_343);
or U990 (N_990,In_273,In_971);
and U991 (N_991,In_12,In_722);
or U992 (N_992,In_522,In_755);
nor U993 (N_993,In_769,In_461);
nor U994 (N_994,In_550,In_29);
xor U995 (N_995,In_470,In_341);
and U996 (N_996,In_804,In_904);
and U997 (N_997,In_56,In_795);
or U998 (N_998,In_683,In_889);
and U999 (N_999,In_239,In_201);
and U1000 (N_1000,N_683,N_691);
or U1001 (N_1001,N_820,N_581);
nand U1002 (N_1002,N_770,N_279);
nand U1003 (N_1003,N_870,N_397);
nor U1004 (N_1004,N_71,N_185);
and U1005 (N_1005,N_917,N_126);
nand U1006 (N_1006,N_408,N_863);
and U1007 (N_1007,N_573,N_218);
and U1008 (N_1008,N_231,N_767);
or U1009 (N_1009,N_757,N_862);
nor U1010 (N_1010,N_455,N_68);
and U1011 (N_1011,N_591,N_109);
or U1012 (N_1012,N_626,N_749);
nor U1013 (N_1013,N_611,N_561);
nor U1014 (N_1014,N_336,N_739);
or U1015 (N_1015,N_528,N_79);
or U1016 (N_1016,N_592,N_969);
or U1017 (N_1017,N_681,N_298);
nand U1018 (N_1018,N_213,N_253);
nand U1019 (N_1019,N_388,N_518);
or U1020 (N_1020,N_857,N_539);
nor U1021 (N_1021,N_814,N_574);
and U1022 (N_1022,N_610,N_278);
nand U1023 (N_1023,N_792,N_785);
nand U1024 (N_1024,N_532,N_210);
nand U1025 (N_1025,N_429,N_4);
nand U1026 (N_1026,N_108,N_311);
nand U1027 (N_1027,N_540,N_215);
nor U1028 (N_1028,N_300,N_329);
or U1029 (N_1029,N_982,N_341);
and U1030 (N_1030,N_503,N_3);
nor U1031 (N_1031,N_477,N_419);
nand U1032 (N_1032,N_986,N_238);
nor U1033 (N_1033,N_209,N_149);
nor U1034 (N_1034,N_122,N_617);
xnor U1035 (N_1035,N_76,N_779);
nor U1036 (N_1036,N_967,N_99);
and U1037 (N_1037,N_956,N_993);
and U1038 (N_1038,N_933,N_346);
nor U1039 (N_1039,N_884,N_551);
nor U1040 (N_1040,N_661,N_54);
nor U1041 (N_1041,N_392,N_506);
nor U1042 (N_1042,N_468,N_698);
and U1043 (N_1043,N_51,N_663);
xor U1044 (N_1044,N_643,N_138);
and U1045 (N_1045,N_112,N_297);
nand U1046 (N_1046,N_671,N_143);
and U1047 (N_1047,N_930,N_886);
nand U1048 (N_1048,N_555,N_47);
nand U1049 (N_1049,N_239,N_564);
nand U1050 (N_1050,N_970,N_685);
nand U1051 (N_1051,N_296,N_858);
or U1052 (N_1052,N_438,N_708);
nor U1053 (N_1053,N_487,N_376);
or U1054 (N_1054,N_189,N_22);
or U1055 (N_1055,N_908,N_235);
nor U1056 (N_1056,N_77,N_976);
nor U1057 (N_1057,N_495,N_905);
nand U1058 (N_1058,N_630,N_474);
or U1059 (N_1059,N_491,N_773);
or U1060 (N_1060,N_451,N_276);
or U1061 (N_1061,N_489,N_403);
or U1062 (N_1062,N_601,N_576);
or U1063 (N_1063,N_326,N_406);
and U1064 (N_1064,N_174,N_263);
or U1065 (N_1065,N_306,N_843);
nand U1066 (N_1066,N_224,N_724);
or U1067 (N_1067,N_614,N_777);
nand U1068 (N_1068,N_851,N_650);
nor U1069 (N_1069,N_281,N_507);
and U1070 (N_1070,N_828,N_699);
and U1071 (N_1071,N_736,N_778);
nand U1072 (N_1072,N_395,N_499);
and U1073 (N_1073,N_742,N_965);
and U1074 (N_1074,N_497,N_319);
or U1075 (N_1075,N_890,N_52);
nand U1076 (N_1076,N_554,N_398);
and U1077 (N_1077,N_712,N_620);
nor U1078 (N_1078,N_330,N_173);
or U1079 (N_1079,N_184,N_415);
nand U1080 (N_1080,N_791,N_286);
and U1081 (N_1081,N_937,N_822);
or U1082 (N_1082,N_120,N_316);
or U1083 (N_1083,N_864,N_715);
nand U1084 (N_1084,N_125,N_135);
nand U1085 (N_1085,N_145,N_478);
nor U1086 (N_1086,N_918,N_457);
or U1087 (N_1087,N_60,N_467);
nor U1088 (N_1088,N_84,N_42);
nor U1089 (N_1089,N_168,N_810);
and U1090 (N_1090,N_705,N_729);
nor U1091 (N_1091,N_277,N_413);
nand U1092 (N_1092,N_394,N_803);
nor U1093 (N_1093,N_565,N_25);
or U1094 (N_1094,N_404,N_385);
nand U1095 (N_1095,N_389,N_517);
nand U1096 (N_1096,N_764,N_290);
nor U1097 (N_1097,N_898,N_377);
xnor U1098 (N_1098,N_202,N_740);
nand U1099 (N_1099,N_492,N_984);
or U1100 (N_1100,N_807,N_575);
and U1101 (N_1101,N_343,N_19);
nor U1102 (N_1102,N_544,N_134);
and U1103 (N_1103,N_267,N_312);
or U1104 (N_1104,N_6,N_14);
nor U1105 (N_1105,N_957,N_934);
nor U1106 (N_1106,N_694,N_131);
and U1107 (N_1107,N_496,N_310);
nand U1108 (N_1108,N_436,N_571);
nor U1109 (N_1109,N_465,N_802);
and U1110 (N_1110,N_883,N_827);
nor U1111 (N_1111,N_966,N_292);
nand U1112 (N_1112,N_721,N_763);
or U1113 (N_1113,N_5,N_693);
nor U1114 (N_1114,N_282,N_473);
or U1115 (N_1115,N_268,N_205);
nand U1116 (N_1116,N_747,N_222);
nor U1117 (N_1117,N_625,N_157);
nand U1118 (N_1118,N_470,N_445);
and U1119 (N_1119,N_686,N_954);
nor U1120 (N_1120,N_680,N_391);
nand U1121 (N_1121,N_417,N_755);
nor U1122 (N_1122,N_10,N_83);
and U1123 (N_1123,N_647,N_488);
and U1124 (N_1124,N_999,N_775);
nand U1125 (N_1125,N_628,N_593);
or U1126 (N_1126,N_874,N_946);
and U1127 (N_1127,N_896,N_16);
nor U1128 (N_1128,N_887,N_771);
or U1129 (N_1129,N_633,N_494);
nand U1130 (N_1130,N_59,N_711);
or U1131 (N_1131,N_962,N_968);
nor U1132 (N_1132,N_677,N_524);
nand U1133 (N_1133,N_483,N_362);
and U1134 (N_1134,N_587,N_247);
and U1135 (N_1135,N_817,N_20);
xor U1136 (N_1136,N_212,N_922);
or U1137 (N_1137,N_270,N_948);
nor U1138 (N_1138,N_550,N_204);
and U1139 (N_1139,N_166,N_261);
or U1140 (N_1140,N_45,N_796);
and U1141 (N_1141,N_955,N_910);
nand U1142 (N_1142,N_912,N_439);
nand U1143 (N_1143,N_180,N_61);
and U1144 (N_1144,N_427,N_746);
and U1145 (N_1145,N_104,N_974);
and U1146 (N_1146,N_370,N_865);
nor U1147 (N_1147,N_196,N_776);
nor U1148 (N_1148,N_615,N_12);
or U1149 (N_1149,N_265,N_878);
or U1150 (N_1150,N_903,N_602);
nor U1151 (N_1151,N_859,N_527);
nand U1152 (N_1152,N_836,N_635);
and U1153 (N_1153,N_97,N_481);
and U1154 (N_1154,N_769,N_242);
nor U1155 (N_1155,N_510,N_246);
nor U1156 (N_1156,N_65,N_752);
and U1157 (N_1157,N_228,N_977);
or U1158 (N_1158,N_605,N_735);
or U1159 (N_1159,N_823,N_325);
nor U1160 (N_1160,N_381,N_283);
or U1161 (N_1161,N_351,N_293);
and U1162 (N_1162,N_502,N_162);
xnor U1163 (N_1163,N_287,N_689);
or U1164 (N_1164,N_280,N_295);
nor U1165 (N_1165,N_207,N_784);
and U1166 (N_1166,N_525,N_37);
nand U1167 (N_1167,N_328,N_501);
nand U1168 (N_1168,N_713,N_257);
nand U1169 (N_1169,N_35,N_841);
or U1170 (N_1170,N_288,N_372);
and U1171 (N_1171,N_0,N_386);
and U1172 (N_1172,N_416,N_687);
or U1173 (N_1173,N_93,N_916);
nand U1174 (N_1174,N_217,N_155);
nand U1175 (N_1175,N_349,N_678);
and U1176 (N_1176,N_98,N_696);
or U1177 (N_1177,N_396,N_367);
nand U1178 (N_1178,N_294,N_938);
nand U1179 (N_1179,N_106,N_923);
or U1180 (N_1180,N_214,N_707);
nand U1181 (N_1181,N_33,N_612);
nor U1182 (N_1182,N_197,N_556);
and U1183 (N_1183,N_873,N_432);
and U1184 (N_1184,N_78,N_774);
and U1185 (N_1185,N_623,N_806);
nand U1186 (N_1186,N_179,N_758);
nand U1187 (N_1187,N_975,N_275);
or U1188 (N_1188,N_485,N_412);
or U1189 (N_1189,N_819,N_359);
and U1190 (N_1190,N_500,N_291);
nand U1191 (N_1191,N_949,N_273);
nand U1192 (N_1192,N_718,N_34);
or U1193 (N_1193,N_9,N_460);
nor U1194 (N_1194,N_100,N_855);
nand U1195 (N_1195,N_659,N_833);
nor U1196 (N_1196,N_94,N_355);
and U1197 (N_1197,N_219,N_759);
nand U1198 (N_1198,N_632,N_240);
and U1199 (N_1199,N_195,N_657);
nor U1200 (N_1200,N_165,N_943);
nor U1201 (N_1201,N_289,N_352);
xnor U1202 (N_1202,N_900,N_43);
nand U1203 (N_1203,N_915,N_842);
and U1204 (N_1204,N_921,N_236);
nor U1205 (N_1205,N_868,N_813);
nand U1206 (N_1206,N_563,N_658);
nor U1207 (N_1207,N_304,N_622);
nand U1208 (N_1208,N_941,N_546);
and U1209 (N_1209,N_461,N_449);
nand U1210 (N_1210,N_375,N_636);
and U1211 (N_1211,N_244,N_118);
or U1212 (N_1212,N_357,N_899);
nor U1213 (N_1213,N_484,N_24);
or U1214 (N_1214,N_644,N_353);
or U1215 (N_1215,N_760,N_92);
nor U1216 (N_1216,N_672,N_904);
nand U1217 (N_1217,N_191,N_728);
and U1218 (N_1218,N_651,N_631);
nand U1219 (N_1219,N_988,N_324);
and U1220 (N_1220,N_660,N_299);
nand U1221 (N_1221,N_285,N_80);
and U1222 (N_1222,N_598,N_251);
nor U1223 (N_1223,N_271,N_688);
nor U1224 (N_1224,N_199,N_766);
nand U1225 (N_1225,N_666,N_725);
xnor U1226 (N_1226,N_137,N_942);
nor U1227 (N_1227,N_256,N_880);
nor U1228 (N_1228,N_545,N_566);
or U1229 (N_1229,N_69,N_882);
nor U1230 (N_1230,N_704,N_454);
and U1231 (N_1231,N_66,N_72);
nor U1232 (N_1232,N_74,N_327);
nor U1233 (N_1233,N_211,N_164);
nor U1234 (N_1234,N_272,N_221);
nor U1235 (N_1235,N_676,N_318);
nor U1236 (N_1236,N_365,N_136);
nand U1237 (N_1237,N_669,N_642);
nor U1238 (N_1238,N_800,N_875);
or U1239 (N_1239,N_453,N_837);
or U1240 (N_1240,N_861,N_992);
or U1241 (N_1241,N_552,N_613);
and U1242 (N_1242,N_241,N_85);
and U1243 (N_1243,N_579,N_714);
and U1244 (N_1244,N_609,N_81);
nor U1245 (N_1245,N_692,N_719);
nor U1246 (N_1246,N_32,N_547);
nand U1247 (N_1247,N_110,N_153);
nand U1248 (N_1248,N_315,N_849);
and U1249 (N_1249,N_490,N_744);
nor U1250 (N_1250,N_382,N_405);
or U1251 (N_1251,N_102,N_682);
nand U1252 (N_1252,N_462,N_600);
nand U1253 (N_1253,N_114,N_424);
or U1254 (N_1254,N_789,N_804);
and U1255 (N_1255,N_369,N_604);
nor U1256 (N_1256,N_876,N_437);
xnor U1257 (N_1257,N_640,N_529);
nand U1258 (N_1258,N_331,N_846);
or U1259 (N_1259,N_535,N_701);
xnor U1260 (N_1260,N_472,N_508);
nor U1261 (N_1261,N_393,N_542);
nand U1262 (N_1262,N_834,N_146);
nand U1263 (N_1263,N_727,N_765);
or U1264 (N_1264,N_818,N_379);
nand U1265 (N_1265,N_139,N_914);
nor U1266 (N_1266,N_232,N_901);
nand U1267 (N_1267,N_50,N_892);
and U1268 (N_1268,N_505,N_509);
and U1269 (N_1269,N_307,N_401);
nor U1270 (N_1270,N_249,N_549);
and U1271 (N_1271,N_538,N_562);
nand U1272 (N_1272,N_730,N_313);
nand U1273 (N_1273,N_321,N_407);
or U1274 (N_1274,N_128,N_426);
or U1275 (N_1275,N_801,N_486);
nor U1276 (N_1276,N_44,N_226);
nor U1277 (N_1277,N_772,N_38);
nor U1278 (N_1278,N_578,N_332);
or U1279 (N_1279,N_754,N_710);
nor U1280 (N_1280,N_891,N_595);
and U1281 (N_1281,N_384,N_374);
and U1282 (N_1282,N_649,N_981);
nor U1283 (N_1283,N_568,N_751);
nor U1284 (N_1284,N_808,N_638);
nor U1285 (N_1285,N_302,N_936);
nand U1286 (N_1286,N_839,N_284);
nor U1287 (N_1287,N_743,N_464);
and U1288 (N_1288,N_932,N_266);
and U1289 (N_1289,N_28,N_963);
or U1290 (N_1290,N_323,N_906);
or U1291 (N_1291,N_414,N_926);
nand U1292 (N_1292,N_62,N_848);
nand U1293 (N_1293,N_952,N_991);
nor U1294 (N_1294,N_201,N_703);
nand U1295 (N_1295,N_459,N_619);
or U1296 (N_1296,N_252,N_373);
or U1297 (N_1297,N_980,N_190);
nand U1298 (N_1298,N_171,N_186);
and U1299 (N_1299,N_230,N_31);
nand U1300 (N_1300,N_867,N_223);
nand U1301 (N_1301,N_334,N_216);
and U1302 (N_1302,N_360,N_151);
or U1303 (N_1303,N_584,N_428);
or U1304 (N_1304,N_21,N_700);
and U1305 (N_1305,N_142,N_193);
nor U1306 (N_1306,N_103,N_96);
or U1307 (N_1307,N_243,N_260);
nor U1308 (N_1308,N_192,N_141);
and U1309 (N_1309,N_183,N_86);
and U1310 (N_1310,N_537,N_964);
or U1311 (N_1311,N_788,N_148);
or U1312 (N_1312,N_795,N_152);
and U1313 (N_1313,N_130,N_987);
or U1314 (N_1314,N_452,N_440);
or U1315 (N_1315,N_673,N_378);
nor U1316 (N_1316,N_902,N_826);
nand U1317 (N_1317,N_732,N_522);
nor U1318 (N_1318,N_668,N_569);
nand U1319 (N_1319,N_198,N_953);
nor U1320 (N_1320,N_175,N_911);
and U1321 (N_1321,N_782,N_410);
or U1322 (N_1322,N_511,N_940);
nor U1323 (N_1323,N_361,N_557);
and U1324 (N_1324,N_971,N_274);
and U1325 (N_1325,N_761,N_741);
xnor U1326 (N_1326,N_637,N_254);
nor U1327 (N_1327,N_667,N_390);
nor U1328 (N_1328,N_11,N_627);
nor U1329 (N_1329,N_748,N_646);
or U1330 (N_1330,N_607,N_177);
nand U1331 (N_1331,N_845,N_140);
nor U1332 (N_1332,N_400,N_41);
or U1333 (N_1333,N_603,N_989);
and U1334 (N_1334,N_53,N_17);
nor U1335 (N_1335,N_513,N_154);
nor U1336 (N_1336,N_624,N_860);
nor U1337 (N_1337,N_726,N_133);
and U1338 (N_1338,N_590,N_82);
or U1339 (N_1339,N_541,N_809);
or U1340 (N_1340,N_29,N_107);
or U1341 (N_1341,N_738,N_919);
or U1342 (N_1342,N_63,N_441);
nand U1343 (N_1343,N_570,N_621);
nor U1344 (N_1344,N_450,N_64);
nor U1345 (N_1345,N_56,N_723);
nor U1346 (N_1346,N_530,N_255);
nand U1347 (N_1347,N_781,N_553);
and U1348 (N_1348,N_816,N_383);
and U1349 (N_1349,N_422,N_655);
or U1350 (N_1350,N_27,N_629);
nor U1351 (N_1351,N_58,N_229);
or U1352 (N_1352,N_342,N_7);
nand U1353 (N_1353,N_664,N_812);
nand U1354 (N_1354,N_706,N_997);
nor U1355 (N_1355,N_36,N_26);
nand U1356 (N_1356,N_589,N_840);
and U1357 (N_1357,N_783,N_15);
and U1358 (N_1358,N_117,N_448);
or U1359 (N_1359,N_423,N_161);
nor U1360 (N_1360,N_690,N_493);
nor U1361 (N_1361,N_674,N_844);
or U1362 (N_1362,N_856,N_158);
and U1363 (N_1363,N_40,N_512);
xor U1364 (N_1364,N_893,N_652);
nand U1365 (N_1365,N_89,N_194);
nor U1366 (N_1366,N_830,N_734);
nand U1367 (N_1367,N_927,N_821);
nand U1368 (N_1368,N_737,N_434);
nand U1369 (N_1369,N_959,N_333);
or U1370 (N_1370,N_794,N_156);
and U1371 (N_1371,N_220,N_945);
nand U1372 (N_1372,N_314,N_656);
nand U1373 (N_1373,N_399,N_994);
xor U1374 (N_1374,N_170,N_805);
xnor U1375 (N_1375,N_866,N_431);
nor U1376 (N_1376,N_894,N_645);
nor U1377 (N_1377,N_648,N_998);
xnor U1378 (N_1378,N_560,N_90);
nand U1379 (N_1379,N_160,N_925);
and U1380 (N_1380,N_269,N_897);
and U1381 (N_1381,N_305,N_420);
nand U1382 (N_1382,N_815,N_924);
or U1383 (N_1383,N_354,N_793);
nor U1384 (N_1384,N_203,N_847);
or U1385 (N_1385,N_973,N_46);
nor U1386 (N_1386,N_159,N_380);
or U1387 (N_1387,N_322,N_88);
nand U1388 (N_1388,N_163,N_18);
nand U1389 (N_1389,N_95,N_476);
nor U1390 (N_1390,N_39,N_717);
and U1391 (N_1391,N_889,N_895);
nor U1392 (N_1392,N_339,N_733);
nand U1393 (N_1393,N_835,N_73);
or U1394 (N_1394,N_829,N_838);
nand U1395 (N_1395,N_580,N_608);
nor U1396 (N_1396,N_750,N_387);
nand U1397 (N_1397,N_475,N_13);
or U1398 (N_1398,N_944,N_504);
nor U1399 (N_1399,N_303,N_606);
and U1400 (N_1400,N_516,N_978);
xnor U1401 (N_1401,N_947,N_662);
or U1402 (N_1402,N_308,N_363);
nand U1403 (N_1403,N_433,N_797);
nand U1404 (N_1404,N_702,N_582);
or U1405 (N_1405,N_345,N_123);
nand U1406 (N_1406,N_526,N_356);
or U1407 (N_1407,N_913,N_983);
and U1408 (N_1408,N_634,N_888);
nor U1409 (N_1409,N_931,N_885);
or U1410 (N_1410,N_172,N_583);
and U1411 (N_1411,N_443,N_435);
nor U1412 (N_1412,N_188,N_597);
xor U1413 (N_1413,N_338,N_653);
or U1414 (N_1414,N_245,N_129);
nor U1415 (N_1415,N_780,N_409);
nor U1416 (N_1416,N_559,N_558);
nand U1417 (N_1417,N_939,N_695);
nor U1418 (N_1418,N_430,N_444);
nand U1419 (N_1419,N_958,N_259);
nor U1420 (N_1420,N_317,N_588);
and U1421 (N_1421,N_167,N_548);
nand U1422 (N_1422,N_950,N_879);
nand U1423 (N_1423,N_679,N_577);
and U1424 (N_1424,N_176,N_534);
nand U1425 (N_1425,N_2,N_418);
nand U1426 (N_1426,N_178,N_596);
nand U1427 (N_1427,N_234,N_786);
nor U1428 (N_1428,N_572,N_8);
and U1429 (N_1429,N_442,N_872);
and U1430 (N_1430,N_831,N_320);
nor U1431 (N_1431,N_850,N_909);
or U1432 (N_1432,N_756,N_101);
or U1433 (N_1433,N_91,N_208);
nor U1434 (N_1434,N_206,N_337);
nand U1435 (N_1435,N_869,N_340);
and U1436 (N_1436,N_832,N_411);
nand U1437 (N_1437,N_990,N_514);
and U1438 (N_1438,N_421,N_87);
nor U1439 (N_1439,N_466,N_144);
and U1440 (N_1440,N_57,N_616);
nor U1441 (N_1441,N_935,N_250);
nand U1442 (N_1442,N_227,N_697);
and U1443 (N_1443,N_402,N_811);
nand U1444 (N_1444,N_985,N_995);
nor U1445 (N_1445,N_790,N_181);
nor U1446 (N_1446,N_979,N_854);
or U1447 (N_1447,N_853,N_799);
or U1448 (N_1448,N_521,N_169);
nand U1449 (N_1449,N_536,N_132);
or U1450 (N_1450,N_347,N_519);
or U1451 (N_1451,N_23,N_787);
nor U1452 (N_1452,N_237,N_105);
or U1453 (N_1453,N_654,N_929);
or U1454 (N_1454,N_745,N_182);
nor U1455 (N_1455,N_150,N_960);
and U1456 (N_1456,N_30,N_147);
or U1457 (N_1457,N_258,N_350);
or U1458 (N_1458,N_684,N_722);
or U1459 (N_1459,N_482,N_49);
and U1460 (N_1460,N_301,N_480);
nor U1461 (N_1461,N_366,N_920);
nand U1462 (N_1462,N_618,N_127);
nor U1463 (N_1463,N_447,N_996);
nor U1464 (N_1464,N_972,N_720);
and U1465 (N_1465,N_825,N_798);
nor U1466 (N_1466,N_498,N_523);
nand U1467 (N_1467,N_124,N_456);
or U1468 (N_1468,N_716,N_187);
nand U1469 (N_1469,N_531,N_335);
nor U1470 (N_1470,N_425,N_928);
nor U1471 (N_1471,N_364,N_225);
nand U1472 (N_1472,N_348,N_675);
nor U1473 (N_1473,N_471,N_371);
nand U1474 (N_1474,N_119,N_753);
and U1475 (N_1475,N_877,N_233);
or U1476 (N_1476,N_262,N_543);
nand U1477 (N_1477,N_824,N_121);
or U1478 (N_1478,N_458,N_871);
nor U1479 (N_1479,N_75,N_533);
nand U1480 (N_1480,N_585,N_762);
and U1481 (N_1481,N_907,N_70);
nand U1482 (N_1482,N_55,N_515);
nand U1483 (N_1483,N_200,N_469);
nor U1484 (N_1484,N_520,N_586);
or U1485 (N_1485,N_567,N_48);
and U1486 (N_1486,N_111,N_113);
or U1487 (N_1487,N_479,N_264);
nor U1488 (N_1488,N_446,N_116);
nor U1489 (N_1489,N_463,N_709);
nand U1490 (N_1490,N_248,N_1);
nor U1491 (N_1491,N_594,N_639);
and U1492 (N_1492,N_358,N_731);
nor U1493 (N_1493,N_344,N_768);
nand U1494 (N_1494,N_951,N_599);
and U1495 (N_1495,N_665,N_670);
and U1496 (N_1496,N_961,N_368);
nor U1497 (N_1497,N_641,N_881);
and U1498 (N_1498,N_309,N_115);
nor U1499 (N_1499,N_67,N_852);
xnor U1500 (N_1500,N_854,N_500);
or U1501 (N_1501,N_282,N_183);
or U1502 (N_1502,N_396,N_54);
nor U1503 (N_1503,N_178,N_938);
nand U1504 (N_1504,N_714,N_713);
nor U1505 (N_1505,N_63,N_684);
or U1506 (N_1506,N_307,N_350);
or U1507 (N_1507,N_382,N_252);
or U1508 (N_1508,N_83,N_678);
nor U1509 (N_1509,N_772,N_839);
nor U1510 (N_1510,N_329,N_573);
and U1511 (N_1511,N_538,N_743);
and U1512 (N_1512,N_195,N_231);
xnor U1513 (N_1513,N_923,N_717);
nand U1514 (N_1514,N_535,N_687);
nand U1515 (N_1515,N_854,N_460);
nor U1516 (N_1516,N_264,N_593);
nand U1517 (N_1517,N_889,N_876);
nand U1518 (N_1518,N_828,N_301);
or U1519 (N_1519,N_922,N_448);
or U1520 (N_1520,N_750,N_557);
and U1521 (N_1521,N_673,N_767);
or U1522 (N_1522,N_887,N_993);
or U1523 (N_1523,N_971,N_676);
and U1524 (N_1524,N_345,N_725);
xnor U1525 (N_1525,N_242,N_109);
nor U1526 (N_1526,N_215,N_209);
nand U1527 (N_1527,N_378,N_703);
xor U1528 (N_1528,N_549,N_588);
and U1529 (N_1529,N_936,N_797);
and U1530 (N_1530,N_733,N_192);
nor U1531 (N_1531,N_694,N_821);
nor U1532 (N_1532,N_862,N_607);
or U1533 (N_1533,N_189,N_243);
nor U1534 (N_1534,N_566,N_280);
nor U1535 (N_1535,N_429,N_576);
and U1536 (N_1536,N_429,N_904);
or U1537 (N_1537,N_441,N_329);
or U1538 (N_1538,N_273,N_625);
nor U1539 (N_1539,N_163,N_169);
nand U1540 (N_1540,N_673,N_698);
nor U1541 (N_1541,N_146,N_843);
nand U1542 (N_1542,N_905,N_264);
nand U1543 (N_1543,N_264,N_774);
or U1544 (N_1544,N_430,N_840);
or U1545 (N_1545,N_593,N_436);
nand U1546 (N_1546,N_567,N_109);
or U1547 (N_1547,N_621,N_67);
and U1548 (N_1548,N_602,N_498);
nand U1549 (N_1549,N_624,N_48);
or U1550 (N_1550,N_916,N_293);
xor U1551 (N_1551,N_670,N_532);
nor U1552 (N_1552,N_241,N_204);
and U1553 (N_1553,N_473,N_244);
or U1554 (N_1554,N_840,N_948);
and U1555 (N_1555,N_231,N_182);
and U1556 (N_1556,N_988,N_468);
nand U1557 (N_1557,N_636,N_155);
or U1558 (N_1558,N_523,N_209);
and U1559 (N_1559,N_73,N_950);
and U1560 (N_1560,N_691,N_84);
or U1561 (N_1561,N_171,N_293);
nand U1562 (N_1562,N_900,N_303);
or U1563 (N_1563,N_499,N_404);
and U1564 (N_1564,N_978,N_706);
or U1565 (N_1565,N_640,N_456);
xor U1566 (N_1566,N_363,N_254);
nand U1567 (N_1567,N_778,N_177);
or U1568 (N_1568,N_815,N_25);
nand U1569 (N_1569,N_195,N_793);
nand U1570 (N_1570,N_912,N_491);
nand U1571 (N_1571,N_795,N_646);
xor U1572 (N_1572,N_236,N_483);
and U1573 (N_1573,N_110,N_456);
or U1574 (N_1574,N_870,N_873);
or U1575 (N_1575,N_83,N_880);
xnor U1576 (N_1576,N_381,N_504);
nor U1577 (N_1577,N_18,N_845);
and U1578 (N_1578,N_385,N_317);
nor U1579 (N_1579,N_895,N_658);
or U1580 (N_1580,N_891,N_180);
nand U1581 (N_1581,N_779,N_235);
or U1582 (N_1582,N_935,N_86);
xor U1583 (N_1583,N_354,N_641);
nand U1584 (N_1584,N_184,N_126);
and U1585 (N_1585,N_539,N_948);
nand U1586 (N_1586,N_282,N_797);
nor U1587 (N_1587,N_753,N_756);
nor U1588 (N_1588,N_56,N_449);
or U1589 (N_1589,N_114,N_32);
or U1590 (N_1590,N_602,N_990);
nand U1591 (N_1591,N_691,N_468);
nor U1592 (N_1592,N_956,N_244);
or U1593 (N_1593,N_600,N_146);
or U1594 (N_1594,N_769,N_751);
nand U1595 (N_1595,N_893,N_48);
or U1596 (N_1596,N_613,N_256);
nand U1597 (N_1597,N_369,N_621);
or U1598 (N_1598,N_541,N_611);
nand U1599 (N_1599,N_471,N_811);
and U1600 (N_1600,N_999,N_216);
and U1601 (N_1601,N_566,N_40);
or U1602 (N_1602,N_335,N_140);
nor U1603 (N_1603,N_974,N_134);
or U1604 (N_1604,N_447,N_985);
or U1605 (N_1605,N_275,N_279);
nand U1606 (N_1606,N_733,N_248);
or U1607 (N_1607,N_771,N_103);
and U1608 (N_1608,N_554,N_92);
or U1609 (N_1609,N_895,N_473);
nor U1610 (N_1610,N_297,N_839);
nand U1611 (N_1611,N_380,N_609);
nand U1612 (N_1612,N_370,N_970);
or U1613 (N_1613,N_579,N_984);
or U1614 (N_1614,N_205,N_207);
nor U1615 (N_1615,N_836,N_123);
nand U1616 (N_1616,N_734,N_947);
or U1617 (N_1617,N_577,N_515);
nand U1618 (N_1618,N_126,N_453);
nand U1619 (N_1619,N_648,N_312);
nor U1620 (N_1620,N_154,N_746);
nand U1621 (N_1621,N_138,N_204);
nor U1622 (N_1622,N_528,N_794);
nor U1623 (N_1623,N_568,N_769);
or U1624 (N_1624,N_599,N_944);
nand U1625 (N_1625,N_472,N_979);
or U1626 (N_1626,N_995,N_446);
and U1627 (N_1627,N_834,N_551);
or U1628 (N_1628,N_177,N_793);
and U1629 (N_1629,N_35,N_61);
xor U1630 (N_1630,N_326,N_707);
nand U1631 (N_1631,N_931,N_760);
nand U1632 (N_1632,N_279,N_284);
and U1633 (N_1633,N_86,N_781);
nand U1634 (N_1634,N_537,N_511);
or U1635 (N_1635,N_275,N_843);
or U1636 (N_1636,N_94,N_716);
and U1637 (N_1637,N_493,N_751);
nor U1638 (N_1638,N_943,N_583);
or U1639 (N_1639,N_997,N_842);
or U1640 (N_1640,N_945,N_927);
and U1641 (N_1641,N_258,N_201);
or U1642 (N_1642,N_939,N_489);
nor U1643 (N_1643,N_976,N_354);
nor U1644 (N_1644,N_289,N_697);
or U1645 (N_1645,N_304,N_653);
or U1646 (N_1646,N_426,N_353);
and U1647 (N_1647,N_832,N_205);
nor U1648 (N_1648,N_863,N_12);
or U1649 (N_1649,N_681,N_96);
nor U1650 (N_1650,N_225,N_932);
and U1651 (N_1651,N_568,N_398);
nor U1652 (N_1652,N_286,N_273);
nor U1653 (N_1653,N_326,N_287);
and U1654 (N_1654,N_718,N_397);
and U1655 (N_1655,N_97,N_27);
and U1656 (N_1656,N_256,N_67);
nand U1657 (N_1657,N_192,N_20);
or U1658 (N_1658,N_822,N_820);
nand U1659 (N_1659,N_96,N_985);
nand U1660 (N_1660,N_383,N_129);
nand U1661 (N_1661,N_164,N_9);
nor U1662 (N_1662,N_630,N_158);
and U1663 (N_1663,N_614,N_297);
or U1664 (N_1664,N_775,N_573);
nor U1665 (N_1665,N_21,N_813);
or U1666 (N_1666,N_720,N_279);
or U1667 (N_1667,N_70,N_840);
nor U1668 (N_1668,N_72,N_344);
nand U1669 (N_1669,N_962,N_662);
or U1670 (N_1670,N_987,N_305);
and U1671 (N_1671,N_480,N_966);
nand U1672 (N_1672,N_45,N_747);
nor U1673 (N_1673,N_752,N_339);
nand U1674 (N_1674,N_361,N_785);
and U1675 (N_1675,N_705,N_981);
or U1676 (N_1676,N_700,N_729);
or U1677 (N_1677,N_898,N_2);
nor U1678 (N_1678,N_879,N_797);
nand U1679 (N_1679,N_732,N_37);
and U1680 (N_1680,N_11,N_385);
nand U1681 (N_1681,N_992,N_454);
or U1682 (N_1682,N_953,N_225);
nor U1683 (N_1683,N_383,N_741);
nor U1684 (N_1684,N_368,N_355);
or U1685 (N_1685,N_356,N_82);
nor U1686 (N_1686,N_120,N_85);
nand U1687 (N_1687,N_172,N_395);
and U1688 (N_1688,N_170,N_479);
nand U1689 (N_1689,N_718,N_980);
or U1690 (N_1690,N_72,N_532);
nand U1691 (N_1691,N_156,N_622);
nand U1692 (N_1692,N_396,N_544);
and U1693 (N_1693,N_359,N_972);
and U1694 (N_1694,N_625,N_726);
nor U1695 (N_1695,N_7,N_321);
nand U1696 (N_1696,N_436,N_492);
or U1697 (N_1697,N_320,N_596);
xor U1698 (N_1698,N_525,N_670);
nand U1699 (N_1699,N_305,N_873);
nand U1700 (N_1700,N_47,N_704);
or U1701 (N_1701,N_552,N_162);
and U1702 (N_1702,N_421,N_635);
or U1703 (N_1703,N_596,N_406);
or U1704 (N_1704,N_955,N_41);
nor U1705 (N_1705,N_804,N_658);
nand U1706 (N_1706,N_831,N_642);
nor U1707 (N_1707,N_331,N_186);
nor U1708 (N_1708,N_566,N_956);
or U1709 (N_1709,N_444,N_771);
or U1710 (N_1710,N_420,N_42);
nand U1711 (N_1711,N_488,N_27);
nand U1712 (N_1712,N_963,N_604);
nor U1713 (N_1713,N_218,N_466);
or U1714 (N_1714,N_326,N_354);
or U1715 (N_1715,N_905,N_723);
and U1716 (N_1716,N_227,N_672);
nor U1717 (N_1717,N_142,N_393);
nor U1718 (N_1718,N_841,N_296);
and U1719 (N_1719,N_756,N_368);
nand U1720 (N_1720,N_904,N_432);
or U1721 (N_1721,N_919,N_720);
or U1722 (N_1722,N_270,N_52);
nor U1723 (N_1723,N_798,N_871);
and U1724 (N_1724,N_856,N_76);
nand U1725 (N_1725,N_262,N_141);
nor U1726 (N_1726,N_322,N_748);
and U1727 (N_1727,N_358,N_259);
and U1728 (N_1728,N_176,N_564);
and U1729 (N_1729,N_114,N_243);
nor U1730 (N_1730,N_837,N_550);
or U1731 (N_1731,N_66,N_799);
nor U1732 (N_1732,N_591,N_355);
or U1733 (N_1733,N_941,N_740);
or U1734 (N_1734,N_848,N_746);
or U1735 (N_1735,N_930,N_787);
or U1736 (N_1736,N_376,N_578);
nand U1737 (N_1737,N_980,N_500);
and U1738 (N_1738,N_796,N_71);
nand U1739 (N_1739,N_970,N_183);
nand U1740 (N_1740,N_82,N_218);
and U1741 (N_1741,N_882,N_806);
nand U1742 (N_1742,N_812,N_954);
and U1743 (N_1743,N_556,N_840);
xor U1744 (N_1744,N_79,N_935);
nor U1745 (N_1745,N_382,N_196);
or U1746 (N_1746,N_122,N_49);
and U1747 (N_1747,N_399,N_843);
nand U1748 (N_1748,N_891,N_259);
nor U1749 (N_1749,N_622,N_379);
nand U1750 (N_1750,N_525,N_285);
nand U1751 (N_1751,N_113,N_896);
or U1752 (N_1752,N_134,N_897);
nor U1753 (N_1753,N_555,N_293);
or U1754 (N_1754,N_393,N_397);
and U1755 (N_1755,N_53,N_208);
or U1756 (N_1756,N_790,N_888);
xor U1757 (N_1757,N_243,N_688);
nand U1758 (N_1758,N_968,N_207);
nand U1759 (N_1759,N_573,N_519);
and U1760 (N_1760,N_26,N_205);
and U1761 (N_1761,N_596,N_704);
nor U1762 (N_1762,N_852,N_358);
and U1763 (N_1763,N_974,N_6);
or U1764 (N_1764,N_792,N_203);
or U1765 (N_1765,N_276,N_305);
or U1766 (N_1766,N_404,N_51);
nand U1767 (N_1767,N_894,N_331);
and U1768 (N_1768,N_513,N_115);
or U1769 (N_1769,N_300,N_51);
or U1770 (N_1770,N_448,N_41);
or U1771 (N_1771,N_997,N_187);
and U1772 (N_1772,N_821,N_272);
or U1773 (N_1773,N_478,N_560);
nand U1774 (N_1774,N_816,N_86);
and U1775 (N_1775,N_249,N_394);
nor U1776 (N_1776,N_176,N_551);
nor U1777 (N_1777,N_266,N_637);
nor U1778 (N_1778,N_382,N_970);
and U1779 (N_1779,N_485,N_885);
nand U1780 (N_1780,N_997,N_563);
or U1781 (N_1781,N_743,N_86);
or U1782 (N_1782,N_129,N_242);
and U1783 (N_1783,N_866,N_643);
xor U1784 (N_1784,N_628,N_79);
and U1785 (N_1785,N_929,N_446);
nand U1786 (N_1786,N_833,N_531);
or U1787 (N_1787,N_103,N_313);
xor U1788 (N_1788,N_487,N_235);
nor U1789 (N_1789,N_297,N_284);
and U1790 (N_1790,N_419,N_375);
or U1791 (N_1791,N_566,N_596);
nand U1792 (N_1792,N_917,N_136);
or U1793 (N_1793,N_885,N_809);
or U1794 (N_1794,N_279,N_21);
or U1795 (N_1795,N_33,N_735);
or U1796 (N_1796,N_913,N_690);
nand U1797 (N_1797,N_88,N_761);
or U1798 (N_1798,N_910,N_269);
or U1799 (N_1799,N_383,N_99);
nor U1800 (N_1800,N_504,N_168);
and U1801 (N_1801,N_495,N_444);
nand U1802 (N_1802,N_231,N_341);
nor U1803 (N_1803,N_961,N_166);
or U1804 (N_1804,N_143,N_782);
and U1805 (N_1805,N_347,N_294);
or U1806 (N_1806,N_558,N_416);
or U1807 (N_1807,N_208,N_404);
and U1808 (N_1808,N_512,N_136);
or U1809 (N_1809,N_409,N_990);
nor U1810 (N_1810,N_219,N_606);
nand U1811 (N_1811,N_430,N_317);
and U1812 (N_1812,N_268,N_313);
or U1813 (N_1813,N_880,N_916);
and U1814 (N_1814,N_932,N_854);
nand U1815 (N_1815,N_666,N_787);
and U1816 (N_1816,N_816,N_144);
nor U1817 (N_1817,N_31,N_653);
and U1818 (N_1818,N_487,N_704);
nor U1819 (N_1819,N_299,N_250);
and U1820 (N_1820,N_477,N_245);
nor U1821 (N_1821,N_673,N_155);
nand U1822 (N_1822,N_17,N_676);
nand U1823 (N_1823,N_797,N_779);
nor U1824 (N_1824,N_159,N_634);
nand U1825 (N_1825,N_374,N_772);
and U1826 (N_1826,N_534,N_927);
or U1827 (N_1827,N_823,N_767);
and U1828 (N_1828,N_389,N_892);
nand U1829 (N_1829,N_96,N_374);
nor U1830 (N_1830,N_420,N_629);
nor U1831 (N_1831,N_960,N_569);
nand U1832 (N_1832,N_431,N_873);
or U1833 (N_1833,N_142,N_539);
or U1834 (N_1834,N_99,N_57);
nor U1835 (N_1835,N_409,N_829);
or U1836 (N_1836,N_753,N_439);
nand U1837 (N_1837,N_372,N_178);
nor U1838 (N_1838,N_195,N_598);
nor U1839 (N_1839,N_165,N_307);
and U1840 (N_1840,N_524,N_0);
and U1841 (N_1841,N_710,N_957);
xor U1842 (N_1842,N_639,N_568);
nor U1843 (N_1843,N_497,N_639);
or U1844 (N_1844,N_905,N_577);
xnor U1845 (N_1845,N_632,N_705);
nor U1846 (N_1846,N_394,N_481);
or U1847 (N_1847,N_121,N_569);
nand U1848 (N_1848,N_757,N_784);
and U1849 (N_1849,N_531,N_706);
nor U1850 (N_1850,N_390,N_613);
nand U1851 (N_1851,N_762,N_90);
or U1852 (N_1852,N_476,N_803);
nand U1853 (N_1853,N_462,N_658);
nand U1854 (N_1854,N_525,N_217);
and U1855 (N_1855,N_777,N_724);
nor U1856 (N_1856,N_249,N_790);
and U1857 (N_1857,N_270,N_47);
or U1858 (N_1858,N_658,N_42);
nand U1859 (N_1859,N_968,N_677);
or U1860 (N_1860,N_251,N_238);
and U1861 (N_1861,N_814,N_886);
or U1862 (N_1862,N_175,N_711);
nor U1863 (N_1863,N_54,N_475);
and U1864 (N_1864,N_92,N_416);
nor U1865 (N_1865,N_497,N_358);
and U1866 (N_1866,N_488,N_507);
and U1867 (N_1867,N_632,N_891);
and U1868 (N_1868,N_149,N_140);
nand U1869 (N_1869,N_316,N_882);
nand U1870 (N_1870,N_93,N_931);
and U1871 (N_1871,N_319,N_308);
and U1872 (N_1872,N_508,N_278);
or U1873 (N_1873,N_482,N_6);
nand U1874 (N_1874,N_553,N_807);
or U1875 (N_1875,N_958,N_839);
or U1876 (N_1876,N_236,N_719);
nand U1877 (N_1877,N_922,N_323);
nand U1878 (N_1878,N_203,N_715);
nand U1879 (N_1879,N_824,N_152);
or U1880 (N_1880,N_872,N_709);
nand U1881 (N_1881,N_908,N_558);
or U1882 (N_1882,N_392,N_919);
nand U1883 (N_1883,N_958,N_482);
and U1884 (N_1884,N_272,N_535);
nor U1885 (N_1885,N_911,N_328);
and U1886 (N_1886,N_928,N_184);
nor U1887 (N_1887,N_247,N_533);
nor U1888 (N_1888,N_535,N_921);
nor U1889 (N_1889,N_3,N_176);
nor U1890 (N_1890,N_601,N_569);
nor U1891 (N_1891,N_290,N_872);
or U1892 (N_1892,N_90,N_577);
or U1893 (N_1893,N_339,N_607);
nor U1894 (N_1894,N_601,N_653);
and U1895 (N_1895,N_380,N_777);
nor U1896 (N_1896,N_540,N_406);
nand U1897 (N_1897,N_64,N_589);
nor U1898 (N_1898,N_617,N_570);
nand U1899 (N_1899,N_87,N_513);
and U1900 (N_1900,N_238,N_174);
and U1901 (N_1901,N_651,N_436);
nor U1902 (N_1902,N_404,N_617);
nor U1903 (N_1903,N_343,N_720);
and U1904 (N_1904,N_951,N_326);
xor U1905 (N_1905,N_960,N_411);
or U1906 (N_1906,N_244,N_953);
and U1907 (N_1907,N_269,N_536);
nor U1908 (N_1908,N_923,N_225);
and U1909 (N_1909,N_507,N_805);
nand U1910 (N_1910,N_820,N_871);
or U1911 (N_1911,N_961,N_699);
and U1912 (N_1912,N_406,N_107);
or U1913 (N_1913,N_344,N_136);
nor U1914 (N_1914,N_822,N_4);
nor U1915 (N_1915,N_466,N_370);
or U1916 (N_1916,N_744,N_322);
or U1917 (N_1917,N_248,N_428);
or U1918 (N_1918,N_133,N_486);
nand U1919 (N_1919,N_780,N_643);
nand U1920 (N_1920,N_271,N_213);
and U1921 (N_1921,N_855,N_335);
nor U1922 (N_1922,N_369,N_855);
or U1923 (N_1923,N_918,N_737);
or U1924 (N_1924,N_210,N_773);
and U1925 (N_1925,N_808,N_272);
and U1926 (N_1926,N_189,N_49);
and U1927 (N_1927,N_362,N_740);
and U1928 (N_1928,N_287,N_324);
nor U1929 (N_1929,N_773,N_477);
nand U1930 (N_1930,N_375,N_908);
or U1931 (N_1931,N_954,N_536);
or U1932 (N_1932,N_378,N_328);
nor U1933 (N_1933,N_171,N_911);
nand U1934 (N_1934,N_622,N_247);
or U1935 (N_1935,N_903,N_112);
nor U1936 (N_1936,N_5,N_808);
or U1937 (N_1937,N_506,N_935);
nor U1938 (N_1938,N_854,N_83);
or U1939 (N_1939,N_793,N_260);
and U1940 (N_1940,N_777,N_814);
nand U1941 (N_1941,N_310,N_938);
nand U1942 (N_1942,N_644,N_537);
nor U1943 (N_1943,N_325,N_145);
or U1944 (N_1944,N_424,N_511);
nor U1945 (N_1945,N_734,N_138);
or U1946 (N_1946,N_123,N_406);
nand U1947 (N_1947,N_998,N_980);
nor U1948 (N_1948,N_391,N_244);
and U1949 (N_1949,N_311,N_486);
nor U1950 (N_1950,N_37,N_553);
nand U1951 (N_1951,N_55,N_32);
nor U1952 (N_1952,N_2,N_712);
or U1953 (N_1953,N_157,N_554);
nand U1954 (N_1954,N_423,N_68);
and U1955 (N_1955,N_388,N_279);
nor U1956 (N_1956,N_980,N_557);
and U1957 (N_1957,N_169,N_54);
or U1958 (N_1958,N_322,N_752);
nand U1959 (N_1959,N_887,N_94);
and U1960 (N_1960,N_678,N_54);
and U1961 (N_1961,N_592,N_897);
nor U1962 (N_1962,N_680,N_854);
or U1963 (N_1963,N_567,N_103);
or U1964 (N_1964,N_573,N_919);
nand U1965 (N_1965,N_812,N_305);
nand U1966 (N_1966,N_488,N_914);
nor U1967 (N_1967,N_944,N_243);
nor U1968 (N_1968,N_739,N_885);
xor U1969 (N_1969,N_127,N_288);
nand U1970 (N_1970,N_402,N_493);
nand U1971 (N_1971,N_536,N_853);
and U1972 (N_1972,N_75,N_248);
nand U1973 (N_1973,N_869,N_597);
and U1974 (N_1974,N_1,N_442);
nor U1975 (N_1975,N_42,N_326);
or U1976 (N_1976,N_734,N_268);
nor U1977 (N_1977,N_38,N_684);
nor U1978 (N_1978,N_718,N_109);
or U1979 (N_1979,N_722,N_688);
nor U1980 (N_1980,N_270,N_587);
nor U1981 (N_1981,N_813,N_149);
and U1982 (N_1982,N_352,N_103);
or U1983 (N_1983,N_329,N_96);
and U1984 (N_1984,N_556,N_254);
nor U1985 (N_1985,N_78,N_803);
or U1986 (N_1986,N_531,N_20);
and U1987 (N_1987,N_645,N_558);
nand U1988 (N_1988,N_628,N_57);
nand U1989 (N_1989,N_155,N_21);
and U1990 (N_1990,N_371,N_332);
nor U1991 (N_1991,N_780,N_308);
and U1992 (N_1992,N_866,N_463);
nand U1993 (N_1993,N_586,N_268);
nand U1994 (N_1994,N_405,N_490);
or U1995 (N_1995,N_989,N_494);
nor U1996 (N_1996,N_608,N_57);
nor U1997 (N_1997,N_811,N_740);
and U1998 (N_1998,N_559,N_198);
and U1999 (N_1999,N_159,N_739);
nand U2000 (N_2000,N_1971,N_1406);
nor U2001 (N_2001,N_1142,N_1478);
or U2002 (N_2002,N_1747,N_1739);
nand U2003 (N_2003,N_1117,N_1540);
nor U2004 (N_2004,N_1087,N_1974);
xor U2005 (N_2005,N_1611,N_1486);
or U2006 (N_2006,N_1066,N_1013);
and U2007 (N_2007,N_1006,N_1377);
nor U2008 (N_2008,N_1815,N_1904);
and U2009 (N_2009,N_1397,N_1362);
nor U2010 (N_2010,N_1476,N_1244);
and U2011 (N_2011,N_1316,N_1820);
or U2012 (N_2012,N_1961,N_1190);
nand U2013 (N_2013,N_1568,N_1559);
or U2014 (N_2014,N_1738,N_1034);
nand U2015 (N_2015,N_1280,N_1854);
nand U2016 (N_2016,N_1274,N_1224);
and U2017 (N_2017,N_1879,N_1832);
nand U2018 (N_2018,N_1749,N_1062);
xnor U2019 (N_2019,N_1933,N_1044);
or U2020 (N_2020,N_1252,N_1425);
or U2021 (N_2021,N_1569,N_1707);
or U2022 (N_2022,N_1038,N_1881);
nor U2023 (N_2023,N_1673,N_1711);
nor U2024 (N_2024,N_1701,N_1657);
nand U2025 (N_2025,N_1418,N_1620);
or U2026 (N_2026,N_1619,N_1090);
or U2027 (N_2027,N_1957,N_1847);
and U2028 (N_2028,N_1850,N_1203);
and U2029 (N_2029,N_1866,N_1295);
nand U2030 (N_2030,N_1774,N_1980);
or U2031 (N_2031,N_1344,N_1465);
and U2032 (N_2032,N_1950,N_1487);
nor U2033 (N_2033,N_1134,N_1480);
nand U2034 (N_2034,N_1470,N_1155);
or U2035 (N_2035,N_1369,N_1951);
and U2036 (N_2036,N_1007,N_1681);
nor U2037 (N_2037,N_1901,N_1777);
and U2038 (N_2038,N_1366,N_1570);
and U2039 (N_2039,N_1511,N_1136);
nor U2040 (N_2040,N_1089,N_1212);
nand U2041 (N_2041,N_1760,N_1589);
nand U2042 (N_2042,N_1693,N_1718);
or U2043 (N_2043,N_1947,N_1011);
or U2044 (N_2044,N_1053,N_1768);
nor U2045 (N_2045,N_1122,N_1084);
and U2046 (N_2046,N_1473,N_1201);
or U2047 (N_2047,N_1451,N_1621);
nand U2048 (N_2048,N_1598,N_1684);
nand U2049 (N_2049,N_1723,N_1085);
or U2050 (N_2050,N_1236,N_1272);
and U2051 (N_2051,N_1293,N_1209);
nand U2052 (N_2052,N_1528,N_1125);
or U2053 (N_2053,N_1311,N_1440);
or U2054 (N_2054,N_1271,N_1938);
or U2055 (N_2055,N_1438,N_1700);
nor U2056 (N_2056,N_1497,N_1735);
or U2057 (N_2057,N_1869,N_1849);
nor U2058 (N_2058,N_1093,N_1148);
or U2059 (N_2059,N_1515,N_1431);
or U2060 (N_2060,N_1112,N_1934);
nand U2061 (N_2061,N_1948,N_1335);
xor U2062 (N_2062,N_1636,N_1900);
nand U2063 (N_2063,N_1027,N_1207);
xnor U2064 (N_2064,N_1048,N_1078);
nand U2065 (N_2065,N_1161,N_1555);
or U2066 (N_2066,N_1283,N_1098);
nand U2067 (N_2067,N_1896,N_1814);
or U2068 (N_2068,N_1870,N_1510);
and U2069 (N_2069,N_1778,N_1593);
nand U2070 (N_2070,N_1249,N_1533);
or U2071 (N_2071,N_1858,N_1223);
nor U2072 (N_2072,N_1743,N_1996);
nand U2073 (N_2073,N_1143,N_1919);
or U2074 (N_2074,N_1821,N_1855);
and U2075 (N_2075,N_1928,N_1604);
nand U2076 (N_2076,N_1075,N_1634);
and U2077 (N_2077,N_1535,N_1705);
nor U2078 (N_2078,N_1285,N_1172);
and U2079 (N_2079,N_1780,N_1068);
or U2080 (N_2080,N_1025,N_1245);
or U2081 (N_2081,N_1643,N_1024);
and U2082 (N_2082,N_1750,N_1724);
and U2083 (N_2083,N_1983,N_1288);
or U2084 (N_2084,N_1583,N_1321);
nand U2085 (N_2085,N_1842,N_1100);
xnor U2086 (N_2086,N_1276,N_1617);
nor U2087 (N_2087,N_1408,N_1697);
xnor U2088 (N_2088,N_1003,N_1446);
and U2089 (N_2089,N_1502,N_1302);
nor U2090 (N_2090,N_1672,N_1175);
xnor U2091 (N_2091,N_1364,N_1887);
or U2092 (N_2092,N_1002,N_1234);
nand U2093 (N_2093,N_1453,N_1520);
or U2094 (N_2094,N_1065,N_1460);
and U2095 (N_2095,N_1686,N_1071);
or U2096 (N_2096,N_1477,N_1770);
and U2097 (N_2097,N_1412,N_1386);
nand U2098 (N_2098,N_1613,N_1167);
and U2099 (N_2099,N_1184,N_1860);
nor U2100 (N_2100,N_1633,N_1096);
nand U2101 (N_2101,N_1602,N_1199);
nand U2102 (N_2102,N_1665,N_1399);
or U2103 (N_2103,N_1905,N_1334);
nand U2104 (N_2104,N_1826,N_1157);
and U2105 (N_2105,N_1978,N_1278);
nand U2106 (N_2106,N_1748,N_1069);
or U2107 (N_2107,N_1456,N_1940);
nand U2108 (N_2108,N_1014,N_1585);
nor U2109 (N_2109,N_1231,N_1466);
or U2110 (N_2110,N_1287,N_1196);
or U2111 (N_2111,N_1927,N_1758);
and U2112 (N_2112,N_1638,N_1691);
nor U2113 (N_2113,N_1198,N_1115);
xor U2114 (N_2114,N_1719,N_1496);
or U2115 (N_2115,N_1594,N_1518);
nor U2116 (N_2116,N_1217,N_1326);
or U2117 (N_2117,N_1865,N_1356);
nor U2118 (N_2118,N_1906,N_1126);
and U2119 (N_2119,N_1902,N_1314);
nor U2120 (N_2120,N_1298,N_1578);
nor U2121 (N_2121,N_1367,N_1177);
or U2122 (N_2122,N_1785,N_1388);
nor U2123 (N_2123,N_1648,N_1267);
or U2124 (N_2124,N_1985,N_1703);
or U2125 (N_2125,N_1233,N_1921);
nor U2126 (N_2126,N_1498,N_1822);
and U2127 (N_2127,N_1668,N_1892);
nand U2128 (N_2128,N_1443,N_1095);
and U2129 (N_2129,N_1725,N_1588);
nor U2130 (N_2130,N_1475,N_1361);
nand U2131 (N_2131,N_1054,N_1519);
and U2132 (N_2132,N_1082,N_1186);
xnor U2133 (N_2133,N_1253,N_1363);
nand U2134 (N_2134,N_1187,N_1998);
and U2135 (N_2135,N_1941,N_1831);
or U2136 (N_2136,N_1883,N_1825);
or U2137 (N_2137,N_1146,N_1575);
or U2138 (N_2138,N_1246,N_1999);
nand U2139 (N_2139,N_1309,N_1227);
and U2140 (N_2140,N_1433,N_1164);
and U2141 (N_2141,N_1899,N_1968);
or U2142 (N_2142,N_1816,N_1370);
nor U2143 (N_2143,N_1337,N_1058);
or U2144 (N_2144,N_1376,N_1057);
and U2145 (N_2145,N_1120,N_1714);
or U2146 (N_2146,N_1525,N_1107);
or U2147 (N_2147,N_1163,N_1827);
or U2148 (N_2148,N_1264,N_1704);
nand U2149 (N_2149,N_1912,N_1424);
xnor U2150 (N_2150,N_1571,N_1208);
nor U2151 (N_2151,N_1189,N_1949);
or U2152 (N_2152,N_1325,N_1618);
and U2153 (N_2153,N_1484,N_1333);
or U2154 (N_2154,N_1566,N_1028);
nand U2155 (N_2155,N_1629,N_1573);
nand U2156 (N_2156,N_1171,N_1759);
xnor U2157 (N_2157,N_1269,N_1894);
nor U2158 (N_2158,N_1586,N_1182);
and U2159 (N_2159,N_1324,N_1835);
or U2160 (N_2160,N_1534,N_1315);
nand U2161 (N_2161,N_1138,N_1137);
nor U2162 (N_2162,N_1371,N_1884);
nand U2163 (N_2163,N_1351,N_1554);
or U2164 (N_2164,N_1103,N_1492);
and U2165 (N_2165,N_1726,N_1527);
nand U2166 (N_2166,N_1606,N_1210);
and U2167 (N_2167,N_1384,N_1124);
nand U2168 (N_2168,N_1811,N_1834);
and U2169 (N_2169,N_1852,N_1505);
or U2170 (N_2170,N_1522,N_1917);
nor U2171 (N_2171,N_1615,N_1308);
or U2172 (N_2172,N_1359,N_1449);
xor U2173 (N_2173,N_1461,N_1872);
nand U2174 (N_2174,N_1523,N_1296);
and U2175 (N_2175,N_1577,N_1320);
or U2176 (N_2176,N_1060,N_1565);
and U2177 (N_2177,N_1517,N_1669);
and U2178 (N_2178,N_1882,N_1414);
or U2179 (N_2179,N_1997,N_1086);
and U2180 (N_2180,N_1385,N_1754);
nand U2181 (N_2181,N_1074,N_1258);
nand U2182 (N_2182,N_1174,N_1863);
or U2183 (N_2183,N_1216,N_1282);
or U2184 (N_2184,N_1592,N_1608);
nor U2185 (N_2185,N_1962,N_1848);
nand U2186 (N_2186,N_1885,N_1402);
xor U2187 (N_2187,N_1340,N_1045);
nor U2188 (N_2188,N_1230,N_1610);
and U2189 (N_2189,N_1330,N_1357);
or U2190 (N_2190,N_1247,N_1539);
nand U2191 (N_2191,N_1886,N_1802);
and U2192 (N_2192,N_1080,N_1303);
and U2193 (N_2193,N_1741,N_1411);
and U2194 (N_2194,N_1448,N_1410);
nand U2195 (N_2195,N_1427,N_1955);
or U2196 (N_2196,N_1445,N_1312);
nor U2197 (N_2197,N_1929,N_1888);
nand U2198 (N_2198,N_1944,N_1818);
and U2199 (N_2199,N_1911,N_1035);
and U2200 (N_2200,N_1685,N_1185);
nor U2201 (N_2201,N_1409,N_1856);
nor U2202 (N_2202,N_1352,N_1463);
or U2203 (N_2203,N_1339,N_1787);
and U2204 (N_2204,N_1183,N_1874);
nor U2205 (N_2205,N_1779,N_1031);
nand U2206 (N_2206,N_1790,N_1471);
nor U2207 (N_2207,N_1772,N_1304);
and U2208 (N_2208,N_1623,N_1455);
or U2209 (N_2209,N_1557,N_1683);
nand U2210 (N_2210,N_1574,N_1717);
and U2211 (N_2211,N_1422,N_1979);
or U2212 (N_2212,N_1846,N_1239);
and U2213 (N_2213,N_1784,N_1404);
nand U2214 (N_2214,N_1291,N_1671);
nor U2215 (N_2215,N_1211,N_1810);
nand U2216 (N_2216,N_1348,N_1942);
and U2217 (N_2217,N_1268,N_1110);
nor U2218 (N_2218,N_1162,N_1823);
and U2219 (N_2219,N_1582,N_1490);
and U2220 (N_2220,N_1173,N_1056);
and U2221 (N_2221,N_1482,N_1839);
nor U2222 (N_2222,N_1988,N_1680);
and U2223 (N_2223,N_1458,N_1392);
nand U2224 (N_2224,N_1088,N_1121);
nand U2225 (N_2225,N_1878,N_1931);
nand U2226 (N_2226,N_1179,N_1029);
or U2227 (N_2227,N_1459,N_1710);
and U2228 (N_2228,N_1301,N_1509);
and U2229 (N_2229,N_1218,N_1713);
nand U2230 (N_2230,N_1964,N_1219);
nor U2231 (N_2231,N_1677,N_1373);
nand U2232 (N_2232,N_1764,N_1444);
nor U2233 (N_2233,N_1052,N_1489);
or U2234 (N_2234,N_1401,N_1795);
nor U2235 (N_2235,N_1970,N_1798);
and U2236 (N_2236,N_1660,N_1903);
and U2237 (N_2237,N_1867,N_1880);
nor U2238 (N_2238,N_1689,N_1639);
nand U2239 (N_2239,N_1506,N_1228);
nor U2240 (N_2240,N_1954,N_1977);
nand U2241 (N_2241,N_1391,N_1061);
or U2242 (N_2242,N_1773,N_1494);
and U2243 (N_2243,N_1552,N_1628);
nor U2244 (N_2244,N_1720,N_1129);
or U2245 (N_2245,N_1144,N_1745);
or U2246 (N_2246,N_1695,N_1488);
nand U2247 (N_2247,N_1439,N_1039);
nor U2248 (N_2248,N_1242,N_1631);
and U2249 (N_2249,N_1192,N_1799);
nand U2250 (N_2250,N_1214,N_1472);
or U2251 (N_2251,N_1877,N_1262);
and U2252 (N_2252,N_1300,N_1389);
and U2253 (N_2253,N_1263,N_1939);
or U2254 (N_2254,N_1116,N_1500);
and U2255 (N_2255,N_1421,N_1259);
and U2256 (N_2256,N_1766,N_1139);
nor U2257 (N_2257,N_1712,N_1393);
nor U2258 (N_2258,N_1358,N_1873);
and U2259 (N_2259,N_1800,N_1170);
nand U2260 (N_2260,N_1765,N_1432);
nor U2261 (N_2261,N_1600,N_1261);
or U2262 (N_2262,N_1319,N_1674);
nand U2263 (N_2263,N_1524,N_1817);
nand U2264 (N_2264,N_1696,N_1804);
nand U2265 (N_2265,N_1730,N_1907);
and U2266 (N_2266,N_1646,N_1803);
nand U2267 (N_2267,N_1687,N_1546);
or U2268 (N_2268,N_1937,N_1666);
or U2269 (N_2269,N_1776,N_1659);
nor U2270 (N_2270,N_1156,N_1215);
or U2271 (N_2271,N_1550,N_1154);
and U2272 (N_2272,N_1197,N_1794);
or U2273 (N_2273,N_1612,N_1769);
nand U2274 (N_2274,N_1036,N_1729);
or U2275 (N_2275,N_1507,N_1828);
and U2276 (N_2276,N_1413,N_1097);
nand U2277 (N_2277,N_1213,N_1273);
nor U2278 (N_2278,N_1694,N_1699);
nand U2279 (N_2279,N_1796,N_1430);
nor U2280 (N_2280,N_1853,N_1226);
or U2281 (N_2281,N_1529,N_1468);
nand U2282 (N_2282,N_1454,N_1436);
and U2283 (N_2283,N_1441,N_1310);
nand U2284 (N_2284,N_1976,N_1596);
nand U2285 (N_2285,N_1915,N_1584);
or U2286 (N_2286,N_1635,N_1450);
or U2287 (N_2287,N_1113,N_1806);
nor U2288 (N_2288,N_1650,N_1407);
nor U2289 (N_2289,N_1992,N_1149);
or U2290 (N_2290,N_1562,N_1530);
and U2291 (N_2291,N_1081,N_1682);
and U2292 (N_2292,N_1783,N_1499);
nand U2293 (N_2293,N_1147,N_1180);
nor U2294 (N_2294,N_1380,N_1336);
or U2295 (N_2295,N_1587,N_1857);
or U2296 (N_2296,N_1923,N_1994);
and U2297 (N_2297,N_1642,N_1109);
or U2298 (N_2298,N_1567,N_1016);
nand U2299 (N_2299,N_1662,N_1512);
or U2300 (N_2300,N_1323,N_1178);
or U2301 (N_2301,N_1995,N_1558);
or U2302 (N_2302,N_1420,N_1322);
nor U2303 (N_2303,N_1419,N_1188);
nor U2304 (N_2304,N_1396,N_1265);
and U2305 (N_2305,N_1479,N_1133);
or U2306 (N_2306,N_1379,N_1819);
nor U2307 (N_2307,N_1083,N_1895);
nand U2308 (N_2308,N_1020,N_1343);
and U2309 (N_2309,N_1292,N_1653);
nor U2310 (N_2310,N_1355,N_1924);
and U2311 (N_2311,N_1289,N_1374);
nor U2312 (N_2312,N_1807,N_1805);
and U2313 (N_2313,N_1248,N_1317);
nor U2314 (N_2314,N_1833,N_1742);
and U2315 (N_2315,N_1047,N_1485);
xnor U2316 (N_2316,N_1953,N_1875);
nor U2317 (N_2317,N_1108,N_1793);
and U2318 (N_2318,N_1624,N_1676);
nand U2319 (N_2319,N_1544,N_1260);
nand U2320 (N_2320,N_1859,N_1946);
nor U2321 (N_2321,N_1381,N_1347);
nor U2322 (N_2322,N_1651,N_1023);
xnor U2323 (N_2323,N_1627,N_1200);
nand U2324 (N_2324,N_1284,N_1042);
nor U2325 (N_2325,N_1597,N_1165);
and U2326 (N_2326,N_1428,N_1092);
xor U2327 (N_2327,N_1046,N_1722);
nor U2328 (N_2328,N_1281,N_1238);
and U2329 (N_2329,N_1152,N_1844);
nand U2330 (N_2330,N_1114,N_1070);
nand U2331 (N_2331,N_1266,N_1063);
and U2332 (N_2332,N_1603,N_1897);
nor U2333 (N_2333,N_1622,N_1375);
or U2334 (N_2334,N_1563,N_1914);
nand U2335 (N_2335,N_1206,N_1508);
and U2336 (N_2336,N_1493,N_1829);
nor U2337 (N_2337,N_1299,N_1667);
and U2338 (N_2338,N_1740,N_1652);
nand U2339 (N_2339,N_1864,N_1128);
or U2340 (N_2340,N_1503,N_1532);
nand U2341 (N_2341,N_1734,N_1781);
and U2342 (N_2342,N_1395,N_1055);
and U2343 (N_2343,N_1590,N_1836);
xnor U2344 (N_2344,N_1982,N_1437);
nand U2345 (N_2345,N_1091,N_1342);
nor U2346 (N_2346,N_1972,N_1580);
xnor U2347 (N_2347,N_1936,N_1797);
nor U2348 (N_2348,N_1991,N_1545);
or U2349 (N_2349,N_1841,N_1607);
or U2350 (N_2350,N_1943,N_1744);
or U2351 (N_2351,N_1969,N_1094);
xnor U2352 (N_2352,N_1050,N_1812);
nor U2353 (N_2353,N_1229,N_1706);
nor U2354 (N_2354,N_1973,N_1032);
nand U2355 (N_2355,N_1464,N_1429);
nor U2356 (N_2356,N_1305,N_1733);
nand U2357 (N_2357,N_1041,N_1987);
or U2358 (N_2358,N_1131,N_1135);
nand U2359 (N_2359,N_1925,N_1751);
nand U2360 (N_2360,N_1033,N_1019);
and U2361 (N_2361,N_1004,N_1762);
nor U2362 (N_2362,N_1101,N_1132);
nor U2363 (N_2363,N_1141,N_1782);
nor U2364 (N_2364,N_1501,N_1076);
nand U2365 (N_2365,N_1159,N_1614);
nand U2366 (N_2366,N_1791,N_1541);
and U2367 (N_2367,N_1556,N_1191);
nor U2368 (N_2368,N_1059,N_1067);
and U2369 (N_2369,N_1015,N_1531);
nor U2370 (N_2370,N_1279,N_1251);
nand U2371 (N_2371,N_1576,N_1889);
or U2372 (N_2372,N_1365,N_1327);
or U2373 (N_2373,N_1256,N_1130);
and U2374 (N_2374,N_1043,N_1656);
nor U2375 (N_2375,N_1329,N_1119);
and U2376 (N_2376,N_1840,N_1018);
nor U2377 (N_2377,N_1469,N_1118);
nor U2378 (N_2378,N_1194,N_1767);
or U2379 (N_2379,N_1990,N_1037);
and U2380 (N_2380,N_1099,N_1548);
nor U2381 (N_2381,N_1504,N_1625);
and U2382 (N_2382,N_1481,N_1959);
nand U2383 (N_2383,N_1513,N_1434);
or U2384 (N_2384,N_1346,N_1294);
or U2385 (N_2385,N_1728,N_1581);
and U2386 (N_2386,N_1158,N_1675);
nand U2387 (N_2387,N_1813,N_1193);
xnor U2388 (N_2388,N_1383,N_1051);
nor U2389 (N_2389,N_1649,N_1290);
and U2390 (N_2390,N_1871,N_1307);
or U2391 (N_2391,N_1561,N_1543);
nor U2392 (N_2392,N_1232,N_1930);
nand U2393 (N_2393,N_1965,N_1516);
or U2394 (N_2394,N_1655,N_1372);
nand U2395 (N_2395,N_1442,N_1368);
nor U2396 (N_2396,N_1564,N_1984);
nor U2397 (N_2397,N_1542,N_1275);
and U2398 (N_2398,N_1474,N_1547);
and U2399 (N_2399,N_1123,N_1876);
and U2400 (N_2400,N_1678,N_1645);
or U2401 (N_2401,N_1553,N_1181);
nor U2402 (N_2402,N_1690,N_1752);
or U2403 (N_2403,N_1626,N_1104);
nand U2404 (N_2404,N_1009,N_1255);
nand U2405 (N_2405,N_1963,N_1663);
nor U2406 (N_2406,N_1435,N_1756);
or U2407 (N_2407,N_1789,N_1851);
and U2408 (N_2408,N_1916,N_1644);
and U2409 (N_2409,N_1106,N_1721);
nand U2410 (N_2410,N_1830,N_1243);
or U2411 (N_2411,N_1140,N_1286);
and U2412 (N_2412,N_1030,N_1416);
xnor U2413 (N_2413,N_1975,N_1022);
and U2414 (N_2414,N_1176,N_1727);
nor U2415 (N_2415,N_1918,N_1240);
and U2416 (N_2416,N_1993,N_1079);
nor U2417 (N_2417,N_1168,N_1483);
xnor U2418 (N_2418,N_1641,N_1632);
and U2419 (N_2419,N_1195,N_1153);
or U2420 (N_2420,N_1012,N_1732);
nor U2421 (N_2421,N_1241,N_1491);
and U2422 (N_2422,N_1328,N_1861);
and U2423 (N_2423,N_1981,N_1935);
nor U2424 (N_2424,N_1609,N_1235);
nor U2425 (N_2425,N_1354,N_1001);
nor U2426 (N_2426,N_1630,N_1757);
or U2427 (N_2427,N_1838,N_1560);
nand U2428 (N_2428,N_1605,N_1306);
and U2429 (N_2429,N_1160,N_1868);
nand U2430 (N_2430,N_1332,N_1415);
and U2431 (N_2431,N_1549,N_1967);
nor U2432 (N_2432,N_1225,N_1843);
or U2433 (N_2433,N_1221,N_1702);
or U2434 (N_2434,N_1792,N_1105);
or U2435 (N_2435,N_1526,N_1394);
xnor U2436 (N_2436,N_1127,N_1989);
nor U2437 (N_2437,N_1824,N_1026);
or U2438 (N_2438,N_1679,N_1688);
and U2439 (N_2439,N_1390,N_1909);
nor U2440 (N_2440,N_1761,N_1893);
and U2441 (N_2441,N_1837,N_1495);
or U2442 (N_2442,N_1205,N_1341);
and U2443 (N_2443,N_1338,N_1716);
nand U2444 (N_2444,N_1908,N_1664);
nand U2445 (N_2445,N_1786,N_1637);
nor U2446 (N_2446,N_1898,N_1077);
xnor U2447 (N_2447,N_1254,N_1462);
and U2448 (N_2448,N_1400,N_1360);
and U2449 (N_2449,N_1890,N_1423);
nand U2450 (N_2450,N_1008,N_1353);
or U2451 (N_2451,N_1920,N_1000);
or U2452 (N_2452,N_1387,N_1616);
nor U2453 (N_2453,N_1064,N_1922);
and U2454 (N_2454,N_1250,N_1452);
or U2455 (N_2455,N_1202,N_1378);
nand U2456 (N_2456,N_1599,N_1102);
nor U2457 (N_2457,N_1788,N_1318);
nor U2458 (N_2458,N_1204,N_1551);
nand U2459 (N_2459,N_1403,N_1417);
nand U2460 (N_2460,N_1715,N_1670);
and U2461 (N_2461,N_1049,N_1382);
or U2462 (N_2462,N_1297,N_1151);
nand U2463 (N_2463,N_1345,N_1538);
and U2464 (N_2464,N_1775,N_1862);
and U2465 (N_2465,N_1960,N_1845);
nor U2466 (N_2466,N_1521,N_1111);
nor U2467 (N_2467,N_1040,N_1222);
nor U2468 (N_2468,N_1591,N_1647);
nor U2469 (N_2469,N_1926,N_1072);
nor U2470 (N_2470,N_1910,N_1601);
nand U2471 (N_2471,N_1572,N_1753);
nor U2472 (N_2472,N_1945,N_1536);
nand U2473 (N_2473,N_1709,N_1447);
nand U2474 (N_2474,N_1808,N_1313);
and U2475 (N_2475,N_1277,N_1801);
and U2476 (N_2476,N_1349,N_1017);
nor U2477 (N_2477,N_1595,N_1579);
nand U2478 (N_2478,N_1654,N_1270);
and U2479 (N_2479,N_1891,N_1932);
nor U2480 (N_2480,N_1698,N_1692);
nand U2481 (N_2481,N_1746,N_1737);
and U2482 (N_2482,N_1010,N_1537);
or U2483 (N_2483,N_1257,N_1956);
nand U2484 (N_2484,N_1467,N_1426);
nor U2485 (N_2485,N_1021,N_1166);
nor U2486 (N_2486,N_1809,N_1457);
nor U2487 (N_2487,N_1913,N_1708);
or U2488 (N_2488,N_1331,N_1220);
nand U2489 (N_2489,N_1150,N_1658);
nor U2490 (N_2490,N_1350,N_1952);
nand U2491 (N_2491,N_1755,N_1661);
and U2492 (N_2492,N_1398,N_1731);
nor U2493 (N_2493,N_1966,N_1237);
and U2494 (N_2494,N_1958,N_1073);
nor U2495 (N_2495,N_1736,N_1145);
nor U2496 (N_2496,N_1005,N_1986);
and U2497 (N_2497,N_1405,N_1514);
or U2498 (N_2498,N_1169,N_1763);
or U2499 (N_2499,N_1771,N_1640);
and U2500 (N_2500,N_1826,N_1370);
or U2501 (N_2501,N_1352,N_1359);
or U2502 (N_2502,N_1546,N_1140);
nor U2503 (N_2503,N_1358,N_1566);
and U2504 (N_2504,N_1746,N_1661);
nor U2505 (N_2505,N_1816,N_1662);
nor U2506 (N_2506,N_1581,N_1696);
nand U2507 (N_2507,N_1614,N_1437);
nor U2508 (N_2508,N_1517,N_1887);
nand U2509 (N_2509,N_1599,N_1325);
or U2510 (N_2510,N_1105,N_1977);
and U2511 (N_2511,N_1762,N_1205);
nand U2512 (N_2512,N_1136,N_1329);
nor U2513 (N_2513,N_1707,N_1644);
nor U2514 (N_2514,N_1030,N_1811);
nand U2515 (N_2515,N_1842,N_1605);
and U2516 (N_2516,N_1954,N_1389);
xor U2517 (N_2517,N_1635,N_1237);
and U2518 (N_2518,N_1101,N_1278);
and U2519 (N_2519,N_1424,N_1773);
nand U2520 (N_2520,N_1067,N_1314);
nand U2521 (N_2521,N_1944,N_1613);
nand U2522 (N_2522,N_1613,N_1428);
xor U2523 (N_2523,N_1706,N_1198);
or U2524 (N_2524,N_1400,N_1066);
and U2525 (N_2525,N_1273,N_1009);
xor U2526 (N_2526,N_1591,N_1054);
nand U2527 (N_2527,N_1274,N_1472);
and U2528 (N_2528,N_1360,N_1522);
nor U2529 (N_2529,N_1465,N_1155);
or U2530 (N_2530,N_1650,N_1076);
and U2531 (N_2531,N_1490,N_1706);
or U2532 (N_2532,N_1140,N_1874);
and U2533 (N_2533,N_1169,N_1627);
nor U2534 (N_2534,N_1985,N_1646);
nand U2535 (N_2535,N_1678,N_1369);
nor U2536 (N_2536,N_1667,N_1638);
and U2537 (N_2537,N_1614,N_1376);
and U2538 (N_2538,N_1426,N_1462);
and U2539 (N_2539,N_1901,N_1887);
nand U2540 (N_2540,N_1788,N_1135);
or U2541 (N_2541,N_1640,N_1242);
or U2542 (N_2542,N_1794,N_1978);
or U2543 (N_2543,N_1585,N_1007);
nor U2544 (N_2544,N_1124,N_1903);
and U2545 (N_2545,N_1949,N_1219);
nor U2546 (N_2546,N_1230,N_1435);
nand U2547 (N_2547,N_1759,N_1011);
nor U2548 (N_2548,N_1875,N_1237);
nor U2549 (N_2549,N_1879,N_1986);
and U2550 (N_2550,N_1350,N_1150);
and U2551 (N_2551,N_1408,N_1923);
or U2552 (N_2552,N_1863,N_1859);
or U2553 (N_2553,N_1163,N_1748);
and U2554 (N_2554,N_1705,N_1541);
or U2555 (N_2555,N_1891,N_1317);
or U2556 (N_2556,N_1108,N_1635);
and U2557 (N_2557,N_1512,N_1868);
and U2558 (N_2558,N_1167,N_1570);
nand U2559 (N_2559,N_1390,N_1502);
nor U2560 (N_2560,N_1675,N_1838);
nor U2561 (N_2561,N_1254,N_1390);
or U2562 (N_2562,N_1967,N_1680);
nor U2563 (N_2563,N_1774,N_1446);
nor U2564 (N_2564,N_1733,N_1307);
or U2565 (N_2565,N_1311,N_1201);
nor U2566 (N_2566,N_1215,N_1786);
or U2567 (N_2567,N_1298,N_1696);
and U2568 (N_2568,N_1940,N_1497);
nand U2569 (N_2569,N_1051,N_1475);
nand U2570 (N_2570,N_1246,N_1577);
nor U2571 (N_2571,N_1626,N_1006);
nand U2572 (N_2572,N_1937,N_1355);
nor U2573 (N_2573,N_1964,N_1950);
nand U2574 (N_2574,N_1560,N_1401);
nand U2575 (N_2575,N_1871,N_1194);
nand U2576 (N_2576,N_1361,N_1994);
nor U2577 (N_2577,N_1458,N_1139);
and U2578 (N_2578,N_1008,N_1821);
nand U2579 (N_2579,N_1278,N_1812);
nand U2580 (N_2580,N_1037,N_1123);
nand U2581 (N_2581,N_1735,N_1107);
nand U2582 (N_2582,N_1128,N_1341);
or U2583 (N_2583,N_1631,N_1360);
nand U2584 (N_2584,N_1231,N_1056);
nor U2585 (N_2585,N_1818,N_1419);
nor U2586 (N_2586,N_1233,N_1466);
or U2587 (N_2587,N_1437,N_1483);
and U2588 (N_2588,N_1271,N_1144);
or U2589 (N_2589,N_1945,N_1558);
nor U2590 (N_2590,N_1212,N_1814);
nand U2591 (N_2591,N_1275,N_1330);
and U2592 (N_2592,N_1310,N_1948);
and U2593 (N_2593,N_1277,N_1864);
and U2594 (N_2594,N_1283,N_1723);
nor U2595 (N_2595,N_1214,N_1786);
nand U2596 (N_2596,N_1752,N_1456);
and U2597 (N_2597,N_1313,N_1174);
xor U2598 (N_2598,N_1967,N_1861);
and U2599 (N_2599,N_1138,N_1006);
nand U2600 (N_2600,N_1485,N_1658);
or U2601 (N_2601,N_1564,N_1239);
and U2602 (N_2602,N_1460,N_1998);
and U2603 (N_2603,N_1688,N_1537);
or U2604 (N_2604,N_1583,N_1974);
nor U2605 (N_2605,N_1023,N_1792);
nand U2606 (N_2606,N_1612,N_1756);
nor U2607 (N_2607,N_1020,N_1105);
and U2608 (N_2608,N_1849,N_1103);
nor U2609 (N_2609,N_1120,N_1863);
nor U2610 (N_2610,N_1891,N_1719);
or U2611 (N_2611,N_1836,N_1983);
nand U2612 (N_2612,N_1220,N_1693);
and U2613 (N_2613,N_1907,N_1627);
or U2614 (N_2614,N_1982,N_1373);
or U2615 (N_2615,N_1926,N_1769);
or U2616 (N_2616,N_1488,N_1140);
and U2617 (N_2617,N_1723,N_1989);
nor U2618 (N_2618,N_1023,N_1863);
nor U2619 (N_2619,N_1491,N_1250);
nor U2620 (N_2620,N_1630,N_1793);
nor U2621 (N_2621,N_1269,N_1157);
nand U2622 (N_2622,N_1493,N_1800);
and U2623 (N_2623,N_1603,N_1569);
and U2624 (N_2624,N_1835,N_1374);
or U2625 (N_2625,N_1643,N_1562);
and U2626 (N_2626,N_1267,N_1811);
or U2627 (N_2627,N_1147,N_1068);
nor U2628 (N_2628,N_1040,N_1502);
nor U2629 (N_2629,N_1291,N_1811);
nor U2630 (N_2630,N_1125,N_1428);
or U2631 (N_2631,N_1471,N_1268);
and U2632 (N_2632,N_1406,N_1787);
and U2633 (N_2633,N_1839,N_1678);
and U2634 (N_2634,N_1059,N_1986);
nand U2635 (N_2635,N_1747,N_1257);
or U2636 (N_2636,N_1045,N_1830);
nor U2637 (N_2637,N_1261,N_1729);
or U2638 (N_2638,N_1558,N_1835);
and U2639 (N_2639,N_1430,N_1976);
and U2640 (N_2640,N_1770,N_1735);
or U2641 (N_2641,N_1209,N_1324);
nor U2642 (N_2642,N_1040,N_1503);
nand U2643 (N_2643,N_1372,N_1231);
or U2644 (N_2644,N_1543,N_1611);
or U2645 (N_2645,N_1213,N_1036);
nor U2646 (N_2646,N_1268,N_1897);
nand U2647 (N_2647,N_1746,N_1903);
or U2648 (N_2648,N_1823,N_1599);
or U2649 (N_2649,N_1375,N_1589);
and U2650 (N_2650,N_1647,N_1731);
and U2651 (N_2651,N_1021,N_1368);
nor U2652 (N_2652,N_1302,N_1983);
nor U2653 (N_2653,N_1254,N_1710);
nor U2654 (N_2654,N_1975,N_1403);
or U2655 (N_2655,N_1158,N_1858);
nand U2656 (N_2656,N_1487,N_1692);
nand U2657 (N_2657,N_1362,N_1907);
and U2658 (N_2658,N_1199,N_1882);
or U2659 (N_2659,N_1157,N_1226);
nor U2660 (N_2660,N_1593,N_1297);
nor U2661 (N_2661,N_1096,N_1048);
nand U2662 (N_2662,N_1449,N_1324);
and U2663 (N_2663,N_1094,N_1480);
nand U2664 (N_2664,N_1037,N_1666);
or U2665 (N_2665,N_1335,N_1972);
or U2666 (N_2666,N_1300,N_1873);
or U2667 (N_2667,N_1448,N_1252);
xor U2668 (N_2668,N_1258,N_1010);
nand U2669 (N_2669,N_1943,N_1612);
nand U2670 (N_2670,N_1252,N_1064);
and U2671 (N_2671,N_1529,N_1159);
nor U2672 (N_2672,N_1827,N_1585);
and U2673 (N_2673,N_1326,N_1645);
nor U2674 (N_2674,N_1485,N_1398);
nand U2675 (N_2675,N_1388,N_1061);
and U2676 (N_2676,N_1820,N_1254);
xor U2677 (N_2677,N_1544,N_1475);
and U2678 (N_2678,N_1811,N_1225);
nor U2679 (N_2679,N_1425,N_1462);
and U2680 (N_2680,N_1412,N_1349);
and U2681 (N_2681,N_1365,N_1304);
nand U2682 (N_2682,N_1670,N_1033);
nor U2683 (N_2683,N_1717,N_1194);
nor U2684 (N_2684,N_1058,N_1363);
and U2685 (N_2685,N_1114,N_1835);
nand U2686 (N_2686,N_1771,N_1569);
or U2687 (N_2687,N_1587,N_1006);
and U2688 (N_2688,N_1851,N_1534);
and U2689 (N_2689,N_1161,N_1610);
or U2690 (N_2690,N_1605,N_1493);
nand U2691 (N_2691,N_1069,N_1405);
and U2692 (N_2692,N_1917,N_1339);
or U2693 (N_2693,N_1185,N_1605);
nand U2694 (N_2694,N_1320,N_1295);
nand U2695 (N_2695,N_1570,N_1464);
nor U2696 (N_2696,N_1162,N_1660);
nor U2697 (N_2697,N_1628,N_1310);
nand U2698 (N_2698,N_1467,N_1197);
nand U2699 (N_2699,N_1521,N_1822);
or U2700 (N_2700,N_1862,N_1522);
nor U2701 (N_2701,N_1233,N_1840);
nand U2702 (N_2702,N_1380,N_1582);
or U2703 (N_2703,N_1200,N_1826);
or U2704 (N_2704,N_1742,N_1908);
nor U2705 (N_2705,N_1010,N_1525);
or U2706 (N_2706,N_1560,N_1801);
or U2707 (N_2707,N_1180,N_1227);
nand U2708 (N_2708,N_1761,N_1520);
and U2709 (N_2709,N_1049,N_1370);
nor U2710 (N_2710,N_1253,N_1626);
nor U2711 (N_2711,N_1331,N_1793);
nor U2712 (N_2712,N_1606,N_1750);
nand U2713 (N_2713,N_1099,N_1135);
or U2714 (N_2714,N_1632,N_1760);
nand U2715 (N_2715,N_1156,N_1130);
or U2716 (N_2716,N_1661,N_1097);
nand U2717 (N_2717,N_1306,N_1876);
nor U2718 (N_2718,N_1259,N_1910);
and U2719 (N_2719,N_1739,N_1079);
nand U2720 (N_2720,N_1310,N_1786);
nand U2721 (N_2721,N_1524,N_1942);
nor U2722 (N_2722,N_1491,N_1079);
nor U2723 (N_2723,N_1873,N_1419);
nor U2724 (N_2724,N_1233,N_1362);
nor U2725 (N_2725,N_1835,N_1260);
and U2726 (N_2726,N_1584,N_1009);
or U2727 (N_2727,N_1190,N_1716);
nand U2728 (N_2728,N_1988,N_1677);
and U2729 (N_2729,N_1661,N_1232);
and U2730 (N_2730,N_1396,N_1615);
nand U2731 (N_2731,N_1528,N_1010);
and U2732 (N_2732,N_1151,N_1418);
and U2733 (N_2733,N_1215,N_1367);
nor U2734 (N_2734,N_1345,N_1631);
nor U2735 (N_2735,N_1948,N_1362);
or U2736 (N_2736,N_1429,N_1512);
and U2737 (N_2737,N_1432,N_1123);
or U2738 (N_2738,N_1820,N_1400);
xnor U2739 (N_2739,N_1832,N_1008);
or U2740 (N_2740,N_1287,N_1913);
nor U2741 (N_2741,N_1691,N_1348);
nand U2742 (N_2742,N_1709,N_1136);
or U2743 (N_2743,N_1182,N_1039);
nor U2744 (N_2744,N_1299,N_1668);
nand U2745 (N_2745,N_1565,N_1985);
nand U2746 (N_2746,N_1800,N_1053);
and U2747 (N_2747,N_1934,N_1517);
and U2748 (N_2748,N_1525,N_1285);
nor U2749 (N_2749,N_1887,N_1040);
xor U2750 (N_2750,N_1886,N_1697);
nand U2751 (N_2751,N_1244,N_1387);
or U2752 (N_2752,N_1329,N_1059);
nand U2753 (N_2753,N_1012,N_1816);
nor U2754 (N_2754,N_1714,N_1506);
nand U2755 (N_2755,N_1967,N_1432);
nand U2756 (N_2756,N_1924,N_1745);
or U2757 (N_2757,N_1495,N_1405);
and U2758 (N_2758,N_1523,N_1200);
or U2759 (N_2759,N_1422,N_1517);
nand U2760 (N_2760,N_1923,N_1261);
or U2761 (N_2761,N_1978,N_1189);
nor U2762 (N_2762,N_1977,N_1832);
nand U2763 (N_2763,N_1377,N_1218);
nand U2764 (N_2764,N_1404,N_1332);
nor U2765 (N_2765,N_1166,N_1302);
and U2766 (N_2766,N_1026,N_1401);
and U2767 (N_2767,N_1050,N_1641);
and U2768 (N_2768,N_1989,N_1791);
or U2769 (N_2769,N_1113,N_1477);
or U2770 (N_2770,N_1156,N_1615);
and U2771 (N_2771,N_1676,N_1467);
nand U2772 (N_2772,N_1516,N_1777);
or U2773 (N_2773,N_1230,N_1805);
and U2774 (N_2774,N_1768,N_1885);
nand U2775 (N_2775,N_1603,N_1570);
nand U2776 (N_2776,N_1899,N_1253);
or U2777 (N_2777,N_1299,N_1277);
or U2778 (N_2778,N_1193,N_1849);
nand U2779 (N_2779,N_1110,N_1628);
or U2780 (N_2780,N_1971,N_1313);
nand U2781 (N_2781,N_1141,N_1113);
or U2782 (N_2782,N_1395,N_1315);
or U2783 (N_2783,N_1781,N_1490);
and U2784 (N_2784,N_1015,N_1326);
or U2785 (N_2785,N_1999,N_1320);
and U2786 (N_2786,N_1937,N_1227);
nand U2787 (N_2787,N_1554,N_1757);
nand U2788 (N_2788,N_1079,N_1254);
nor U2789 (N_2789,N_1938,N_1664);
nor U2790 (N_2790,N_1270,N_1518);
and U2791 (N_2791,N_1212,N_1896);
and U2792 (N_2792,N_1197,N_1086);
and U2793 (N_2793,N_1967,N_1633);
nand U2794 (N_2794,N_1002,N_1965);
nand U2795 (N_2795,N_1109,N_1714);
and U2796 (N_2796,N_1891,N_1495);
nor U2797 (N_2797,N_1606,N_1239);
or U2798 (N_2798,N_1131,N_1239);
nor U2799 (N_2799,N_1267,N_1028);
nand U2800 (N_2800,N_1224,N_1006);
nor U2801 (N_2801,N_1011,N_1185);
nand U2802 (N_2802,N_1781,N_1119);
nand U2803 (N_2803,N_1081,N_1739);
and U2804 (N_2804,N_1922,N_1709);
and U2805 (N_2805,N_1366,N_1129);
and U2806 (N_2806,N_1201,N_1132);
nand U2807 (N_2807,N_1538,N_1572);
and U2808 (N_2808,N_1239,N_1557);
nor U2809 (N_2809,N_1064,N_1486);
nand U2810 (N_2810,N_1967,N_1560);
nor U2811 (N_2811,N_1158,N_1582);
and U2812 (N_2812,N_1949,N_1381);
or U2813 (N_2813,N_1938,N_1479);
nor U2814 (N_2814,N_1847,N_1017);
and U2815 (N_2815,N_1197,N_1712);
or U2816 (N_2816,N_1512,N_1884);
or U2817 (N_2817,N_1279,N_1611);
or U2818 (N_2818,N_1679,N_1430);
and U2819 (N_2819,N_1672,N_1595);
nand U2820 (N_2820,N_1580,N_1302);
nor U2821 (N_2821,N_1762,N_1448);
nor U2822 (N_2822,N_1526,N_1509);
nand U2823 (N_2823,N_1151,N_1940);
and U2824 (N_2824,N_1099,N_1839);
nand U2825 (N_2825,N_1958,N_1149);
nor U2826 (N_2826,N_1357,N_1133);
nor U2827 (N_2827,N_1221,N_1600);
nand U2828 (N_2828,N_1090,N_1774);
nor U2829 (N_2829,N_1193,N_1907);
nor U2830 (N_2830,N_1449,N_1742);
or U2831 (N_2831,N_1886,N_1814);
nand U2832 (N_2832,N_1899,N_1422);
nand U2833 (N_2833,N_1047,N_1660);
nand U2834 (N_2834,N_1212,N_1947);
nand U2835 (N_2835,N_1619,N_1650);
nand U2836 (N_2836,N_1525,N_1635);
or U2837 (N_2837,N_1596,N_1000);
or U2838 (N_2838,N_1533,N_1872);
nand U2839 (N_2839,N_1479,N_1179);
nand U2840 (N_2840,N_1248,N_1272);
or U2841 (N_2841,N_1413,N_1975);
and U2842 (N_2842,N_1441,N_1565);
or U2843 (N_2843,N_1519,N_1483);
and U2844 (N_2844,N_1172,N_1028);
nand U2845 (N_2845,N_1123,N_1809);
and U2846 (N_2846,N_1465,N_1675);
or U2847 (N_2847,N_1573,N_1299);
or U2848 (N_2848,N_1548,N_1758);
nor U2849 (N_2849,N_1896,N_1872);
or U2850 (N_2850,N_1882,N_1564);
nor U2851 (N_2851,N_1378,N_1770);
nor U2852 (N_2852,N_1928,N_1013);
or U2853 (N_2853,N_1066,N_1844);
or U2854 (N_2854,N_1388,N_1157);
and U2855 (N_2855,N_1567,N_1213);
nor U2856 (N_2856,N_1743,N_1942);
and U2857 (N_2857,N_1949,N_1896);
and U2858 (N_2858,N_1566,N_1092);
or U2859 (N_2859,N_1978,N_1601);
and U2860 (N_2860,N_1182,N_1790);
nor U2861 (N_2861,N_1631,N_1912);
or U2862 (N_2862,N_1250,N_1941);
nand U2863 (N_2863,N_1665,N_1551);
nor U2864 (N_2864,N_1522,N_1040);
or U2865 (N_2865,N_1222,N_1958);
and U2866 (N_2866,N_1787,N_1262);
nor U2867 (N_2867,N_1602,N_1977);
or U2868 (N_2868,N_1978,N_1453);
nand U2869 (N_2869,N_1294,N_1016);
and U2870 (N_2870,N_1505,N_1187);
or U2871 (N_2871,N_1107,N_1464);
or U2872 (N_2872,N_1664,N_1317);
nand U2873 (N_2873,N_1944,N_1585);
or U2874 (N_2874,N_1799,N_1840);
or U2875 (N_2875,N_1637,N_1639);
and U2876 (N_2876,N_1389,N_1008);
nand U2877 (N_2877,N_1874,N_1624);
nand U2878 (N_2878,N_1464,N_1811);
nand U2879 (N_2879,N_1882,N_1629);
or U2880 (N_2880,N_1133,N_1706);
nand U2881 (N_2881,N_1511,N_1057);
xor U2882 (N_2882,N_1069,N_1214);
or U2883 (N_2883,N_1019,N_1963);
xor U2884 (N_2884,N_1505,N_1763);
or U2885 (N_2885,N_1628,N_1430);
or U2886 (N_2886,N_1835,N_1575);
nor U2887 (N_2887,N_1818,N_1774);
nor U2888 (N_2888,N_1437,N_1782);
and U2889 (N_2889,N_1696,N_1020);
and U2890 (N_2890,N_1721,N_1713);
xnor U2891 (N_2891,N_1243,N_1247);
nand U2892 (N_2892,N_1422,N_1969);
nor U2893 (N_2893,N_1161,N_1253);
or U2894 (N_2894,N_1966,N_1807);
nand U2895 (N_2895,N_1170,N_1671);
and U2896 (N_2896,N_1687,N_1296);
or U2897 (N_2897,N_1288,N_1658);
and U2898 (N_2898,N_1334,N_1534);
and U2899 (N_2899,N_1768,N_1025);
and U2900 (N_2900,N_1670,N_1912);
nand U2901 (N_2901,N_1307,N_1851);
nor U2902 (N_2902,N_1081,N_1500);
or U2903 (N_2903,N_1042,N_1883);
nand U2904 (N_2904,N_1852,N_1738);
and U2905 (N_2905,N_1340,N_1223);
nor U2906 (N_2906,N_1005,N_1222);
or U2907 (N_2907,N_1467,N_1024);
and U2908 (N_2908,N_1480,N_1448);
and U2909 (N_2909,N_1741,N_1047);
and U2910 (N_2910,N_1128,N_1977);
nand U2911 (N_2911,N_1319,N_1467);
nor U2912 (N_2912,N_1994,N_1039);
or U2913 (N_2913,N_1523,N_1453);
nor U2914 (N_2914,N_1332,N_1335);
nor U2915 (N_2915,N_1712,N_1806);
or U2916 (N_2916,N_1171,N_1062);
nor U2917 (N_2917,N_1790,N_1257);
nand U2918 (N_2918,N_1687,N_1713);
or U2919 (N_2919,N_1534,N_1462);
nand U2920 (N_2920,N_1204,N_1626);
nor U2921 (N_2921,N_1063,N_1773);
nor U2922 (N_2922,N_1536,N_1466);
and U2923 (N_2923,N_1431,N_1151);
nor U2924 (N_2924,N_1375,N_1352);
and U2925 (N_2925,N_1758,N_1845);
or U2926 (N_2926,N_1498,N_1538);
or U2927 (N_2927,N_1465,N_1623);
nand U2928 (N_2928,N_1568,N_1902);
or U2929 (N_2929,N_1405,N_1336);
or U2930 (N_2930,N_1111,N_1822);
and U2931 (N_2931,N_1351,N_1172);
or U2932 (N_2932,N_1031,N_1432);
nand U2933 (N_2933,N_1949,N_1777);
xor U2934 (N_2934,N_1485,N_1172);
and U2935 (N_2935,N_1299,N_1122);
or U2936 (N_2936,N_1572,N_1305);
or U2937 (N_2937,N_1025,N_1816);
nor U2938 (N_2938,N_1400,N_1620);
nor U2939 (N_2939,N_1261,N_1143);
and U2940 (N_2940,N_1876,N_1561);
nor U2941 (N_2941,N_1069,N_1464);
xor U2942 (N_2942,N_1940,N_1636);
and U2943 (N_2943,N_1777,N_1510);
and U2944 (N_2944,N_1271,N_1368);
or U2945 (N_2945,N_1491,N_1226);
nor U2946 (N_2946,N_1709,N_1611);
nand U2947 (N_2947,N_1788,N_1218);
nand U2948 (N_2948,N_1930,N_1913);
nor U2949 (N_2949,N_1041,N_1762);
nor U2950 (N_2950,N_1870,N_1082);
nor U2951 (N_2951,N_1800,N_1225);
nand U2952 (N_2952,N_1940,N_1003);
nand U2953 (N_2953,N_1976,N_1254);
nand U2954 (N_2954,N_1847,N_1470);
nand U2955 (N_2955,N_1501,N_1248);
nand U2956 (N_2956,N_1193,N_1873);
nor U2957 (N_2957,N_1374,N_1565);
nand U2958 (N_2958,N_1104,N_1300);
nand U2959 (N_2959,N_1301,N_1923);
or U2960 (N_2960,N_1232,N_1105);
and U2961 (N_2961,N_1001,N_1959);
and U2962 (N_2962,N_1343,N_1960);
or U2963 (N_2963,N_1356,N_1111);
and U2964 (N_2964,N_1974,N_1562);
nand U2965 (N_2965,N_1546,N_1231);
or U2966 (N_2966,N_1560,N_1379);
nand U2967 (N_2967,N_1073,N_1481);
or U2968 (N_2968,N_1559,N_1601);
nand U2969 (N_2969,N_1333,N_1139);
and U2970 (N_2970,N_1474,N_1859);
and U2971 (N_2971,N_1322,N_1500);
and U2972 (N_2972,N_1796,N_1823);
or U2973 (N_2973,N_1016,N_1928);
nor U2974 (N_2974,N_1759,N_1376);
and U2975 (N_2975,N_1260,N_1726);
nand U2976 (N_2976,N_1740,N_1865);
nand U2977 (N_2977,N_1538,N_1194);
and U2978 (N_2978,N_1376,N_1260);
xnor U2979 (N_2979,N_1092,N_1395);
nand U2980 (N_2980,N_1967,N_1119);
nor U2981 (N_2981,N_1022,N_1190);
nor U2982 (N_2982,N_1865,N_1598);
or U2983 (N_2983,N_1079,N_1877);
or U2984 (N_2984,N_1374,N_1874);
and U2985 (N_2985,N_1686,N_1369);
nor U2986 (N_2986,N_1755,N_1432);
or U2987 (N_2987,N_1113,N_1786);
nand U2988 (N_2988,N_1309,N_1027);
nand U2989 (N_2989,N_1688,N_1596);
and U2990 (N_2990,N_1647,N_1221);
nor U2991 (N_2991,N_1979,N_1002);
or U2992 (N_2992,N_1653,N_1936);
and U2993 (N_2993,N_1273,N_1013);
and U2994 (N_2994,N_1394,N_1720);
or U2995 (N_2995,N_1501,N_1598);
or U2996 (N_2996,N_1400,N_1822);
and U2997 (N_2997,N_1020,N_1000);
nand U2998 (N_2998,N_1800,N_1265);
xnor U2999 (N_2999,N_1977,N_1975);
xnor U3000 (N_3000,N_2349,N_2692);
nor U3001 (N_3001,N_2250,N_2574);
and U3002 (N_3002,N_2750,N_2303);
and U3003 (N_3003,N_2737,N_2573);
nor U3004 (N_3004,N_2264,N_2643);
and U3005 (N_3005,N_2175,N_2465);
nor U3006 (N_3006,N_2145,N_2523);
or U3007 (N_3007,N_2867,N_2851);
nand U3008 (N_3008,N_2232,N_2255);
nor U3009 (N_3009,N_2583,N_2334);
nor U3010 (N_3010,N_2901,N_2990);
nand U3011 (N_3011,N_2393,N_2512);
nor U3012 (N_3012,N_2212,N_2454);
or U3013 (N_3013,N_2998,N_2056);
and U3014 (N_3014,N_2722,N_2738);
nor U3015 (N_3015,N_2272,N_2730);
nand U3016 (N_3016,N_2732,N_2556);
and U3017 (N_3017,N_2922,N_2505);
or U3018 (N_3018,N_2532,N_2872);
or U3019 (N_3019,N_2527,N_2641);
xnor U3020 (N_3020,N_2391,N_2161);
or U3021 (N_3021,N_2499,N_2447);
or U3022 (N_3022,N_2311,N_2474);
or U3023 (N_3023,N_2430,N_2126);
nor U3024 (N_3024,N_2899,N_2216);
or U3025 (N_3025,N_2453,N_2858);
nor U3026 (N_3026,N_2804,N_2617);
nand U3027 (N_3027,N_2397,N_2824);
nor U3028 (N_3028,N_2847,N_2050);
or U3029 (N_3029,N_2408,N_2038);
and U3030 (N_3030,N_2670,N_2096);
or U3031 (N_3031,N_2071,N_2261);
nand U3032 (N_3032,N_2906,N_2830);
nor U3033 (N_3033,N_2375,N_2542);
nand U3034 (N_3034,N_2884,N_2840);
nor U3035 (N_3035,N_2543,N_2023);
xor U3036 (N_3036,N_2213,N_2995);
nand U3037 (N_3037,N_2195,N_2024);
nand U3038 (N_3038,N_2235,N_2073);
and U3039 (N_3039,N_2686,N_2339);
nand U3040 (N_3040,N_2580,N_2194);
and U3041 (N_3041,N_2258,N_2870);
nor U3042 (N_3042,N_2887,N_2040);
nor U3043 (N_3043,N_2151,N_2618);
or U3044 (N_3044,N_2657,N_2306);
and U3045 (N_3045,N_2874,N_2090);
nor U3046 (N_3046,N_2985,N_2383);
nand U3047 (N_3047,N_2828,N_2677);
or U3048 (N_3048,N_2350,N_2415);
or U3049 (N_3049,N_2114,N_2822);
nand U3050 (N_3050,N_2109,N_2329);
nor U3051 (N_3051,N_2513,N_2490);
nand U3052 (N_3052,N_2136,N_2260);
nand U3053 (N_3053,N_2941,N_2243);
or U3054 (N_3054,N_2936,N_2110);
and U3055 (N_3055,N_2275,N_2278);
or U3056 (N_3056,N_2914,N_2797);
xor U3057 (N_3057,N_2077,N_2736);
nor U3058 (N_3058,N_2060,N_2094);
and U3059 (N_3059,N_2575,N_2705);
and U3060 (N_3060,N_2374,N_2353);
nand U3061 (N_3061,N_2898,N_2456);
nand U3062 (N_3062,N_2507,N_2020);
nor U3063 (N_3063,N_2860,N_2596);
nand U3064 (N_3064,N_2927,N_2209);
nor U3065 (N_3065,N_2504,N_2771);
nand U3066 (N_3066,N_2398,N_2116);
nand U3067 (N_3067,N_2183,N_2880);
nand U3068 (N_3068,N_2577,N_2103);
and U3069 (N_3069,N_2855,N_2091);
or U3070 (N_3070,N_2939,N_2702);
or U3071 (N_3071,N_2099,N_2917);
nor U3072 (N_3072,N_2912,N_2081);
and U3073 (N_3073,N_2761,N_2361);
and U3074 (N_3074,N_2545,N_2200);
nor U3075 (N_3075,N_2530,N_2274);
nor U3076 (N_3076,N_2399,N_2609);
or U3077 (N_3077,N_2957,N_2895);
and U3078 (N_3078,N_2841,N_2389);
nor U3079 (N_3079,N_2741,N_2902);
nand U3080 (N_3080,N_2432,N_2286);
or U3081 (N_3081,N_2291,N_2006);
nor U3082 (N_3082,N_2352,N_2777);
and U3083 (N_3083,N_2614,N_2446);
nand U3084 (N_3084,N_2612,N_2137);
nand U3085 (N_3085,N_2324,N_2564);
nand U3086 (N_3086,N_2593,N_2052);
or U3087 (N_3087,N_2214,N_2239);
and U3088 (N_3088,N_2540,N_2146);
nor U3089 (N_3089,N_2655,N_2791);
nor U3090 (N_3090,N_2699,N_2016);
nor U3091 (N_3091,N_2069,N_2220);
or U3092 (N_3092,N_2034,N_2503);
and U3093 (N_3093,N_2431,N_2179);
and U3094 (N_3094,N_2696,N_2994);
xnor U3095 (N_3095,N_2178,N_2581);
nor U3096 (N_3096,N_2520,N_2188);
or U3097 (N_3097,N_2392,N_2767);
or U3098 (N_3098,N_2054,N_2967);
or U3099 (N_3099,N_2719,N_2700);
or U3100 (N_3100,N_2043,N_2066);
and U3101 (N_3101,N_2658,N_2422);
nor U3102 (N_3102,N_2229,N_2904);
nand U3103 (N_3103,N_2506,N_2913);
xor U3104 (N_3104,N_2369,N_2916);
and U3105 (N_3105,N_2687,N_2438);
or U3106 (N_3106,N_2565,N_2315);
or U3107 (N_3107,N_2418,N_2186);
xnor U3108 (N_3108,N_2231,N_2153);
or U3109 (N_3109,N_2603,N_2343);
nor U3110 (N_3110,N_2570,N_2550);
xnor U3111 (N_3111,N_2846,N_2442);
xor U3112 (N_3112,N_2783,N_2591);
or U3113 (N_3113,N_2005,N_2210);
nor U3114 (N_3114,N_2367,N_2176);
nand U3115 (N_3115,N_2204,N_2265);
nand U3116 (N_3116,N_2063,N_2764);
nand U3117 (N_3117,N_2553,N_2225);
nor U3118 (N_3118,N_2423,N_2362);
or U3119 (N_3119,N_2585,N_2218);
nand U3120 (N_3120,N_2511,N_2586);
and U3121 (N_3121,N_2592,N_2160);
nand U3122 (N_3122,N_2835,N_2800);
and U3123 (N_3123,N_2781,N_2890);
nand U3124 (N_3124,N_2509,N_2246);
and U3125 (N_3125,N_2486,N_2171);
nor U3126 (N_3126,N_2597,N_2604);
nor U3127 (N_3127,N_2241,N_2107);
and U3128 (N_3128,N_2245,N_2120);
and U3129 (N_3129,N_2296,N_2372);
and U3130 (N_3130,N_2944,N_2298);
nand U3131 (N_3131,N_2785,N_2067);
nor U3132 (N_3132,N_2413,N_2108);
nor U3133 (N_3133,N_2388,N_2460);
and U3134 (N_3134,N_2875,N_2027);
and U3135 (N_3135,N_2009,N_2610);
nand U3136 (N_3136,N_2285,N_2811);
nor U3137 (N_3137,N_2684,N_2607);
nor U3138 (N_3138,N_2792,N_2414);
nand U3139 (N_3139,N_2975,N_2247);
or U3140 (N_3140,N_2588,N_2314);
and U3141 (N_3141,N_2908,N_2206);
nor U3142 (N_3142,N_2680,N_2058);
nand U3143 (N_3143,N_2668,N_2763);
nand U3144 (N_3144,N_2497,N_2991);
nand U3145 (N_3145,N_2467,N_2313);
and U3146 (N_3146,N_2862,N_2358);
or U3147 (N_3147,N_2886,N_2873);
nor U3148 (N_3148,N_2669,N_2778);
or U3149 (N_3149,N_2379,N_2814);
nor U3150 (N_3150,N_2159,N_2227);
nor U3151 (N_3151,N_2605,N_2333);
nor U3152 (N_3152,N_2646,N_2576);
and U3153 (N_3153,N_2582,N_2952);
nand U3154 (N_3154,N_2093,N_2428);
or U3155 (N_3155,N_2436,N_2953);
and U3156 (N_3156,N_2017,N_2253);
nor U3157 (N_3157,N_2788,N_2911);
and U3158 (N_3158,N_2674,N_2130);
and U3159 (N_3159,N_2373,N_2405);
and U3160 (N_3160,N_2602,N_2988);
xor U3161 (N_3161,N_2861,N_2080);
or U3162 (N_3162,N_2776,N_2173);
and U3163 (N_3163,N_2184,N_2878);
nor U3164 (N_3164,N_2008,N_2134);
or U3165 (N_3165,N_2749,N_2595);
nand U3166 (N_3166,N_2671,N_2335);
nand U3167 (N_3167,N_2106,N_2528);
or U3168 (N_3168,N_2224,N_2457);
nor U3169 (N_3169,N_2885,N_2572);
nor U3170 (N_3170,N_2562,N_2059);
xnor U3171 (N_3171,N_2336,N_2928);
or U3172 (N_3172,N_2407,N_2004);
nor U3173 (N_3173,N_2135,N_2088);
nand U3174 (N_3174,N_2471,N_2404);
nor U3175 (N_3175,N_2197,N_2117);
nor U3176 (N_3176,N_2337,N_2795);
or U3177 (N_3177,N_2755,N_2932);
or U3178 (N_3178,N_2466,N_2794);
or U3179 (N_3179,N_2089,N_2555);
nand U3180 (N_3180,N_2746,N_2829);
nand U3181 (N_3181,N_2376,N_2715);
and U3182 (N_3182,N_2538,N_2964);
and U3183 (N_3183,N_2305,N_2297);
and U3184 (N_3184,N_2561,N_2396);
and U3185 (N_3185,N_2843,N_2226);
or U3186 (N_3186,N_2720,N_2185);
nand U3187 (N_3187,N_2889,N_2891);
and U3188 (N_3188,N_2481,N_2918);
and U3189 (N_3189,N_2013,N_2723);
and U3190 (N_3190,N_2728,N_2429);
nor U3191 (N_3191,N_2650,N_2546);
nor U3192 (N_3192,N_2676,N_2790);
and U3193 (N_3193,N_2571,N_2635);
or U3194 (N_3194,N_2892,N_2782);
xnor U3195 (N_3195,N_2772,N_2667);
nand U3196 (N_3196,N_2271,N_2775);
nand U3197 (N_3197,N_2193,N_2118);
nor U3198 (N_3198,N_2266,N_2933);
nor U3199 (N_3199,N_2999,N_2122);
and U3200 (N_3200,N_2981,N_2385);
and U3201 (N_3201,N_2045,N_2087);
and U3202 (N_3202,N_2086,N_2425);
nor U3203 (N_3203,N_2476,N_2625);
or U3204 (N_3204,N_2132,N_2019);
and U3205 (N_3205,N_2718,N_2128);
xor U3206 (N_3206,N_2238,N_2690);
nor U3207 (N_3207,N_2064,N_2745);
nor U3208 (N_3208,N_2987,N_2100);
nand U3209 (N_3209,N_2281,N_2802);
nand U3210 (N_3210,N_2208,N_2934);
nand U3211 (N_3211,N_2410,N_2003);
or U3212 (N_3212,N_2269,N_2524);
and U3213 (N_3213,N_2021,N_2535);
or U3214 (N_3214,N_2234,N_2919);
or U3215 (N_3215,N_2356,N_2445);
or U3216 (N_3216,N_2864,N_2638);
nor U3217 (N_3217,N_2807,N_2784);
and U3218 (N_3218,N_2252,N_2223);
or U3219 (N_3219,N_2112,N_2307);
nor U3220 (N_3220,N_2289,N_2882);
or U3221 (N_3221,N_2833,N_2986);
or U3222 (N_3222,N_2863,N_2611);
nor U3223 (N_3223,N_2139,N_2150);
and U3224 (N_3224,N_2868,N_2158);
and U3225 (N_3225,N_2327,N_2222);
or U3226 (N_3226,N_2706,N_2810);
and U3227 (N_3227,N_2963,N_2945);
nand U3228 (N_3228,N_2549,N_2584);
nand U3229 (N_3229,N_2849,N_2664);
and U3230 (N_3230,N_2689,N_2850);
nor U3231 (N_3231,N_2133,N_2978);
nor U3232 (N_3232,N_2165,N_2039);
nand U3233 (N_3233,N_2636,N_2390);
nor U3234 (N_3234,N_2735,N_2464);
and U3235 (N_3235,N_2368,N_2237);
or U3236 (N_3236,N_2249,N_2779);
and U3237 (N_3237,N_2685,N_2082);
nand U3238 (N_3238,N_2248,N_2300);
or U3239 (N_3239,N_2030,N_2155);
and U3240 (N_3240,N_2470,N_2263);
nor U3241 (N_3241,N_2979,N_2798);
nor U3242 (N_3242,N_2703,N_2473);
nor U3243 (N_3243,N_2923,N_2493);
nor U3244 (N_3244,N_2113,N_2192);
nand U3245 (N_3245,N_2515,N_2381);
nor U3246 (N_3246,N_2925,N_2697);
and U3247 (N_3247,N_2345,N_2616);
and U3248 (N_3248,N_2101,N_2085);
nand U3249 (N_3249,N_2837,N_2187);
or U3250 (N_3250,N_2451,N_2731);
nand U3251 (N_3251,N_2037,N_2724);
or U3252 (N_3252,N_2725,N_2644);
nor U3253 (N_3253,N_2156,N_2753);
and U3254 (N_3254,N_2522,N_2386);
nor U3255 (N_3255,N_2627,N_2443);
nor U3256 (N_3256,N_2105,N_2487);
xnor U3257 (N_3257,N_2817,N_2548);
xor U3258 (N_3258,N_2962,N_2519);
and U3259 (N_3259,N_2931,N_2201);
nor U3260 (N_3260,N_2104,N_2531);
or U3261 (N_3261,N_2097,N_2510);
or U3262 (N_3262,N_2083,N_2848);
and U3263 (N_3263,N_2463,N_2707);
nand U3264 (N_3264,N_2025,N_2529);
and U3265 (N_3265,N_2310,N_2541);
and U3266 (N_3266,N_2808,N_2946);
nor U3267 (N_3267,N_2818,N_2279);
or U3268 (N_3268,N_2384,N_2163);
and U3269 (N_3269,N_2293,N_2240);
nand U3270 (N_3270,N_2836,N_2256);
or U3271 (N_3271,N_2357,N_2558);
or U3272 (N_3272,N_2951,N_2041);
or U3273 (N_3273,N_2640,N_2320);
or U3274 (N_3274,N_2970,N_2733);
and U3275 (N_3275,N_2370,N_2325);
or U3276 (N_3276,N_2960,N_2626);
and U3277 (N_3277,N_2949,N_2992);
and U3278 (N_3278,N_2439,N_2434);
nor U3279 (N_3279,N_2773,N_2806);
and U3280 (N_3280,N_2055,N_2965);
nor U3281 (N_3281,N_2950,N_2092);
nand U3282 (N_3282,N_2228,N_2714);
or U3283 (N_3283,N_2031,N_2075);
nor U3284 (N_3284,N_2483,N_2517);
xor U3285 (N_3285,N_2681,N_2799);
nand U3286 (N_3286,N_2477,N_2198);
or U3287 (N_3287,N_2654,N_2959);
nor U3288 (N_3288,N_2495,N_2012);
or U3289 (N_3289,N_2624,N_2461);
nand U3290 (N_3290,N_2935,N_2061);
nor U3291 (N_3291,N_2141,N_2629);
or U3292 (N_3292,N_2569,N_2380);
nor U3293 (N_3293,N_2876,N_2170);
and U3294 (N_3294,N_2652,N_2757);
nor U3295 (N_3295,N_2257,N_2955);
or U3296 (N_3296,N_2202,N_2268);
and U3297 (N_3297,N_2734,N_2827);
nor U3298 (N_3298,N_2956,N_2172);
or U3299 (N_3299,N_2857,N_2930);
or U3300 (N_3300,N_2653,N_2400);
and U3301 (N_3301,N_2717,N_2309);
nor U3302 (N_3302,N_2416,N_2823);
and U3303 (N_3303,N_2974,N_2844);
nor U3304 (N_3304,N_2666,N_2539);
nor U3305 (N_3305,N_2437,N_2996);
xnor U3306 (N_3306,N_2364,N_2102);
or U3307 (N_3307,N_2015,N_2754);
xor U3308 (N_3308,N_2929,N_2623);
or U3309 (N_3309,N_2351,N_2319);
or U3310 (N_3310,N_2149,N_2270);
nand U3311 (N_3311,N_2651,N_2694);
and U3312 (N_3312,N_2682,N_2328);
and U3313 (N_3313,N_2182,N_2018);
nor U3314 (N_3314,N_2450,N_2663);
nor U3315 (N_3315,N_2290,N_2154);
and U3316 (N_3316,N_2683,N_2566);
nand U3317 (N_3317,N_2633,N_2712);
and U3318 (N_3318,N_2809,N_2805);
or U3319 (N_3319,N_2752,N_2262);
and U3320 (N_3320,N_2125,N_2815);
nand U3321 (N_3321,N_2982,N_2711);
nand U3322 (N_3322,N_2710,N_2007);
or U3323 (N_3323,N_2924,N_2634);
and U3324 (N_3324,N_2441,N_2747);
or U3325 (N_3325,N_2331,N_2205);
nand U3326 (N_3326,N_2244,N_2793);
xor U3327 (N_3327,N_2518,N_2148);
and U3328 (N_3328,N_2427,N_2387);
nor U3329 (N_3329,N_2199,N_2395);
nand U3330 (N_3330,N_2332,N_2675);
nand U3331 (N_3331,N_2971,N_2462);
nor U3332 (N_3332,N_2283,N_2288);
nand U3333 (N_3333,N_2533,N_2940);
and U3334 (N_3334,N_2869,N_2508);
and U3335 (N_3335,N_2742,N_2559);
nand U3336 (N_3336,N_2406,N_2409);
nand U3337 (N_3337,N_2346,N_2131);
or U3338 (N_3338,N_2338,N_2937);
nor U3339 (N_3339,N_2412,N_2028);
and U3340 (N_3340,N_2853,N_2174);
or U3341 (N_3341,N_2276,N_2537);
nand U3342 (N_3342,N_2280,N_2299);
or U3343 (N_3343,N_2177,N_2302);
nor U3344 (N_3344,N_2267,N_2014);
nor U3345 (N_3345,N_2900,N_2852);
or U3346 (N_3346,N_2993,N_2947);
or U3347 (N_3347,N_2579,N_2147);
and U3348 (N_3348,N_2044,N_2312);
nor U3349 (N_3349,N_2648,N_2502);
nand U3350 (N_3350,N_2046,N_2424);
nor U3351 (N_3351,N_2854,N_2812);
or U3352 (N_3352,N_2448,N_2219);
and U3353 (N_3353,N_2084,N_2047);
and U3354 (N_3354,N_2976,N_2000);
nor U3355 (N_3355,N_2766,N_2938);
nor U3356 (N_3356,N_2078,N_2709);
and U3357 (N_3357,N_2726,N_2825);
nor U3358 (N_3358,N_2287,N_2284);
or U3359 (N_3359,N_2661,N_2679);
nand U3360 (N_3360,N_2521,N_2613);
nor U3361 (N_3361,N_2273,N_2316);
or U3362 (N_3362,N_2968,N_2758);
nand U3363 (N_3363,N_2589,N_2032);
nand U3364 (N_3364,N_2123,N_2926);
and U3365 (N_3365,N_2639,N_2943);
or U3366 (N_3366,N_2888,N_2601);
nand U3367 (N_3367,N_2124,N_2563);
nand U3368 (N_3368,N_2157,N_2164);
and U3369 (N_3369,N_2484,N_2347);
and U3370 (N_3370,N_2421,N_2479);
nand U3371 (N_3371,N_2762,N_2905);
and U3372 (N_3372,N_2656,N_2739);
and U3373 (N_3373,N_2866,N_2637);
nand U3374 (N_3374,N_2485,N_2578);
or U3375 (N_3375,N_2459,N_2010);
and U3376 (N_3376,N_2002,N_2631);
and U3377 (N_3377,N_2254,N_2366);
nand U3378 (N_3378,N_2525,N_2673);
or U3379 (N_3379,N_2475,N_2662);
or U3380 (N_3380,N_2909,N_2062);
xnor U3381 (N_3381,N_2534,N_2033);
nor U3382 (N_3382,N_2615,N_2468);
nand U3383 (N_3383,N_2127,N_2594);
and U3384 (N_3384,N_2233,N_2590);
and U3385 (N_3385,N_2355,N_2167);
and U3386 (N_3386,N_2743,N_2645);
nand U3387 (N_3387,N_2879,N_2304);
or U3388 (N_3388,N_2619,N_2954);
or U3389 (N_3389,N_2942,N_2897);
and U3390 (N_3390,N_2472,N_2189);
and U3391 (N_3391,N_2259,N_2251);
nor U3392 (N_3392,N_2560,N_2877);
and U3393 (N_3393,N_2526,N_2342);
nand U3394 (N_3394,N_2688,N_2277);
or U3395 (N_3395,N_2984,N_2360);
or U3396 (N_3396,N_2865,N_2098);
nor U3397 (N_3397,N_2660,N_2547);
or U3398 (N_3398,N_2042,N_2378);
and U3399 (N_3399,N_2301,N_2318);
or U3400 (N_3400,N_2983,N_2621);
nand U3401 (N_3401,N_2444,N_2910);
nand U3402 (N_3402,N_2420,N_2191);
and U3403 (N_3403,N_2842,N_2138);
nor U3404 (N_3404,N_2972,N_2215);
or U3405 (N_3405,N_2980,N_2751);
and U3406 (N_3406,N_2469,N_2704);
or U3407 (N_3407,N_2359,N_2903);
or U3408 (N_3408,N_2449,N_2121);
or U3409 (N_3409,N_2744,N_2452);
or U3410 (N_3410,N_2948,N_2691);
nor U3411 (N_3411,N_2647,N_2458);
nor U3412 (N_3412,N_2433,N_2029);
nand U3413 (N_3413,N_2966,N_2317);
nand U3414 (N_3414,N_2169,N_2881);
or U3415 (N_3415,N_2419,N_2494);
and U3416 (N_3416,N_2819,N_2321);
and U3417 (N_3417,N_2768,N_2838);
or U3418 (N_3418,N_2190,N_2587);
and U3419 (N_3419,N_2893,N_2813);
or U3420 (N_3420,N_2363,N_2382);
nor U3421 (N_3421,N_2140,N_2856);
nor U3422 (N_3422,N_2816,N_2217);
nand U3423 (N_3423,N_2035,N_2871);
nand U3424 (N_3424,N_2894,N_2834);
and U3425 (N_3425,N_2920,N_2440);
nor U3426 (N_3426,N_2011,N_2567);
nor U3427 (N_3427,N_2072,N_2721);
and U3428 (N_3428,N_2482,N_2552);
or U3429 (N_3429,N_2780,N_2230);
xor U3430 (N_3430,N_2770,N_2606);
xnor U3431 (N_3431,N_2142,N_2065);
nor U3432 (N_3432,N_2119,N_2501);
and U3433 (N_3433,N_2211,N_2701);
nor U3434 (N_3434,N_2649,N_2354);
nand U3435 (N_3435,N_2969,N_2115);
and U3436 (N_3436,N_2492,N_2070);
nand U3437 (N_3437,N_2292,N_2074);
and U3438 (N_3438,N_2774,N_2491);
nand U3439 (N_3439,N_2756,N_2435);
and U3440 (N_3440,N_2129,N_2236);
and U3441 (N_3441,N_2196,N_2095);
nor U3442 (N_3442,N_2557,N_2480);
nand U3443 (N_3443,N_2402,N_2308);
and U3444 (N_3444,N_2678,N_2977);
nor U3445 (N_3445,N_2371,N_2989);
nand U3446 (N_3446,N_2144,N_2551);
nand U3447 (N_3447,N_2598,N_2068);
or U3448 (N_3448,N_2665,N_2348);
or U3449 (N_3449,N_2554,N_2789);
nand U3450 (N_3450,N_2053,N_2973);
nand U3451 (N_3451,N_2915,N_2426);
nand U3452 (N_3452,N_2496,N_2727);
and U3453 (N_3453,N_2997,N_2831);
nand U3454 (N_3454,N_2516,N_2203);
or U3455 (N_3455,N_2111,N_2401);
and U3456 (N_3456,N_2760,N_2455);
nand U3457 (N_3457,N_2608,N_2026);
or U3458 (N_3458,N_2411,N_2417);
nor U3459 (N_3459,N_2143,N_2659);
nor U3460 (N_3460,N_2330,N_2620);
nand U3461 (N_3461,N_2821,N_2180);
nand U3462 (N_3462,N_2498,N_2832);
or U3463 (N_3463,N_2672,N_2036);
nor U3464 (N_3464,N_2907,N_2883);
xnor U3465 (N_3465,N_2921,N_2796);
and U3466 (N_3466,N_2786,N_2207);
or U3467 (N_3467,N_2489,N_2168);
and U3468 (N_3468,N_2740,N_2748);
nor U3469 (N_3469,N_2322,N_2787);
and U3470 (N_3470,N_2152,N_2820);
and U3471 (N_3471,N_2695,N_2403);
nor U3472 (N_3472,N_2765,N_2057);
nor U3473 (N_3473,N_2632,N_2051);
nor U3474 (N_3474,N_2488,N_2630);
or U3475 (N_3475,N_2622,N_2162);
nor U3476 (N_3476,N_2708,N_2394);
nand U3477 (N_3477,N_2377,N_2323);
nand U3478 (N_3478,N_2599,N_2826);
and U3479 (N_3479,N_2166,N_2845);
nand U3480 (N_3480,N_2803,N_2544);
xnor U3481 (N_3481,N_2295,N_2769);
nand U3482 (N_3482,N_2958,N_2628);
or U3483 (N_3483,N_2500,N_2242);
nor U3484 (N_3484,N_2282,N_2079);
and U3485 (N_3485,N_2642,N_2365);
nor U3486 (N_3486,N_2514,N_2181);
nand U3487 (N_3487,N_2048,N_2716);
nor U3488 (N_3488,N_2340,N_2961);
or U3489 (N_3489,N_2693,N_2839);
or U3490 (N_3490,N_2896,N_2478);
nand U3491 (N_3491,N_2568,N_2049);
and U3492 (N_3492,N_2759,N_2344);
or U3493 (N_3493,N_2001,N_2600);
or U3494 (N_3494,N_2729,N_2536);
nand U3495 (N_3495,N_2076,N_2022);
or U3496 (N_3496,N_2294,N_2801);
and U3497 (N_3497,N_2326,N_2859);
nand U3498 (N_3498,N_2221,N_2698);
nor U3499 (N_3499,N_2713,N_2341);
nor U3500 (N_3500,N_2844,N_2784);
and U3501 (N_3501,N_2212,N_2147);
nor U3502 (N_3502,N_2491,N_2792);
or U3503 (N_3503,N_2545,N_2191);
nor U3504 (N_3504,N_2509,N_2945);
nor U3505 (N_3505,N_2371,N_2596);
nand U3506 (N_3506,N_2203,N_2220);
and U3507 (N_3507,N_2846,N_2894);
nor U3508 (N_3508,N_2439,N_2572);
nor U3509 (N_3509,N_2412,N_2943);
nor U3510 (N_3510,N_2750,N_2343);
xnor U3511 (N_3511,N_2036,N_2904);
and U3512 (N_3512,N_2802,N_2771);
nand U3513 (N_3513,N_2992,N_2917);
or U3514 (N_3514,N_2751,N_2513);
xnor U3515 (N_3515,N_2481,N_2456);
or U3516 (N_3516,N_2671,N_2175);
or U3517 (N_3517,N_2014,N_2606);
or U3518 (N_3518,N_2162,N_2986);
xnor U3519 (N_3519,N_2677,N_2507);
and U3520 (N_3520,N_2115,N_2752);
nor U3521 (N_3521,N_2604,N_2484);
nor U3522 (N_3522,N_2218,N_2835);
or U3523 (N_3523,N_2931,N_2646);
nand U3524 (N_3524,N_2064,N_2784);
nand U3525 (N_3525,N_2592,N_2882);
or U3526 (N_3526,N_2288,N_2573);
nand U3527 (N_3527,N_2779,N_2121);
and U3528 (N_3528,N_2982,N_2039);
nand U3529 (N_3529,N_2871,N_2761);
nor U3530 (N_3530,N_2489,N_2152);
and U3531 (N_3531,N_2663,N_2399);
and U3532 (N_3532,N_2207,N_2351);
nand U3533 (N_3533,N_2607,N_2521);
nor U3534 (N_3534,N_2733,N_2720);
and U3535 (N_3535,N_2895,N_2520);
nand U3536 (N_3536,N_2605,N_2538);
nand U3537 (N_3537,N_2860,N_2520);
nand U3538 (N_3538,N_2787,N_2391);
or U3539 (N_3539,N_2053,N_2016);
nor U3540 (N_3540,N_2287,N_2033);
and U3541 (N_3541,N_2577,N_2437);
and U3542 (N_3542,N_2260,N_2518);
nor U3543 (N_3543,N_2510,N_2849);
or U3544 (N_3544,N_2282,N_2377);
or U3545 (N_3545,N_2047,N_2794);
nor U3546 (N_3546,N_2383,N_2394);
nor U3547 (N_3547,N_2393,N_2732);
or U3548 (N_3548,N_2926,N_2719);
nand U3549 (N_3549,N_2825,N_2872);
and U3550 (N_3550,N_2893,N_2962);
nand U3551 (N_3551,N_2524,N_2240);
and U3552 (N_3552,N_2101,N_2878);
or U3553 (N_3553,N_2080,N_2008);
nor U3554 (N_3554,N_2452,N_2571);
or U3555 (N_3555,N_2668,N_2090);
nand U3556 (N_3556,N_2873,N_2325);
or U3557 (N_3557,N_2471,N_2255);
nor U3558 (N_3558,N_2863,N_2571);
and U3559 (N_3559,N_2113,N_2668);
nand U3560 (N_3560,N_2890,N_2281);
nand U3561 (N_3561,N_2976,N_2536);
or U3562 (N_3562,N_2734,N_2053);
nor U3563 (N_3563,N_2418,N_2594);
or U3564 (N_3564,N_2646,N_2670);
or U3565 (N_3565,N_2825,N_2006);
nor U3566 (N_3566,N_2465,N_2328);
or U3567 (N_3567,N_2995,N_2504);
or U3568 (N_3568,N_2649,N_2522);
nand U3569 (N_3569,N_2613,N_2325);
nor U3570 (N_3570,N_2506,N_2364);
and U3571 (N_3571,N_2439,N_2738);
nand U3572 (N_3572,N_2128,N_2770);
nand U3573 (N_3573,N_2535,N_2946);
or U3574 (N_3574,N_2705,N_2821);
nand U3575 (N_3575,N_2879,N_2197);
nand U3576 (N_3576,N_2926,N_2568);
nor U3577 (N_3577,N_2565,N_2557);
nand U3578 (N_3578,N_2129,N_2253);
or U3579 (N_3579,N_2256,N_2324);
xnor U3580 (N_3580,N_2131,N_2591);
or U3581 (N_3581,N_2922,N_2253);
or U3582 (N_3582,N_2176,N_2414);
or U3583 (N_3583,N_2405,N_2519);
xor U3584 (N_3584,N_2178,N_2835);
nand U3585 (N_3585,N_2631,N_2951);
and U3586 (N_3586,N_2403,N_2486);
or U3587 (N_3587,N_2451,N_2886);
or U3588 (N_3588,N_2352,N_2599);
nand U3589 (N_3589,N_2865,N_2888);
nor U3590 (N_3590,N_2436,N_2506);
nor U3591 (N_3591,N_2908,N_2493);
or U3592 (N_3592,N_2634,N_2249);
nor U3593 (N_3593,N_2200,N_2810);
nor U3594 (N_3594,N_2422,N_2474);
nor U3595 (N_3595,N_2071,N_2000);
nor U3596 (N_3596,N_2763,N_2247);
nor U3597 (N_3597,N_2126,N_2659);
and U3598 (N_3598,N_2855,N_2557);
nand U3599 (N_3599,N_2301,N_2971);
and U3600 (N_3600,N_2192,N_2481);
nor U3601 (N_3601,N_2274,N_2603);
and U3602 (N_3602,N_2150,N_2198);
or U3603 (N_3603,N_2642,N_2245);
xnor U3604 (N_3604,N_2538,N_2097);
or U3605 (N_3605,N_2189,N_2805);
and U3606 (N_3606,N_2371,N_2247);
xnor U3607 (N_3607,N_2411,N_2134);
nand U3608 (N_3608,N_2011,N_2354);
nand U3609 (N_3609,N_2339,N_2404);
and U3610 (N_3610,N_2456,N_2876);
xor U3611 (N_3611,N_2884,N_2747);
nor U3612 (N_3612,N_2896,N_2091);
or U3613 (N_3613,N_2563,N_2916);
nor U3614 (N_3614,N_2509,N_2056);
and U3615 (N_3615,N_2570,N_2067);
and U3616 (N_3616,N_2307,N_2815);
or U3617 (N_3617,N_2810,N_2035);
nand U3618 (N_3618,N_2732,N_2182);
nor U3619 (N_3619,N_2045,N_2102);
nand U3620 (N_3620,N_2659,N_2708);
nand U3621 (N_3621,N_2616,N_2957);
nor U3622 (N_3622,N_2510,N_2768);
or U3623 (N_3623,N_2932,N_2536);
and U3624 (N_3624,N_2419,N_2973);
or U3625 (N_3625,N_2964,N_2896);
or U3626 (N_3626,N_2260,N_2720);
nand U3627 (N_3627,N_2470,N_2336);
nor U3628 (N_3628,N_2928,N_2982);
nand U3629 (N_3629,N_2368,N_2458);
nor U3630 (N_3630,N_2023,N_2900);
xnor U3631 (N_3631,N_2809,N_2708);
xnor U3632 (N_3632,N_2814,N_2448);
nor U3633 (N_3633,N_2617,N_2474);
and U3634 (N_3634,N_2684,N_2613);
and U3635 (N_3635,N_2584,N_2410);
nor U3636 (N_3636,N_2361,N_2302);
or U3637 (N_3637,N_2851,N_2043);
and U3638 (N_3638,N_2211,N_2466);
and U3639 (N_3639,N_2373,N_2817);
nand U3640 (N_3640,N_2773,N_2741);
nor U3641 (N_3641,N_2964,N_2246);
or U3642 (N_3642,N_2671,N_2249);
nor U3643 (N_3643,N_2017,N_2349);
and U3644 (N_3644,N_2900,N_2819);
xnor U3645 (N_3645,N_2151,N_2555);
nor U3646 (N_3646,N_2388,N_2837);
or U3647 (N_3647,N_2760,N_2498);
or U3648 (N_3648,N_2464,N_2855);
xor U3649 (N_3649,N_2478,N_2021);
and U3650 (N_3650,N_2510,N_2714);
nor U3651 (N_3651,N_2594,N_2520);
nand U3652 (N_3652,N_2416,N_2422);
nand U3653 (N_3653,N_2323,N_2467);
nor U3654 (N_3654,N_2959,N_2308);
xor U3655 (N_3655,N_2030,N_2138);
nor U3656 (N_3656,N_2216,N_2029);
nor U3657 (N_3657,N_2558,N_2402);
nand U3658 (N_3658,N_2054,N_2583);
nor U3659 (N_3659,N_2757,N_2355);
and U3660 (N_3660,N_2865,N_2814);
or U3661 (N_3661,N_2984,N_2676);
and U3662 (N_3662,N_2355,N_2001);
or U3663 (N_3663,N_2484,N_2088);
and U3664 (N_3664,N_2713,N_2646);
nor U3665 (N_3665,N_2520,N_2226);
nor U3666 (N_3666,N_2712,N_2696);
nand U3667 (N_3667,N_2702,N_2647);
nand U3668 (N_3668,N_2254,N_2942);
nand U3669 (N_3669,N_2500,N_2508);
and U3670 (N_3670,N_2394,N_2150);
or U3671 (N_3671,N_2937,N_2242);
nand U3672 (N_3672,N_2967,N_2959);
and U3673 (N_3673,N_2372,N_2651);
nand U3674 (N_3674,N_2656,N_2391);
nor U3675 (N_3675,N_2039,N_2950);
or U3676 (N_3676,N_2095,N_2067);
nor U3677 (N_3677,N_2524,N_2737);
or U3678 (N_3678,N_2186,N_2746);
nand U3679 (N_3679,N_2687,N_2008);
nor U3680 (N_3680,N_2818,N_2278);
and U3681 (N_3681,N_2728,N_2583);
or U3682 (N_3682,N_2284,N_2633);
and U3683 (N_3683,N_2162,N_2168);
nor U3684 (N_3684,N_2628,N_2605);
nand U3685 (N_3685,N_2718,N_2176);
nor U3686 (N_3686,N_2707,N_2635);
nor U3687 (N_3687,N_2010,N_2643);
or U3688 (N_3688,N_2548,N_2224);
or U3689 (N_3689,N_2099,N_2913);
xnor U3690 (N_3690,N_2008,N_2883);
or U3691 (N_3691,N_2132,N_2792);
and U3692 (N_3692,N_2852,N_2818);
nand U3693 (N_3693,N_2257,N_2732);
and U3694 (N_3694,N_2749,N_2044);
nand U3695 (N_3695,N_2376,N_2510);
or U3696 (N_3696,N_2270,N_2084);
xnor U3697 (N_3697,N_2968,N_2819);
or U3698 (N_3698,N_2795,N_2901);
nand U3699 (N_3699,N_2900,N_2135);
nor U3700 (N_3700,N_2552,N_2945);
nand U3701 (N_3701,N_2089,N_2682);
or U3702 (N_3702,N_2924,N_2777);
nand U3703 (N_3703,N_2005,N_2739);
nor U3704 (N_3704,N_2522,N_2933);
nor U3705 (N_3705,N_2582,N_2842);
nand U3706 (N_3706,N_2132,N_2308);
nand U3707 (N_3707,N_2391,N_2297);
nor U3708 (N_3708,N_2648,N_2171);
or U3709 (N_3709,N_2375,N_2819);
and U3710 (N_3710,N_2212,N_2921);
nand U3711 (N_3711,N_2099,N_2461);
or U3712 (N_3712,N_2649,N_2964);
and U3713 (N_3713,N_2127,N_2178);
or U3714 (N_3714,N_2113,N_2107);
or U3715 (N_3715,N_2912,N_2548);
nor U3716 (N_3716,N_2519,N_2011);
nand U3717 (N_3717,N_2506,N_2347);
xnor U3718 (N_3718,N_2236,N_2751);
nand U3719 (N_3719,N_2851,N_2633);
or U3720 (N_3720,N_2277,N_2670);
or U3721 (N_3721,N_2858,N_2518);
nor U3722 (N_3722,N_2428,N_2101);
or U3723 (N_3723,N_2550,N_2536);
or U3724 (N_3724,N_2648,N_2207);
or U3725 (N_3725,N_2855,N_2190);
nor U3726 (N_3726,N_2227,N_2875);
nand U3727 (N_3727,N_2040,N_2431);
nand U3728 (N_3728,N_2399,N_2504);
nand U3729 (N_3729,N_2843,N_2076);
nand U3730 (N_3730,N_2186,N_2772);
nor U3731 (N_3731,N_2040,N_2816);
nand U3732 (N_3732,N_2446,N_2702);
nand U3733 (N_3733,N_2256,N_2584);
nor U3734 (N_3734,N_2815,N_2829);
or U3735 (N_3735,N_2106,N_2810);
nor U3736 (N_3736,N_2061,N_2609);
nor U3737 (N_3737,N_2073,N_2728);
nand U3738 (N_3738,N_2949,N_2790);
or U3739 (N_3739,N_2694,N_2492);
nor U3740 (N_3740,N_2845,N_2721);
or U3741 (N_3741,N_2936,N_2594);
nor U3742 (N_3742,N_2867,N_2392);
nand U3743 (N_3743,N_2780,N_2898);
or U3744 (N_3744,N_2943,N_2636);
nand U3745 (N_3745,N_2595,N_2014);
nor U3746 (N_3746,N_2726,N_2922);
nand U3747 (N_3747,N_2761,N_2244);
or U3748 (N_3748,N_2451,N_2745);
nor U3749 (N_3749,N_2595,N_2006);
or U3750 (N_3750,N_2225,N_2712);
nand U3751 (N_3751,N_2122,N_2471);
nor U3752 (N_3752,N_2990,N_2669);
or U3753 (N_3753,N_2297,N_2278);
nor U3754 (N_3754,N_2303,N_2200);
xor U3755 (N_3755,N_2843,N_2577);
nand U3756 (N_3756,N_2390,N_2338);
nor U3757 (N_3757,N_2662,N_2347);
nand U3758 (N_3758,N_2011,N_2418);
nor U3759 (N_3759,N_2143,N_2947);
nor U3760 (N_3760,N_2747,N_2830);
nor U3761 (N_3761,N_2085,N_2726);
or U3762 (N_3762,N_2630,N_2899);
nor U3763 (N_3763,N_2072,N_2319);
or U3764 (N_3764,N_2561,N_2318);
or U3765 (N_3765,N_2621,N_2073);
nor U3766 (N_3766,N_2647,N_2305);
or U3767 (N_3767,N_2002,N_2336);
or U3768 (N_3768,N_2167,N_2954);
or U3769 (N_3769,N_2367,N_2446);
and U3770 (N_3770,N_2318,N_2860);
nor U3771 (N_3771,N_2500,N_2445);
and U3772 (N_3772,N_2674,N_2212);
nand U3773 (N_3773,N_2154,N_2933);
nor U3774 (N_3774,N_2052,N_2456);
and U3775 (N_3775,N_2276,N_2258);
and U3776 (N_3776,N_2702,N_2771);
nor U3777 (N_3777,N_2253,N_2467);
and U3778 (N_3778,N_2309,N_2791);
nand U3779 (N_3779,N_2974,N_2007);
nand U3780 (N_3780,N_2462,N_2344);
and U3781 (N_3781,N_2081,N_2871);
and U3782 (N_3782,N_2453,N_2329);
nor U3783 (N_3783,N_2530,N_2907);
nor U3784 (N_3784,N_2723,N_2171);
or U3785 (N_3785,N_2475,N_2354);
and U3786 (N_3786,N_2439,N_2479);
nor U3787 (N_3787,N_2789,N_2629);
nand U3788 (N_3788,N_2572,N_2236);
nor U3789 (N_3789,N_2195,N_2788);
and U3790 (N_3790,N_2887,N_2594);
nor U3791 (N_3791,N_2995,N_2135);
nor U3792 (N_3792,N_2902,N_2777);
or U3793 (N_3793,N_2083,N_2589);
or U3794 (N_3794,N_2617,N_2619);
or U3795 (N_3795,N_2261,N_2491);
or U3796 (N_3796,N_2480,N_2256);
nand U3797 (N_3797,N_2096,N_2163);
and U3798 (N_3798,N_2204,N_2547);
and U3799 (N_3799,N_2716,N_2266);
nand U3800 (N_3800,N_2852,N_2555);
and U3801 (N_3801,N_2401,N_2860);
nand U3802 (N_3802,N_2695,N_2802);
and U3803 (N_3803,N_2425,N_2770);
and U3804 (N_3804,N_2818,N_2013);
nand U3805 (N_3805,N_2672,N_2711);
nand U3806 (N_3806,N_2348,N_2440);
nand U3807 (N_3807,N_2974,N_2650);
xor U3808 (N_3808,N_2454,N_2912);
or U3809 (N_3809,N_2399,N_2859);
nor U3810 (N_3810,N_2160,N_2343);
or U3811 (N_3811,N_2841,N_2489);
or U3812 (N_3812,N_2551,N_2650);
nor U3813 (N_3813,N_2468,N_2248);
and U3814 (N_3814,N_2530,N_2519);
nand U3815 (N_3815,N_2732,N_2055);
or U3816 (N_3816,N_2846,N_2736);
or U3817 (N_3817,N_2461,N_2410);
nor U3818 (N_3818,N_2907,N_2641);
nor U3819 (N_3819,N_2988,N_2607);
nand U3820 (N_3820,N_2222,N_2943);
and U3821 (N_3821,N_2467,N_2769);
or U3822 (N_3822,N_2117,N_2835);
nor U3823 (N_3823,N_2305,N_2025);
nor U3824 (N_3824,N_2324,N_2649);
and U3825 (N_3825,N_2743,N_2936);
or U3826 (N_3826,N_2018,N_2906);
nand U3827 (N_3827,N_2172,N_2645);
nand U3828 (N_3828,N_2990,N_2045);
or U3829 (N_3829,N_2922,N_2901);
nor U3830 (N_3830,N_2763,N_2495);
nor U3831 (N_3831,N_2951,N_2822);
nor U3832 (N_3832,N_2370,N_2838);
or U3833 (N_3833,N_2376,N_2166);
nor U3834 (N_3834,N_2998,N_2048);
and U3835 (N_3835,N_2161,N_2207);
and U3836 (N_3836,N_2335,N_2523);
and U3837 (N_3837,N_2841,N_2895);
nor U3838 (N_3838,N_2717,N_2385);
or U3839 (N_3839,N_2753,N_2526);
nor U3840 (N_3840,N_2297,N_2969);
and U3841 (N_3841,N_2484,N_2212);
xor U3842 (N_3842,N_2377,N_2564);
or U3843 (N_3843,N_2652,N_2569);
and U3844 (N_3844,N_2616,N_2481);
or U3845 (N_3845,N_2105,N_2679);
xor U3846 (N_3846,N_2489,N_2917);
xor U3847 (N_3847,N_2210,N_2727);
and U3848 (N_3848,N_2816,N_2036);
and U3849 (N_3849,N_2442,N_2142);
nor U3850 (N_3850,N_2857,N_2722);
or U3851 (N_3851,N_2011,N_2939);
or U3852 (N_3852,N_2943,N_2427);
nor U3853 (N_3853,N_2353,N_2058);
nor U3854 (N_3854,N_2269,N_2438);
and U3855 (N_3855,N_2118,N_2391);
nand U3856 (N_3856,N_2543,N_2196);
and U3857 (N_3857,N_2756,N_2293);
and U3858 (N_3858,N_2726,N_2958);
nor U3859 (N_3859,N_2510,N_2012);
nor U3860 (N_3860,N_2894,N_2447);
nor U3861 (N_3861,N_2462,N_2879);
nand U3862 (N_3862,N_2096,N_2259);
and U3863 (N_3863,N_2982,N_2323);
and U3864 (N_3864,N_2385,N_2996);
nor U3865 (N_3865,N_2721,N_2095);
or U3866 (N_3866,N_2491,N_2083);
or U3867 (N_3867,N_2686,N_2385);
and U3868 (N_3868,N_2440,N_2417);
xor U3869 (N_3869,N_2707,N_2173);
and U3870 (N_3870,N_2743,N_2971);
nand U3871 (N_3871,N_2106,N_2847);
nor U3872 (N_3872,N_2680,N_2767);
and U3873 (N_3873,N_2912,N_2780);
nor U3874 (N_3874,N_2420,N_2075);
nand U3875 (N_3875,N_2191,N_2396);
and U3876 (N_3876,N_2064,N_2261);
or U3877 (N_3877,N_2634,N_2780);
nor U3878 (N_3878,N_2560,N_2508);
or U3879 (N_3879,N_2922,N_2630);
and U3880 (N_3880,N_2659,N_2709);
or U3881 (N_3881,N_2559,N_2288);
or U3882 (N_3882,N_2979,N_2762);
and U3883 (N_3883,N_2906,N_2601);
or U3884 (N_3884,N_2120,N_2232);
and U3885 (N_3885,N_2581,N_2966);
and U3886 (N_3886,N_2458,N_2063);
or U3887 (N_3887,N_2332,N_2709);
and U3888 (N_3888,N_2453,N_2429);
nor U3889 (N_3889,N_2571,N_2773);
and U3890 (N_3890,N_2506,N_2080);
or U3891 (N_3891,N_2078,N_2862);
or U3892 (N_3892,N_2011,N_2392);
or U3893 (N_3893,N_2258,N_2283);
and U3894 (N_3894,N_2083,N_2960);
nor U3895 (N_3895,N_2414,N_2322);
and U3896 (N_3896,N_2560,N_2880);
and U3897 (N_3897,N_2681,N_2327);
nor U3898 (N_3898,N_2550,N_2288);
and U3899 (N_3899,N_2242,N_2767);
or U3900 (N_3900,N_2704,N_2719);
nor U3901 (N_3901,N_2455,N_2205);
or U3902 (N_3902,N_2464,N_2194);
nand U3903 (N_3903,N_2798,N_2867);
nor U3904 (N_3904,N_2935,N_2283);
and U3905 (N_3905,N_2310,N_2258);
and U3906 (N_3906,N_2169,N_2957);
and U3907 (N_3907,N_2290,N_2089);
nor U3908 (N_3908,N_2983,N_2936);
and U3909 (N_3909,N_2429,N_2451);
or U3910 (N_3910,N_2991,N_2182);
and U3911 (N_3911,N_2992,N_2525);
and U3912 (N_3912,N_2338,N_2773);
and U3913 (N_3913,N_2350,N_2588);
nor U3914 (N_3914,N_2083,N_2922);
nor U3915 (N_3915,N_2942,N_2030);
and U3916 (N_3916,N_2342,N_2500);
nor U3917 (N_3917,N_2532,N_2684);
and U3918 (N_3918,N_2190,N_2576);
nor U3919 (N_3919,N_2354,N_2811);
nor U3920 (N_3920,N_2937,N_2553);
nor U3921 (N_3921,N_2565,N_2288);
and U3922 (N_3922,N_2708,N_2384);
nand U3923 (N_3923,N_2506,N_2868);
nor U3924 (N_3924,N_2696,N_2569);
nand U3925 (N_3925,N_2964,N_2572);
nor U3926 (N_3926,N_2434,N_2513);
and U3927 (N_3927,N_2786,N_2687);
or U3928 (N_3928,N_2032,N_2215);
nor U3929 (N_3929,N_2175,N_2689);
nand U3930 (N_3930,N_2359,N_2229);
or U3931 (N_3931,N_2444,N_2115);
or U3932 (N_3932,N_2167,N_2726);
or U3933 (N_3933,N_2105,N_2971);
or U3934 (N_3934,N_2311,N_2459);
nand U3935 (N_3935,N_2081,N_2355);
nand U3936 (N_3936,N_2086,N_2720);
or U3937 (N_3937,N_2161,N_2153);
and U3938 (N_3938,N_2824,N_2833);
or U3939 (N_3939,N_2167,N_2130);
or U3940 (N_3940,N_2799,N_2746);
or U3941 (N_3941,N_2651,N_2095);
and U3942 (N_3942,N_2327,N_2826);
nand U3943 (N_3943,N_2009,N_2513);
or U3944 (N_3944,N_2571,N_2281);
nor U3945 (N_3945,N_2678,N_2759);
or U3946 (N_3946,N_2979,N_2777);
and U3947 (N_3947,N_2374,N_2670);
nor U3948 (N_3948,N_2296,N_2652);
or U3949 (N_3949,N_2883,N_2874);
and U3950 (N_3950,N_2511,N_2421);
nor U3951 (N_3951,N_2021,N_2723);
nand U3952 (N_3952,N_2573,N_2226);
and U3953 (N_3953,N_2212,N_2789);
nand U3954 (N_3954,N_2008,N_2809);
and U3955 (N_3955,N_2404,N_2825);
nand U3956 (N_3956,N_2950,N_2854);
nand U3957 (N_3957,N_2335,N_2733);
xor U3958 (N_3958,N_2247,N_2770);
nor U3959 (N_3959,N_2422,N_2957);
nor U3960 (N_3960,N_2103,N_2656);
nand U3961 (N_3961,N_2779,N_2185);
nand U3962 (N_3962,N_2577,N_2584);
or U3963 (N_3963,N_2426,N_2765);
or U3964 (N_3964,N_2969,N_2474);
xor U3965 (N_3965,N_2572,N_2142);
nor U3966 (N_3966,N_2475,N_2729);
and U3967 (N_3967,N_2663,N_2971);
nor U3968 (N_3968,N_2635,N_2319);
and U3969 (N_3969,N_2946,N_2304);
nor U3970 (N_3970,N_2652,N_2278);
and U3971 (N_3971,N_2170,N_2127);
nor U3972 (N_3972,N_2529,N_2810);
nand U3973 (N_3973,N_2795,N_2956);
and U3974 (N_3974,N_2244,N_2862);
and U3975 (N_3975,N_2782,N_2745);
or U3976 (N_3976,N_2111,N_2278);
nand U3977 (N_3977,N_2042,N_2934);
nor U3978 (N_3978,N_2244,N_2875);
nand U3979 (N_3979,N_2186,N_2026);
or U3980 (N_3980,N_2693,N_2194);
or U3981 (N_3981,N_2665,N_2986);
nand U3982 (N_3982,N_2106,N_2675);
nor U3983 (N_3983,N_2741,N_2399);
and U3984 (N_3984,N_2713,N_2709);
nor U3985 (N_3985,N_2448,N_2530);
nand U3986 (N_3986,N_2659,N_2777);
or U3987 (N_3987,N_2418,N_2198);
nor U3988 (N_3988,N_2873,N_2137);
or U3989 (N_3989,N_2008,N_2839);
nand U3990 (N_3990,N_2660,N_2112);
or U3991 (N_3991,N_2498,N_2391);
and U3992 (N_3992,N_2151,N_2631);
or U3993 (N_3993,N_2513,N_2857);
nand U3994 (N_3994,N_2553,N_2828);
nor U3995 (N_3995,N_2124,N_2555);
or U3996 (N_3996,N_2319,N_2015);
nor U3997 (N_3997,N_2979,N_2358);
or U3998 (N_3998,N_2594,N_2509);
nand U3999 (N_3999,N_2480,N_2343);
and U4000 (N_4000,N_3944,N_3580);
and U4001 (N_4001,N_3581,N_3904);
nand U4002 (N_4002,N_3279,N_3495);
or U4003 (N_4003,N_3011,N_3171);
nor U4004 (N_4004,N_3801,N_3808);
nor U4005 (N_4005,N_3515,N_3217);
nor U4006 (N_4006,N_3162,N_3697);
nor U4007 (N_4007,N_3490,N_3377);
and U4008 (N_4008,N_3274,N_3401);
nor U4009 (N_4009,N_3565,N_3951);
nand U4010 (N_4010,N_3151,N_3586);
nand U4011 (N_4011,N_3044,N_3080);
and U4012 (N_4012,N_3215,N_3441);
nor U4013 (N_4013,N_3692,N_3295);
nand U4014 (N_4014,N_3887,N_3329);
and U4015 (N_4015,N_3566,N_3110);
and U4016 (N_4016,N_3559,N_3334);
and U4017 (N_4017,N_3804,N_3033);
or U4018 (N_4018,N_3353,N_3280);
nor U4019 (N_4019,N_3270,N_3042);
and U4020 (N_4020,N_3406,N_3731);
and U4021 (N_4021,N_3462,N_3831);
nor U4022 (N_4022,N_3198,N_3165);
nor U4023 (N_4023,N_3619,N_3319);
and U4024 (N_4024,N_3449,N_3035);
or U4025 (N_4025,N_3138,N_3448);
or U4026 (N_4026,N_3857,N_3900);
and U4027 (N_4027,N_3679,N_3119);
nor U4028 (N_4028,N_3598,N_3469);
and U4029 (N_4029,N_3558,N_3840);
or U4030 (N_4030,N_3133,N_3820);
nor U4031 (N_4031,N_3242,N_3592);
nand U4032 (N_4032,N_3127,N_3243);
nand U4033 (N_4033,N_3968,N_3388);
nor U4034 (N_4034,N_3611,N_3267);
nand U4035 (N_4035,N_3288,N_3910);
or U4036 (N_4036,N_3043,N_3491);
and U4037 (N_4037,N_3766,N_3934);
or U4038 (N_4038,N_3958,N_3902);
nand U4039 (N_4039,N_3878,N_3071);
or U4040 (N_4040,N_3427,N_3949);
and U4041 (N_4041,N_3460,N_3023);
nor U4042 (N_4042,N_3529,N_3988);
or U4043 (N_4043,N_3528,N_3301);
and U4044 (N_4044,N_3678,N_3300);
nor U4045 (N_4045,N_3028,N_3153);
or U4046 (N_4046,N_3214,N_3473);
nor U4047 (N_4047,N_3913,N_3053);
or U4048 (N_4048,N_3596,N_3352);
xor U4049 (N_4049,N_3056,N_3336);
nor U4050 (N_4050,N_3889,N_3257);
and U4051 (N_4051,N_3081,N_3255);
or U4052 (N_4052,N_3411,N_3224);
nand U4053 (N_4053,N_3973,N_3942);
and U4054 (N_4054,N_3754,N_3677);
and U4055 (N_4055,N_3239,N_3435);
nand U4056 (N_4056,N_3501,N_3893);
nand U4057 (N_4057,N_3374,N_3982);
and U4058 (N_4058,N_3745,N_3045);
nor U4059 (N_4059,N_3254,N_3649);
or U4060 (N_4060,N_3147,N_3899);
nor U4061 (N_4061,N_3548,N_3380);
or U4062 (N_4062,N_3666,N_3739);
nor U4063 (N_4063,N_3854,N_3720);
nand U4064 (N_4064,N_3476,N_3143);
and U4065 (N_4065,N_3313,N_3376);
and U4066 (N_4066,N_3123,N_3773);
nand U4067 (N_4067,N_3195,N_3231);
or U4068 (N_4068,N_3767,N_3048);
nor U4069 (N_4069,N_3419,N_3432);
nand U4070 (N_4070,N_3519,N_3991);
and U4071 (N_4071,N_3707,N_3833);
nand U4072 (N_4072,N_3895,N_3971);
and U4073 (N_4073,N_3832,N_3729);
and U4074 (N_4074,N_3121,N_3131);
or U4075 (N_4075,N_3703,N_3140);
and U4076 (N_4076,N_3068,N_3571);
and U4077 (N_4077,N_3675,N_3695);
nand U4078 (N_4078,N_3278,N_3488);
or U4079 (N_4079,N_3463,N_3281);
nor U4080 (N_4080,N_3225,N_3472);
nand U4081 (N_4081,N_3095,N_3437);
or U4082 (N_4082,N_3136,N_3498);
nor U4083 (N_4083,N_3796,N_3644);
or U4084 (N_4084,N_3593,N_3293);
and U4085 (N_4085,N_3087,N_3628);
and U4086 (N_4086,N_3404,N_3927);
and U4087 (N_4087,N_3622,N_3892);
and U4088 (N_4088,N_3470,N_3689);
or U4089 (N_4089,N_3260,N_3015);
nor U4090 (N_4090,N_3330,N_3715);
and U4091 (N_4091,N_3637,N_3829);
nand U4092 (N_4092,N_3502,N_3538);
nand U4093 (N_4093,N_3497,N_3828);
and U4094 (N_4094,N_3054,N_3010);
and U4095 (N_4095,N_3757,N_3367);
and U4096 (N_4096,N_3451,N_3640);
nand U4097 (N_4097,N_3183,N_3290);
and U4098 (N_4098,N_3063,N_3345);
nor U4099 (N_4099,N_3768,N_3306);
and U4100 (N_4100,N_3641,N_3111);
and U4101 (N_4101,N_3438,N_3393);
or U4102 (N_4102,N_3713,N_3207);
and U4103 (N_4103,N_3762,N_3935);
nand U4104 (N_4104,N_3024,N_3163);
nor U4105 (N_4105,N_3174,N_3952);
or U4106 (N_4106,N_3977,N_3030);
or U4107 (N_4107,N_3761,N_3685);
and U4108 (N_4108,N_3608,N_3817);
nand U4109 (N_4109,N_3219,N_3702);
or U4110 (N_4110,N_3753,N_3712);
nor U4111 (N_4111,N_3969,N_3776);
and U4112 (N_4112,N_3499,N_3326);
and U4113 (N_4113,N_3803,N_3510);
or U4114 (N_4114,N_3021,N_3132);
or U4115 (N_4115,N_3069,N_3237);
nand U4116 (N_4116,N_3836,N_3057);
and U4117 (N_4117,N_3590,N_3305);
and U4118 (N_4118,N_3047,N_3112);
or U4119 (N_4119,N_3858,N_3425);
nand U4120 (N_4120,N_3218,N_3582);
and U4121 (N_4121,N_3778,N_3576);
and U4122 (N_4122,N_3972,N_3447);
and U4123 (N_4123,N_3009,N_3025);
or U4124 (N_4124,N_3845,N_3418);
and U4125 (N_4125,N_3667,N_3724);
or U4126 (N_4126,N_3603,N_3318);
or U4127 (N_4127,N_3083,N_3959);
and U4128 (N_4128,N_3660,N_3312);
nand U4129 (N_4129,N_3126,N_3698);
nand U4130 (N_4130,N_3152,N_3302);
or U4131 (N_4131,N_3355,N_3478);
and U4132 (N_4132,N_3560,N_3384);
nand U4133 (N_4133,N_3019,N_3671);
nor U4134 (N_4134,N_3458,N_3208);
nand U4135 (N_4135,N_3760,N_3005);
and U4136 (N_4136,N_3524,N_3549);
nor U4137 (N_4137,N_3533,N_3777);
xnor U4138 (N_4138,N_3752,N_3924);
and U4139 (N_4139,N_3849,N_3545);
nand U4140 (N_4140,N_3688,N_3718);
nand U4141 (N_4141,N_3366,N_3125);
and U4142 (N_4142,N_3815,N_3442);
or U4143 (N_4143,N_3813,N_3719);
or U4144 (N_4144,N_3308,N_3706);
nand U4145 (N_4145,N_3950,N_3074);
and U4146 (N_4146,N_3879,N_3122);
and U4147 (N_4147,N_3585,N_3625);
and U4148 (N_4148,N_3908,N_3477);
nand U4149 (N_4149,N_3169,N_3128);
or U4150 (N_4150,N_3109,N_3541);
and U4151 (N_4151,N_3161,N_3452);
nor U4152 (N_4152,N_3787,N_3861);
nor U4153 (N_4153,N_3755,N_3555);
nand U4154 (N_4154,N_3975,N_3534);
and U4155 (N_4155,N_3097,N_3691);
and U4156 (N_4156,N_3405,N_3454);
and U4157 (N_4157,N_3299,N_3134);
or U4158 (N_4158,N_3956,N_3064);
and U4159 (N_4159,N_3396,N_3853);
nor U4160 (N_4160,N_3633,N_3626);
or U4161 (N_4161,N_3962,N_3874);
nand U4162 (N_4162,N_3417,N_3589);
or U4163 (N_4163,N_3526,N_3618);
nand U4164 (N_4164,N_3520,N_3711);
nor U4165 (N_4165,N_3155,N_3430);
nand U4166 (N_4166,N_3184,N_3967);
nor U4167 (N_4167,N_3294,N_3717);
nand U4168 (N_4168,N_3769,N_3226);
nor U4169 (N_4169,N_3725,N_3016);
and U4170 (N_4170,N_3164,N_3827);
nor U4171 (N_4171,N_3487,N_3645);
or U4172 (N_4172,N_3575,N_3550);
or U4173 (N_4173,N_3403,N_3323);
nand U4174 (N_4174,N_3407,N_3118);
or U4175 (N_4175,N_3500,N_3130);
nor U4176 (N_4176,N_3450,N_3765);
nor U4177 (N_4177,N_3894,N_3408);
xnor U4178 (N_4178,N_3573,N_3794);
nand U4179 (N_4179,N_3093,N_3716);
nand U4180 (N_4180,N_3456,N_3834);
nand U4181 (N_4181,N_3875,N_3014);
nor U4182 (N_4182,N_3993,N_3912);
xor U4183 (N_4183,N_3465,N_3751);
or U4184 (N_4184,N_3253,N_3117);
xor U4185 (N_4185,N_3343,N_3012);
nor U4186 (N_4186,N_3189,N_3039);
nand U4187 (N_4187,N_3824,N_3995);
and U4188 (N_4188,N_3263,N_3201);
nor U4189 (N_4189,N_3399,N_3606);
and U4190 (N_4190,N_3346,N_3873);
nand U4191 (N_4191,N_3966,N_3429);
nand U4192 (N_4192,N_3536,N_3202);
nand U4193 (N_4193,N_3819,N_3175);
nor U4194 (N_4194,N_3599,N_3615);
and U4195 (N_4195,N_3997,N_3604);
nor U4196 (N_4196,N_3646,N_3735);
nand U4197 (N_4197,N_3996,N_3461);
nor U4198 (N_4198,N_3483,N_3386);
nor U4199 (N_4199,N_3938,N_3259);
or U4200 (N_4200,N_3075,N_3287);
or U4201 (N_4201,N_3106,N_3372);
nor U4202 (N_4202,N_3786,N_3310);
nand U4203 (N_4203,N_3321,N_3082);
nand U4204 (N_4204,N_3433,N_3286);
nor U4205 (N_4205,N_3236,N_3837);
and U4206 (N_4206,N_3516,N_3459);
nor U4207 (N_4207,N_3770,N_3180);
nand U4208 (N_4208,N_3320,N_3061);
nor U4209 (N_4209,N_3701,N_3464);
and U4210 (N_4210,N_3865,N_3394);
nand U4211 (N_4211,N_3493,N_3998);
and U4212 (N_4212,N_3289,N_3296);
nor U4213 (N_4213,N_3758,N_3839);
and U4214 (N_4214,N_3922,N_3283);
or U4215 (N_4215,N_3105,N_3978);
nor U4216 (N_4216,N_3381,N_3228);
and U4217 (N_4217,N_3869,N_3791);
nand U4218 (N_4218,N_3727,N_3793);
nor U4219 (N_4219,N_3232,N_3291);
xor U4220 (N_4220,N_3414,N_3932);
xnor U4221 (N_4221,N_3365,N_3256);
and U4222 (N_4222,N_3234,N_3521);
and U4223 (N_4223,N_3213,N_3693);
nor U4224 (N_4224,N_3335,N_3850);
and U4225 (N_4225,N_3535,N_3020);
nand U4226 (N_4226,N_3036,N_3398);
or U4227 (N_4227,N_3509,N_3049);
nand U4228 (N_4228,N_3065,N_3588);
xor U4229 (N_4229,N_3665,N_3624);
xor U4230 (N_4230,N_3444,N_3395);
and U4231 (N_4231,N_3282,N_3659);
nand U4232 (N_4232,N_3587,N_3055);
nand U4233 (N_4233,N_3657,N_3480);
nand U4234 (N_4234,N_3870,N_3965);
and U4235 (N_4235,N_3426,N_3652);
nor U4236 (N_4236,N_3371,N_3440);
nor U4237 (N_4237,N_3943,N_3272);
or U4238 (N_4238,N_3514,N_3780);
and U4239 (N_4239,N_3271,N_3347);
nor U4240 (N_4240,N_3732,N_3979);
or U4241 (N_4241,N_3188,N_3656);
nor U4242 (N_4242,N_3101,N_3527);
nand U4243 (N_4243,N_3107,N_3750);
nor U4244 (N_4244,N_3613,N_3268);
nand U4245 (N_4245,N_3494,N_3360);
nor U4246 (N_4246,N_3662,N_3547);
and U4247 (N_4247,N_3882,N_3210);
nor U4248 (N_4248,N_3792,N_3199);
nand U4249 (N_4249,N_3331,N_3930);
or U4250 (N_4250,N_3554,N_3643);
or U4251 (N_4251,N_3981,N_3743);
nand U4252 (N_4252,N_3532,N_3062);
nand U4253 (N_4253,N_3051,N_3116);
or U4254 (N_4254,N_3034,N_3492);
nor U4255 (N_4255,N_3681,N_3031);
nand U4256 (N_4256,N_3091,N_3484);
or U4257 (N_4257,N_3986,N_3976);
or U4258 (N_4258,N_3723,N_3562);
nor U4259 (N_4259,N_3772,N_3142);
nand U4260 (N_4260,N_3314,N_3385);
and U4261 (N_4261,N_3928,N_3358);
xor U4262 (N_4262,N_3249,N_3884);
nand U4263 (N_4263,N_3872,N_3680);
nor U4264 (N_4264,N_3221,N_3961);
nand U4265 (N_4265,N_3058,N_3916);
xnor U4266 (N_4266,N_3173,N_3759);
or U4267 (N_4267,N_3052,N_3368);
and U4268 (N_4268,N_3744,N_3084);
or U4269 (N_4269,N_3160,N_3145);
or U4270 (N_4270,N_3946,N_3471);
or U4271 (N_4271,N_3424,N_3954);
or U4272 (N_4272,N_3333,N_3413);
and U4273 (N_4273,N_3992,N_3223);
or U4274 (N_4274,N_3983,N_3915);
or U4275 (N_4275,N_3307,N_3038);
and U4276 (N_4276,N_3844,N_3327);
and U4277 (N_4277,N_3923,N_3522);
and U4278 (N_4278,N_3356,N_3322);
and U4279 (N_4279,N_3265,N_3919);
nand U4280 (N_4280,N_3542,N_3600);
and U4281 (N_4281,N_3439,N_3809);
or U4282 (N_4282,N_3994,N_3149);
and U4283 (N_4283,N_3668,N_3027);
and U4284 (N_4284,N_3614,N_3505);
nor U4285 (N_4285,N_3632,N_3569);
nor U4286 (N_4286,N_3338,N_3672);
nor U4287 (N_4287,N_3383,N_3673);
nor U4288 (N_4288,N_3621,N_3220);
nand U4289 (N_4289,N_3911,N_3003);
nand U4290 (N_4290,N_3017,N_3830);
or U4291 (N_4291,N_3742,N_3475);
and U4292 (N_4292,N_3709,N_3496);
nor U4293 (N_4293,N_3181,N_3059);
nand U4294 (N_4294,N_3653,N_3141);
or U4295 (N_4295,N_3273,N_3847);
nor U4296 (N_4296,N_3848,N_3191);
nand U4297 (N_4297,N_3937,N_3888);
and U4298 (N_4298,N_3664,N_3342);
nor U4299 (N_4299,N_3185,N_3103);
and U4300 (N_4300,N_3316,N_3802);
and U4301 (N_4301,N_3594,N_3906);
and U4302 (N_4302,N_3203,N_3948);
and U4303 (N_4303,N_3654,N_3568);
nand U4304 (N_4304,N_3194,N_3806);
nand U4305 (N_4305,N_3387,N_3229);
or U4306 (N_4306,N_3325,N_3708);
and U4307 (N_4307,N_3859,N_3192);
and U4308 (N_4308,N_3357,N_3085);
or U4309 (N_4309,N_3567,N_3563);
and U4310 (N_4310,N_3193,N_3157);
nand U4311 (N_4311,N_3073,N_3985);
or U4312 (N_4312,N_3783,N_3482);
and U4313 (N_4313,N_3749,N_3108);
or U4314 (N_4314,N_3907,N_3896);
or U4315 (N_4315,N_3670,N_3690);
and U4316 (N_4316,N_3006,N_3856);
or U4317 (N_4317,N_3209,N_3797);
nor U4318 (N_4318,N_3705,N_3206);
nand U4319 (N_4319,N_3546,N_3078);
nor U4320 (N_4320,N_3196,N_3349);
nor U4321 (N_4321,N_3481,N_3092);
and U4322 (N_4322,N_3066,N_3763);
or U4323 (N_4323,N_3790,N_3304);
nand U4324 (N_4324,N_3001,N_3655);
and U4325 (N_4325,N_3741,N_3574);
and U4326 (N_4326,N_3642,N_3651);
nand U4327 (N_4327,N_3422,N_3317);
nor U4328 (N_4328,N_3072,N_3244);
nor U4329 (N_4329,N_3553,N_3798);
nand U4330 (N_4330,N_3018,N_3026);
or U4331 (N_4331,N_3258,N_3771);
nand U4332 (N_4332,N_3129,N_3747);
nor U4333 (N_4333,N_3379,N_3098);
or U4334 (N_4334,N_3369,N_3262);
or U4335 (N_4335,N_3617,N_3315);
nand U4336 (N_4336,N_3583,N_3512);
nand U4337 (N_4337,N_3647,N_3455);
or U4338 (N_4338,N_3764,N_3612);
or U4339 (N_4339,N_3363,N_3389);
nand U4340 (N_4340,N_3537,N_3235);
nor U4341 (N_4341,N_3150,N_3963);
nand U4342 (N_4342,N_3168,N_3577);
or U4343 (N_4343,N_3543,N_3479);
or U4344 (N_4344,N_3862,N_3000);
and U4345 (N_4345,N_3987,N_3453);
nor U4346 (N_4346,N_3811,N_3443);
and U4347 (N_4347,N_3851,N_3205);
and U4348 (N_4348,N_3860,N_3113);
and U4349 (N_4349,N_3104,N_3400);
and U4350 (N_4350,N_3457,N_3980);
nor U4351 (N_4351,N_3636,N_3261);
and U4352 (N_4352,N_3227,N_3931);
or U4353 (N_4353,N_3816,N_3953);
or U4354 (N_4354,N_3167,N_3503);
nor U4355 (N_4355,N_3552,N_3818);
nand U4356 (N_4356,N_3821,N_3897);
and U4357 (N_4357,N_3517,N_3086);
nor U4358 (N_4358,N_3914,N_3089);
nand U4359 (N_4359,N_3324,N_3686);
nand U4360 (N_4360,N_3863,N_3008);
nand U4361 (N_4361,N_3037,N_3623);
and U4362 (N_4362,N_3868,N_3252);
or U4363 (N_4363,N_3079,N_3876);
or U4364 (N_4364,N_3823,N_3309);
nor U4365 (N_4365,N_3135,N_3661);
nor U4366 (N_4366,N_3341,N_3245);
xor U4367 (N_4367,N_3090,N_3578);
or U4368 (N_4368,N_3362,N_3784);
and U4369 (N_4369,N_3076,N_3197);
or U4370 (N_4370,N_3428,N_3721);
xor U4371 (N_4371,N_3211,N_3781);
or U4372 (N_4372,N_3391,N_3311);
nand U4373 (N_4373,N_3022,N_3124);
nor U4374 (N_4374,N_3826,N_3351);
nand U4375 (N_4375,N_3373,N_3648);
nor U4376 (N_4376,N_3246,N_3240);
and U4377 (N_4377,N_3704,N_3250);
nand U4378 (N_4378,N_3926,N_3556);
or U4379 (N_4379,N_3572,N_3190);
and U4380 (N_4380,N_3468,N_3740);
and U4381 (N_4381,N_3285,N_3957);
or U4382 (N_4382,N_3722,N_3891);
and U4383 (N_4383,N_3340,N_3867);
or U4384 (N_4384,N_3835,N_3222);
and U4385 (N_4385,N_3531,N_3788);
or U4386 (N_4386,N_3939,N_3013);
nand U4387 (N_4387,N_3990,N_3630);
nand U4388 (N_4388,N_3597,N_3842);
and U4389 (N_4389,N_3251,N_3775);
nand U4390 (N_4390,N_3040,N_3810);
or U4391 (N_4391,N_3843,N_3276);
nand U4392 (N_4392,N_3390,N_3694);
nand U4393 (N_4393,N_3375,N_3779);
nand U4394 (N_4394,N_3805,N_3638);
or U4395 (N_4395,N_3485,N_3841);
nand U4396 (N_4396,N_3204,N_3736);
and U4397 (N_4397,N_3789,N_3855);
nand U4398 (N_4398,N_3539,N_3627);
nor U4399 (N_4399,N_3933,N_3852);
and U4400 (N_4400,N_3941,N_3148);
xnor U4401 (N_4401,N_3674,N_3067);
or U4402 (N_4402,N_3917,N_3871);
nand U4403 (N_4403,N_3466,N_3506);
nand U4404 (N_4404,N_3814,N_3004);
nor U4405 (N_4405,N_3088,N_3178);
and U4406 (N_4406,N_3561,N_3467);
nor U4407 (N_4407,N_3909,N_3898);
nand U4408 (N_4408,N_3738,N_3639);
nand U4409 (N_4409,N_3518,N_3050);
nand U4410 (N_4410,N_3007,N_3504);
or U4411 (N_4411,N_3344,N_3328);
nand U4412 (N_4412,N_3507,N_3436);
nand U4413 (N_4413,N_3513,N_3115);
and U4414 (N_4414,N_3540,N_3881);
nor U4415 (N_4415,N_3370,N_3795);
nor U4416 (N_4416,N_3866,N_3298);
nor U4417 (N_4417,N_3339,N_3756);
or U4418 (N_4418,N_3176,N_3846);
or U4419 (N_4419,N_3431,N_3029);
xor U4420 (N_4420,N_3822,N_3486);
nor U4421 (N_4421,N_3423,N_3629);
or U4422 (N_4422,N_3989,N_3557);
and U4423 (N_4423,N_3297,N_3269);
nand U4424 (N_4424,N_3100,N_3392);
and U4425 (N_4425,N_3359,N_3570);
or U4426 (N_4426,N_3825,N_3864);
nand U4427 (N_4427,N_3415,N_3676);
nand U4428 (N_4428,N_3591,N_3489);
xor U4429 (N_4429,N_3730,N_3102);
nand U4430 (N_4430,N_3292,N_3683);
nor U4431 (N_4431,N_3905,N_3446);
nand U4432 (N_4432,N_3060,N_3154);
or U4433 (N_4433,N_3807,N_3146);
nor U4434 (N_4434,N_3970,N_3099);
nor U4435 (N_4435,N_3041,N_3350);
nor U4436 (N_4436,N_3266,N_3920);
nor U4437 (N_4437,N_3434,N_3880);
nand U4438 (N_4438,N_3610,N_3378);
nand U4439 (N_4439,N_3886,N_3710);
nor U4440 (N_4440,N_3523,N_3800);
and U4441 (N_4441,N_3337,N_3734);
nor U4442 (N_4442,N_3579,N_3564);
or U4443 (N_4443,N_3921,N_3658);
nand U4444 (N_4444,N_3120,N_3233);
or U4445 (N_4445,N_3883,N_3412);
nand U4446 (N_4446,N_3544,N_3631);
or U4447 (N_4447,N_3364,N_3669);
nand U4448 (N_4448,N_3277,N_3156);
nor U4449 (N_4449,N_3663,N_3696);
or U4450 (N_4450,N_3602,N_3177);
or U4451 (N_4451,N_3172,N_3416);
or U4452 (N_4452,N_3774,N_3737);
or U4453 (N_4453,N_3179,N_3947);
nor U4454 (N_4454,N_3885,N_3508);
and U4455 (N_4455,N_3170,N_3940);
and U4456 (N_4456,N_3607,N_3890);
nand U4457 (N_4457,N_3182,N_3595);
nor U4458 (N_4458,N_3726,N_3159);
nor U4459 (N_4459,N_3901,N_3748);
nor U4460 (N_4460,N_3918,N_3421);
nand U4461 (N_4461,N_3166,N_3158);
and U4462 (N_4462,N_3955,N_3332);
or U4463 (N_4463,N_3096,N_3782);
xor U4464 (N_4464,N_3746,N_3699);
nor U4465 (N_4465,N_3728,N_3984);
nor U4466 (N_4466,N_3397,N_3284);
and U4467 (N_4467,N_3999,N_3903);
nand U4468 (N_4468,N_3812,N_3046);
and U4469 (N_4469,N_3929,N_3248);
xnor U4470 (N_4470,N_3354,N_3303);
or U4471 (N_4471,N_3094,N_3650);
or U4472 (N_4472,N_3238,N_3936);
or U4473 (N_4473,N_3114,N_3525);
nor U4474 (N_4474,N_3925,N_3002);
nand U4475 (N_4475,N_3687,N_3200);
nand U4476 (N_4476,N_3799,N_3620);
nor U4477 (N_4477,N_3964,N_3077);
nand U4478 (N_4478,N_3635,N_3960);
and U4479 (N_4479,N_3684,N_3609);
and U4480 (N_4480,N_3616,N_3700);
or U4481 (N_4481,N_3144,N_3186);
or U4482 (N_4482,N_3601,N_3838);
nor U4483 (N_4483,N_3445,N_3137);
nor U4484 (N_4484,N_3584,N_3634);
or U4485 (N_4485,N_3247,N_3070);
nand U4486 (N_4486,N_3409,N_3511);
and U4487 (N_4487,N_3974,N_3785);
nor U4488 (N_4488,N_3945,N_3474);
nor U4489 (N_4489,N_3241,N_3733);
or U4490 (N_4490,N_3382,N_3187);
or U4491 (N_4491,N_3420,N_3264);
nor U4492 (N_4492,N_3139,N_3410);
nor U4493 (N_4493,N_3530,N_3032);
nor U4494 (N_4494,N_3212,N_3682);
nor U4495 (N_4495,N_3551,N_3348);
or U4496 (N_4496,N_3714,N_3877);
nor U4497 (N_4497,N_3361,N_3402);
nor U4498 (N_4498,N_3216,N_3605);
or U4499 (N_4499,N_3230,N_3275);
or U4500 (N_4500,N_3539,N_3725);
or U4501 (N_4501,N_3503,N_3931);
nand U4502 (N_4502,N_3761,N_3416);
nand U4503 (N_4503,N_3165,N_3268);
nand U4504 (N_4504,N_3332,N_3705);
nor U4505 (N_4505,N_3338,N_3215);
and U4506 (N_4506,N_3505,N_3283);
or U4507 (N_4507,N_3185,N_3622);
or U4508 (N_4508,N_3889,N_3210);
nand U4509 (N_4509,N_3490,N_3874);
or U4510 (N_4510,N_3697,N_3597);
nor U4511 (N_4511,N_3735,N_3849);
nor U4512 (N_4512,N_3547,N_3524);
nand U4513 (N_4513,N_3463,N_3346);
xor U4514 (N_4514,N_3466,N_3887);
nand U4515 (N_4515,N_3418,N_3642);
or U4516 (N_4516,N_3784,N_3408);
nor U4517 (N_4517,N_3622,N_3058);
nor U4518 (N_4518,N_3055,N_3385);
nand U4519 (N_4519,N_3026,N_3520);
and U4520 (N_4520,N_3499,N_3026);
or U4521 (N_4521,N_3869,N_3247);
nor U4522 (N_4522,N_3162,N_3733);
and U4523 (N_4523,N_3200,N_3294);
or U4524 (N_4524,N_3213,N_3168);
or U4525 (N_4525,N_3900,N_3148);
or U4526 (N_4526,N_3649,N_3476);
nand U4527 (N_4527,N_3069,N_3301);
nand U4528 (N_4528,N_3564,N_3219);
xor U4529 (N_4529,N_3835,N_3568);
and U4530 (N_4530,N_3483,N_3879);
nand U4531 (N_4531,N_3927,N_3857);
nor U4532 (N_4532,N_3096,N_3304);
nor U4533 (N_4533,N_3280,N_3990);
nor U4534 (N_4534,N_3139,N_3869);
nor U4535 (N_4535,N_3447,N_3384);
or U4536 (N_4536,N_3253,N_3755);
xnor U4537 (N_4537,N_3865,N_3993);
or U4538 (N_4538,N_3098,N_3369);
and U4539 (N_4539,N_3515,N_3617);
and U4540 (N_4540,N_3833,N_3339);
nor U4541 (N_4541,N_3864,N_3804);
nand U4542 (N_4542,N_3053,N_3984);
nor U4543 (N_4543,N_3394,N_3748);
or U4544 (N_4544,N_3490,N_3281);
nor U4545 (N_4545,N_3539,N_3857);
and U4546 (N_4546,N_3489,N_3231);
or U4547 (N_4547,N_3022,N_3641);
and U4548 (N_4548,N_3865,N_3150);
and U4549 (N_4549,N_3270,N_3332);
nand U4550 (N_4550,N_3591,N_3769);
xnor U4551 (N_4551,N_3096,N_3764);
and U4552 (N_4552,N_3859,N_3457);
nand U4553 (N_4553,N_3110,N_3950);
nand U4554 (N_4554,N_3632,N_3030);
nor U4555 (N_4555,N_3220,N_3120);
or U4556 (N_4556,N_3691,N_3914);
nand U4557 (N_4557,N_3516,N_3790);
nor U4558 (N_4558,N_3527,N_3260);
and U4559 (N_4559,N_3874,N_3997);
nand U4560 (N_4560,N_3862,N_3649);
or U4561 (N_4561,N_3204,N_3624);
nand U4562 (N_4562,N_3144,N_3061);
or U4563 (N_4563,N_3222,N_3706);
nor U4564 (N_4564,N_3177,N_3762);
nor U4565 (N_4565,N_3917,N_3313);
or U4566 (N_4566,N_3675,N_3864);
or U4567 (N_4567,N_3929,N_3340);
or U4568 (N_4568,N_3266,N_3238);
and U4569 (N_4569,N_3284,N_3079);
or U4570 (N_4570,N_3694,N_3065);
nor U4571 (N_4571,N_3333,N_3568);
nand U4572 (N_4572,N_3027,N_3003);
or U4573 (N_4573,N_3166,N_3391);
or U4574 (N_4574,N_3256,N_3631);
nand U4575 (N_4575,N_3240,N_3477);
nor U4576 (N_4576,N_3790,N_3882);
and U4577 (N_4577,N_3863,N_3746);
nand U4578 (N_4578,N_3790,N_3892);
and U4579 (N_4579,N_3561,N_3503);
nand U4580 (N_4580,N_3893,N_3626);
or U4581 (N_4581,N_3880,N_3252);
and U4582 (N_4582,N_3258,N_3475);
and U4583 (N_4583,N_3619,N_3818);
xnor U4584 (N_4584,N_3846,N_3485);
or U4585 (N_4585,N_3628,N_3381);
nor U4586 (N_4586,N_3292,N_3817);
or U4587 (N_4587,N_3283,N_3634);
nand U4588 (N_4588,N_3417,N_3210);
nor U4589 (N_4589,N_3085,N_3979);
nand U4590 (N_4590,N_3744,N_3530);
nor U4591 (N_4591,N_3130,N_3568);
nand U4592 (N_4592,N_3880,N_3329);
nor U4593 (N_4593,N_3746,N_3382);
or U4594 (N_4594,N_3291,N_3725);
or U4595 (N_4595,N_3984,N_3454);
or U4596 (N_4596,N_3908,N_3957);
nand U4597 (N_4597,N_3769,N_3636);
and U4598 (N_4598,N_3394,N_3837);
nor U4599 (N_4599,N_3814,N_3879);
and U4600 (N_4600,N_3620,N_3270);
and U4601 (N_4601,N_3855,N_3841);
xnor U4602 (N_4602,N_3925,N_3888);
and U4603 (N_4603,N_3221,N_3126);
and U4604 (N_4604,N_3195,N_3907);
or U4605 (N_4605,N_3146,N_3067);
and U4606 (N_4606,N_3902,N_3199);
nor U4607 (N_4607,N_3815,N_3437);
nand U4608 (N_4608,N_3622,N_3554);
nand U4609 (N_4609,N_3070,N_3534);
or U4610 (N_4610,N_3702,N_3072);
and U4611 (N_4611,N_3889,N_3556);
nand U4612 (N_4612,N_3043,N_3344);
nand U4613 (N_4613,N_3794,N_3125);
nor U4614 (N_4614,N_3172,N_3165);
or U4615 (N_4615,N_3043,N_3157);
nor U4616 (N_4616,N_3895,N_3399);
or U4617 (N_4617,N_3538,N_3752);
and U4618 (N_4618,N_3790,N_3509);
nand U4619 (N_4619,N_3962,N_3787);
nor U4620 (N_4620,N_3112,N_3073);
or U4621 (N_4621,N_3200,N_3520);
nor U4622 (N_4622,N_3251,N_3707);
and U4623 (N_4623,N_3304,N_3464);
nand U4624 (N_4624,N_3504,N_3063);
nand U4625 (N_4625,N_3680,N_3975);
nand U4626 (N_4626,N_3484,N_3624);
nor U4627 (N_4627,N_3842,N_3592);
nor U4628 (N_4628,N_3112,N_3736);
or U4629 (N_4629,N_3382,N_3909);
nand U4630 (N_4630,N_3081,N_3507);
or U4631 (N_4631,N_3865,N_3035);
nand U4632 (N_4632,N_3813,N_3455);
nand U4633 (N_4633,N_3278,N_3463);
and U4634 (N_4634,N_3101,N_3981);
nand U4635 (N_4635,N_3418,N_3086);
nor U4636 (N_4636,N_3686,N_3960);
or U4637 (N_4637,N_3535,N_3012);
nor U4638 (N_4638,N_3258,N_3807);
or U4639 (N_4639,N_3249,N_3905);
nand U4640 (N_4640,N_3081,N_3923);
nand U4641 (N_4641,N_3591,N_3881);
nor U4642 (N_4642,N_3445,N_3716);
or U4643 (N_4643,N_3886,N_3364);
nor U4644 (N_4644,N_3998,N_3045);
or U4645 (N_4645,N_3791,N_3631);
and U4646 (N_4646,N_3621,N_3739);
nor U4647 (N_4647,N_3071,N_3029);
nor U4648 (N_4648,N_3407,N_3402);
and U4649 (N_4649,N_3295,N_3161);
nor U4650 (N_4650,N_3313,N_3907);
and U4651 (N_4651,N_3490,N_3388);
and U4652 (N_4652,N_3350,N_3971);
nand U4653 (N_4653,N_3364,N_3209);
xnor U4654 (N_4654,N_3048,N_3455);
nand U4655 (N_4655,N_3891,N_3159);
nand U4656 (N_4656,N_3541,N_3283);
nor U4657 (N_4657,N_3343,N_3280);
and U4658 (N_4658,N_3829,N_3542);
nand U4659 (N_4659,N_3604,N_3920);
and U4660 (N_4660,N_3294,N_3290);
nor U4661 (N_4661,N_3651,N_3585);
or U4662 (N_4662,N_3324,N_3845);
or U4663 (N_4663,N_3281,N_3341);
and U4664 (N_4664,N_3874,N_3272);
nor U4665 (N_4665,N_3253,N_3500);
nor U4666 (N_4666,N_3884,N_3287);
and U4667 (N_4667,N_3292,N_3045);
nor U4668 (N_4668,N_3631,N_3520);
or U4669 (N_4669,N_3985,N_3460);
nor U4670 (N_4670,N_3542,N_3559);
or U4671 (N_4671,N_3989,N_3826);
and U4672 (N_4672,N_3452,N_3927);
and U4673 (N_4673,N_3219,N_3307);
and U4674 (N_4674,N_3891,N_3768);
nor U4675 (N_4675,N_3789,N_3092);
xor U4676 (N_4676,N_3958,N_3500);
nor U4677 (N_4677,N_3688,N_3236);
or U4678 (N_4678,N_3057,N_3450);
and U4679 (N_4679,N_3441,N_3179);
and U4680 (N_4680,N_3742,N_3277);
nor U4681 (N_4681,N_3083,N_3806);
and U4682 (N_4682,N_3881,N_3224);
and U4683 (N_4683,N_3178,N_3968);
and U4684 (N_4684,N_3638,N_3795);
and U4685 (N_4685,N_3831,N_3056);
and U4686 (N_4686,N_3072,N_3369);
nor U4687 (N_4687,N_3539,N_3433);
xor U4688 (N_4688,N_3111,N_3099);
or U4689 (N_4689,N_3595,N_3618);
nor U4690 (N_4690,N_3778,N_3188);
xnor U4691 (N_4691,N_3609,N_3740);
nor U4692 (N_4692,N_3296,N_3993);
or U4693 (N_4693,N_3167,N_3348);
and U4694 (N_4694,N_3724,N_3043);
and U4695 (N_4695,N_3227,N_3314);
nand U4696 (N_4696,N_3344,N_3069);
nand U4697 (N_4697,N_3421,N_3209);
and U4698 (N_4698,N_3395,N_3634);
nand U4699 (N_4699,N_3045,N_3090);
or U4700 (N_4700,N_3001,N_3988);
or U4701 (N_4701,N_3953,N_3118);
nand U4702 (N_4702,N_3887,N_3809);
and U4703 (N_4703,N_3414,N_3135);
nor U4704 (N_4704,N_3408,N_3656);
nor U4705 (N_4705,N_3654,N_3586);
or U4706 (N_4706,N_3809,N_3830);
nand U4707 (N_4707,N_3885,N_3121);
nand U4708 (N_4708,N_3443,N_3057);
nand U4709 (N_4709,N_3325,N_3962);
and U4710 (N_4710,N_3149,N_3620);
or U4711 (N_4711,N_3613,N_3381);
nor U4712 (N_4712,N_3779,N_3886);
or U4713 (N_4713,N_3571,N_3654);
nand U4714 (N_4714,N_3779,N_3506);
nor U4715 (N_4715,N_3251,N_3439);
and U4716 (N_4716,N_3223,N_3855);
nand U4717 (N_4717,N_3862,N_3285);
nand U4718 (N_4718,N_3001,N_3486);
nor U4719 (N_4719,N_3695,N_3863);
or U4720 (N_4720,N_3257,N_3007);
nor U4721 (N_4721,N_3152,N_3937);
and U4722 (N_4722,N_3609,N_3314);
nor U4723 (N_4723,N_3784,N_3190);
and U4724 (N_4724,N_3139,N_3975);
and U4725 (N_4725,N_3373,N_3857);
and U4726 (N_4726,N_3689,N_3463);
nor U4727 (N_4727,N_3952,N_3835);
and U4728 (N_4728,N_3291,N_3734);
and U4729 (N_4729,N_3752,N_3941);
xor U4730 (N_4730,N_3103,N_3879);
nor U4731 (N_4731,N_3993,N_3335);
or U4732 (N_4732,N_3295,N_3215);
and U4733 (N_4733,N_3189,N_3962);
nor U4734 (N_4734,N_3056,N_3885);
and U4735 (N_4735,N_3908,N_3744);
nor U4736 (N_4736,N_3066,N_3809);
and U4737 (N_4737,N_3151,N_3324);
or U4738 (N_4738,N_3167,N_3408);
nor U4739 (N_4739,N_3198,N_3510);
nand U4740 (N_4740,N_3107,N_3117);
nor U4741 (N_4741,N_3047,N_3063);
or U4742 (N_4742,N_3155,N_3903);
or U4743 (N_4743,N_3219,N_3587);
or U4744 (N_4744,N_3770,N_3397);
or U4745 (N_4745,N_3731,N_3509);
or U4746 (N_4746,N_3153,N_3295);
nand U4747 (N_4747,N_3374,N_3931);
nor U4748 (N_4748,N_3302,N_3335);
nor U4749 (N_4749,N_3098,N_3399);
or U4750 (N_4750,N_3347,N_3232);
or U4751 (N_4751,N_3440,N_3840);
or U4752 (N_4752,N_3619,N_3019);
nor U4753 (N_4753,N_3930,N_3443);
nand U4754 (N_4754,N_3042,N_3079);
nor U4755 (N_4755,N_3880,N_3962);
nand U4756 (N_4756,N_3806,N_3784);
and U4757 (N_4757,N_3296,N_3548);
nor U4758 (N_4758,N_3871,N_3890);
nor U4759 (N_4759,N_3438,N_3789);
nand U4760 (N_4760,N_3913,N_3081);
nor U4761 (N_4761,N_3551,N_3460);
and U4762 (N_4762,N_3118,N_3894);
or U4763 (N_4763,N_3758,N_3980);
or U4764 (N_4764,N_3077,N_3867);
or U4765 (N_4765,N_3033,N_3670);
or U4766 (N_4766,N_3376,N_3096);
or U4767 (N_4767,N_3926,N_3320);
nor U4768 (N_4768,N_3971,N_3006);
or U4769 (N_4769,N_3366,N_3759);
nand U4770 (N_4770,N_3640,N_3159);
nand U4771 (N_4771,N_3440,N_3909);
nor U4772 (N_4772,N_3205,N_3181);
nand U4773 (N_4773,N_3295,N_3847);
nor U4774 (N_4774,N_3559,N_3741);
nand U4775 (N_4775,N_3242,N_3611);
and U4776 (N_4776,N_3105,N_3565);
nand U4777 (N_4777,N_3808,N_3476);
and U4778 (N_4778,N_3288,N_3689);
nand U4779 (N_4779,N_3933,N_3250);
or U4780 (N_4780,N_3664,N_3086);
or U4781 (N_4781,N_3889,N_3141);
and U4782 (N_4782,N_3864,N_3624);
nor U4783 (N_4783,N_3836,N_3222);
and U4784 (N_4784,N_3226,N_3807);
nand U4785 (N_4785,N_3211,N_3308);
nor U4786 (N_4786,N_3351,N_3719);
nor U4787 (N_4787,N_3540,N_3031);
or U4788 (N_4788,N_3206,N_3589);
nand U4789 (N_4789,N_3552,N_3415);
or U4790 (N_4790,N_3662,N_3302);
nand U4791 (N_4791,N_3628,N_3241);
nand U4792 (N_4792,N_3335,N_3715);
nand U4793 (N_4793,N_3983,N_3953);
nand U4794 (N_4794,N_3403,N_3805);
nor U4795 (N_4795,N_3557,N_3890);
and U4796 (N_4796,N_3077,N_3287);
nor U4797 (N_4797,N_3232,N_3975);
and U4798 (N_4798,N_3582,N_3321);
nor U4799 (N_4799,N_3883,N_3661);
nand U4800 (N_4800,N_3806,N_3329);
and U4801 (N_4801,N_3096,N_3552);
nand U4802 (N_4802,N_3112,N_3794);
or U4803 (N_4803,N_3530,N_3226);
and U4804 (N_4804,N_3095,N_3950);
nand U4805 (N_4805,N_3169,N_3393);
nand U4806 (N_4806,N_3951,N_3896);
nand U4807 (N_4807,N_3072,N_3564);
and U4808 (N_4808,N_3510,N_3391);
nor U4809 (N_4809,N_3281,N_3259);
and U4810 (N_4810,N_3990,N_3298);
nand U4811 (N_4811,N_3715,N_3044);
nand U4812 (N_4812,N_3748,N_3745);
nand U4813 (N_4813,N_3284,N_3825);
nand U4814 (N_4814,N_3686,N_3025);
or U4815 (N_4815,N_3593,N_3360);
nor U4816 (N_4816,N_3471,N_3435);
or U4817 (N_4817,N_3932,N_3227);
nand U4818 (N_4818,N_3264,N_3758);
nand U4819 (N_4819,N_3648,N_3233);
or U4820 (N_4820,N_3481,N_3455);
or U4821 (N_4821,N_3543,N_3131);
and U4822 (N_4822,N_3469,N_3060);
or U4823 (N_4823,N_3877,N_3624);
and U4824 (N_4824,N_3315,N_3037);
and U4825 (N_4825,N_3109,N_3962);
nor U4826 (N_4826,N_3098,N_3312);
nand U4827 (N_4827,N_3727,N_3439);
and U4828 (N_4828,N_3662,N_3812);
or U4829 (N_4829,N_3308,N_3881);
and U4830 (N_4830,N_3500,N_3991);
or U4831 (N_4831,N_3883,N_3660);
or U4832 (N_4832,N_3769,N_3929);
nor U4833 (N_4833,N_3864,N_3235);
nor U4834 (N_4834,N_3191,N_3416);
and U4835 (N_4835,N_3252,N_3711);
and U4836 (N_4836,N_3663,N_3351);
and U4837 (N_4837,N_3000,N_3145);
or U4838 (N_4838,N_3737,N_3015);
nand U4839 (N_4839,N_3742,N_3405);
xor U4840 (N_4840,N_3703,N_3688);
and U4841 (N_4841,N_3909,N_3872);
nor U4842 (N_4842,N_3144,N_3234);
and U4843 (N_4843,N_3079,N_3880);
and U4844 (N_4844,N_3017,N_3272);
nor U4845 (N_4845,N_3508,N_3932);
or U4846 (N_4846,N_3159,N_3393);
nor U4847 (N_4847,N_3103,N_3262);
and U4848 (N_4848,N_3372,N_3904);
or U4849 (N_4849,N_3135,N_3977);
and U4850 (N_4850,N_3463,N_3644);
or U4851 (N_4851,N_3704,N_3963);
or U4852 (N_4852,N_3623,N_3327);
nor U4853 (N_4853,N_3955,N_3005);
or U4854 (N_4854,N_3927,N_3905);
nand U4855 (N_4855,N_3601,N_3777);
and U4856 (N_4856,N_3711,N_3981);
and U4857 (N_4857,N_3030,N_3870);
nor U4858 (N_4858,N_3311,N_3025);
nand U4859 (N_4859,N_3687,N_3287);
and U4860 (N_4860,N_3433,N_3467);
and U4861 (N_4861,N_3655,N_3232);
or U4862 (N_4862,N_3024,N_3203);
or U4863 (N_4863,N_3312,N_3492);
nand U4864 (N_4864,N_3504,N_3520);
nand U4865 (N_4865,N_3869,N_3937);
nor U4866 (N_4866,N_3720,N_3941);
and U4867 (N_4867,N_3662,N_3612);
and U4868 (N_4868,N_3639,N_3842);
nand U4869 (N_4869,N_3452,N_3898);
and U4870 (N_4870,N_3583,N_3595);
nand U4871 (N_4871,N_3631,N_3704);
nand U4872 (N_4872,N_3998,N_3599);
nor U4873 (N_4873,N_3508,N_3386);
nor U4874 (N_4874,N_3228,N_3732);
or U4875 (N_4875,N_3145,N_3095);
nand U4876 (N_4876,N_3808,N_3625);
nor U4877 (N_4877,N_3837,N_3616);
nand U4878 (N_4878,N_3586,N_3159);
and U4879 (N_4879,N_3060,N_3840);
and U4880 (N_4880,N_3981,N_3905);
nand U4881 (N_4881,N_3322,N_3022);
xnor U4882 (N_4882,N_3787,N_3869);
nand U4883 (N_4883,N_3322,N_3348);
nor U4884 (N_4884,N_3377,N_3529);
nand U4885 (N_4885,N_3634,N_3313);
nor U4886 (N_4886,N_3317,N_3917);
nor U4887 (N_4887,N_3328,N_3213);
or U4888 (N_4888,N_3168,N_3617);
nand U4889 (N_4889,N_3921,N_3478);
and U4890 (N_4890,N_3006,N_3703);
nor U4891 (N_4891,N_3596,N_3016);
nand U4892 (N_4892,N_3266,N_3371);
nand U4893 (N_4893,N_3616,N_3771);
and U4894 (N_4894,N_3603,N_3927);
nor U4895 (N_4895,N_3961,N_3959);
nand U4896 (N_4896,N_3585,N_3574);
or U4897 (N_4897,N_3235,N_3743);
nor U4898 (N_4898,N_3471,N_3532);
or U4899 (N_4899,N_3240,N_3173);
or U4900 (N_4900,N_3824,N_3315);
or U4901 (N_4901,N_3144,N_3790);
nand U4902 (N_4902,N_3134,N_3214);
nor U4903 (N_4903,N_3638,N_3959);
or U4904 (N_4904,N_3220,N_3664);
and U4905 (N_4905,N_3426,N_3140);
and U4906 (N_4906,N_3809,N_3063);
nor U4907 (N_4907,N_3840,N_3548);
and U4908 (N_4908,N_3153,N_3224);
or U4909 (N_4909,N_3918,N_3908);
and U4910 (N_4910,N_3856,N_3944);
nor U4911 (N_4911,N_3622,N_3907);
or U4912 (N_4912,N_3145,N_3884);
nand U4913 (N_4913,N_3326,N_3769);
or U4914 (N_4914,N_3359,N_3914);
and U4915 (N_4915,N_3173,N_3465);
nand U4916 (N_4916,N_3532,N_3952);
nand U4917 (N_4917,N_3238,N_3696);
nand U4918 (N_4918,N_3245,N_3908);
and U4919 (N_4919,N_3631,N_3963);
nand U4920 (N_4920,N_3369,N_3855);
nand U4921 (N_4921,N_3460,N_3041);
and U4922 (N_4922,N_3269,N_3408);
nor U4923 (N_4923,N_3309,N_3630);
or U4924 (N_4924,N_3045,N_3423);
nor U4925 (N_4925,N_3975,N_3074);
nor U4926 (N_4926,N_3179,N_3910);
nand U4927 (N_4927,N_3342,N_3148);
nand U4928 (N_4928,N_3741,N_3696);
nor U4929 (N_4929,N_3722,N_3946);
nand U4930 (N_4930,N_3241,N_3678);
nor U4931 (N_4931,N_3728,N_3395);
nor U4932 (N_4932,N_3844,N_3473);
nor U4933 (N_4933,N_3067,N_3054);
or U4934 (N_4934,N_3531,N_3725);
or U4935 (N_4935,N_3789,N_3477);
nand U4936 (N_4936,N_3173,N_3075);
nor U4937 (N_4937,N_3565,N_3506);
nor U4938 (N_4938,N_3030,N_3825);
nand U4939 (N_4939,N_3131,N_3975);
or U4940 (N_4940,N_3771,N_3106);
nand U4941 (N_4941,N_3914,N_3271);
or U4942 (N_4942,N_3927,N_3041);
nand U4943 (N_4943,N_3905,N_3217);
or U4944 (N_4944,N_3495,N_3379);
or U4945 (N_4945,N_3787,N_3515);
nor U4946 (N_4946,N_3901,N_3381);
nand U4947 (N_4947,N_3894,N_3836);
nand U4948 (N_4948,N_3975,N_3507);
nor U4949 (N_4949,N_3428,N_3246);
nand U4950 (N_4950,N_3524,N_3470);
nor U4951 (N_4951,N_3305,N_3010);
and U4952 (N_4952,N_3071,N_3942);
or U4953 (N_4953,N_3294,N_3848);
and U4954 (N_4954,N_3555,N_3735);
nand U4955 (N_4955,N_3486,N_3053);
or U4956 (N_4956,N_3763,N_3072);
and U4957 (N_4957,N_3835,N_3153);
or U4958 (N_4958,N_3400,N_3990);
nor U4959 (N_4959,N_3199,N_3499);
nor U4960 (N_4960,N_3724,N_3242);
or U4961 (N_4961,N_3723,N_3786);
and U4962 (N_4962,N_3167,N_3122);
or U4963 (N_4963,N_3024,N_3016);
nand U4964 (N_4964,N_3906,N_3850);
xnor U4965 (N_4965,N_3283,N_3338);
xnor U4966 (N_4966,N_3745,N_3881);
nor U4967 (N_4967,N_3841,N_3643);
nand U4968 (N_4968,N_3904,N_3689);
nand U4969 (N_4969,N_3075,N_3370);
xnor U4970 (N_4970,N_3848,N_3355);
or U4971 (N_4971,N_3382,N_3498);
or U4972 (N_4972,N_3000,N_3261);
and U4973 (N_4973,N_3237,N_3574);
or U4974 (N_4974,N_3057,N_3193);
nor U4975 (N_4975,N_3539,N_3531);
nand U4976 (N_4976,N_3452,N_3925);
xnor U4977 (N_4977,N_3822,N_3786);
nor U4978 (N_4978,N_3231,N_3862);
nor U4979 (N_4979,N_3708,N_3913);
nand U4980 (N_4980,N_3233,N_3403);
and U4981 (N_4981,N_3784,N_3849);
nand U4982 (N_4982,N_3194,N_3226);
nand U4983 (N_4983,N_3376,N_3493);
nand U4984 (N_4984,N_3867,N_3838);
and U4985 (N_4985,N_3924,N_3009);
xor U4986 (N_4986,N_3222,N_3293);
nor U4987 (N_4987,N_3351,N_3191);
or U4988 (N_4988,N_3515,N_3050);
nor U4989 (N_4989,N_3651,N_3031);
and U4990 (N_4990,N_3513,N_3587);
nand U4991 (N_4991,N_3535,N_3710);
or U4992 (N_4992,N_3614,N_3270);
or U4993 (N_4993,N_3172,N_3226);
and U4994 (N_4994,N_3673,N_3217);
nand U4995 (N_4995,N_3423,N_3214);
or U4996 (N_4996,N_3545,N_3734);
nand U4997 (N_4997,N_3546,N_3055);
or U4998 (N_4998,N_3185,N_3059);
nand U4999 (N_4999,N_3291,N_3700);
nand U5000 (N_5000,N_4236,N_4669);
or U5001 (N_5001,N_4361,N_4511);
or U5002 (N_5002,N_4542,N_4420);
nor U5003 (N_5003,N_4196,N_4890);
nand U5004 (N_5004,N_4691,N_4775);
and U5005 (N_5005,N_4421,N_4166);
nand U5006 (N_5006,N_4144,N_4168);
nor U5007 (N_5007,N_4972,N_4872);
nor U5008 (N_5008,N_4475,N_4367);
nand U5009 (N_5009,N_4540,N_4637);
or U5010 (N_5010,N_4129,N_4635);
nor U5011 (N_5011,N_4779,N_4650);
or U5012 (N_5012,N_4114,N_4215);
or U5013 (N_5013,N_4656,N_4892);
nor U5014 (N_5014,N_4014,N_4247);
and U5015 (N_5015,N_4823,N_4921);
and U5016 (N_5016,N_4906,N_4132);
nor U5017 (N_5017,N_4104,N_4251);
nand U5018 (N_5018,N_4235,N_4182);
nor U5019 (N_5019,N_4122,N_4573);
and U5020 (N_5020,N_4894,N_4191);
and U5021 (N_5021,N_4507,N_4744);
and U5022 (N_5022,N_4581,N_4075);
nor U5023 (N_5023,N_4792,N_4926);
and U5024 (N_5024,N_4451,N_4042);
or U5025 (N_5025,N_4924,N_4037);
or U5026 (N_5026,N_4081,N_4268);
nor U5027 (N_5027,N_4636,N_4722);
nor U5028 (N_5028,N_4445,N_4315);
nand U5029 (N_5029,N_4529,N_4790);
xnor U5030 (N_5030,N_4167,N_4534);
or U5031 (N_5031,N_4801,N_4040);
or U5032 (N_5032,N_4738,N_4219);
or U5033 (N_5033,N_4305,N_4718);
and U5034 (N_5034,N_4474,N_4039);
or U5035 (N_5035,N_4883,N_4611);
xor U5036 (N_5036,N_4527,N_4918);
nand U5037 (N_5037,N_4772,N_4446);
or U5038 (N_5038,N_4108,N_4661);
and U5039 (N_5039,N_4958,N_4754);
and U5040 (N_5040,N_4087,N_4130);
or U5041 (N_5041,N_4632,N_4804);
and U5042 (N_5042,N_4616,N_4332);
or U5043 (N_5043,N_4406,N_4165);
and U5044 (N_5044,N_4214,N_4536);
nand U5045 (N_5045,N_4175,N_4047);
and U5046 (N_5046,N_4648,N_4645);
xor U5047 (N_5047,N_4362,N_4677);
nor U5048 (N_5048,N_4568,N_4461);
and U5049 (N_5049,N_4008,N_4671);
nand U5050 (N_5050,N_4503,N_4580);
and U5051 (N_5051,N_4389,N_4567);
and U5052 (N_5052,N_4909,N_4286);
nand U5053 (N_5053,N_4350,N_4470);
and U5054 (N_5054,N_4942,N_4410);
and U5055 (N_5055,N_4030,N_4387);
nand U5056 (N_5056,N_4417,N_4543);
and U5057 (N_5057,N_4293,N_4907);
nor U5058 (N_5058,N_4370,N_4755);
and U5059 (N_5059,N_4485,N_4549);
nand U5060 (N_5060,N_4774,N_4939);
and U5061 (N_5061,N_4223,N_4875);
or U5062 (N_5062,N_4452,N_4569);
and U5063 (N_5063,N_4244,N_4433);
nand U5064 (N_5064,N_4643,N_4579);
or U5065 (N_5065,N_4237,N_4811);
nand U5066 (N_5066,N_4148,N_4245);
nor U5067 (N_5067,N_4859,N_4145);
and U5068 (N_5068,N_4173,N_4592);
nor U5069 (N_5069,N_4630,N_4816);
and U5070 (N_5070,N_4262,N_4937);
and U5071 (N_5071,N_4491,N_4654);
nor U5072 (N_5072,N_4267,N_4437);
or U5073 (N_5073,N_4283,N_4711);
nor U5074 (N_5074,N_4947,N_4732);
or U5075 (N_5075,N_4572,N_4723);
nand U5076 (N_5076,N_4506,N_4831);
or U5077 (N_5077,N_4970,N_4399);
nor U5078 (N_5078,N_4988,N_4094);
nor U5079 (N_5079,N_4646,N_4441);
and U5080 (N_5080,N_4374,N_4464);
nand U5081 (N_5081,N_4062,N_4742);
or U5082 (N_5082,N_4061,N_4422);
nor U5083 (N_5083,N_4992,N_4734);
and U5084 (N_5084,N_4398,N_4885);
nor U5085 (N_5085,N_4856,N_4931);
nand U5086 (N_5086,N_4591,N_4471);
and U5087 (N_5087,N_4176,N_4318);
or U5088 (N_5088,N_4986,N_4477);
or U5089 (N_5089,N_4996,N_4002);
nand U5090 (N_5090,N_4815,N_4209);
xnor U5091 (N_5091,N_4714,N_4074);
or U5092 (N_5092,N_4917,N_4783);
nand U5093 (N_5093,N_4152,N_4207);
nand U5094 (N_5094,N_4045,N_4408);
nand U5095 (N_5095,N_4863,N_4858);
and U5096 (N_5096,N_4509,N_4384);
or U5097 (N_5097,N_4462,N_4941);
and U5098 (N_5098,N_4659,N_4871);
nor U5099 (N_5099,N_4673,N_4955);
nand U5100 (N_5100,N_4463,N_4302);
or U5101 (N_5101,N_4431,N_4403);
or U5102 (N_5102,N_4344,N_4032);
or U5103 (N_5103,N_4838,N_4480);
nand U5104 (N_5104,N_4442,N_4997);
nor U5105 (N_5105,N_4716,N_4914);
nand U5106 (N_5106,N_4253,N_4840);
or U5107 (N_5107,N_4880,N_4513);
or U5108 (N_5108,N_4261,N_4192);
or U5109 (N_5109,N_4205,N_4901);
and U5110 (N_5110,N_4467,N_4934);
nand U5111 (N_5111,N_4720,N_4899);
and U5112 (N_5112,N_4920,N_4246);
and U5113 (N_5113,N_4701,N_4472);
nor U5114 (N_5114,N_4757,N_4686);
nor U5115 (N_5115,N_4874,N_4147);
and U5116 (N_5116,N_4563,N_4769);
or U5117 (N_5117,N_4853,N_4036);
nand U5118 (N_5118,N_4404,N_4436);
and U5119 (N_5119,N_4021,N_4758);
nand U5120 (N_5120,N_4134,N_4183);
nor U5121 (N_5121,N_4836,N_4311);
nor U5122 (N_5122,N_4230,N_4832);
nand U5123 (N_5123,N_4903,N_4574);
nor U5124 (N_5124,N_4983,N_4954);
nand U5125 (N_5125,N_4109,N_4658);
and U5126 (N_5126,N_4019,N_4493);
and U5127 (N_5127,N_4626,N_4297);
nand U5128 (N_5128,N_4935,N_4843);
and U5129 (N_5129,N_4557,N_4323);
or U5130 (N_5130,N_4796,N_4256);
nand U5131 (N_5131,N_4748,N_4618);
nand U5132 (N_5132,N_4963,N_4140);
nor U5133 (N_5133,N_4867,N_4522);
nand U5134 (N_5134,N_4946,N_4953);
nand U5135 (N_5135,N_4495,N_4112);
nor U5136 (N_5136,N_4208,N_4976);
and U5137 (N_5137,N_4123,N_4975);
or U5138 (N_5138,N_4204,N_4566);
nand U5139 (N_5139,N_4900,N_4575);
nor U5140 (N_5140,N_4020,N_4961);
and U5141 (N_5141,N_4107,N_4465);
or U5142 (N_5142,N_4492,N_4077);
and U5143 (N_5143,N_4582,N_4049);
nand U5144 (N_5144,N_4510,N_4153);
or U5145 (N_5145,N_4951,N_4106);
and U5146 (N_5146,N_4809,N_4065);
or U5147 (N_5147,N_4400,N_4226);
and U5148 (N_5148,N_4829,N_4541);
nand U5149 (N_5149,N_4232,N_4990);
and U5150 (N_5150,N_4562,N_4960);
or U5151 (N_5151,N_4760,N_4034);
nor U5152 (N_5152,N_4613,N_4199);
nor U5153 (N_5153,N_4080,N_4338);
nand U5154 (N_5154,N_4078,N_4310);
or U5155 (N_5155,N_4179,N_4340);
or U5156 (N_5156,N_4979,N_4101);
nor U5157 (N_5157,N_4807,N_4897);
or U5158 (N_5158,N_4644,N_4317);
nor U5159 (N_5159,N_4424,N_4469);
or U5160 (N_5160,N_4103,N_4526);
nor U5161 (N_5161,N_4670,N_4396);
or U5162 (N_5162,N_4304,N_4088);
or U5163 (N_5163,N_4322,N_4967);
or U5164 (N_5164,N_4368,N_4365);
nor U5165 (N_5165,N_4624,N_4847);
nand U5166 (N_5166,N_4177,N_4915);
or U5167 (N_5167,N_4057,N_4759);
or U5168 (N_5168,N_4762,N_4458);
nor U5169 (N_5169,N_4561,N_4546);
nand U5170 (N_5170,N_4352,N_4124);
nor U5171 (N_5171,N_4161,N_4678);
and U5172 (N_5172,N_4444,N_4764);
nand U5173 (N_5173,N_4303,N_4597);
or U5174 (N_5174,N_4985,N_4483);
nor U5175 (N_5175,N_4877,N_4415);
or U5176 (N_5176,N_4265,N_4457);
nand U5177 (N_5177,N_4274,N_4733);
and U5178 (N_5178,N_4258,N_4058);
nand U5179 (N_5179,N_4489,N_4601);
nand U5180 (N_5180,N_4910,N_4887);
nor U5181 (N_5181,N_4625,N_4620);
nand U5182 (N_5182,N_4993,N_4602);
or U5183 (N_5183,N_4827,N_4824);
or U5184 (N_5184,N_4127,N_4373);
and U5185 (N_5185,N_4280,N_4537);
xor U5186 (N_5186,N_4133,N_4518);
nor U5187 (N_5187,N_4347,N_4922);
and U5188 (N_5188,N_4429,N_4281);
nand U5189 (N_5189,N_4113,N_4060);
or U5190 (N_5190,N_4725,N_4105);
nand U5191 (N_5191,N_4089,N_4348);
nor U5192 (N_5192,N_4928,N_4750);
and U5193 (N_5193,N_4216,N_4353);
and U5194 (N_5194,N_4929,N_4959);
nand U5195 (N_5195,N_4412,N_4413);
or U5196 (N_5196,N_4156,N_4565);
nor U5197 (N_5197,N_4595,N_4968);
nand U5198 (N_5198,N_4936,N_4666);
nor U5199 (N_5199,N_4427,N_4741);
nor U5200 (N_5200,N_4018,N_4589);
or U5201 (N_5201,N_4099,N_4912);
or U5202 (N_5202,N_4726,N_4693);
nand U5203 (N_5203,N_4502,N_4110);
nand U5204 (N_5204,N_4320,N_4041);
or U5205 (N_5205,N_4453,N_4137);
or U5206 (N_5206,N_4713,N_4243);
and U5207 (N_5207,N_4210,N_4025);
nand U5208 (N_5208,N_4789,N_4944);
and U5209 (N_5209,N_4505,N_4870);
nor U5210 (N_5210,N_4957,N_4916);
nand U5211 (N_5211,N_4770,N_4893);
and U5212 (N_5212,N_4411,N_4206);
or U5213 (N_5213,N_4615,N_4767);
or U5214 (N_5214,N_4100,N_4539);
nor U5215 (N_5215,N_4481,N_4096);
or U5216 (N_5216,N_4418,N_4095);
or U5217 (N_5217,N_4519,N_4696);
and U5218 (N_5218,N_4288,N_4221);
and U5219 (N_5219,N_4982,N_4649);
nand U5220 (N_5220,N_4084,N_4584);
nor U5221 (N_5221,N_4397,N_4271);
nand U5222 (N_5222,N_4605,N_4702);
and U5223 (N_5223,N_4301,N_4015);
nand U5224 (N_5224,N_4826,N_4694);
and U5225 (N_5225,N_4242,N_4357);
nand U5226 (N_5226,N_4814,N_4409);
nor U5227 (N_5227,N_4687,N_4476);
nand U5228 (N_5228,N_4146,N_4068);
nor U5229 (N_5229,N_4977,N_4706);
or U5230 (N_5230,N_4980,N_4170);
and U5231 (N_5231,N_4059,N_4187);
or U5232 (N_5232,N_4608,N_4312);
or U5233 (N_5233,N_4593,N_4841);
nor U5234 (N_5234,N_4544,N_4285);
or U5235 (N_5235,N_4860,N_4520);
and U5236 (N_5236,N_4321,N_4548);
nor U5237 (N_5237,N_4781,N_4195);
nand U5238 (N_5238,N_4430,N_4052);
nor U5239 (N_5239,N_4309,N_4331);
nor U5240 (N_5240,N_4555,N_4333);
and U5241 (N_5241,N_4576,N_4496);
xnor U5242 (N_5242,N_4642,N_4468);
or U5243 (N_5243,N_4023,N_4048);
and U5244 (N_5244,N_4545,N_4825);
and U5245 (N_5245,N_4228,N_4707);
nand U5246 (N_5246,N_4805,N_4525);
nand U5247 (N_5247,N_4500,N_4006);
nor U5248 (N_5248,N_4692,N_4369);
and U5249 (N_5249,N_4940,N_4538);
nor U5250 (N_5250,N_4290,N_4984);
or U5251 (N_5251,N_4342,N_4813);
or U5252 (N_5252,N_4499,N_4448);
xor U5253 (N_5253,N_4402,N_4276);
nor U5254 (N_5254,N_4695,N_4684);
and U5255 (N_5255,N_4126,N_4911);
or U5256 (N_5256,N_4751,N_4621);
or U5257 (N_5257,N_4160,N_4000);
nand U5258 (N_5258,N_4459,N_4745);
xor U5259 (N_5259,N_4966,N_4394);
nand U5260 (N_5260,N_4440,N_4401);
or U5261 (N_5261,N_4780,N_4260);
or U5262 (N_5262,N_4371,N_4033);
and U5263 (N_5263,N_4820,N_4363);
nor U5264 (N_5264,N_4439,N_4837);
nor U5265 (N_5265,N_4007,N_4512);
nand U5266 (N_5266,N_4482,N_4270);
or U5267 (N_5267,N_4001,N_4822);
nand U5268 (N_5268,N_4391,N_4700);
nand U5269 (N_5269,N_4135,N_4460);
nand U5270 (N_5270,N_4913,N_4866);
nand U5271 (N_5271,N_4050,N_4610);
nor U5272 (N_5272,N_4514,N_4447);
or U5273 (N_5273,N_4895,N_4623);
and U5274 (N_5274,N_4638,N_4416);
and U5275 (N_5275,N_4255,N_4819);
nor U5276 (N_5276,N_4521,N_4359);
nor U5277 (N_5277,N_4619,N_4728);
nand U5278 (N_5278,N_4299,N_4668);
nor U5279 (N_5279,N_4393,N_4690);
or U5280 (N_5280,N_4231,N_4806);
xnor U5281 (N_5281,N_4056,N_4987);
nand U5282 (N_5282,N_4834,N_4349);
or U5283 (N_5283,N_4307,N_4143);
nor U5284 (N_5284,N_4115,N_4587);
and U5285 (N_5285,N_4553,N_4679);
nor U5286 (N_5286,N_4011,N_4335);
nand U5287 (N_5287,N_4717,N_4375);
nand U5288 (N_5288,N_4981,N_4259);
nor U5289 (N_5289,N_4812,N_4155);
nand U5290 (N_5290,N_4128,N_4746);
or U5291 (N_5291,N_4709,N_4009);
nand U5292 (N_5292,N_4224,N_4434);
and U5293 (N_5293,N_4324,N_4719);
nor U5294 (N_5294,N_4688,N_4795);
or U5295 (N_5295,N_4116,N_4184);
or U5296 (N_5296,N_4842,N_4343);
or U5297 (N_5297,N_4200,N_4395);
and U5298 (N_5298,N_4927,N_4329);
nor U5299 (N_5299,N_4308,N_4341);
and U5300 (N_5300,N_4064,N_4454);
and U5301 (N_5301,N_4425,N_4292);
or U5302 (N_5302,N_4802,N_4817);
or U5303 (N_5303,N_4428,N_4849);
nand U5304 (N_5304,N_4850,N_4662);
xor U5305 (N_5305,N_4225,N_4423);
and U5306 (N_5306,N_4186,N_4594);
and U5307 (N_5307,N_4898,N_4596);
nor U5308 (N_5308,N_4385,N_4891);
and U5309 (N_5309,N_4752,N_4777);
nor U5310 (N_5310,N_4697,N_4676);
nor U5311 (N_5311,N_4821,N_4055);
or U5312 (N_5312,N_4180,N_4358);
nand U5313 (N_5313,N_4250,N_4142);
nand U5314 (N_5314,N_4054,N_4945);
and U5315 (N_5315,N_4449,N_4739);
and U5316 (N_5316,N_4355,N_4252);
and U5317 (N_5317,N_4046,N_4508);
or U5318 (N_5318,N_4053,N_4157);
and U5319 (N_5319,N_4473,N_4229);
or U5320 (N_5320,N_4730,N_4995);
nand U5321 (N_5321,N_4278,N_4194);
nor U5322 (N_5322,N_4158,N_4392);
and U5323 (N_5323,N_4786,N_4295);
xnor U5324 (N_5324,N_4346,N_4703);
nand U5325 (N_5325,N_4016,N_4450);
nor U5326 (N_5326,N_4532,N_4269);
nor U5327 (N_5327,N_4634,N_4889);
or U5328 (N_5328,N_4377,N_4031);
or U5329 (N_5329,N_4138,N_4390);
nand U5330 (N_5330,N_4354,N_4071);
and U5331 (N_5331,N_4379,N_4178);
nand U5332 (N_5332,N_4908,N_4943);
or U5333 (N_5333,N_4086,N_4664);
nand U5334 (N_5334,N_4003,N_4063);
nand U5335 (N_5335,N_4139,N_4326);
and U5336 (N_5336,N_4498,N_4846);
nand U5337 (N_5337,N_4197,N_4699);
or U5338 (N_5338,N_4217,N_4043);
nand U5339 (N_5339,N_4782,N_4600);
and U5340 (N_5340,N_4486,N_4848);
and U5341 (N_5341,N_4533,N_4851);
or U5342 (N_5342,N_4724,N_4298);
or U5343 (N_5343,N_4066,N_4213);
and U5344 (N_5344,N_4855,N_4351);
or U5345 (N_5345,N_4991,N_4141);
nor U5346 (N_5346,N_4073,N_4766);
nor U5347 (N_5347,N_4097,N_4273);
and U5348 (N_5348,N_4749,N_4121);
and U5349 (N_5349,N_4729,N_4873);
nand U5350 (N_5350,N_4793,N_4254);
or U5351 (N_5351,N_4484,N_4070);
and U5352 (N_5352,N_4609,N_4810);
nand U5353 (N_5353,N_4028,N_4325);
and U5354 (N_5354,N_4263,N_4628);
nand U5355 (N_5355,N_4845,N_4202);
or U5356 (N_5356,N_4092,N_4698);
nor U5357 (N_5357,N_4120,N_4535);
nor U5358 (N_5358,N_4784,N_4882);
nand U5359 (N_5359,N_4013,N_4136);
nor U5360 (N_5360,N_4300,N_4282);
or U5361 (N_5361,N_4524,N_4586);
nand U5362 (N_5362,N_4785,N_4466);
nand U5363 (N_5363,N_4218,N_4098);
nand U5364 (N_5364,N_4435,N_4736);
or U5365 (N_5365,N_4778,N_4296);
nand U5366 (N_5366,N_4558,N_4614);
nand U5367 (N_5367,N_4159,N_4721);
xnor U5368 (N_5368,N_4680,N_4577);
or U5369 (N_5369,N_4211,N_4497);
nor U5370 (N_5370,N_4559,N_4854);
nand U5371 (N_5371,N_4833,N_4487);
nor U5372 (N_5372,N_4798,N_4768);
or U5373 (N_5373,N_4163,N_4456);
nand U5374 (N_5374,N_4345,N_4038);
nor U5375 (N_5375,N_4740,N_4012);
and U5376 (N_5376,N_4999,N_4174);
or U5377 (N_5377,N_4169,N_4264);
or U5378 (N_5378,N_4027,N_4923);
nand U5379 (N_5379,N_4334,N_4381);
and U5380 (N_5380,N_4675,N_4715);
or U5381 (N_5381,N_4076,N_4753);
or U5382 (N_5382,N_4378,N_4603);
nor U5383 (N_5383,N_4154,N_4896);
or U5384 (N_5384,N_4249,N_4005);
and U5385 (N_5385,N_4082,N_4682);
or U5386 (N_5386,N_4306,N_4667);
and U5387 (N_5387,N_4240,N_4069);
and U5388 (N_5388,N_4571,N_4657);
xor U5389 (N_5389,N_4599,N_4093);
nand U5390 (N_5390,N_4171,N_4090);
nor U5391 (N_5391,N_4633,N_4627);
and U5392 (N_5392,N_4079,N_4663);
nor U5393 (N_5393,N_4904,N_4026);
nor U5394 (N_5394,N_4949,N_4029);
xor U5395 (N_5395,N_4930,N_4653);
nand U5396 (N_5396,N_4952,N_4731);
xor U5397 (N_5397,N_4844,N_4797);
or U5398 (N_5398,N_4426,N_4248);
nand U5399 (N_5399,N_4414,N_4287);
or U5400 (N_5400,N_4380,N_4865);
or U5401 (N_5401,N_4672,N_4083);
or U5402 (N_5402,N_4564,N_4443);
and U5403 (N_5403,N_4570,N_4554);
nor U5404 (N_5404,N_4488,N_4327);
nor U5405 (N_5405,N_4291,N_4072);
and U5406 (N_5406,N_4655,N_4652);
and U5407 (N_5407,N_4761,N_4364);
and U5408 (N_5408,N_4978,N_4530);
and U5409 (N_5409,N_4902,N_4631);
and U5410 (N_5410,N_4660,N_4617);
and U5411 (N_5411,N_4085,N_4583);
or U5412 (N_5412,N_4188,N_4998);
and U5413 (N_5413,N_4438,N_4515);
and U5414 (N_5414,N_4337,N_4239);
nand U5415 (N_5415,N_4330,N_4788);
nand U5416 (N_5416,N_4227,N_4585);
nor U5417 (N_5417,N_4547,N_4550);
or U5418 (N_5418,N_4886,N_4004);
and U5419 (N_5419,N_4193,N_4639);
or U5420 (N_5420,N_4683,N_4257);
nor U5421 (N_5421,N_4932,N_4791);
or U5422 (N_5422,N_4091,N_4973);
or U5423 (N_5423,N_4919,N_4172);
nor U5424 (N_5424,N_4017,N_4888);
nor U5425 (N_5425,N_4531,N_4878);
or U5426 (N_5426,N_4284,N_4241);
or U5427 (N_5427,N_4969,N_4776);
or U5428 (N_5428,N_4607,N_4800);
and U5429 (N_5429,N_4523,N_4971);
xnor U5430 (N_5430,N_4839,N_4314);
nor U5431 (N_5431,N_4111,N_4386);
or U5432 (N_5432,N_4516,N_4035);
or U5433 (N_5433,N_4765,N_4234);
or U5434 (N_5434,N_4794,N_4950);
nand U5435 (N_5435,N_4504,N_4151);
nor U5436 (N_5436,N_4517,N_4289);
or U5437 (N_5437,N_4102,N_4862);
and U5438 (N_5438,N_4962,N_4198);
nor U5439 (N_5439,N_4024,N_4861);
nand U5440 (N_5440,N_4705,N_4852);
nor U5441 (N_5441,N_4328,N_4201);
nor U5442 (N_5442,N_4876,N_4879);
nor U5443 (N_5443,N_4220,N_4356);
nand U5444 (N_5444,N_4803,N_4336);
and U5445 (N_5445,N_4162,N_4674);
and U5446 (N_5446,N_4490,N_4604);
nor U5447 (N_5447,N_4681,N_4022);
nand U5448 (N_5448,N_4010,N_4828);
nand U5449 (N_5449,N_4933,N_4737);
or U5450 (N_5450,N_4407,N_4388);
or U5451 (N_5451,N_4560,N_4598);
and U5452 (N_5452,N_4708,N_4405);
or U5453 (N_5453,N_4857,N_4956);
nor U5454 (N_5454,N_4612,N_4808);
nor U5455 (N_5455,N_4647,N_4313);
nor U5456 (N_5456,N_4884,N_4383);
and U5457 (N_5457,N_4131,N_4455);
and U5458 (N_5458,N_4051,N_4763);
nor U5459 (N_5459,N_4277,N_4881);
or U5460 (N_5460,N_4704,N_4588);
or U5461 (N_5461,N_4419,N_4372);
nand U5462 (N_5462,N_4743,N_4771);
or U5463 (N_5463,N_4606,N_4640);
nand U5464 (N_5464,N_4622,N_4773);
and U5465 (N_5465,N_4864,N_4279);
nor U5466 (N_5466,N_4044,N_4119);
or U5467 (N_5467,N_4989,N_4835);
nand U5468 (N_5468,N_4727,N_4366);
nand U5469 (N_5469,N_4189,N_4925);
and U5470 (N_5470,N_4868,N_4272);
nand U5471 (N_5471,N_4275,N_4222);
or U5472 (N_5472,N_4818,N_4551);
or U5473 (N_5473,N_4149,N_4787);
or U5474 (N_5474,N_4266,N_4578);
nor U5475 (N_5475,N_4181,N_4799);
or U5476 (N_5476,N_4641,N_4869);
or U5477 (N_5477,N_4590,N_4552);
nand U5478 (N_5478,N_4665,N_4629);
nand U5479 (N_5479,N_4756,N_4747);
nand U5480 (N_5480,N_4150,N_4067);
xnor U5481 (N_5481,N_4319,N_4501);
or U5482 (N_5482,N_4238,N_4974);
nor U5483 (N_5483,N_4185,N_4964);
nor U5484 (N_5484,N_4233,N_4938);
nand U5485 (N_5485,N_4316,N_4190);
nor U5486 (N_5486,N_4118,N_4710);
nand U5487 (N_5487,N_4556,N_4339);
nor U5488 (N_5488,N_4376,N_4164);
nor U5489 (N_5489,N_4203,N_4651);
and U5490 (N_5490,N_4294,N_4905);
nor U5491 (N_5491,N_4360,N_4689);
and U5492 (N_5492,N_4994,N_4830);
nand U5493 (N_5493,N_4494,N_4479);
and U5494 (N_5494,N_4528,N_4117);
or U5495 (N_5495,N_4948,N_4212);
or U5496 (N_5496,N_4382,N_4432);
or U5497 (N_5497,N_4685,N_4478);
nand U5498 (N_5498,N_4712,N_4965);
and U5499 (N_5499,N_4735,N_4125);
or U5500 (N_5500,N_4458,N_4540);
nor U5501 (N_5501,N_4109,N_4955);
or U5502 (N_5502,N_4467,N_4015);
nand U5503 (N_5503,N_4303,N_4061);
and U5504 (N_5504,N_4807,N_4842);
nor U5505 (N_5505,N_4821,N_4249);
nor U5506 (N_5506,N_4828,N_4630);
nand U5507 (N_5507,N_4254,N_4609);
or U5508 (N_5508,N_4549,N_4719);
or U5509 (N_5509,N_4557,N_4733);
or U5510 (N_5510,N_4921,N_4673);
nand U5511 (N_5511,N_4951,N_4604);
or U5512 (N_5512,N_4066,N_4087);
nand U5513 (N_5513,N_4637,N_4148);
or U5514 (N_5514,N_4621,N_4784);
or U5515 (N_5515,N_4936,N_4601);
and U5516 (N_5516,N_4662,N_4411);
nand U5517 (N_5517,N_4886,N_4937);
and U5518 (N_5518,N_4720,N_4304);
and U5519 (N_5519,N_4161,N_4090);
and U5520 (N_5520,N_4223,N_4851);
or U5521 (N_5521,N_4987,N_4146);
and U5522 (N_5522,N_4451,N_4241);
nand U5523 (N_5523,N_4321,N_4279);
nor U5524 (N_5524,N_4705,N_4247);
or U5525 (N_5525,N_4518,N_4493);
and U5526 (N_5526,N_4065,N_4499);
and U5527 (N_5527,N_4181,N_4310);
and U5528 (N_5528,N_4409,N_4875);
nor U5529 (N_5529,N_4774,N_4653);
or U5530 (N_5530,N_4816,N_4392);
nand U5531 (N_5531,N_4325,N_4793);
or U5532 (N_5532,N_4036,N_4623);
or U5533 (N_5533,N_4822,N_4930);
nand U5534 (N_5534,N_4413,N_4518);
nand U5535 (N_5535,N_4385,N_4403);
or U5536 (N_5536,N_4369,N_4093);
nand U5537 (N_5537,N_4797,N_4924);
and U5538 (N_5538,N_4072,N_4793);
or U5539 (N_5539,N_4503,N_4063);
and U5540 (N_5540,N_4396,N_4052);
or U5541 (N_5541,N_4105,N_4576);
nand U5542 (N_5542,N_4034,N_4467);
nor U5543 (N_5543,N_4884,N_4501);
and U5544 (N_5544,N_4620,N_4642);
and U5545 (N_5545,N_4470,N_4844);
and U5546 (N_5546,N_4934,N_4919);
nand U5547 (N_5547,N_4723,N_4569);
or U5548 (N_5548,N_4119,N_4033);
nand U5549 (N_5549,N_4246,N_4938);
or U5550 (N_5550,N_4394,N_4057);
nand U5551 (N_5551,N_4694,N_4494);
and U5552 (N_5552,N_4011,N_4262);
xnor U5553 (N_5553,N_4398,N_4633);
nand U5554 (N_5554,N_4508,N_4015);
or U5555 (N_5555,N_4520,N_4340);
nand U5556 (N_5556,N_4307,N_4331);
nor U5557 (N_5557,N_4660,N_4891);
nand U5558 (N_5558,N_4202,N_4507);
or U5559 (N_5559,N_4374,N_4602);
nor U5560 (N_5560,N_4031,N_4110);
nand U5561 (N_5561,N_4210,N_4125);
and U5562 (N_5562,N_4284,N_4653);
nand U5563 (N_5563,N_4092,N_4708);
nor U5564 (N_5564,N_4627,N_4844);
nand U5565 (N_5565,N_4792,N_4617);
nand U5566 (N_5566,N_4899,N_4194);
nor U5567 (N_5567,N_4575,N_4771);
nand U5568 (N_5568,N_4156,N_4102);
and U5569 (N_5569,N_4820,N_4699);
and U5570 (N_5570,N_4330,N_4955);
and U5571 (N_5571,N_4615,N_4749);
nand U5572 (N_5572,N_4458,N_4989);
nor U5573 (N_5573,N_4033,N_4662);
nand U5574 (N_5574,N_4408,N_4680);
nor U5575 (N_5575,N_4102,N_4838);
nand U5576 (N_5576,N_4090,N_4253);
nor U5577 (N_5577,N_4425,N_4532);
nand U5578 (N_5578,N_4983,N_4719);
or U5579 (N_5579,N_4846,N_4945);
nand U5580 (N_5580,N_4148,N_4103);
and U5581 (N_5581,N_4598,N_4106);
or U5582 (N_5582,N_4597,N_4136);
and U5583 (N_5583,N_4030,N_4792);
or U5584 (N_5584,N_4068,N_4995);
nand U5585 (N_5585,N_4119,N_4730);
nor U5586 (N_5586,N_4186,N_4781);
and U5587 (N_5587,N_4433,N_4538);
and U5588 (N_5588,N_4315,N_4401);
or U5589 (N_5589,N_4400,N_4587);
nor U5590 (N_5590,N_4428,N_4758);
and U5591 (N_5591,N_4100,N_4976);
nand U5592 (N_5592,N_4997,N_4469);
or U5593 (N_5593,N_4388,N_4202);
nand U5594 (N_5594,N_4633,N_4843);
nand U5595 (N_5595,N_4710,N_4353);
and U5596 (N_5596,N_4076,N_4507);
or U5597 (N_5597,N_4631,N_4889);
nor U5598 (N_5598,N_4577,N_4271);
nand U5599 (N_5599,N_4190,N_4894);
nor U5600 (N_5600,N_4095,N_4780);
and U5601 (N_5601,N_4927,N_4041);
or U5602 (N_5602,N_4295,N_4227);
or U5603 (N_5603,N_4630,N_4868);
nor U5604 (N_5604,N_4629,N_4149);
and U5605 (N_5605,N_4378,N_4453);
nand U5606 (N_5606,N_4518,N_4017);
nand U5607 (N_5607,N_4362,N_4114);
nor U5608 (N_5608,N_4645,N_4290);
nor U5609 (N_5609,N_4039,N_4295);
nor U5610 (N_5610,N_4412,N_4931);
and U5611 (N_5611,N_4636,N_4269);
or U5612 (N_5612,N_4093,N_4414);
or U5613 (N_5613,N_4540,N_4528);
and U5614 (N_5614,N_4818,N_4302);
or U5615 (N_5615,N_4557,N_4218);
nand U5616 (N_5616,N_4523,N_4399);
nand U5617 (N_5617,N_4711,N_4720);
nor U5618 (N_5618,N_4541,N_4360);
nand U5619 (N_5619,N_4888,N_4307);
or U5620 (N_5620,N_4152,N_4830);
nand U5621 (N_5621,N_4579,N_4312);
or U5622 (N_5622,N_4663,N_4285);
nand U5623 (N_5623,N_4958,N_4136);
nor U5624 (N_5624,N_4776,N_4015);
nor U5625 (N_5625,N_4999,N_4251);
nand U5626 (N_5626,N_4293,N_4895);
nand U5627 (N_5627,N_4237,N_4016);
or U5628 (N_5628,N_4660,N_4812);
nand U5629 (N_5629,N_4505,N_4532);
nor U5630 (N_5630,N_4490,N_4569);
nand U5631 (N_5631,N_4661,N_4076);
nor U5632 (N_5632,N_4475,N_4687);
or U5633 (N_5633,N_4973,N_4755);
or U5634 (N_5634,N_4250,N_4548);
and U5635 (N_5635,N_4653,N_4892);
nor U5636 (N_5636,N_4402,N_4498);
nor U5637 (N_5637,N_4576,N_4299);
and U5638 (N_5638,N_4181,N_4449);
and U5639 (N_5639,N_4319,N_4347);
nor U5640 (N_5640,N_4425,N_4089);
and U5641 (N_5641,N_4116,N_4646);
nand U5642 (N_5642,N_4133,N_4980);
nand U5643 (N_5643,N_4815,N_4754);
or U5644 (N_5644,N_4516,N_4419);
and U5645 (N_5645,N_4247,N_4523);
and U5646 (N_5646,N_4922,N_4173);
or U5647 (N_5647,N_4202,N_4869);
nand U5648 (N_5648,N_4405,N_4159);
nor U5649 (N_5649,N_4244,N_4505);
nand U5650 (N_5650,N_4512,N_4880);
nor U5651 (N_5651,N_4120,N_4098);
nor U5652 (N_5652,N_4340,N_4446);
or U5653 (N_5653,N_4117,N_4067);
nand U5654 (N_5654,N_4274,N_4508);
nor U5655 (N_5655,N_4683,N_4294);
nor U5656 (N_5656,N_4141,N_4208);
nand U5657 (N_5657,N_4659,N_4555);
nor U5658 (N_5658,N_4729,N_4173);
and U5659 (N_5659,N_4631,N_4892);
and U5660 (N_5660,N_4124,N_4891);
or U5661 (N_5661,N_4532,N_4473);
nand U5662 (N_5662,N_4530,N_4144);
or U5663 (N_5663,N_4678,N_4638);
and U5664 (N_5664,N_4323,N_4520);
nor U5665 (N_5665,N_4702,N_4504);
nor U5666 (N_5666,N_4951,N_4575);
xor U5667 (N_5667,N_4737,N_4085);
nor U5668 (N_5668,N_4519,N_4943);
and U5669 (N_5669,N_4530,N_4477);
or U5670 (N_5670,N_4566,N_4023);
or U5671 (N_5671,N_4605,N_4879);
nand U5672 (N_5672,N_4615,N_4368);
nand U5673 (N_5673,N_4347,N_4483);
or U5674 (N_5674,N_4773,N_4009);
and U5675 (N_5675,N_4289,N_4419);
or U5676 (N_5676,N_4607,N_4827);
or U5677 (N_5677,N_4337,N_4724);
nand U5678 (N_5678,N_4281,N_4066);
nand U5679 (N_5679,N_4654,N_4790);
nor U5680 (N_5680,N_4026,N_4659);
nor U5681 (N_5681,N_4522,N_4031);
nor U5682 (N_5682,N_4512,N_4249);
and U5683 (N_5683,N_4161,N_4348);
nor U5684 (N_5684,N_4935,N_4451);
nor U5685 (N_5685,N_4090,N_4139);
or U5686 (N_5686,N_4178,N_4846);
and U5687 (N_5687,N_4617,N_4210);
nand U5688 (N_5688,N_4553,N_4537);
or U5689 (N_5689,N_4611,N_4997);
or U5690 (N_5690,N_4694,N_4096);
and U5691 (N_5691,N_4922,N_4669);
nand U5692 (N_5692,N_4727,N_4317);
nor U5693 (N_5693,N_4626,N_4535);
and U5694 (N_5694,N_4381,N_4148);
and U5695 (N_5695,N_4134,N_4591);
nand U5696 (N_5696,N_4883,N_4817);
nand U5697 (N_5697,N_4718,N_4179);
or U5698 (N_5698,N_4168,N_4218);
nor U5699 (N_5699,N_4313,N_4515);
nand U5700 (N_5700,N_4794,N_4961);
and U5701 (N_5701,N_4419,N_4772);
and U5702 (N_5702,N_4563,N_4587);
nor U5703 (N_5703,N_4765,N_4799);
nand U5704 (N_5704,N_4340,N_4022);
nand U5705 (N_5705,N_4719,N_4138);
or U5706 (N_5706,N_4126,N_4617);
nor U5707 (N_5707,N_4623,N_4103);
or U5708 (N_5708,N_4149,N_4274);
or U5709 (N_5709,N_4017,N_4829);
nor U5710 (N_5710,N_4855,N_4676);
nor U5711 (N_5711,N_4324,N_4343);
nand U5712 (N_5712,N_4380,N_4062);
or U5713 (N_5713,N_4965,N_4503);
nor U5714 (N_5714,N_4105,N_4135);
nand U5715 (N_5715,N_4575,N_4194);
nand U5716 (N_5716,N_4050,N_4832);
nand U5717 (N_5717,N_4260,N_4658);
xnor U5718 (N_5718,N_4795,N_4140);
and U5719 (N_5719,N_4723,N_4963);
nand U5720 (N_5720,N_4766,N_4977);
nand U5721 (N_5721,N_4607,N_4183);
or U5722 (N_5722,N_4526,N_4045);
nand U5723 (N_5723,N_4489,N_4605);
nor U5724 (N_5724,N_4848,N_4246);
and U5725 (N_5725,N_4656,N_4718);
or U5726 (N_5726,N_4609,N_4897);
and U5727 (N_5727,N_4358,N_4984);
and U5728 (N_5728,N_4791,N_4647);
nand U5729 (N_5729,N_4274,N_4791);
and U5730 (N_5730,N_4965,N_4788);
or U5731 (N_5731,N_4931,N_4590);
or U5732 (N_5732,N_4814,N_4549);
or U5733 (N_5733,N_4674,N_4417);
and U5734 (N_5734,N_4683,N_4088);
nor U5735 (N_5735,N_4320,N_4899);
or U5736 (N_5736,N_4150,N_4430);
or U5737 (N_5737,N_4300,N_4782);
or U5738 (N_5738,N_4257,N_4422);
nand U5739 (N_5739,N_4252,N_4733);
or U5740 (N_5740,N_4335,N_4161);
nand U5741 (N_5741,N_4697,N_4462);
nor U5742 (N_5742,N_4036,N_4297);
nor U5743 (N_5743,N_4941,N_4530);
or U5744 (N_5744,N_4746,N_4797);
nand U5745 (N_5745,N_4686,N_4901);
or U5746 (N_5746,N_4746,N_4547);
or U5747 (N_5747,N_4776,N_4429);
or U5748 (N_5748,N_4408,N_4687);
or U5749 (N_5749,N_4231,N_4851);
or U5750 (N_5750,N_4164,N_4356);
nor U5751 (N_5751,N_4629,N_4843);
or U5752 (N_5752,N_4678,N_4188);
nand U5753 (N_5753,N_4744,N_4351);
nor U5754 (N_5754,N_4571,N_4694);
nand U5755 (N_5755,N_4371,N_4218);
nor U5756 (N_5756,N_4942,N_4586);
nand U5757 (N_5757,N_4601,N_4151);
or U5758 (N_5758,N_4852,N_4427);
and U5759 (N_5759,N_4256,N_4395);
and U5760 (N_5760,N_4137,N_4558);
or U5761 (N_5761,N_4906,N_4243);
nand U5762 (N_5762,N_4737,N_4261);
or U5763 (N_5763,N_4013,N_4823);
and U5764 (N_5764,N_4670,N_4676);
and U5765 (N_5765,N_4477,N_4714);
nor U5766 (N_5766,N_4962,N_4369);
nand U5767 (N_5767,N_4183,N_4236);
nor U5768 (N_5768,N_4467,N_4633);
and U5769 (N_5769,N_4960,N_4262);
or U5770 (N_5770,N_4998,N_4521);
or U5771 (N_5771,N_4111,N_4005);
nand U5772 (N_5772,N_4479,N_4318);
and U5773 (N_5773,N_4756,N_4007);
nand U5774 (N_5774,N_4457,N_4479);
or U5775 (N_5775,N_4301,N_4755);
nor U5776 (N_5776,N_4246,N_4811);
nor U5777 (N_5777,N_4952,N_4368);
or U5778 (N_5778,N_4717,N_4560);
nand U5779 (N_5779,N_4392,N_4041);
nand U5780 (N_5780,N_4160,N_4517);
and U5781 (N_5781,N_4527,N_4673);
or U5782 (N_5782,N_4771,N_4148);
nand U5783 (N_5783,N_4697,N_4300);
and U5784 (N_5784,N_4233,N_4034);
and U5785 (N_5785,N_4386,N_4977);
nor U5786 (N_5786,N_4629,N_4325);
nand U5787 (N_5787,N_4532,N_4760);
and U5788 (N_5788,N_4286,N_4689);
or U5789 (N_5789,N_4516,N_4903);
and U5790 (N_5790,N_4560,N_4646);
nand U5791 (N_5791,N_4492,N_4974);
xnor U5792 (N_5792,N_4457,N_4384);
nand U5793 (N_5793,N_4607,N_4549);
or U5794 (N_5794,N_4679,N_4382);
or U5795 (N_5795,N_4848,N_4855);
nand U5796 (N_5796,N_4004,N_4882);
or U5797 (N_5797,N_4624,N_4439);
nand U5798 (N_5798,N_4141,N_4602);
and U5799 (N_5799,N_4489,N_4296);
and U5800 (N_5800,N_4641,N_4599);
or U5801 (N_5801,N_4594,N_4268);
and U5802 (N_5802,N_4041,N_4440);
and U5803 (N_5803,N_4855,N_4086);
nand U5804 (N_5804,N_4508,N_4721);
nand U5805 (N_5805,N_4171,N_4567);
and U5806 (N_5806,N_4444,N_4199);
and U5807 (N_5807,N_4147,N_4490);
or U5808 (N_5808,N_4160,N_4612);
or U5809 (N_5809,N_4039,N_4963);
and U5810 (N_5810,N_4672,N_4387);
or U5811 (N_5811,N_4578,N_4448);
or U5812 (N_5812,N_4480,N_4546);
or U5813 (N_5813,N_4515,N_4208);
or U5814 (N_5814,N_4397,N_4597);
or U5815 (N_5815,N_4429,N_4363);
and U5816 (N_5816,N_4925,N_4734);
xor U5817 (N_5817,N_4969,N_4296);
and U5818 (N_5818,N_4453,N_4740);
or U5819 (N_5819,N_4457,N_4539);
xnor U5820 (N_5820,N_4733,N_4671);
or U5821 (N_5821,N_4583,N_4499);
nand U5822 (N_5822,N_4477,N_4284);
or U5823 (N_5823,N_4304,N_4610);
and U5824 (N_5824,N_4737,N_4283);
xnor U5825 (N_5825,N_4350,N_4208);
nor U5826 (N_5826,N_4485,N_4395);
nor U5827 (N_5827,N_4678,N_4198);
and U5828 (N_5828,N_4533,N_4264);
and U5829 (N_5829,N_4672,N_4973);
nand U5830 (N_5830,N_4133,N_4495);
nor U5831 (N_5831,N_4285,N_4498);
and U5832 (N_5832,N_4094,N_4303);
and U5833 (N_5833,N_4019,N_4837);
nand U5834 (N_5834,N_4655,N_4716);
and U5835 (N_5835,N_4440,N_4582);
or U5836 (N_5836,N_4940,N_4956);
nor U5837 (N_5837,N_4368,N_4410);
nor U5838 (N_5838,N_4121,N_4679);
nand U5839 (N_5839,N_4378,N_4493);
nand U5840 (N_5840,N_4998,N_4324);
or U5841 (N_5841,N_4634,N_4893);
or U5842 (N_5842,N_4405,N_4031);
nor U5843 (N_5843,N_4058,N_4806);
and U5844 (N_5844,N_4511,N_4374);
nor U5845 (N_5845,N_4244,N_4533);
and U5846 (N_5846,N_4151,N_4693);
and U5847 (N_5847,N_4129,N_4431);
nand U5848 (N_5848,N_4345,N_4487);
and U5849 (N_5849,N_4039,N_4837);
nand U5850 (N_5850,N_4040,N_4649);
or U5851 (N_5851,N_4106,N_4564);
and U5852 (N_5852,N_4457,N_4669);
nand U5853 (N_5853,N_4782,N_4075);
nor U5854 (N_5854,N_4927,N_4251);
nand U5855 (N_5855,N_4588,N_4068);
nor U5856 (N_5856,N_4862,N_4443);
nand U5857 (N_5857,N_4584,N_4455);
or U5858 (N_5858,N_4992,N_4654);
and U5859 (N_5859,N_4264,N_4568);
nor U5860 (N_5860,N_4151,N_4626);
nand U5861 (N_5861,N_4162,N_4421);
and U5862 (N_5862,N_4163,N_4087);
nor U5863 (N_5863,N_4576,N_4520);
nor U5864 (N_5864,N_4722,N_4831);
and U5865 (N_5865,N_4331,N_4621);
xor U5866 (N_5866,N_4217,N_4461);
or U5867 (N_5867,N_4256,N_4878);
nand U5868 (N_5868,N_4368,N_4422);
or U5869 (N_5869,N_4192,N_4056);
and U5870 (N_5870,N_4261,N_4098);
nor U5871 (N_5871,N_4836,N_4714);
and U5872 (N_5872,N_4608,N_4381);
nand U5873 (N_5873,N_4155,N_4672);
nand U5874 (N_5874,N_4998,N_4938);
nor U5875 (N_5875,N_4440,N_4389);
or U5876 (N_5876,N_4317,N_4487);
or U5877 (N_5877,N_4268,N_4832);
xor U5878 (N_5878,N_4189,N_4637);
or U5879 (N_5879,N_4529,N_4272);
nand U5880 (N_5880,N_4108,N_4589);
nand U5881 (N_5881,N_4518,N_4556);
nor U5882 (N_5882,N_4117,N_4593);
nor U5883 (N_5883,N_4836,N_4839);
nand U5884 (N_5884,N_4813,N_4339);
nand U5885 (N_5885,N_4490,N_4698);
and U5886 (N_5886,N_4556,N_4361);
nor U5887 (N_5887,N_4795,N_4871);
or U5888 (N_5888,N_4190,N_4736);
and U5889 (N_5889,N_4659,N_4315);
or U5890 (N_5890,N_4129,N_4706);
nand U5891 (N_5891,N_4918,N_4300);
or U5892 (N_5892,N_4315,N_4089);
and U5893 (N_5893,N_4434,N_4798);
nor U5894 (N_5894,N_4075,N_4244);
or U5895 (N_5895,N_4830,N_4719);
or U5896 (N_5896,N_4015,N_4726);
nor U5897 (N_5897,N_4670,N_4297);
nor U5898 (N_5898,N_4998,N_4774);
xnor U5899 (N_5899,N_4419,N_4607);
nand U5900 (N_5900,N_4875,N_4531);
and U5901 (N_5901,N_4398,N_4675);
nand U5902 (N_5902,N_4337,N_4681);
nor U5903 (N_5903,N_4452,N_4092);
or U5904 (N_5904,N_4769,N_4802);
nor U5905 (N_5905,N_4118,N_4733);
nor U5906 (N_5906,N_4696,N_4772);
xor U5907 (N_5907,N_4200,N_4270);
xor U5908 (N_5908,N_4591,N_4194);
and U5909 (N_5909,N_4758,N_4081);
or U5910 (N_5910,N_4027,N_4645);
xor U5911 (N_5911,N_4881,N_4800);
nor U5912 (N_5912,N_4183,N_4751);
or U5913 (N_5913,N_4552,N_4675);
nor U5914 (N_5914,N_4571,N_4850);
or U5915 (N_5915,N_4418,N_4402);
or U5916 (N_5916,N_4771,N_4228);
nor U5917 (N_5917,N_4362,N_4920);
or U5918 (N_5918,N_4836,N_4596);
nand U5919 (N_5919,N_4909,N_4740);
nor U5920 (N_5920,N_4569,N_4765);
nand U5921 (N_5921,N_4837,N_4224);
and U5922 (N_5922,N_4943,N_4799);
nand U5923 (N_5923,N_4522,N_4854);
or U5924 (N_5924,N_4689,N_4786);
and U5925 (N_5925,N_4465,N_4862);
nor U5926 (N_5926,N_4439,N_4937);
and U5927 (N_5927,N_4550,N_4981);
or U5928 (N_5928,N_4392,N_4025);
and U5929 (N_5929,N_4642,N_4993);
nor U5930 (N_5930,N_4065,N_4781);
xor U5931 (N_5931,N_4137,N_4580);
and U5932 (N_5932,N_4213,N_4227);
and U5933 (N_5933,N_4069,N_4102);
nor U5934 (N_5934,N_4727,N_4135);
nor U5935 (N_5935,N_4136,N_4977);
nor U5936 (N_5936,N_4474,N_4206);
or U5937 (N_5937,N_4434,N_4402);
and U5938 (N_5938,N_4760,N_4027);
nor U5939 (N_5939,N_4372,N_4641);
nand U5940 (N_5940,N_4033,N_4485);
and U5941 (N_5941,N_4398,N_4836);
nor U5942 (N_5942,N_4191,N_4998);
or U5943 (N_5943,N_4344,N_4228);
and U5944 (N_5944,N_4252,N_4262);
or U5945 (N_5945,N_4896,N_4614);
nor U5946 (N_5946,N_4763,N_4401);
nand U5947 (N_5947,N_4651,N_4202);
or U5948 (N_5948,N_4163,N_4314);
or U5949 (N_5949,N_4580,N_4179);
and U5950 (N_5950,N_4905,N_4156);
nor U5951 (N_5951,N_4675,N_4664);
and U5952 (N_5952,N_4808,N_4565);
nand U5953 (N_5953,N_4477,N_4777);
nand U5954 (N_5954,N_4532,N_4319);
nor U5955 (N_5955,N_4848,N_4271);
and U5956 (N_5956,N_4925,N_4716);
nor U5957 (N_5957,N_4651,N_4165);
nand U5958 (N_5958,N_4170,N_4057);
nor U5959 (N_5959,N_4137,N_4838);
nor U5960 (N_5960,N_4224,N_4025);
nor U5961 (N_5961,N_4471,N_4848);
nor U5962 (N_5962,N_4449,N_4256);
nand U5963 (N_5963,N_4376,N_4048);
nor U5964 (N_5964,N_4050,N_4270);
and U5965 (N_5965,N_4227,N_4484);
and U5966 (N_5966,N_4687,N_4815);
or U5967 (N_5967,N_4272,N_4739);
nor U5968 (N_5968,N_4263,N_4299);
or U5969 (N_5969,N_4421,N_4932);
nor U5970 (N_5970,N_4817,N_4882);
nor U5971 (N_5971,N_4875,N_4459);
nor U5972 (N_5972,N_4368,N_4869);
or U5973 (N_5973,N_4942,N_4222);
nor U5974 (N_5974,N_4130,N_4301);
nand U5975 (N_5975,N_4986,N_4772);
nand U5976 (N_5976,N_4057,N_4603);
and U5977 (N_5977,N_4721,N_4486);
nand U5978 (N_5978,N_4418,N_4343);
nor U5979 (N_5979,N_4578,N_4676);
and U5980 (N_5980,N_4637,N_4463);
nor U5981 (N_5981,N_4457,N_4102);
nand U5982 (N_5982,N_4899,N_4121);
and U5983 (N_5983,N_4984,N_4613);
or U5984 (N_5984,N_4384,N_4350);
nor U5985 (N_5985,N_4222,N_4268);
or U5986 (N_5986,N_4652,N_4133);
nand U5987 (N_5987,N_4942,N_4328);
nor U5988 (N_5988,N_4110,N_4605);
nor U5989 (N_5989,N_4727,N_4350);
nand U5990 (N_5990,N_4767,N_4362);
and U5991 (N_5991,N_4076,N_4579);
and U5992 (N_5992,N_4921,N_4223);
and U5993 (N_5993,N_4719,N_4833);
and U5994 (N_5994,N_4127,N_4097);
nand U5995 (N_5995,N_4085,N_4003);
or U5996 (N_5996,N_4323,N_4356);
or U5997 (N_5997,N_4301,N_4786);
and U5998 (N_5998,N_4606,N_4380);
and U5999 (N_5999,N_4318,N_4026);
nand U6000 (N_6000,N_5445,N_5259);
or U6001 (N_6001,N_5470,N_5262);
and U6002 (N_6002,N_5731,N_5324);
and U6003 (N_6003,N_5148,N_5986);
and U6004 (N_6004,N_5448,N_5431);
and U6005 (N_6005,N_5608,N_5564);
nor U6006 (N_6006,N_5839,N_5573);
and U6007 (N_6007,N_5648,N_5076);
and U6008 (N_6008,N_5131,N_5689);
and U6009 (N_6009,N_5124,N_5897);
nor U6010 (N_6010,N_5908,N_5070);
nand U6011 (N_6011,N_5949,N_5581);
nand U6012 (N_6012,N_5342,N_5900);
nand U6013 (N_6013,N_5368,N_5770);
nand U6014 (N_6014,N_5674,N_5275);
and U6015 (N_6015,N_5941,N_5746);
or U6016 (N_6016,N_5842,N_5354);
xor U6017 (N_6017,N_5576,N_5558);
nand U6018 (N_6018,N_5319,N_5232);
xnor U6019 (N_6019,N_5539,N_5025);
nor U6020 (N_6020,N_5910,N_5359);
nor U6021 (N_6021,N_5312,N_5433);
and U6022 (N_6022,N_5589,N_5379);
nand U6023 (N_6023,N_5765,N_5351);
or U6024 (N_6024,N_5384,N_5942);
and U6025 (N_6025,N_5236,N_5988);
nor U6026 (N_6026,N_5940,N_5929);
and U6027 (N_6027,N_5487,N_5622);
nand U6028 (N_6028,N_5420,N_5626);
nor U6029 (N_6029,N_5041,N_5902);
nand U6030 (N_6030,N_5550,N_5206);
nand U6031 (N_6031,N_5009,N_5017);
nor U6032 (N_6032,N_5584,N_5453);
nand U6033 (N_6033,N_5887,N_5611);
nand U6034 (N_6034,N_5752,N_5464);
and U6035 (N_6035,N_5185,N_5593);
nand U6036 (N_6036,N_5040,N_5273);
nor U6037 (N_6037,N_5653,N_5142);
or U6038 (N_6038,N_5775,N_5216);
nor U6039 (N_6039,N_5382,N_5679);
or U6040 (N_6040,N_5305,N_5754);
and U6041 (N_6041,N_5636,N_5526);
and U6042 (N_6042,N_5082,N_5256);
or U6043 (N_6043,N_5514,N_5792);
or U6044 (N_6044,N_5089,N_5184);
nand U6045 (N_6045,N_5187,N_5178);
nor U6046 (N_6046,N_5429,N_5906);
or U6047 (N_6047,N_5575,N_5660);
nor U6048 (N_6048,N_5771,N_5594);
nor U6049 (N_6049,N_5591,N_5747);
nor U6050 (N_6050,N_5323,N_5479);
or U6051 (N_6051,N_5534,N_5117);
and U6052 (N_6052,N_5779,N_5834);
or U6053 (N_6053,N_5450,N_5045);
nor U6054 (N_6054,N_5123,N_5046);
nor U6055 (N_6055,N_5716,N_5537);
and U6056 (N_6056,N_5592,N_5270);
and U6057 (N_6057,N_5953,N_5791);
nor U6058 (N_6058,N_5212,N_5952);
or U6059 (N_6059,N_5349,N_5203);
or U6060 (N_6060,N_5145,N_5451);
nand U6061 (N_6061,N_5794,N_5821);
or U6062 (N_6062,N_5449,N_5664);
and U6063 (N_6063,N_5296,N_5536);
nand U6064 (N_6064,N_5501,N_5582);
nand U6065 (N_6065,N_5700,N_5086);
nor U6066 (N_6066,N_5935,N_5238);
nand U6067 (N_6067,N_5036,N_5790);
nor U6068 (N_6068,N_5098,N_5859);
nand U6069 (N_6069,N_5743,N_5111);
and U6070 (N_6070,N_5641,N_5390);
nor U6071 (N_6071,N_5056,N_5924);
and U6072 (N_6072,N_5494,N_5866);
or U6073 (N_6073,N_5326,N_5353);
and U6074 (N_6074,N_5049,N_5201);
and U6075 (N_6075,N_5764,N_5288);
nand U6076 (N_6076,N_5901,N_5394);
nand U6077 (N_6077,N_5110,N_5960);
and U6078 (N_6078,N_5987,N_5402);
nor U6079 (N_6079,N_5345,N_5826);
and U6080 (N_6080,N_5852,N_5998);
nand U6081 (N_6081,N_5688,N_5886);
or U6082 (N_6082,N_5180,N_5217);
or U6083 (N_6083,N_5478,N_5297);
and U6084 (N_6084,N_5334,N_5175);
nor U6085 (N_6085,N_5726,N_5419);
nor U6086 (N_6086,N_5856,N_5512);
and U6087 (N_6087,N_5704,N_5029);
nand U6088 (N_6088,N_5410,N_5461);
nand U6089 (N_6089,N_5643,N_5515);
nand U6090 (N_6090,N_5965,N_5154);
and U6091 (N_6091,N_5223,N_5999);
nand U6092 (N_6092,N_5411,N_5915);
nor U6093 (N_6093,N_5918,N_5724);
and U6094 (N_6094,N_5804,N_5773);
and U6095 (N_6095,N_5244,N_5993);
and U6096 (N_6096,N_5605,N_5417);
and U6097 (N_6097,N_5369,N_5905);
and U6098 (N_6098,N_5427,N_5251);
and U6099 (N_6099,N_5899,N_5841);
or U6100 (N_6100,N_5613,N_5944);
nor U6101 (N_6101,N_5883,N_5248);
and U6102 (N_6102,N_5126,N_5090);
or U6103 (N_6103,N_5541,N_5545);
nor U6104 (N_6104,N_5492,N_5817);
nor U6105 (N_6105,N_5882,N_5308);
nand U6106 (N_6106,N_5454,N_5340);
nand U6107 (N_6107,N_5936,N_5970);
xor U6108 (N_6108,N_5559,N_5493);
xor U6109 (N_6109,N_5631,N_5426);
and U6110 (N_6110,N_5723,N_5188);
nor U6111 (N_6111,N_5759,N_5415);
and U6112 (N_6112,N_5022,N_5521);
nand U6113 (N_6113,N_5332,N_5809);
nand U6114 (N_6114,N_5051,N_5365);
or U6115 (N_6115,N_5511,N_5532);
nand U6116 (N_6116,N_5242,N_5985);
nand U6117 (N_6117,N_5624,N_5829);
nand U6118 (N_6118,N_5425,N_5371);
nand U6119 (N_6119,N_5566,N_5362);
nor U6120 (N_6120,N_5815,N_5416);
nand U6121 (N_6121,N_5037,N_5476);
nand U6122 (N_6122,N_5896,N_5447);
and U6123 (N_6123,N_5489,N_5661);
and U6124 (N_6124,N_5926,N_5604);
and U6125 (N_6125,N_5577,N_5781);
nor U6126 (N_6126,N_5586,N_5686);
nand U6127 (N_6127,N_5505,N_5128);
nor U6128 (N_6128,N_5615,N_5482);
and U6129 (N_6129,N_5498,N_5623);
nor U6130 (N_6130,N_5343,N_5705);
xor U6131 (N_6131,N_5682,N_5182);
nor U6132 (N_6132,N_5920,N_5260);
nand U6133 (N_6133,N_5300,N_5321);
and U6134 (N_6134,N_5278,N_5619);
nor U6135 (N_6135,N_5285,N_5233);
or U6136 (N_6136,N_5913,N_5093);
nor U6137 (N_6137,N_5435,N_5668);
and U6138 (N_6138,N_5655,N_5676);
and U6139 (N_6139,N_5540,N_5062);
and U6140 (N_6140,N_5782,N_5071);
or U6141 (N_6141,N_5956,N_5504);
or U6142 (N_6142,N_5745,N_5396);
or U6143 (N_6143,N_5838,N_5711);
or U6144 (N_6144,N_5143,N_5028);
and U6145 (N_6145,N_5799,N_5966);
nand U6146 (N_6146,N_5927,N_5120);
or U6147 (N_6147,N_5702,N_5292);
and U6148 (N_6148,N_5879,N_5614);
nand U6149 (N_6149,N_5397,N_5951);
xor U6150 (N_6150,N_5084,N_5921);
nor U6151 (N_6151,N_5173,N_5968);
and U6152 (N_6152,N_5833,N_5736);
nand U6153 (N_6153,N_5876,N_5717);
nand U6154 (N_6154,N_5789,N_5563);
or U6155 (N_6155,N_5508,N_5207);
or U6156 (N_6156,N_5346,N_5325);
and U6157 (N_6157,N_5116,N_5159);
and U6158 (N_6158,N_5347,N_5685);
nand U6159 (N_6159,N_5122,N_5950);
nor U6160 (N_6160,N_5165,N_5467);
nor U6161 (N_6161,N_5246,N_5818);
and U6162 (N_6162,N_5778,N_5691);
nor U6163 (N_6163,N_5979,N_5585);
nor U6164 (N_6164,N_5129,N_5708);
or U6165 (N_6165,N_5038,N_5665);
or U6166 (N_6166,N_5571,N_5113);
nand U6167 (N_6167,N_5058,N_5130);
or U6168 (N_6168,N_5831,N_5327);
nor U6169 (N_6169,N_5119,N_5205);
and U6170 (N_6170,N_5853,N_5072);
nand U6171 (N_6171,N_5083,N_5506);
nor U6172 (N_6172,N_5272,N_5339);
or U6173 (N_6173,N_5471,N_5567);
and U6174 (N_6174,N_5578,N_5599);
nand U6175 (N_6175,N_5336,N_5580);
and U6176 (N_6176,N_5398,N_5197);
and U6177 (N_6177,N_5224,N_5925);
nand U6178 (N_6178,N_5836,N_5301);
or U6179 (N_6179,N_5155,N_5463);
nor U6180 (N_6180,N_5307,N_5881);
or U6181 (N_6181,N_5500,N_5177);
and U6182 (N_6182,N_5280,N_5858);
xnor U6183 (N_6183,N_5277,N_5549);
xor U6184 (N_6184,N_5378,N_5135);
nor U6185 (N_6185,N_5065,N_5483);
or U6186 (N_6186,N_5452,N_5081);
nor U6187 (N_6187,N_5338,N_5517);
and U6188 (N_6188,N_5672,N_5257);
or U6189 (N_6189,N_5698,N_5245);
nand U6190 (N_6190,N_5769,N_5004);
nor U6191 (N_6191,N_5560,N_5255);
and U6192 (N_6192,N_5172,N_5048);
or U6193 (N_6193,N_5068,N_5847);
and U6194 (N_6194,N_5673,N_5687);
and U6195 (N_6195,N_5772,N_5074);
and U6196 (N_6196,N_5738,N_5033);
and U6197 (N_6197,N_5003,N_5010);
nand U6198 (N_6198,N_5218,N_5019);
nand U6199 (N_6199,N_5737,N_5706);
and U6200 (N_6200,N_5638,N_5803);
and U6201 (N_6201,N_5819,N_5957);
nor U6202 (N_6202,N_5432,N_5850);
nand U6203 (N_6203,N_5984,N_5796);
or U6204 (N_6204,N_5458,N_5335);
and U6205 (N_6205,N_5080,N_5392);
nand U6206 (N_6206,N_5042,N_5802);
xor U6207 (N_6207,N_5366,N_5097);
and U6208 (N_6208,N_5755,N_5488);
or U6209 (N_6209,N_5525,N_5055);
nor U6210 (N_6210,N_5034,N_5136);
or U6211 (N_6211,N_5917,N_5767);
nor U6212 (N_6212,N_5250,N_5800);
and U6213 (N_6213,N_5075,N_5663);
nor U6214 (N_6214,N_5945,N_5894);
nand U6215 (N_6215,N_5441,N_5027);
xor U6216 (N_6216,N_5228,N_5955);
nand U6217 (N_6217,N_5480,N_5108);
or U6218 (N_6218,N_5287,N_5712);
nand U6219 (N_6219,N_5215,N_5844);
nand U6220 (N_6220,N_5374,N_5720);
nand U6221 (N_6221,N_5403,N_5088);
nor U6222 (N_6222,N_5628,N_5587);
and U6223 (N_6223,N_5967,N_5104);
nor U6224 (N_6224,N_5995,N_5385);
nor U6225 (N_6225,N_5649,N_5780);
or U6226 (N_6226,N_5529,N_5372);
or U6227 (N_6227,N_5867,N_5138);
and U6228 (N_6228,N_5533,N_5404);
or U6229 (N_6229,N_5409,N_5472);
and U6230 (N_6230,N_5652,N_5981);
nand U6231 (N_6231,N_5570,N_5620);
or U6232 (N_6232,N_5520,N_5057);
nand U6233 (N_6233,N_5428,N_5199);
or U6234 (N_6234,N_5094,N_5118);
and U6235 (N_6235,N_5013,N_5391);
and U6236 (N_6236,N_5078,N_5364);
or U6237 (N_6237,N_5715,N_5721);
and U6238 (N_6238,N_5189,N_5101);
or U6239 (N_6239,N_5561,N_5141);
nor U6240 (N_6240,N_5934,N_5820);
nand U6241 (N_6241,N_5309,N_5741);
or U6242 (N_6242,N_5732,N_5888);
and U6243 (N_6243,N_5763,N_5024);
xnor U6244 (N_6244,N_5002,N_5825);
nor U6245 (N_6245,N_5837,N_5909);
or U6246 (N_6246,N_5827,N_5699);
and U6247 (N_6247,N_5583,N_5485);
and U6248 (N_6248,N_5174,N_5835);
or U6249 (N_6249,N_5510,N_5516);
and U6250 (N_6250,N_5171,N_5812);
or U6251 (N_6251,N_5760,N_5304);
or U6252 (N_6252,N_5210,N_5313);
nand U6253 (N_6253,N_5252,N_5121);
nor U6254 (N_6254,N_5279,N_5328);
nand U6255 (N_6255,N_5880,N_5161);
xnor U6256 (N_6256,N_5748,N_5061);
or U6257 (N_6257,N_5857,N_5787);
nand U6258 (N_6258,N_5658,N_5258);
and U6259 (N_6259,N_5437,N_5457);
nand U6260 (N_6260,N_5728,N_5241);
nor U6261 (N_6261,N_5133,N_5840);
nor U6262 (N_6262,N_5209,N_5310);
nor U6263 (N_6263,N_5314,N_5994);
nand U6264 (N_6264,N_5502,N_5848);
nand U6265 (N_6265,N_5635,N_5933);
and U6266 (N_6266,N_5612,N_5168);
nor U6267 (N_6267,N_5389,N_5295);
and U6268 (N_6268,N_5753,N_5127);
and U6269 (N_6269,N_5008,N_5430);
nand U6270 (N_6270,N_5793,N_5546);
nor U6271 (N_6271,N_5713,N_5317);
nor U6272 (N_6272,N_5481,N_5776);
nand U6273 (N_6273,N_5269,N_5509);
nand U6274 (N_6274,N_5522,N_5642);
or U6275 (N_6275,N_5647,N_5693);
and U6276 (N_6276,N_5337,N_5400);
nand U6277 (N_6277,N_5367,N_5361);
and U6278 (N_6278,N_5291,N_5616);
nor U6279 (N_6279,N_5650,N_5811);
nand U6280 (N_6280,N_5692,N_5109);
nand U6281 (N_6281,N_5873,N_5018);
or U6282 (N_6282,N_5456,N_5972);
nor U6283 (N_6283,N_5551,N_5609);
nand U6284 (N_6284,N_5446,N_5497);
nand U6285 (N_6285,N_5438,N_5229);
and U6286 (N_6286,N_5962,N_5633);
nor U6287 (N_6287,N_5376,N_5423);
or U6288 (N_6288,N_5595,N_5749);
nand U6289 (N_6289,N_5169,N_5610);
and U6290 (N_6290,N_5221,N_5077);
nor U6291 (N_6291,N_5315,N_5156);
and U6292 (N_6292,N_5158,N_5845);
or U6293 (N_6293,N_5484,N_5303);
nand U6294 (N_6294,N_5102,N_5200);
nor U6295 (N_6295,N_5703,N_5134);
and U6296 (N_6296,N_5087,N_5320);
nor U6297 (N_6297,N_5044,N_5322);
or U6298 (N_6298,N_5877,N_5271);
nand U6299 (N_6299,N_5667,N_5442);
and U6300 (N_6300,N_5606,N_5937);
nor U6301 (N_6301,N_5670,N_5196);
or U6302 (N_6302,N_5341,N_5634);
or U6303 (N_6303,N_5474,N_5629);
nor U6304 (N_6304,N_5878,N_5035);
nor U6305 (N_6305,N_5598,N_5542);
or U6306 (N_6306,N_5662,N_5299);
xor U6307 (N_6307,N_5774,N_5651);
nor U6308 (N_6308,N_5331,N_5192);
or U6309 (N_6309,N_5047,N_5434);
or U6310 (N_6310,N_5734,N_5152);
and U6311 (N_6311,N_5179,N_5290);
nand U6312 (N_6312,N_5729,N_5344);
nor U6313 (N_6313,N_5557,N_5399);
nor U6314 (N_6314,N_5459,N_5574);
nand U6315 (N_6315,N_5475,N_5473);
nor U6316 (N_6316,N_5701,N_5640);
nor U6317 (N_6317,N_5181,N_5973);
nand U6318 (N_6318,N_5235,N_5824);
nor U6319 (N_6319,N_5875,N_5601);
and U6320 (N_6320,N_5043,N_5054);
nor U6321 (N_6321,N_5418,N_5239);
or U6322 (N_6322,N_5766,N_5730);
nand U6323 (N_6323,N_5727,N_5719);
xor U6324 (N_6324,N_5751,N_5012);
and U6325 (N_6325,N_5243,N_5637);
and U6326 (N_6326,N_5978,N_5225);
and U6327 (N_6327,N_5617,N_5190);
nand U6328 (N_6328,N_5079,N_5067);
or U6329 (N_6329,N_5524,N_5455);
or U6330 (N_6330,N_5348,N_5193);
nor U6331 (N_6331,N_5247,N_5176);
nand U6332 (N_6332,N_5722,N_5026);
and U6333 (N_6333,N_5572,N_5414);
nor U6334 (N_6334,N_5535,N_5860);
or U6335 (N_6335,N_5100,N_5519);
nand U6336 (N_6336,N_5554,N_5618);
nand U6337 (N_6337,N_5132,N_5518);
and U6338 (N_6338,N_5961,N_5164);
and U6339 (N_6339,N_5096,N_5030);
and U6340 (N_6340,N_5370,N_5281);
nor U6341 (N_6341,N_5237,N_5646);
or U6342 (N_6342,N_5846,N_5816);
and U6343 (N_6343,N_5253,N_5191);
or U6344 (N_6344,N_5356,N_5408);
and U6345 (N_6345,N_5862,N_5675);
nor U6346 (N_6346,N_5666,N_5073);
xor U6347 (N_6347,N_5393,N_5115);
and U6348 (N_6348,N_5477,N_5264);
and U6349 (N_6349,N_5316,N_5632);
xnor U6350 (N_6350,N_5267,N_5625);
or U6351 (N_6351,N_5869,N_5007);
nand U6352 (N_6352,N_5997,N_5146);
and U6353 (N_6353,N_5690,N_5311);
nand U6354 (N_6354,N_5163,N_5263);
or U6355 (N_6355,N_5744,N_5865);
nor U6356 (N_6356,N_5680,N_5777);
nand U6357 (N_6357,N_5735,N_5219);
and U6358 (N_6358,N_5014,N_5740);
nor U6359 (N_6359,N_5671,N_5465);
nand U6360 (N_6360,N_5588,N_5996);
nor U6361 (N_6361,N_5932,N_5443);
and U6362 (N_6362,N_5709,N_5421);
and U6363 (N_6363,N_5870,N_5579);
nor U6364 (N_6364,N_5931,N_5496);
and U6365 (N_6365,N_5383,N_5565);
or U6366 (N_6366,N_5656,N_5405);
nand U6367 (N_6367,N_5553,N_5552);
nor U6368 (N_6368,N_5669,N_5783);
and U6369 (N_6369,N_5387,N_5202);
or U6370 (N_6370,N_5099,N_5293);
and U6371 (N_6371,N_5556,N_5329);
nor U6372 (N_6372,N_5460,N_5406);
nor U6373 (N_6373,N_5923,N_5137);
nand U6374 (N_6374,N_5964,N_5659);
and U6375 (N_6375,N_5360,N_5424);
and U6376 (N_6376,N_5851,N_5718);
and U6377 (N_6377,N_5639,N_5306);
and U6378 (N_6378,N_5801,N_5725);
nand U6379 (N_6379,N_5352,N_5021);
nor U6380 (N_6380,N_5644,N_5091);
and U6381 (N_6381,N_5469,N_5696);
and U6382 (N_6382,N_5654,N_5092);
nor U6383 (N_6383,N_5872,N_5627);
or U6384 (N_6384,N_5015,N_5555);
nand U6385 (N_6385,N_5948,N_5160);
nand U6386 (N_6386,N_5681,N_5756);
and U6387 (N_6387,N_5969,N_5903);
nor U6388 (N_6388,N_5381,N_5914);
nand U6389 (N_6389,N_5195,N_5375);
nor U6390 (N_6390,N_5885,N_5707);
and U6391 (N_6391,N_5889,N_5714);
nor U6392 (N_6392,N_5742,N_5147);
nor U6393 (N_6393,N_5095,N_5710);
nor U6394 (N_6394,N_5125,N_5600);
and U6395 (N_6395,N_5602,N_5513);
and U6396 (N_6396,N_5757,N_5788);
nand U6397 (N_6397,N_5153,N_5495);
nand U6398 (N_6398,N_5254,N_5211);
nand U6399 (N_6399,N_5060,N_5005);
nand U6400 (N_6400,N_5050,N_5330);
nor U6401 (N_6401,N_5294,N_5499);
nor U6402 (N_6402,N_5983,N_5758);
nand U6403 (N_6403,N_5198,N_5597);
or U6404 (N_6404,N_5543,N_5798);
nor U6405 (N_6405,N_5444,N_5982);
or U6406 (N_6406,N_5064,N_5892);
and U6407 (N_6407,N_5440,N_5805);
or U6408 (N_6408,N_5204,N_5170);
or U6409 (N_6409,N_5468,N_5874);
nor U6410 (N_6410,N_5466,N_5830);
or U6411 (N_6411,N_5603,N_5750);
nor U6412 (N_6412,N_5797,N_5286);
nand U6413 (N_6413,N_5808,N_5854);
xnor U6414 (N_6414,N_5388,N_5868);
nand U6415 (N_6415,N_5226,N_5208);
or U6416 (N_6416,N_5568,N_5943);
nor U6417 (N_6417,N_5971,N_5531);
nand U6418 (N_6418,N_5491,N_5462);
and U6419 (N_6419,N_5282,N_5318);
or U6420 (N_6420,N_5103,N_5490);
and U6421 (N_6421,N_5785,N_5106);
nand U6422 (N_6422,N_5144,N_5954);
and U6423 (N_6423,N_5363,N_5538);
or U6424 (N_6424,N_5938,N_5032);
and U6425 (N_6425,N_5001,N_5052);
or U6426 (N_6426,N_5380,N_5166);
nor U6427 (N_6427,N_5059,N_5544);
nor U6428 (N_6428,N_5507,N_5992);
or U6429 (N_6429,N_5140,N_5621);
xnor U6430 (N_6430,N_5283,N_5828);
and U6431 (N_6431,N_5039,N_5694);
nor U6432 (N_6432,N_5151,N_5063);
nand U6433 (N_6433,N_5884,N_5990);
nand U6434 (N_6434,N_5657,N_5768);
and U6435 (N_6435,N_5358,N_5503);
nand U6436 (N_6436,N_5395,N_5898);
nand U6437 (N_6437,N_5000,N_5864);
or U6438 (N_6438,N_5919,N_5107);
nor U6439 (N_6439,N_5523,N_5922);
or U6440 (N_6440,N_5486,N_5806);
or U6441 (N_6441,N_5861,N_5333);
nand U6442 (N_6442,N_5904,N_5183);
and U6443 (N_6443,N_5912,N_5810);
nor U6444 (N_6444,N_5413,N_5976);
or U6445 (N_6445,N_5112,N_5843);
and U6446 (N_6446,N_5907,N_5849);
nand U6447 (N_6447,N_5222,N_5020);
nor U6448 (N_6448,N_5373,N_5194);
and U6449 (N_6449,N_5016,N_5011);
or U6450 (N_6450,N_5157,N_5284);
xor U6451 (N_6451,N_5678,N_5234);
and U6452 (N_6452,N_5590,N_5871);
nand U6453 (N_6453,N_5268,N_5562);
nor U6454 (N_6454,N_5139,N_5249);
nor U6455 (N_6455,N_5814,N_5946);
nand U6456 (N_6456,N_5947,N_5911);
nand U6457 (N_6457,N_5377,N_5289);
nor U6458 (N_6458,N_5085,N_5930);
xor U6459 (N_6459,N_5053,N_5220);
xor U6460 (N_6460,N_5677,N_5213);
and U6461 (N_6461,N_5916,N_5066);
or U6462 (N_6462,N_5422,N_5527);
and U6463 (N_6463,N_5980,N_5963);
nor U6464 (N_6464,N_5162,N_5893);
nor U6465 (N_6465,N_5891,N_5031);
and U6466 (N_6466,N_5298,N_5214);
nand U6467 (N_6467,N_5928,N_5230);
or U6468 (N_6468,N_5350,N_5436);
and U6469 (N_6469,N_5784,N_5302);
nand U6470 (N_6470,N_5528,N_5974);
nor U6471 (N_6471,N_5240,N_5683);
xor U6472 (N_6472,N_5813,N_5547);
nand U6473 (N_6473,N_5786,N_5975);
or U6474 (N_6474,N_5939,N_5733);
and U6475 (N_6475,N_5167,N_5977);
and U6476 (N_6476,N_5261,N_5989);
and U6477 (N_6477,N_5991,N_5006);
or U6478 (N_6478,N_5863,N_5761);
nand U6479 (N_6479,N_5265,N_5231);
nand U6480 (N_6480,N_5274,N_5276);
nor U6481 (N_6481,N_5890,N_5114);
nand U6482 (N_6482,N_5959,N_5823);
nand U6483 (N_6483,N_5407,N_5596);
nand U6484 (N_6484,N_5355,N_5069);
and U6485 (N_6485,N_5684,N_5412);
nand U6486 (N_6486,N_5386,N_5832);
and U6487 (N_6487,N_5645,N_5855);
nand U6488 (N_6488,N_5630,N_5807);
xor U6489 (N_6489,N_5607,N_5227);
nand U6490 (N_6490,N_5548,N_5795);
or U6491 (N_6491,N_5401,N_5149);
and U6492 (N_6492,N_5150,N_5695);
nand U6493 (N_6493,N_5186,N_5697);
or U6494 (N_6494,N_5895,N_5266);
and U6495 (N_6495,N_5958,N_5569);
nand U6496 (N_6496,N_5762,N_5439);
nor U6497 (N_6497,N_5357,N_5822);
nor U6498 (N_6498,N_5105,N_5530);
nor U6499 (N_6499,N_5739,N_5023);
or U6500 (N_6500,N_5136,N_5087);
or U6501 (N_6501,N_5287,N_5139);
and U6502 (N_6502,N_5936,N_5043);
nor U6503 (N_6503,N_5611,N_5759);
nand U6504 (N_6504,N_5520,N_5778);
nor U6505 (N_6505,N_5468,N_5419);
nand U6506 (N_6506,N_5148,N_5746);
nand U6507 (N_6507,N_5621,N_5496);
nand U6508 (N_6508,N_5542,N_5931);
nand U6509 (N_6509,N_5055,N_5693);
and U6510 (N_6510,N_5138,N_5648);
nor U6511 (N_6511,N_5913,N_5697);
nor U6512 (N_6512,N_5762,N_5704);
and U6513 (N_6513,N_5763,N_5348);
or U6514 (N_6514,N_5805,N_5015);
xor U6515 (N_6515,N_5771,N_5587);
and U6516 (N_6516,N_5039,N_5456);
nor U6517 (N_6517,N_5685,N_5539);
or U6518 (N_6518,N_5329,N_5170);
xor U6519 (N_6519,N_5573,N_5619);
and U6520 (N_6520,N_5505,N_5981);
nor U6521 (N_6521,N_5410,N_5214);
or U6522 (N_6522,N_5760,N_5839);
and U6523 (N_6523,N_5519,N_5275);
nor U6524 (N_6524,N_5814,N_5197);
xor U6525 (N_6525,N_5714,N_5702);
or U6526 (N_6526,N_5765,N_5803);
and U6527 (N_6527,N_5493,N_5383);
or U6528 (N_6528,N_5818,N_5201);
or U6529 (N_6529,N_5819,N_5075);
nor U6530 (N_6530,N_5823,N_5789);
xnor U6531 (N_6531,N_5440,N_5281);
and U6532 (N_6532,N_5130,N_5265);
and U6533 (N_6533,N_5145,N_5634);
nor U6534 (N_6534,N_5156,N_5186);
nor U6535 (N_6535,N_5058,N_5932);
and U6536 (N_6536,N_5087,N_5109);
nor U6537 (N_6537,N_5382,N_5415);
or U6538 (N_6538,N_5766,N_5639);
or U6539 (N_6539,N_5515,N_5560);
nor U6540 (N_6540,N_5122,N_5395);
and U6541 (N_6541,N_5591,N_5806);
nor U6542 (N_6542,N_5061,N_5122);
nor U6543 (N_6543,N_5661,N_5653);
or U6544 (N_6544,N_5654,N_5530);
nor U6545 (N_6545,N_5731,N_5135);
nand U6546 (N_6546,N_5510,N_5863);
or U6547 (N_6547,N_5202,N_5643);
nor U6548 (N_6548,N_5391,N_5170);
and U6549 (N_6549,N_5460,N_5242);
or U6550 (N_6550,N_5778,N_5522);
xnor U6551 (N_6551,N_5669,N_5672);
nor U6552 (N_6552,N_5014,N_5728);
nand U6553 (N_6553,N_5189,N_5379);
and U6554 (N_6554,N_5607,N_5256);
nor U6555 (N_6555,N_5296,N_5061);
or U6556 (N_6556,N_5831,N_5267);
and U6557 (N_6557,N_5030,N_5352);
nand U6558 (N_6558,N_5808,N_5765);
and U6559 (N_6559,N_5270,N_5881);
nor U6560 (N_6560,N_5022,N_5553);
and U6561 (N_6561,N_5883,N_5060);
and U6562 (N_6562,N_5274,N_5642);
nor U6563 (N_6563,N_5587,N_5699);
nand U6564 (N_6564,N_5956,N_5594);
or U6565 (N_6565,N_5869,N_5673);
nor U6566 (N_6566,N_5601,N_5531);
nor U6567 (N_6567,N_5700,N_5313);
and U6568 (N_6568,N_5547,N_5212);
and U6569 (N_6569,N_5657,N_5339);
nand U6570 (N_6570,N_5061,N_5046);
nand U6571 (N_6571,N_5479,N_5449);
nor U6572 (N_6572,N_5940,N_5320);
or U6573 (N_6573,N_5546,N_5082);
xnor U6574 (N_6574,N_5618,N_5251);
nand U6575 (N_6575,N_5871,N_5683);
and U6576 (N_6576,N_5312,N_5210);
nor U6577 (N_6577,N_5257,N_5393);
or U6578 (N_6578,N_5771,N_5297);
or U6579 (N_6579,N_5251,N_5848);
and U6580 (N_6580,N_5092,N_5959);
nor U6581 (N_6581,N_5192,N_5156);
and U6582 (N_6582,N_5085,N_5346);
nor U6583 (N_6583,N_5084,N_5448);
xnor U6584 (N_6584,N_5318,N_5846);
or U6585 (N_6585,N_5549,N_5314);
nand U6586 (N_6586,N_5951,N_5579);
and U6587 (N_6587,N_5598,N_5733);
nand U6588 (N_6588,N_5043,N_5562);
nor U6589 (N_6589,N_5446,N_5244);
or U6590 (N_6590,N_5182,N_5885);
nand U6591 (N_6591,N_5282,N_5502);
and U6592 (N_6592,N_5886,N_5231);
nor U6593 (N_6593,N_5002,N_5994);
nor U6594 (N_6594,N_5960,N_5209);
or U6595 (N_6595,N_5823,N_5658);
or U6596 (N_6596,N_5751,N_5990);
nand U6597 (N_6597,N_5217,N_5617);
and U6598 (N_6598,N_5545,N_5503);
or U6599 (N_6599,N_5574,N_5618);
nand U6600 (N_6600,N_5965,N_5726);
xor U6601 (N_6601,N_5447,N_5609);
and U6602 (N_6602,N_5712,N_5995);
and U6603 (N_6603,N_5755,N_5376);
or U6604 (N_6604,N_5450,N_5642);
and U6605 (N_6605,N_5976,N_5627);
nand U6606 (N_6606,N_5927,N_5254);
nor U6607 (N_6607,N_5383,N_5618);
and U6608 (N_6608,N_5613,N_5000);
nor U6609 (N_6609,N_5985,N_5357);
or U6610 (N_6610,N_5892,N_5862);
or U6611 (N_6611,N_5734,N_5519);
nand U6612 (N_6612,N_5626,N_5410);
xor U6613 (N_6613,N_5646,N_5748);
nand U6614 (N_6614,N_5991,N_5321);
nand U6615 (N_6615,N_5176,N_5000);
or U6616 (N_6616,N_5463,N_5077);
nand U6617 (N_6617,N_5285,N_5068);
nor U6618 (N_6618,N_5742,N_5838);
nand U6619 (N_6619,N_5681,N_5511);
and U6620 (N_6620,N_5223,N_5254);
nand U6621 (N_6621,N_5098,N_5496);
nor U6622 (N_6622,N_5871,N_5048);
nor U6623 (N_6623,N_5834,N_5899);
and U6624 (N_6624,N_5085,N_5125);
nor U6625 (N_6625,N_5452,N_5852);
or U6626 (N_6626,N_5779,N_5150);
and U6627 (N_6627,N_5979,N_5605);
nand U6628 (N_6628,N_5287,N_5900);
nor U6629 (N_6629,N_5497,N_5646);
and U6630 (N_6630,N_5774,N_5805);
nor U6631 (N_6631,N_5467,N_5355);
and U6632 (N_6632,N_5364,N_5359);
and U6633 (N_6633,N_5371,N_5318);
and U6634 (N_6634,N_5598,N_5718);
and U6635 (N_6635,N_5037,N_5684);
nand U6636 (N_6636,N_5834,N_5393);
or U6637 (N_6637,N_5591,N_5617);
nand U6638 (N_6638,N_5785,N_5161);
nor U6639 (N_6639,N_5823,N_5075);
or U6640 (N_6640,N_5630,N_5174);
and U6641 (N_6641,N_5484,N_5643);
or U6642 (N_6642,N_5194,N_5575);
nand U6643 (N_6643,N_5069,N_5461);
and U6644 (N_6644,N_5376,N_5790);
nor U6645 (N_6645,N_5003,N_5898);
nand U6646 (N_6646,N_5578,N_5162);
and U6647 (N_6647,N_5157,N_5378);
xnor U6648 (N_6648,N_5245,N_5221);
nand U6649 (N_6649,N_5026,N_5322);
nand U6650 (N_6650,N_5004,N_5068);
or U6651 (N_6651,N_5559,N_5142);
or U6652 (N_6652,N_5590,N_5369);
nand U6653 (N_6653,N_5390,N_5630);
and U6654 (N_6654,N_5329,N_5186);
and U6655 (N_6655,N_5479,N_5547);
nor U6656 (N_6656,N_5703,N_5466);
and U6657 (N_6657,N_5261,N_5707);
nand U6658 (N_6658,N_5313,N_5247);
nand U6659 (N_6659,N_5420,N_5270);
and U6660 (N_6660,N_5474,N_5770);
xor U6661 (N_6661,N_5554,N_5230);
nand U6662 (N_6662,N_5421,N_5711);
or U6663 (N_6663,N_5506,N_5801);
nand U6664 (N_6664,N_5914,N_5221);
or U6665 (N_6665,N_5061,N_5853);
and U6666 (N_6666,N_5215,N_5576);
and U6667 (N_6667,N_5102,N_5318);
or U6668 (N_6668,N_5926,N_5216);
nor U6669 (N_6669,N_5831,N_5837);
or U6670 (N_6670,N_5571,N_5448);
nor U6671 (N_6671,N_5321,N_5207);
and U6672 (N_6672,N_5169,N_5285);
and U6673 (N_6673,N_5209,N_5828);
or U6674 (N_6674,N_5801,N_5628);
or U6675 (N_6675,N_5398,N_5790);
or U6676 (N_6676,N_5561,N_5893);
or U6677 (N_6677,N_5840,N_5428);
nor U6678 (N_6678,N_5487,N_5263);
nor U6679 (N_6679,N_5523,N_5007);
nand U6680 (N_6680,N_5372,N_5135);
and U6681 (N_6681,N_5471,N_5873);
nand U6682 (N_6682,N_5852,N_5670);
nand U6683 (N_6683,N_5971,N_5783);
or U6684 (N_6684,N_5654,N_5301);
nand U6685 (N_6685,N_5190,N_5883);
nand U6686 (N_6686,N_5217,N_5686);
or U6687 (N_6687,N_5128,N_5845);
or U6688 (N_6688,N_5916,N_5096);
or U6689 (N_6689,N_5793,N_5970);
or U6690 (N_6690,N_5483,N_5449);
or U6691 (N_6691,N_5931,N_5111);
nor U6692 (N_6692,N_5174,N_5260);
nand U6693 (N_6693,N_5574,N_5748);
xor U6694 (N_6694,N_5691,N_5190);
nor U6695 (N_6695,N_5582,N_5994);
and U6696 (N_6696,N_5229,N_5770);
or U6697 (N_6697,N_5630,N_5001);
or U6698 (N_6698,N_5478,N_5422);
nand U6699 (N_6699,N_5786,N_5373);
nor U6700 (N_6700,N_5469,N_5552);
nor U6701 (N_6701,N_5097,N_5358);
nor U6702 (N_6702,N_5669,N_5448);
or U6703 (N_6703,N_5668,N_5346);
nor U6704 (N_6704,N_5000,N_5132);
or U6705 (N_6705,N_5283,N_5096);
nand U6706 (N_6706,N_5791,N_5525);
and U6707 (N_6707,N_5340,N_5997);
or U6708 (N_6708,N_5191,N_5972);
or U6709 (N_6709,N_5667,N_5730);
nand U6710 (N_6710,N_5693,N_5493);
or U6711 (N_6711,N_5617,N_5431);
and U6712 (N_6712,N_5241,N_5442);
nand U6713 (N_6713,N_5755,N_5656);
nand U6714 (N_6714,N_5960,N_5046);
nor U6715 (N_6715,N_5646,N_5157);
nand U6716 (N_6716,N_5840,N_5450);
and U6717 (N_6717,N_5988,N_5451);
nand U6718 (N_6718,N_5174,N_5532);
and U6719 (N_6719,N_5288,N_5987);
and U6720 (N_6720,N_5342,N_5430);
or U6721 (N_6721,N_5433,N_5220);
nor U6722 (N_6722,N_5914,N_5670);
and U6723 (N_6723,N_5125,N_5348);
nand U6724 (N_6724,N_5980,N_5760);
and U6725 (N_6725,N_5685,N_5789);
nand U6726 (N_6726,N_5049,N_5060);
or U6727 (N_6727,N_5505,N_5486);
nand U6728 (N_6728,N_5498,N_5508);
nor U6729 (N_6729,N_5473,N_5404);
nor U6730 (N_6730,N_5930,N_5608);
and U6731 (N_6731,N_5930,N_5071);
and U6732 (N_6732,N_5019,N_5005);
nand U6733 (N_6733,N_5297,N_5981);
or U6734 (N_6734,N_5518,N_5492);
nor U6735 (N_6735,N_5721,N_5474);
nand U6736 (N_6736,N_5899,N_5496);
or U6737 (N_6737,N_5188,N_5633);
or U6738 (N_6738,N_5850,N_5283);
and U6739 (N_6739,N_5348,N_5204);
nor U6740 (N_6740,N_5828,N_5043);
nor U6741 (N_6741,N_5470,N_5577);
or U6742 (N_6742,N_5426,N_5630);
nand U6743 (N_6743,N_5415,N_5947);
nor U6744 (N_6744,N_5728,N_5029);
nand U6745 (N_6745,N_5780,N_5526);
or U6746 (N_6746,N_5443,N_5221);
and U6747 (N_6747,N_5161,N_5989);
nand U6748 (N_6748,N_5820,N_5275);
and U6749 (N_6749,N_5929,N_5568);
xnor U6750 (N_6750,N_5238,N_5961);
nor U6751 (N_6751,N_5798,N_5049);
and U6752 (N_6752,N_5189,N_5050);
nor U6753 (N_6753,N_5692,N_5581);
nand U6754 (N_6754,N_5279,N_5472);
nand U6755 (N_6755,N_5236,N_5484);
nand U6756 (N_6756,N_5331,N_5099);
nand U6757 (N_6757,N_5662,N_5645);
or U6758 (N_6758,N_5926,N_5698);
nor U6759 (N_6759,N_5398,N_5734);
nor U6760 (N_6760,N_5745,N_5408);
nand U6761 (N_6761,N_5292,N_5440);
nor U6762 (N_6762,N_5537,N_5810);
nor U6763 (N_6763,N_5893,N_5716);
or U6764 (N_6764,N_5410,N_5968);
or U6765 (N_6765,N_5305,N_5814);
nor U6766 (N_6766,N_5431,N_5782);
nor U6767 (N_6767,N_5126,N_5658);
and U6768 (N_6768,N_5602,N_5774);
nor U6769 (N_6769,N_5988,N_5943);
xor U6770 (N_6770,N_5418,N_5154);
nand U6771 (N_6771,N_5493,N_5675);
nor U6772 (N_6772,N_5603,N_5525);
or U6773 (N_6773,N_5181,N_5295);
nor U6774 (N_6774,N_5516,N_5171);
or U6775 (N_6775,N_5707,N_5753);
and U6776 (N_6776,N_5596,N_5648);
nor U6777 (N_6777,N_5942,N_5113);
or U6778 (N_6778,N_5949,N_5894);
nor U6779 (N_6779,N_5765,N_5605);
nand U6780 (N_6780,N_5791,N_5492);
and U6781 (N_6781,N_5430,N_5252);
or U6782 (N_6782,N_5772,N_5661);
nor U6783 (N_6783,N_5295,N_5200);
and U6784 (N_6784,N_5770,N_5710);
and U6785 (N_6785,N_5582,N_5977);
nand U6786 (N_6786,N_5429,N_5247);
nor U6787 (N_6787,N_5127,N_5782);
and U6788 (N_6788,N_5072,N_5366);
nor U6789 (N_6789,N_5515,N_5460);
and U6790 (N_6790,N_5588,N_5624);
xor U6791 (N_6791,N_5519,N_5295);
nand U6792 (N_6792,N_5496,N_5176);
nand U6793 (N_6793,N_5762,N_5349);
or U6794 (N_6794,N_5828,N_5505);
nand U6795 (N_6795,N_5552,N_5291);
or U6796 (N_6796,N_5620,N_5769);
nand U6797 (N_6797,N_5975,N_5448);
and U6798 (N_6798,N_5454,N_5956);
nand U6799 (N_6799,N_5653,N_5855);
or U6800 (N_6800,N_5695,N_5968);
and U6801 (N_6801,N_5130,N_5698);
nor U6802 (N_6802,N_5892,N_5058);
and U6803 (N_6803,N_5039,N_5113);
nor U6804 (N_6804,N_5030,N_5450);
or U6805 (N_6805,N_5915,N_5967);
and U6806 (N_6806,N_5235,N_5505);
nand U6807 (N_6807,N_5193,N_5591);
nand U6808 (N_6808,N_5114,N_5716);
nand U6809 (N_6809,N_5640,N_5309);
nor U6810 (N_6810,N_5135,N_5516);
nor U6811 (N_6811,N_5241,N_5501);
or U6812 (N_6812,N_5110,N_5996);
nor U6813 (N_6813,N_5147,N_5081);
and U6814 (N_6814,N_5182,N_5782);
or U6815 (N_6815,N_5274,N_5914);
and U6816 (N_6816,N_5992,N_5236);
nand U6817 (N_6817,N_5168,N_5359);
or U6818 (N_6818,N_5029,N_5523);
nor U6819 (N_6819,N_5845,N_5794);
or U6820 (N_6820,N_5204,N_5360);
and U6821 (N_6821,N_5490,N_5982);
nor U6822 (N_6822,N_5489,N_5790);
or U6823 (N_6823,N_5804,N_5562);
nand U6824 (N_6824,N_5881,N_5692);
nor U6825 (N_6825,N_5911,N_5254);
or U6826 (N_6826,N_5668,N_5761);
and U6827 (N_6827,N_5851,N_5168);
nand U6828 (N_6828,N_5859,N_5122);
nor U6829 (N_6829,N_5604,N_5294);
or U6830 (N_6830,N_5015,N_5512);
nor U6831 (N_6831,N_5137,N_5801);
nand U6832 (N_6832,N_5083,N_5144);
nor U6833 (N_6833,N_5224,N_5143);
or U6834 (N_6834,N_5522,N_5010);
and U6835 (N_6835,N_5717,N_5092);
nor U6836 (N_6836,N_5995,N_5750);
nor U6837 (N_6837,N_5334,N_5458);
or U6838 (N_6838,N_5593,N_5658);
nor U6839 (N_6839,N_5075,N_5427);
and U6840 (N_6840,N_5463,N_5037);
or U6841 (N_6841,N_5808,N_5344);
nand U6842 (N_6842,N_5298,N_5363);
nor U6843 (N_6843,N_5596,N_5385);
nor U6844 (N_6844,N_5872,N_5601);
nand U6845 (N_6845,N_5759,N_5273);
or U6846 (N_6846,N_5743,N_5954);
nor U6847 (N_6847,N_5366,N_5021);
or U6848 (N_6848,N_5714,N_5603);
or U6849 (N_6849,N_5973,N_5406);
and U6850 (N_6850,N_5053,N_5173);
xnor U6851 (N_6851,N_5230,N_5046);
xnor U6852 (N_6852,N_5987,N_5341);
and U6853 (N_6853,N_5315,N_5312);
and U6854 (N_6854,N_5367,N_5001);
and U6855 (N_6855,N_5203,N_5544);
nand U6856 (N_6856,N_5892,N_5122);
nand U6857 (N_6857,N_5915,N_5020);
nor U6858 (N_6858,N_5017,N_5914);
or U6859 (N_6859,N_5675,N_5075);
nor U6860 (N_6860,N_5021,N_5495);
nand U6861 (N_6861,N_5558,N_5923);
nor U6862 (N_6862,N_5932,N_5153);
or U6863 (N_6863,N_5008,N_5496);
nand U6864 (N_6864,N_5743,N_5391);
or U6865 (N_6865,N_5583,N_5283);
nand U6866 (N_6866,N_5878,N_5210);
and U6867 (N_6867,N_5317,N_5262);
nor U6868 (N_6868,N_5802,N_5017);
nand U6869 (N_6869,N_5317,N_5839);
or U6870 (N_6870,N_5438,N_5828);
or U6871 (N_6871,N_5001,N_5063);
nor U6872 (N_6872,N_5402,N_5671);
nor U6873 (N_6873,N_5207,N_5841);
and U6874 (N_6874,N_5341,N_5852);
nand U6875 (N_6875,N_5078,N_5173);
or U6876 (N_6876,N_5517,N_5566);
xnor U6877 (N_6877,N_5540,N_5689);
or U6878 (N_6878,N_5449,N_5892);
and U6879 (N_6879,N_5759,N_5249);
nand U6880 (N_6880,N_5811,N_5046);
or U6881 (N_6881,N_5467,N_5821);
nand U6882 (N_6882,N_5070,N_5331);
and U6883 (N_6883,N_5363,N_5573);
and U6884 (N_6884,N_5859,N_5887);
or U6885 (N_6885,N_5261,N_5746);
or U6886 (N_6886,N_5064,N_5967);
nor U6887 (N_6887,N_5553,N_5694);
or U6888 (N_6888,N_5619,N_5225);
nor U6889 (N_6889,N_5425,N_5507);
nor U6890 (N_6890,N_5310,N_5115);
and U6891 (N_6891,N_5633,N_5470);
or U6892 (N_6892,N_5361,N_5748);
and U6893 (N_6893,N_5491,N_5939);
nand U6894 (N_6894,N_5558,N_5491);
nand U6895 (N_6895,N_5986,N_5726);
nand U6896 (N_6896,N_5646,N_5033);
or U6897 (N_6897,N_5180,N_5982);
and U6898 (N_6898,N_5640,N_5885);
nor U6899 (N_6899,N_5407,N_5183);
and U6900 (N_6900,N_5819,N_5710);
and U6901 (N_6901,N_5974,N_5437);
and U6902 (N_6902,N_5068,N_5933);
and U6903 (N_6903,N_5539,N_5549);
nand U6904 (N_6904,N_5965,N_5271);
and U6905 (N_6905,N_5193,N_5873);
or U6906 (N_6906,N_5480,N_5940);
nand U6907 (N_6907,N_5740,N_5038);
and U6908 (N_6908,N_5147,N_5837);
nor U6909 (N_6909,N_5637,N_5635);
nor U6910 (N_6910,N_5666,N_5985);
and U6911 (N_6911,N_5541,N_5088);
or U6912 (N_6912,N_5495,N_5208);
nor U6913 (N_6913,N_5015,N_5850);
nand U6914 (N_6914,N_5705,N_5461);
nand U6915 (N_6915,N_5625,N_5793);
and U6916 (N_6916,N_5893,N_5273);
nor U6917 (N_6917,N_5063,N_5137);
xnor U6918 (N_6918,N_5663,N_5296);
nor U6919 (N_6919,N_5597,N_5980);
nor U6920 (N_6920,N_5502,N_5793);
nor U6921 (N_6921,N_5502,N_5924);
nor U6922 (N_6922,N_5641,N_5816);
xnor U6923 (N_6923,N_5672,N_5046);
nand U6924 (N_6924,N_5230,N_5140);
nand U6925 (N_6925,N_5442,N_5078);
nand U6926 (N_6926,N_5776,N_5939);
nor U6927 (N_6927,N_5420,N_5384);
nand U6928 (N_6928,N_5218,N_5486);
xor U6929 (N_6929,N_5087,N_5734);
nand U6930 (N_6930,N_5804,N_5097);
nor U6931 (N_6931,N_5433,N_5496);
and U6932 (N_6932,N_5188,N_5282);
or U6933 (N_6933,N_5588,N_5435);
nand U6934 (N_6934,N_5398,N_5769);
or U6935 (N_6935,N_5543,N_5686);
nand U6936 (N_6936,N_5038,N_5272);
or U6937 (N_6937,N_5932,N_5597);
or U6938 (N_6938,N_5153,N_5081);
xor U6939 (N_6939,N_5693,N_5762);
nand U6940 (N_6940,N_5875,N_5342);
nand U6941 (N_6941,N_5195,N_5151);
or U6942 (N_6942,N_5015,N_5030);
nor U6943 (N_6943,N_5225,N_5397);
nor U6944 (N_6944,N_5747,N_5300);
or U6945 (N_6945,N_5029,N_5629);
nor U6946 (N_6946,N_5750,N_5551);
and U6947 (N_6947,N_5033,N_5258);
and U6948 (N_6948,N_5090,N_5312);
and U6949 (N_6949,N_5322,N_5919);
and U6950 (N_6950,N_5533,N_5381);
or U6951 (N_6951,N_5514,N_5660);
and U6952 (N_6952,N_5667,N_5301);
nand U6953 (N_6953,N_5218,N_5738);
nor U6954 (N_6954,N_5514,N_5067);
and U6955 (N_6955,N_5957,N_5878);
and U6956 (N_6956,N_5789,N_5835);
nor U6957 (N_6957,N_5589,N_5177);
or U6958 (N_6958,N_5441,N_5974);
nand U6959 (N_6959,N_5583,N_5319);
and U6960 (N_6960,N_5503,N_5105);
nor U6961 (N_6961,N_5357,N_5352);
nor U6962 (N_6962,N_5087,N_5824);
nor U6963 (N_6963,N_5621,N_5545);
or U6964 (N_6964,N_5927,N_5390);
nor U6965 (N_6965,N_5613,N_5770);
nor U6966 (N_6966,N_5285,N_5074);
and U6967 (N_6967,N_5833,N_5349);
nor U6968 (N_6968,N_5736,N_5091);
nand U6969 (N_6969,N_5008,N_5801);
and U6970 (N_6970,N_5436,N_5006);
nand U6971 (N_6971,N_5461,N_5036);
or U6972 (N_6972,N_5060,N_5429);
nand U6973 (N_6973,N_5498,N_5963);
nand U6974 (N_6974,N_5554,N_5528);
and U6975 (N_6975,N_5564,N_5817);
or U6976 (N_6976,N_5633,N_5408);
nor U6977 (N_6977,N_5749,N_5438);
nand U6978 (N_6978,N_5919,N_5272);
nor U6979 (N_6979,N_5193,N_5316);
nor U6980 (N_6980,N_5998,N_5975);
nand U6981 (N_6981,N_5385,N_5789);
nand U6982 (N_6982,N_5036,N_5622);
nand U6983 (N_6983,N_5092,N_5963);
nor U6984 (N_6984,N_5887,N_5685);
and U6985 (N_6985,N_5852,N_5303);
and U6986 (N_6986,N_5545,N_5079);
nor U6987 (N_6987,N_5553,N_5596);
nand U6988 (N_6988,N_5512,N_5597);
or U6989 (N_6989,N_5364,N_5628);
or U6990 (N_6990,N_5738,N_5481);
nand U6991 (N_6991,N_5946,N_5787);
or U6992 (N_6992,N_5218,N_5542);
or U6993 (N_6993,N_5408,N_5121);
nor U6994 (N_6994,N_5539,N_5405);
nand U6995 (N_6995,N_5775,N_5608);
or U6996 (N_6996,N_5866,N_5759);
and U6997 (N_6997,N_5818,N_5609);
nand U6998 (N_6998,N_5220,N_5706);
nand U6999 (N_6999,N_5528,N_5045);
or U7000 (N_7000,N_6290,N_6682);
xor U7001 (N_7001,N_6973,N_6007);
or U7002 (N_7002,N_6302,N_6338);
or U7003 (N_7003,N_6035,N_6868);
nand U7004 (N_7004,N_6760,N_6714);
nor U7005 (N_7005,N_6529,N_6228);
nor U7006 (N_7006,N_6762,N_6523);
nor U7007 (N_7007,N_6698,N_6309);
nor U7008 (N_7008,N_6721,N_6586);
and U7009 (N_7009,N_6447,N_6713);
xor U7010 (N_7010,N_6872,N_6498);
or U7011 (N_7011,N_6922,N_6083);
nor U7012 (N_7012,N_6568,N_6364);
nor U7013 (N_7013,N_6237,N_6177);
nand U7014 (N_7014,N_6494,N_6268);
or U7015 (N_7015,N_6927,N_6312);
or U7016 (N_7016,N_6640,N_6335);
nand U7017 (N_7017,N_6340,N_6054);
xnor U7018 (N_7018,N_6984,N_6960);
nor U7019 (N_7019,N_6056,N_6088);
nand U7020 (N_7020,N_6019,N_6047);
nor U7021 (N_7021,N_6604,N_6483);
nand U7022 (N_7022,N_6784,N_6883);
or U7023 (N_7023,N_6358,N_6427);
nor U7024 (N_7024,N_6255,N_6296);
nand U7025 (N_7025,N_6457,N_6856);
nor U7026 (N_7026,N_6365,N_6459);
nand U7027 (N_7027,N_6754,N_6172);
or U7028 (N_7028,N_6025,N_6802);
or U7029 (N_7029,N_6272,N_6072);
or U7030 (N_7030,N_6474,N_6890);
nand U7031 (N_7031,N_6432,N_6077);
or U7032 (N_7032,N_6398,N_6433);
or U7033 (N_7033,N_6169,N_6504);
nand U7034 (N_7034,N_6545,N_6234);
nor U7035 (N_7035,N_6672,N_6435);
nand U7036 (N_7036,N_6751,N_6059);
nand U7037 (N_7037,N_6253,N_6493);
nand U7038 (N_7038,N_6310,N_6111);
or U7039 (N_7039,N_6330,N_6264);
nand U7040 (N_7040,N_6082,N_6178);
nor U7041 (N_7041,N_6099,N_6933);
nand U7042 (N_7042,N_6243,N_6384);
nand U7043 (N_7043,N_6598,N_6185);
and U7044 (N_7044,N_6959,N_6674);
nand U7045 (N_7045,N_6909,N_6858);
nand U7046 (N_7046,N_6133,N_6347);
or U7047 (N_7047,N_6569,N_6775);
and U7048 (N_7048,N_6198,N_6859);
nor U7049 (N_7049,N_6747,N_6192);
or U7050 (N_7050,N_6334,N_6295);
or U7051 (N_7051,N_6084,N_6062);
or U7052 (N_7052,N_6900,N_6438);
nand U7053 (N_7053,N_6375,N_6625);
or U7054 (N_7054,N_6102,N_6526);
nand U7055 (N_7055,N_6009,N_6583);
nor U7056 (N_7056,N_6824,N_6894);
nand U7057 (N_7057,N_6490,N_6506);
nor U7058 (N_7058,N_6739,N_6238);
or U7059 (N_7059,N_6124,N_6594);
nor U7060 (N_7060,N_6120,N_6694);
or U7061 (N_7061,N_6817,N_6143);
nand U7062 (N_7062,N_6336,N_6635);
nor U7063 (N_7063,N_6241,N_6910);
and U7064 (N_7064,N_6857,N_6259);
nand U7065 (N_7065,N_6434,N_6027);
nor U7066 (N_7066,N_6053,N_6738);
nor U7067 (N_7067,N_6578,N_6958);
and U7068 (N_7068,N_6285,N_6566);
and U7069 (N_7069,N_6743,N_6430);
and U7070 (N_7070,N_6977,N_6725);
xor U7071 (N_7071,N_6477,N_6556);
nor U7072 (N_7072,N_6943,N_6193);
or U7073 (N_7073,N_6125,N_6573);
and U7074 (N_7074,N_6863,N_6669);
nand U7075 (N_7075,N_6683,N_6303);
and U7076 (N_7076,N_6826,N_6632);
nand U7077 (N_7077,N_6429,N_6597);
nor U7078 (N_7078,N_6500,N_6626);
nand U7079 (N_7079,N_6878,N_6881);
and U7080 (N_7080,N_6151,N_6542);
and U7081 (N_7081,N_6936,N_6983);
or U7082 (N_7082,N_6650,N_6337);
nor U7083 (N_7083,N_6965,N_6339);
nor U7084 (N_7084,N_6724,N_6610);
nor U7085 (N_7085,N_6828,N_6677);
xnor U7086 (N_7086,N_6733,N_6456);
nand U7087 (N_7087,N_6399,N_6746);
nor U7088 (N_7088,N_6263,N_6596);
nand U7089 (N_7089,N_6759,N_6908);
and U7090 (N_7090,N_6048,N_6546);
or U7091 (N_7091,N_6046,N_6293);
nand U7092 (N_7092,N_6767,N_6024);
and U7093 (N_7093,N_6488,N_6101);
nand U7094 (N_7094,N_6051,N_6508);
nor U7095 (N_7095,N_6834,N_6843);
and U7096 (N_7096,N_6662,N_6836);
nor U7097 (N_7097,N_6658,N_6605);
nor U7098 (N_7098,N_6362,N_6095);
or U7099 (N_7099,N_6023,N_6100);
nand U7100 (N_7100,N_6663,N_6865);
xor U7101 (N_7101,N_6168,N_6531);
nor U7102 (N_7102,N_6446,N_6415);
or U7103 (N_7103,N_6551,N_6107);
and U7104 (N_7104,N_6142,N_6793);
or U7105 (N_7105,N_6182,N_6219);
nand U7106 (N_7106,N_6113,N_6952);
nand U7107 (N_7107,N_6458,N_6014);
nand U7108 (N_7108,N_6948,N_6460);
or U7109 (N_7109,N_6854,N_6829);
nor U7110 (N_7110,N_6643,N_6882);
nor U7111 (N_7111,N_6855,N_6587);
nor U7112 (N_7112,N_6096,N_6607);
nand U7113 (N_7113,N_6777,N_6078);
or U7114 (N_7114,N_6540,N_6913);
or U7115 (N_7115,N_6252,N_6314);
or U7116 (N_7116,N_6215,N_6208);
nor U7117 (N_7117,N_6031,N_6425);
or U7118 (N_7118,N_6875,N_6299);
nor U7119 (N_7119,N_6935,N_6440);
nand U7120 (N_7120,N_6067,N_6842);
nand U7121 (N_7121,N_6181,N_6139);
nand U7122 (N_7122,N_6507,N_6667);
nand U7123 (N_7123,N_6956,N_6442);
and U7124 (N_7124,N_6788,N_6911);
nand U7125 (N_7125,N_6514,N_6115);
nor U7126 (N_7126,N_6161,N_6939);
nand U7127 (N_7127,N_6557,N_6317);
nor U7128 (N_7128,N_6304,N_6975);
nor U7129 (N_7129,N_6528,N_6837);
nand U7130 (N_7130,N_6307,N_6419);
and U7131 (N_7131,N_6247,N_6515);
nor U7132 (N_7132,N_6116,N_6558);
and U7133 (N_7133,N_6416,N_6403);
and U7134 (N_7134,N_6678,N_6866);
or U7135 (N_7135,N_6397,N_6267);
nand U7136 (N_7136,N_6361,N_6798);
nor U7137 (N_7137,N_6851,N_6286);
or U7138 (N_7138,N_6225,N_6945);
and U7139 (N_7139,N_6703,N_6928);
nor U7140 (N_7140,N_6121,N_6352);
nor U7141 (N_7141,N_6519,N_6070);
or U7142 (N_7142,N_6390,N_6776);
nor U7143 (N_7143,N_6484,N_6501);
xnor U7144 (N_7144,N_6748,N_6249);
or U7145 (N_7145,N_6951,N_6206);
and U7146 (N_7146,N_6565,N_6489);
nor U7147 (N_7147,N_6963,N_6942);
nand U7148 (N_7148,N_6585,N_6173);
nor U7149 (N_7149,N_6131,N_6768);
nor U7150 (N_7150,N_6153,N_6183);
and U7151 (N_7151,N_6414,N_6822);
and U7152 (N_7152,N_6057,N_6261);
and U7153 (N_7153,N_6778,N_6245);
or U7154 (N_7154,N_6726,N_6862);
nand U7155 (N_7155,N_6395,N_6118);
or U7156 (N_7156,N_6970,N_6847);
nor U7157 (N_7157,N_6021,N_6902);
nand U7158 (N_7158,N_6205,N_6394);
or U7159 (N_7159,N_6938,N_6861);
or U7160 (N_7160,N_6972,N_6316);
nand U7161 (N_7161,N_6015,N_6325);
or U7162 (N_7162,N_6979,N_6187);
nor U7163 (N_7163,N_6284,N_6171);
nor U7164 (N_7164,N_6112,N_6982);
and U7165 (N_7165,N_6831,N_6368);
nor U7166 (N_7166,N_6033,N_6967);
nand U7167 (N_7167,N_6321,N_6158);
nor U7168 (N_7168,N_6010,N_6510);
nand U7169 (N_7169,N_6553,N_6745);
and U7170 (N_7170,N_6688,N_6888);
nor U7171 (N_7171,N_6923,N_6475);
or U7172 (N_7172,N_6676,N_6671);
nor U7173 (N_7173,N_6539,N_6097);
or U7174 (N_7174,N_6164,N_6165);
nor U7175 (N_7175,N_6505,N_6379);
nand U7176 (N_7176,N_6797,N_6496);
or U7177 (N_7177,N_6114,N_6396);
nor U7178 (N_7178,N_6222,N_6693);
and U7179 (N_7179,N_6552,N_6659);
and U7180 (N_7180,N_6106,N_6123);
and U7181 (N_7181,N_6685,N_6921);
or U7182 (N_7182,N_6471,N_6647);
nand U7183 (N_7183,N_6319,N_6606);
nor U7184 (N_7184,N_6410,N_6812);
nand U7185 (N_7185,N_6146,N_6816);
nor U7186 (N_7186,N_6697,N_6481);
or U7187 (N_7187,N_6820,N_6346);
nand U7188 (N_7188,N_6473,N_6796);
or U7189 (N_7189,N_6289,N_6660);
nor U7190 (N_7190,N_6479,N_6765);
nand U7191 (N_7191,N_6002,N_6609);
or U7192 (N_7192,N_6452,N_6841);
or U7193 (N_7193,N_6279,N_6648);
nor U7194 (N_7194,N_6149,N_6453);
and U7195 (N_7195,N_6320,N_6277);
nor U7196 (N_7196,N_6377,N_6719);
xor U7197 (N_7197,N_6495,N_6673);
and U7198 (N_7198,N_6305,N_6850);
nand U7199 (N_7199,N_6246,N_6930);
nor U7200 (N_7200,N_6052,N_6076);
nor U7201 (N_7201,N_6603,N_6957);
nor U7202 (N_7202,N_6265,N_6845);
and U7203 (N_7203,N_6702,N_6532);
nand U7204 (N_7204,N_6562,N_6709);
nor U7205 (N_7205,N_6439,N_6406);
and U7206 (N_7206,N_6590,N_6092);
and U7207 (N_7207,N_6896,N_6794);
nor U7208 (N_7208,N_6260,N_6230);
or U7209 (N_7209,N_6373,N_6492);
or U7210 (N_7210,N_6791,N_6617);
nor U7211 (N_7211,N_6188,N_6345);
and U7212 (N_7212,N_6654,N_6050);
nand U7213 (N_7213,N_6852,N_6233);
and U7214 (N_7214,N_6961,N_6413);
xor U7215 (N_7215,N_6710,N_6000);
nand U7216 (N_7216,N_6184,N_6524);
nor U7217 (N_7217,N_6758,N_6122);
and U7218 (N_7218,N_6140,N_6387);
or U7219 (N_7219,N_6004,N_6386);
or U7220 (N_7220,N_6281,N_6848);
nand U7221 (N_7221,N_6653,N_6701);
xnor U7222 (N_7222,N_6200,N_6686);
and U7223 (N_7223,N_6044,N_6810);
or U7224 (N_7224,N_6091,N_6809);
and U7225 (N_7225,N_6250,N_6844);
and U7226 (N_7226,N_6194,N_6175);
or U7227 (N_7227,N_6769,N_6461);
nor U7228 (N_7228,N_6503,N_6469);
nand U7229 (N_7229,N_6782,N_6343);
and U7230 (N_7230,N_6311,N_6916);
nor U7231 (N_7231,N_6991,N_6136);
or U7232 (N_7232,N_6370,N_6600);
nor U7233 (N_7233,N_6360,N_6231);
nor U7234 (N_7234,N_6825,N_6197);
xnor U7235 (N_7235,N_6656,N_6341);
nor U7236 (N_7236,N_6393,N_6235);
or U7237 (N_7237,N_6986,N_6818);
or U7238 (N_7238,N_6012,N_6744);
nand U7239 (N_7239,N_6502,N_6167);
or U7240 (N_7240,N_6363,N_6616);
nand U7241 (N_7241,N_6813,N_6891);
or U7242 (N_7242,N_6795,N_6417);
and U7243 (N_7243,N_6711,N_6918);
nor U7244 (N_7244,N_6451,N_6944);
or U7245 (N_7245,N_6287,N_6884);
and U7246 (N_7246,N_6814,N_6186);
and U7247 (N_7247,N_6431,N_6661);
or U7248 (N_7248,N_6132,N_6899);
nor U7249 (N_7249,N_6723,N_6405);
nand U7250 (N_7250,N_6691,N_6482);
and U7251 (N_7251,N_6800,N_6491);
or U7252 (N_7252,N_6421,N_6889);
nor U7253 (N_7253,N_6592,N_6497);
and U7254 (N_7254,N_6581,N_6849);
or U7255 (N_7255,N_6548,N_6038);
and U7256 (N_7256,N_6380,N_6630);
and U7257 (N_7257,N_6846,N_6547);
and U7258 (N_7258,N_6664,N_6564);
nor U7259 (N_7259,N_6251,N_6214);
or U7260 (N_7260,N_6271,N_6137);
or U7261 (N_7261,N_6412,N_6093);
nor U7262 (N_7262,N_6041,N_6533);
and U7263 (N_7263,N_6623,N_6645);
and U7264 (N_7264,N_6203,N_6919);
nor U7265 (N_7265,N_6207,N_6344);
nand U7266 (N_7266,N_6020,N_6869);
nand U7267 (N_7267,N_6236,N_6955);
nor U7268 (N_7268,N_6638,N_6620);
or U7269 (N_7269,N_6997,N_6378);
nand U7270 (N_7270,N_6032,N_6332);
and U7271 (N_7271,N_6803,N_6879);
and U7272 (N_7272,N_6134,N_6191);
nor U7273 (N_7273,N_6366,N_6915);
nand U7274 (N_7274,N_6001,N_6049);
nand U7275 (N_7275,N_6369,N_6127);
nand U7276 (N_7276,N_6280,N_6144);
nor U7277 (N_7277,N_6478,N_6098);
nor U7278 (N_7278,N_6179,N_6657);
or U7279 (N_7279,N_6717,N_6633);
nand U7280 (N_7280,N_6966,N_6907);
and U7281 (N_7281,N_6750,N_6783);
nand U7282 (N_7282,N_6486,N_6209);
nand U7283 (N_7283,N_6718,N_6629);
nor U7284 (N_7284,N_6740,N_6058);
nand U7285 (N_7285,N_6400,N_6670);
or U7286 (N_7286,N_6003,N_6727);
nand U7287 (N_7287,N_6608,N_6081);
nand U7288 (N_7288,N_6799,N_6512);
nor U7289 (N_7289,N_6270,N_6407);
xor U7290 (N_7290,N_6971,N_6126);
or U7291 (N_7291,N_6210,N_6934);
nor U7292 (N_7292,N_6065,N_6367);
or U7293 (N_7293,N_6521,N_6599);
nand U7294 (N_7294,N_6242,N_6994);
nand U7295 (N_7295,N_6728,N_6833);
nor U7296 (N_7296,N_6068,N_6327);
and U7297 (N_7297,N_6627,N_6066);
nor U7298 (N_7298,N_6516,N_6079);
and U7299 (N_7299,N_6073,N_6064);
nor U7300 (N_7300,N_6163,N_6555);
nand U7301 (N_7301,N_6860,N_6220);
or U7302 (N_7302,N_6454,N_6870);
or U7303 (N_7303,N_6008,N_6463);
or U7304 (N_7304,N_6696,N_6351);
nor U7305 (N_7305,N_6389,N_6763);
nand U7306 (N_7306,N_6428,N_6914);
nand U7307 (N_7307,N_6619,N_6631);
nand U7308 (N_7308,N_6213,N_6628);
and U7309 (N_7309,N_6706,N_6043);
nand U7310 (N_7310,N_6785,N_6217);
xor U7311 (N_7311,N_6353,N_6274);
nand U7312 (N_7312,N_6771,N_6535);
and U7313 (N_7313,N_6018,N_6392);
nand U7314 (N_7314,N_6313,N_6968);
and U7315 (N_7315,N_6781,N_6680);
nor U7316 (N_7316,N_6254,N_6318);
nor U7317 (N_7317,N_6355,N_6275);
or U7318 (N_7318,N_6615,N_6730);
and U7319 (N_7319,N_6448,N_6117);
nor U7320 (N_7320,N_6612,N_6584);
and U7321 (N_7321,N_6611,N_6823);
nand U7322 (N_7322,N_6753,N_6042);
and U7323 (N_7323,N_6080,N_6690);
or U7324 (N_7324,N_6641,N_6525);
nor U7325 (N_7325,N_6988,N_6244);
nand U7326 (N_7326,N_6487,N_6324);
xnor U7327 (N_7327,N_6017,N_6772);
nand U7328 (N_7328,N_6655,N_6601);
xnor U7329 (N_7329,N_6905,N_6450);
nand U7330 (N_7330,N_6195,N_6917);
nor U7331 (N_7331,N_6969,N_6283);
and U7332 (N_7332,N_6110,N_6383);
nor U7333 (N_7333,N_6155,N_6774);
nand U7334 (N_7334,N_6349,N_6887);
nand U7335 (N_7335,N_6639,N_6522);
or U7336 (N_7336,N_6815,N_6513);
nor U7337 (N_7337,N_6326,N_6135);
nor U7338 (N_7338,N_6692,N_6105);
nor U7339 (N_7339,N_6040,N_6835);
xnor U7340 (N_7340,N_6731,N_6550);
and U7341 (N_7341,N_6897,N_6912);
nand U7342 (N_7342,N_6480,N_6278);
and U7343 (N_7343,N_6227,N_6257);
nor U7344 (N_7344,N_6806,N_6821);
nor U7345 (N_7345,N_6687,N_6734);
or U7346 (N_7346,N_6987,N_6853);
xor U7347 (N_7347,N_6148,N_6315);
xnor U7348 (N_7348,N_6162,N_6722);
or U7349 (N_7349,N_6877,N_6946);
nand U7350 (N_7350,N_6582,N_6224);
and U7351 (N_7351,N_6374,N_6104);
or U7352 (N_7352,N_6468,N_6011);
nor U7353 (N_7353,N_6749,N_6294);
or U7354 (N_7354,N_6575,N_6306);
nor U7355 (N_7355,N_6580,N_6176);
nand U7356 (N_7356,N_6786,N_6892);
or U7357 (N_7357,N_6618,N_6770);
nand U7358 (N_7358,N_6204,N_6929);
nand U7359 (N_7359,N_6593,N_6560);
and U7360 (N_7360,N_6174,N_6013);
nor U7361 (N_7361,N_6467,N_6402);
xnor U7362 (N_7362,N_6559,N_6086);
or U7363 (N_7363,N_6992,N_6445);
and U7364 (N_7364,N_6998,N_6472);
or U7365 (N_7365,N_6561,N_6649);
and U7366 (N_7366,N_6549,N_6357);
and U7367 (N_7367,N_6291,N_6060);
or U7368 (N_7368,N_6885,N_6090);
nand U7369 (N_7369,N_6223,N_6895);
and U7370 (N_7370,N_6761,N_6699);
nand U7371 (N_7371,N_6792,N_6634);
nand U7372 (N_7372,N_6554,N_6537);
nor U7373 (N_7373,N_6328,N_6376);
and U7374 (N_7374,N_6061,N_6621);
or U7375 (N_7375,N_6150,N_6704);
xnor U7376 (N_7376,N_6371,N_6530);
nand U7377 (N_7377,N_6423,N_6348);
nor U7378 (N_7378,N_6485,N_6665);
xnor U7379 (N_7379,N_6016,N_6103);
nand U7380 (N_7380,N_6045,N_6873);
xor U7381 (N_7381,N_6180,N_6156);
nor U7382 (N_7382,N_6229,N_6301);
xnor U7383 (N_7383,N_6297,N_6381);
or U7384 (N_7384,N_6563,N_6602);
nor U7385 (N_7385,N_6470,N_6128);
nor U7386 (N_7386,N_6737,N_6801);
nand U7387 (N_7387,N_6920,N_6350);
and U7388 (N_7388,N_6830,N_6570);
nand U7389 (N_7389,N_6756,N_6981);
or U7390 (N_7390,N_6591,N_6511);
nor U7391 (N_7391,N_6941,N_6901);
nand U7392 (N_7392,N_6995,N_6752);
or U7393 (N_7393,N_6577,N_6039);
or U7394 (N_7394,N_6441,N_6411);
and U7395 (N_7395,N_6962,N_6466);
nor U7396 (N_7396,N_6006,N_6108);
and U7397 (N_7397,N_6166,N_6520);
or U7398 (N_7398,N_6642,N_6420);
nor U7399 (N_7399,N_6517,N_6273);
nand U7400 (N_7400,N_6069,N_6544);
and U7401 (N_7401,N_6443,N_6898);
nor U7402 (N_7402,N_6707,N_6201);
nand U7403 (N_7403,N_6571,N_6949);
or U7404 (N_7404,N_6708,N_6666);
nand U7405 (N_7405,N_6147,N_6893);
and U7406 (N_7406,N_6644,N_6700);
or U7407 (N_7407,N_6886,N_6534);
or U7408 (N_7408,N_6266,N_6160);
nor U7409 (N_7409,N_6668,N_6567);
or U7410 (N_7410,N_6388,N_6418);
nor U7411 (N_7411,N_6138,N_6819);
or U7412 (N_7412,N_6298,N_6543);
and U7413 (N_7413,N_6282,N_6904);
nor U7414 (N_7414,N_6329,N_6636);
nand U7415 (N_7415,N_6509,N_6755);
nor U7416 (N_7416,N_6455,N_6705);
or U7417 (N_7417,N_6356,N_6880);
nand U7418 (N_7418,N_6087,N_6141);
and U7419 (N_7419,N_6712,N_6401);
or U7420 (N_7420,N_6808,N_6154);
and U7421 (N_7421,N_6614,N_6874);
and U7422 (N_7422,N_6903,N_6940);
or U7423 (N_7423,N_6288,N_6292);
nand U7424 (N_7424,N_6840,N_6333);
nor U7425 (N_7425,N_6331,N_6071);
nor U7426 (N_7426,N_6408,N_6646);
or U7427 (N_7427,N_6212,N_6766);
nor U7428 (N_7428,N_6063,N_6741);
nand U7429 (N_7429,N_6576,N_6437);
nor U7430 (N_7430,N_6867,N_6354);
or U7431 (N_7431,N_6742,N_6804);
and U7432 (N_7432,N_6218,N_6240);
and U7433 (N_7433,N_6109,N_6735);
or U7434 (N_7434,N_6476,N_6159);
and U7435 (N_7435,N_6906,N_6684);
or U7436 (N_7436,N_6681,N_6436);
and U7437 (N_7437,N_6444,N_6409);
nand U7438 (N_7438,N_6216,N_6239);
nor U7439 (N_7439,N_6716,N_6202);
and U7440 (N_7440,N_6675,N_6022);
or U7441 (N_7441,N_6588,N_6871);
nor U7442 (N_7442,N_6464,N_6342);
or U7443 (N_7443,N_6805,N_6258);
nand U7444 (N_7444,N_6989,N_6613);
or U7445 (N_7445,N_6732,N_6790);
nand U7446 (N_7446,N_6404,N_6827);
or U7447 (N_7447,N_6075,N_6026);
nand U7448 (N_7448,N_6926,N_6449);
xnor U7449 (N_7449,N_6579,N_6838);
nor U7450 (N_7450,N_6322,N_6157);
or U7451 (N_7451,N_6269,N_6232);
nand U7452 (N_7452,N_6689,N_6839);
nand U7453 (N_7453,N_6145,N_6925);
nor U7454 (N_7454,N_6189,N_6947);
or U7455 (N_7455,N_6953,N_6499);
nor U7456 (N_7456,N_6864,N_6773);
nor U7457 (N_7457,N_6536,N_6256);
nand U7458 (N_7458,N_6129,N_6465);
nand U7459 (N_7459,N_6382,N_6211);
or U7460 (N_7460,N_6811,N_6119);
nand U7461 (N_7461,N_6652,N_6391);
nand U7462 (N_7462,N_6832,N_6999);
or U7463 (N_7463,N_6152,N_6993);
or U7464 (N_7464,N_6937,N_6085);
nor U7465 (N_7465,N_6780,N_6572);
nand U7466 (N_7466,N_6037,N_6226);
nor U7467 (N_7467,N_6990,N_6190);
nand U7468 (N_7468,N_6622,N_6931);
nor U7469 (N_7469,N_6055,N_6764);
nand U7470 (N_7470,N_6323,N_6300);
and U7471 (N_7471,N_6695,N_6924);
xor U7472 (N_7472,N_6736,N_6262);
or U7473 (N_7473,N_6787,N_6574);
or U7474 (N_7474,N_6005,N_6980);
nand U7475 (N_7475,N_6462,N_6199);
nand U7476 (N_7476,N_6541,N_6974);
nor U7477 (N_7477,N_6130,N_6089);
nor U7478 (N_7478,N_6424,N_6679);
nor U7479 (N_7479,N_6308,N_6996);
nor U7480 (N_7480,N_6538,N_6372);
nand U7481 (N_7481,N_6094,N_6964);
xnor U7482 (N_7482,N_6422,N_6950);
nor U7483 (N_7483,N_6954,N_6359);
nand U7484 (N_7484,N_6276,N_6624);
and U7485 (N_7485,N_6876,N_6637);
or U7486 (N_7486,N_6651,N_6985);
nor U7487 (N_7487,N_6196,N_6030);
or U7488 (N_7488,N_6029,N_6527);
nand U7489 (N_7489,N_6807,N_6932);
or U7490 (N_7490,N_6595,N_6221);
nor U7491 (N_7491,N_6715,N_6757);
and U7492 (N_7492,N_6028,N_6034);
and U7493 (N_7493,N_6976,N_6074);
nand U7494 (N_7494,N_6518,N_6720);
or U7495 (N_7495,N_6729,N_6789);
and U7496 (N_7496,N_6978,N_6385);
or U7497 (N_7497,N_6779,N_6170);
or U7498 (N_7498,N_6248,N_6036);
or U7499 (N_7499,N_6589,N_6426);
nand U7500 (N_7500,N_6471,N_6380);
nor U7501 (N_7501,N_6344,N_6036);
nand U7502 (N_7502,N_6667,N_6999);
nor U7503 (N_7503,N_6748,N_6642);
and U7504 (N_7504,N_6016,N_6184);
or U7505 (N_7505,N_6291,N_6001);
and U7506 (N_7506,N_6059,N_6417);
nand U7507 (N_7507,N_6990,N_6405);
and U7508 (N_7508,N_6229,N_6681);
and U7509 (N_7509,N_6750,N_6838);
nand U7510 (N_7510,N_6943,N_6049);
nor U7511 (N_7511,N_6646,N_6005);
and U7512 (N_7512,N_6219,N_6411);
and U7513 (N_7513,N_6324,N_6498);
and U7514 (N_7514,N_6191,N_6947);
nor U7515 (N_7515,N_6908,N_6297);
nand U7516 (N_7516,N_6944,N_6355);
or U7517 (N_7517,N_6478,N_6984);
nor U7518 (N_7518,N_6653,N_6001);
and U7519 (N_7519,N_6741,N_6607);
or U7520 (N_7520,N_6014,N_6759);
or U7521 (N_7521,N_6288,N_6193);
and U7522 (N_7522,N_6154,N_6324);
or U7523 (N_7523,N_6978,N_6483);
nor U7524 (N_7524,N_6606,N_6886);
nand U7525 (N_7525,N_6763,N_6845);
or U7526 (N_7526,N_6209,N_6218);
or U7527 (N_7527,N_6096,N_6778);
and U7528 (N_7528,N_6839,N_6446);
xnor U7529 (N_7529,N_6563,N_6125);
nand U7530 (N_7530,N_6292,N_6386);
nand U7531 (N_7531,N_6001,N_6041);
and U7532 (N_7532,N_6457,N_6454);
nand U7533 (N_7533,N_6304,N_6558);
nor U7534 (N_7534,N_6784,N_6164);
nor U7535 (N_7535,N_6593,N_6309);
or U7536 (N_7536,N_6253,N_6912);
and U7537 (N_7537,N_6432,N_6562);
or U7538 (N_7538,N_6448,N_6161);
nor U7539 (N_7539,N_6390,N_6349);
nor U7540 (N_7540,N_6229,N_6985);
nand U7541 (N_7541,N_6861,N_6231);
and U7542 (N_7542,N_6920,N_6211);
and U7543 (N_7543,N_6628,N_6306);
and U7544 (N_7544,N_6726,N_6756);
nand U7545 (N_7545,N_6741,N_6676);
nor U7546 (N_7546,N_6681,N_6353);
or U7547 (N_7547,N_6089,N_6913);
nor U7548 (N_7548,N_6760,N_6955);
xnor U7549 (N_7549,N_6251,N_6257);
nand U7550 (N_7550,N_6050,N_6202);
nand U7551 (N_7551,N_6651,N_6765);
or U7552 (N_7552,N_6884,N_6038);
nor U7553 (N_7553,N_6436,N_6785);
or U7554 (N_7554,N_6226,N_6459);
and U7555 (N_7555,N_6035,N_6933);
or U7556 (N_7556,N_6550,N_6411);
or U7557 (N_7557,N_6052,N_6213);
and U7558 (N_7558,N_6388,N_6532);
nor U7559 (N_7559,N_6550,N_6078);
or U7560 (N_7560,N_6325,N_6199);
and U7561 (N_7561,N_6768,N_6126);
or U7562 (N_7562,N_6148,N_6854);
nand U7563 (N_7563,N_6574,N_6287);
and U7564 (N_7564,N_6360,N_6583);
and U7565 (N_7565,N_6025,N_6275);
nand U7566 (N_7566,N_6209,N_6017);
or U7567 (N_7567,N_6174,N_6015);
or U7568 (N_7568,N_6357,N_6516);
and U7569 (N_7569,N_6549,N_6800);
and U7570 (N_7570,N_6538,N_6956);
or U7571 (N_7571,N_6230,N_6923);
and U7572 (N_7572,N_6371,N_6736);
nand U7573 (N_7573,N_6286,N_6462);
and U7574 (N_7574,N_6979,N_6621);
or U7575 (N_7575,N_6891,N_6766);
nor U7576 (N_7576,N_6455,N_6170);
and U7577 (N_7577,N_6468,N_6351);
xnor U7578 (N_7578,N_6846,N_6478);
and U7579 (N_7579,N_6808,N_6315);
nand U7580 (N_7580,N_6021,N_6880);
xnor U7581 (N_7581,N_6507,N_6733);
or U7582 (N_7582,N_6790,N_6221);
and U7583 (N_7583,N_6602,N_6933);
or U7584 (N_7584,N_6735,N_6459);
xor U7585 (N_7585,N_6247,N_6459);
nand U7586 (N_7586,N_6465,N_6438);
nor U7587 (N_7587,N_6275,N_6770);
and U7588 (N_7588,N_6228,N_6054);
nor U7589 (N_7589,N_6059,N_6385);
nand U7590 (N_7590,N_6653,N_6320);
nand U7591 (N_7591,N_6894,N_6867);
and U7592 (N_7592,N_6903,N_6719);
nand U7593 (N_7593,N_6392,N_6205);
nor U7594 (N_7594,N_6990,N_6183);
nor U7595 (N_7595,N_6346,N_6066);
nand U7596 (N_7596,N_6714,N_6392);
nand U7597 (N_7597,N_6348,N_6884);
or U7598 (N_7598,N_6357,N_6241);
or U7599 (N_7599,N_6948,N_6251);
nor U7600 (N_7600,N_6647,N_6554);
nor U7601 (N_7601,N_6246,N_6109);
nand U7602 (N_7602,N_6107,N_6043);
or U7603 (N_7603,N_6970,N_6341);
or U7604 (N_7604,N_6195,N_6387);
and U7605 (N_7605,N_6746,N_6117);
nand U7606 (N_7606,N_6249,N_6325);
and U7607 (N_7607,N_6107,N_6831);
and U7608 (N_7608,N_6433,N_6140);
nor U7609 (N_7609,N_6344,N_6176);
nand U7610 (N_7610,N_6797,N_6626);
or U7611 (N_7611,N_6089,N_6272);
and U7612 (N_7612,N_6485,N_6275);
and U7613 (N_7613,N_6124,N_6751);
or U7614 (N_7614,N_6053,N_6049);
or U7615 (N_7615,N_6703,N_6179);
and U7616 (N_7616,N_6905,N_6328);
and U7617 (N_7617,N_6145,N_6444);
xnor U7618 (N_7618,N_6713,N_6676);
and U7619 (N_7619,N_6559,N_6910);
nand U7620 (N_7620,N_6149,N_6702);
or U7621 (N_7621,N_6785,N_6051);
nor U7622 (N_7622,N_6253,N_6899);
or U7623 (N_7623,N_6107,N_6036);
nand U7624 (N_7624,N_6489,N_6435);
nor U7625 (N_7625,N_6988,N_6138);
or U7626 (N_7626,N_6056,N_6176);
nor U7627 (N_7627,N_6898,N_6152);
nor U7628 (N_7628,N_6661,N_6321);
nor U7629 (N_7629,N_6141,N_6239);
and U7630 (N_7630,N_6103,N_6779);
nor U7631 (N_7631,N_6430,N_6342);
nand U7632 (N_7632,N_6098,N_6628);
and U7633 (N_7633,N_6005,N_6126);
or U7634 (N_7634,N_6969,N_6625);
nand U7635 (N_7635,N_6639,N_6752);
or U7636 (N_7636,N_6916,N_6919);
nand U7637 (N_7637,N_6670,N_6565);
or U7638 (N_7638,N_6940,N_6242);
nor U7639 (N_7639,N_6445,N_6431);
or U7640 (N_7640,N_6443,N_6751);
or U7641 (N_7641,N_6698,N_6857);
nand U7642 (N_7642,N_6067,N_6168);
and U7643 (N_7643,N_6042,N_6857);
or U7644 (N_7644,N_6490,N_6279);
nand U7645 (N_7645,N_6156,N_6368);
nand U7646 (N_7646,N_6772,N_6475);
nor U7647 (N_7647,N_6972,N_6492);
xor U7648 (N_7648,N_6124,N_6442);
and U7649 (N_7649,N_6737,N_6958);
nand U7650 (N_7650,N_6909,N_6926);
nand U7651 (N_7651,N_6463,N_6565);
nor U7652 (N_7652,N_6553,N_6008);
and U7653 (N_7653,N_6952,N_6646);
nand U7654 (N_7654,N_6264,N_6624);
or U7655 (N_7655,N_6727,N_6105);
nor U7656 (N_7656,N_6480,N_6510);
nand U7657 (N_7657,N_6461,N_6283);
nand U7658 (N_7658,N_6735,N_6096);
or U7659 (N_7659,N_6103,N_6345);
nor U7660 (N_7660,N_6216,N_6382);
nor U7661 (N_7661,N_6169,N_6764);
or U7662 (N_7662,N_6739,N_6244);
nand U7663 (N_7663,N_6859,N_6684);
nor U7664 (N_7664,N_6834,N_6416);
and U7665 (N_7665,N_6575,N_6309);
nor U7666 (N_7666,N_6035,N_6795);
and U7667 (N_7667,N_6760,N_6569);
or U7668 (N_7668,N_6192,N_6149);
and U7669 (N_7669,N_6399,N_6935);
or U7670 (N_7670,N_6857,N_6525);
nor U7671 (N_7671,N_6348,N_6201);
or U7672 (N_7672,N_6238,N_6412);
or U7673 (N_7673,N_6759,N_6949);
and U7674 (N_7674,N_6077,N_6337);
nand U7675 (N_7675,N_6600,N_6591);
nor U7676 (N_7676,N_6586,N_6911);
nand U7677 (N_7677,N_6572,N_6827);
nand U7678 (N_7678,N_6472,N_6260);
nand U7679 (N_7679,N_6401,N_6010);
or U7680 (N_7680,N_6891,N_6926);
nand U7681 (N_7681,N_6835,N_6254);
or U7682 (N_7682,N_6169,N_6916);
and U7683 (N_7683,N_6191,N_6507);
nand U7684 (N_7684,N_6059,N_6159);
nor U7685 (N_7685,N_6134,N_6752);
or U7686 (N_7686,N_6539,N_6521);
nand U7687 (N_7687,N_6873,N_6805);
nor U7688 (N_7688,N_6379,N_6812);
and U7689 (N_7689,N_6200,N_6512);
nand U7690 (N_7690,N_6934,N_6036);
nand U7691 (N_7691,N_6702,N_6666);
nand U7692 (N_7692,N_6037,N_6143);
and U7693 (N_7693,N_6883,N_6735);
and U7694 (N_7694,N_6155,N_6060);
nor U7695 (N_7695,N_6541,N_6085);
nand U7696 (N_7696,N_6127,N_6187);
and U7697 (N_7697,N_6874,N_6722);
nor U7698 (N_7698,N_6487,N_6500);
or U7699 (N_7699,N_6576,N_6729);
nand U7700 (N_7700,N_6485,N_6484);
or U7701 (N_7701,N_6973,N_6684);
or U7702 (N_7702,N_6953,N_6370);
nand U7703 (N_7703,N_6172,N_6474);
and U7704 (N_7704,N_6496,N_6795);
and U7705 (N_7705,N_6245,N_6121);
or U7706 (N_7706,N_6720,N_6823);
or U7707 (N_7707,N_6049,N_6199);
and U7708 (N_7708,N_6949,N_6341);
and U7709 (N_7709,N_6017,N_6704);
or U7710 (N_7710,N_6181,N_6853);
or U7711 (N_7711,N_6232,N_6450);
nor U7712 (N_7712,N_6255,N_6807);
and U7713 (N_7713,N_6306,N_6144);
or U7714 (N_7714,N_6456,N_6101);
and U7715 (N_7715,N_6691,N_6480);
nand U7716 (N_7716,N_6056,N_6943);
and U7717 (N_7717,N_6702,N_6586);
or U7718 (N_7718,N_6753,N_6250);
and U7719 (N_7719,N_6651,N_6039);
nand U7720 (N_7720,N_6996,N_6324);
nand U7721 (N_7721,N_6430,N_6958);
nor U7722 (N_7722,N_6079,N_6650);
nor U7723 (N_7723,N_6416,N_6942);
or U7724 (N_7724,N_6363,N_6415);
xnor U7725 (N_7725,N_6048,N_6902);
or U7726 (N_7726,N_6517,N_6218);
and U7727 (N_7727,N_6692,N_6918);
and U7728 (N_7728,N_6240,N_6084);
or U7729 (N_7729,N_6760,N_6620);
nand U7730 (N_7730,N_6758,N_6401);
or U7731 (N_7731,N_6270,N_6131);
or U7732 (N_7732,N_6512,N_6666);
or U7733 (N_7733,N_6884,N_6983);
nor U7734 (N_7734,N_6913,N_6123);
and U7735 (N_7735,N_6587,N_6173);
nand U7736 (N_7736,N_6904,N_6746);
or U7737 (N_7737,N_6760,N_6191);
and U7738 (N_7738,N_6938,N_6755);
nand U7739 (N_7739,N_6090,N_6010);
and U7740 (N_7740,N_6225,N_6513);
or U7741 (N_7741,N_6043,N_6527);
nor U7742 (N_7742,N_6086,N_6972);
or U7743 (N_7743,N_6844,N_6255);
xor U7744 (N_7744,N_6538,N_6766);
and U7745 (N_7745,N_6888,N_6972);
nor U7746 (N_7746,N_6155,N_6292);
and U7747 (N_7747,N_6027,N_6303);
nor U7748 (N_7748,N_6269,N_6352);
or U7749 (N_7749,N_6912,N_6053);
nand U7750 (N_7750,N_6033,N_6437);
nand U7751 (N_7751,N_6784,N_6948);
and U7752 (N_7752,N_6575,N_6714);
and U7753 (N_7753,N_6402,N_6379);
or U7754 (N_7754,N_6096,N_6520);
and U7755 (N_7755,N_6345,N_6956);
nor U7756 (N_7756,N_6294,N_6627);
nand U7757 (N_7757,N_6323,N_6198);
nor U7758 (N_7758,N_6469,N_6564);
or U7759 (N_7759,N_6248,N_6385);
nor U7760 (N_7760,N_6305,N_6855);
and U7761 (N_7761,N_6937,N_6910);
and U7762 (N_7762,N_6184,N_6477);
or U7763 (N_7763,N_6182,N_6644);
or U7764 (N_7764,N_6792,N_6452);
nor U7765 (N_7765,N_6947,N_6887);
nand U7766 (N_7766,N_6420,N_6429);
and U7767 (N_7767,N_6311,N_6623);
nor U7768 (N_7768,N_6139,N_6196);
nand U7769 (N_7769,N_6706,N_6422);
or U7770 (N_7770,N_6097,N_6122);
nor U7771 (N_7771,N_6271,N_6999);
and U7772 (N_7772,N_6639,N_6540);
nand U7773 (N_7773,N_6225,N_6974);
xnor U7774 (N_7774,N_6417,N_6915);
nor U7775 (N_7775,N_6272,N_6129);
xor U7776 (N_7776,N_6097,N_6590);
and U7777 (N_7777,N_6078,N_6227);
nand U7778 (N_7778,N_6456,N_6572);
nand U7779 (N_7779,N_6875,N_6255);
or U7780 (N_7780,N_6286,N_6853);
or U7781 (N_7781,N_6242,N_6302);
nand U7782 (N_7782,N_6726,N_6940);
nor U7783 (N_7783,N_6735,N_6196);
nor U7784 (N_7784,N_6934,N_6318);
or U7785 (N_7785,N_6117,N_6167);
and U7786 (N_7786,N_6160,N_6096);
and U7787 (N_7787,N_6630,N_6005);
nor U7788 (N_7788,N_6112,N_6666);
and U7789 (N_7789,N_6279,N_6629);
or U7790 (N_7790,N_6566,N_6091);
xnor U7791 (N_7791,N_6512,N_6285);
nor U7792 (N_7792,N_6456,N_6054);
or U7793 (N_7793,N_6041,N_6150);
nand U7794 (N_7794,N_6412,N_6443);
and U7795 (N_7795,N_6914,N_6021);
and U7796 (N_7796,N_6239,N_6150);
or U7797 (N_7797,N_6192,N_6892);
nor U7798 (N_7798,N_6136,N_6077);
and U7799 (N_7799,N_6754,N_6680);
nor U7800 (N_7800,N_6589,N_6621);
or U7801 (N_7801,N_6782,N_6763);
nand U7802 (N_7802,N_6491,N_6638);
nor U7803 (N_7803,N_6956,N_6002);
or U7804 (N_7804,N_6380,N_6505);
and U7805 (N_7805,N_6955,N_6727);
and U7806 (N_7806,N_6725,N_6236);
nand U7807 (N_7807,N_6637,N_6765);
nand U7808 (N_7808,N_6245,N_6461);
nand U7809 (N_7809,N_6156,N_6195);
nand U7810 (N_7810,N_6721,N_6349);
and U7811 (N_7811,N_6426,N_6077);
or U7812 (N_7812,N_6988,N_6654);
or U7813 (N_7813,N_6286,N_6434);
nand U7814 (N_7814,N_6720,N_6153);
or U7815 (N_7815,N_6313,N_6943);
and U7816 (N_7816,N_6875,N_6032);
nor U7817 (N_7817,N_6625,N_6306);
and U7818 (N_7818,N_6357,N_6199);
nor U7819 (N_7819,N_6862,N_6422);
nand U7820 (N_7820,N_6010,N_6155);
nand U7821 (N_7821,N_6447,N_6423);
nor U7822 (N_7822,N_6915,N_6577);
and U7823 (N_7823,N_6809,N_6180);
or U7824 (N_7824,N_6032,N_6592);
or U7825 (N_7825,N_6112,N_6373);
and U7826 (N_7826,N_6381,N_6733);
nand U7827 (N_7827,N_6744,N_6729);
and U7828 (N_7828,N_6140,N_6184);
or U7829 (N_7829,N_6617,N_6483);
nor U7830 (N_7830,N_6834,N_6742);
and U7831 (N_7831,N_6872,N_6678);
nand U7832 (N_7832,N_6837,N_6326);
or U7833 (N_7833,N_6990,N_6059);
or U7834 (N_7834,N_6204,N_6042);
or U7835 (N_7835,N_6610,N_6925);
xnor U7836 (N_7836,N_6236,N_6662);
or U7837 (N_7837,N_6467,N_6959);
xor U7838 (N_7838,N_6463,N_6013);
and U7839 (N_7839,N_6056,N_6706);
xnor U7840 (N_7840,N_6704,N_6822);
or U7841 (N_7841,N_6459,N_6438);
and U7842 (N_7842,N_6494,N_6768);
nand U7843 (N_7843,N_6990,N_6412);
or U7844 (N_7844,N_6864,N_6306);
nor U7845 (N_7845,N_6870,N_6349);
and U7846 (N_7846,N_6920,N_6037);
nor U7847 (N_7847,N_6811,N_6445);
nand U7848 (N_7848,N_6720,N_6219);
or U7849 (N_7849,N_6087,N_6709);
or U7850 (N_7850,N_6403,N_6652);
nor U7851 (N_7851,N_6191,N_6340);
and U7852 (N_7852,N_6397,N_6403);
nor U7853 (N_7853,N_6018,N_6697);
and U7854 (N_7854,N_6895,N_6971);
nor U7855 (N_7855,N_6975,N_6785);
nor U7856 (N_7856,N_6115,N_6365);
nor U7857 (N_7857,N_6704,N_6083);
nor U7858 (N_7858,N_6410,N_6458);
nand U7859 (N_7859,N_6141,N_6221);
nand U7860 (N_7860,N_6894,N_6883);
or U7861 (N_7861,N_6089,N_6412);
nor U7862 (N_7862,N_6141,N_6594);
nand U7863 (N_7863,N_6643,N_6645);
and U7864 (N_7864,N_6055,N_6736);
and U7865 (N_7865,N_6582,N_6453);
or U7866 (N_7866,N_6767,N_6267);
nand U7867 (N_7867,N_6776,N_6965);
nand U7868 (N_7868,N_6285,N_6028);
and U7869 (N_7869,N_6154,N_6282);
and U7870 (N_7870,N_6769,N_6730);
nor U7871 (N_7871,N_6537,N_6035);
or U7872 (N_7872,N_6763,N_6076);
or U7873 (N_7873,N_6363,N_6306);
or U7874 (N_7874,N_6234,N_6435);
nor U7875 (N_7875,N_6888,N_6563);
nand U7876 (N_7876,N_6902,N_6957);
or U7877 (N_7877,N_6542,N_6504);
and U7878 (N_7878,N_6965,N_6527);
nand U7879 (N_7879,N_6467,N_6834);
nor U7880 (N_7880,N_6509,N_6194);
nor U7881 (N_7881,N_6573,N_6165);
or U7882 (N_7882,N_6966,N_6763);
nand U7883 (N_7883,N_6097,N_6959);
nor U7884 (N_7884,N_6750,N_6510);
nor U7885 (N_7885,N_6891,N_6086);
nand U7886 (N_7886,N_6800,N_6332);
nor U7887 (N_7887,N_6557,N_6623);
nor U7888 (N_7888,N_6683,N_6072);
nor U7889 (N_7889,N_6063,N_6610);
and U7890 (N_7890,N_6261,N_6924);
nor U7891 (N_7891,N_6464,N_6924);
nand U7892 (N_7892,N_6656,N_6547);
nor U7893 (N_7893,N_6442,N_6701);
or U7894 (N_7894,N_6683,N_6599);
nand U7895 (N_7895,N_6627,N_6729);
nand U7896 (N_7896,N_6953,N_6528);
nor U7897 (N_7897,N_6455,N_6930);
and U7898 (N_7898,N_6965,N_6132);
and U7899 (N_7899,N_6998,N_6645);
or U7900 (N_7900,N_6600,N_6140);
nor U7901 (N_7901,N_6069,N_6150);
and U7902 (N_7902,N_6901,N_6987);
nand U7903 (N_7903,N_6698,N_6255);
or U7904 (N_7904,N_6809,N_6552);
or U7905 (N_7905,N_6188,N_6145);
or U7906 (N_7906,N_6592,N_6084);
xor U7907 (N_7907,N_6200,N_6809);
or U7908 (N_7908,N_6403,N_6139);
or U7909 (N_7909,N_6467,N_6512);
nor U7910 (N_7910,N_6773,N_6622);
nor U7911 (N_7911,N_6849,N_6248);
or U7912 (N_7912,N_6649,N_6644);
nor U7913 (N_7913,N_6741,N_6082);
and U7914 (N_7914,N_6478,N_6586);
and U7915 (N_7915,N_6498,N_6742);
nand U7916 (N_7916,N_6995,N_6684);
nand U7917 (N_7917,N_6268,N_6397);
nor U7918 (N_7918,N_6684,N_6858);
nand U7919 (N_7919,N_6974,N_6285);
nand U7920 (N_7920,N_6339,N_6009);
nand U7921 (N_7921,N_6503,N_6851);
and U7922 (N_7922,N_6789,N_6484);
or U7923 (N_7923,N_6457,N_6442);
and U7924 (N_7924,N_6890,N_6771);
nor U7925 (N_7925,N_6967,N_6599);
nand U7926 (N_7926,N_6005,N_6973);
nand U7927 (N_7927,N_6416,N_6700);
and U7928 (N_7928,N_6450,N_6128);
and U7929 (N_7929,N_6484,N_6094);
nand U7930 (N_7930,N_6193,N_6933);
nor U7931 (N_7931,N_6220,N_6411);
and U7932 (N_7932,N_6776,N_6728);
nand U7933 (N_7933,N_6416,N_6899);
or U7934 (N_7934,N_6182,N_6826);
or U7935 (N_7935,N_6446,N_6947);
or U7936 (N_7936,N_6187,N_6688);
nand U7937 (N_7937,N_6155,N_6343);
nand U7938 (N_7938,N_6589,N_6523);
or U7939 (N_7939,N_6502,N_6407);
or U7940 (N_7940,N_6707,N_6694);
and U7941 (N_7941,N_6823,N_6241);
nand U7942 (N_7942,N_6581,N_6211);
nand U7943 (N_7943,N_6453,N_6590);
and U7944 (N_7944,N_6043,N_6228);
nand U7945 (N_7945,N_6128,N_6086);
or U7946 (N_7946,N_6383,N_6458);
nor U7947 (N_7947,N_6671,N_6497);
nor U7948 (N_7948,N_6445,N_6519);
and U7949 (N_7949,N_6695,N_6539);
and U7950 (N_7950,N_6632,N_6713);
nor U7951 (N_7951,N_6098,N_6049);
nor U7952 (N_7952,N_6097,N_6736);
or U7953 (N_7953,N_6363,N_6445);
or U7954 (N_7954,N_6978,N_6133);
nand U7955 (N_7955,N_6923,N_6575);
nand U7956 (N_7956,N_6232,N_6071);
nor U7957 (N_7957,N_6188,N_6968);
nand U7958 (N_7958,N_6390,N_6904);
or U7959 (N_7959,N_6221,N_6858);
and U7960 (N_7960,N_6122,N_6137);
nor U7961 (N_7961,N_6844,N_6362);
and U7962 (N_7962,N_6580,N_6151);
nor U7963 (N_7963,N_6247,N_6372);
nand U7964 (N_7964,N_6462,N_6368);
or U7965 (N_7965,N_6017,N_6326);
nand U7966 (N_7966,N_6194,N_6989);
and U7967 (N_7967,N_6692,N_6912);
and U7968 (N_7968,N_6026,N_6500);
nand U7969 (N_7969,N_6757,N_6425);
and U7970 (N_7970,N_6985,N_6087);
and U7971 (N_7971,N_6939,N_6284);
nor U7972 (N_7972,N_6991,N_6836);
nand U7973 (N_7973,N_6317,N_6596);
and U7974 (N_7974,N_6397,N_6656);
nand U7975 (N_7975,N_6785,N_6769);
nand U7976 (N_7976,N_6997,N_6978);
or U7977 (N_7977,N_6111,N_6667);
or U7978 (N_7978,N_6656,N_6031);
nor U7979 (N_7979,N_6164,N_6279);
nand U7980 (N_7980,N_6776,N_6758);
or U7981 (N_7981,N_6927,N_6760);
or U7982 (N_7982,N_6933,N_6218);
nor U7983 (N_7983,N_6941,N_6344);
or U7984 (N_7984,N_6010,N_6705);
nor U7985 (N_7985,N_6243,N_6152);
and U7986 (N_7986,N_6488,N_6053);
nor U7987 (N_7987,N_6002,N_6390);
or U7988 (N_7988,N_6200,N_6519);
nand U7989 (N_7989,N_6099,N_6101);
and U7990 (N_7990,N_6315,N_6614);
nand U7991 (N_7991,N_6582,N_6553);
or U7992 (N_7992,N_6909,N_6189);
nor U7993 (N_7993,N_6663,N_6030);
nor U7994 (N_7994,N_6545,N_6001);
nand U7995 (N_7995,N_6054,N_6135);
and U7996 (N_7996,N_6963,N_6953);
or U7997 (N_7997,N_6979,N_6441);
and U7998 (N_7998,N_6309,N_6437);
and U7999 (N_7999,N_6698,N_6462);
nand U8000 (N_8000,N_7902,N_7707);
and U8001 (N_8001,N_7561,N_7468);
or U8002 (N_8002,N_7673,N_7688);
nor U8003 (N_8003,N_7007,N_7927);
and U8004 (N_8004,N_7363,N_7849);
or U8005 (N_8005,N_7440,N_7784);
nand U8006 (N_8006,N_7329,N_7254);
or U8007 (N_8007,N_7985,N_7162);
nand U8008 (N_8008,N_7103,N_7471);
or U8009 (N_8009,N_7180,N_7819);
or U8010 (N_8010,N_7810,N_7716);
and U8011 (N_8011,N_7624,N_7799);
or U8012 (N_8012,N_7487,N_7637);
and U8013 (N_8013,N_7474,N_7120);
and U8014 (N_8014,N_7404,N_7731);
nor U8015 (N_8015,N_7623,N_7496);
nand U8016 (N_8016,N_7663,N_7840);
nand U8017 (N_8017,N_7607,N_7224);
nor U8018 (N_8018,N_7122,N_7820);
nand U8019 (N_8019,N_7344,N_7386);
nand U8020 (N_8020,N_7172,N_7929);
nor U8021 (N_8021,N_7141,N_7916);
and U8022 (N_8022,N_7566,N_7093);
nand U8023 (N_8023,N_7888,N_7877);
and U8024 (N_8024,N_7159,N_7101);
and U8025 (N_8025,N_7951,N_7578);
and U8026 (N_8026,N_7678,N_7942);
nor U8027 (N_8027,N_7040,N_7744);
or U8028 (N_8028,N_7538,N_7156);
or U8029 (N_8029,N_7096,N_7456);
or U8030 (N_8030,N_7537,N_7695);
and U8031 (N_8031,N_7668,N_7639);
xor U8032 (N_8032,N_7477,N_7323);
or U8033 (N_8033,N_7937,N_7331);
and U8034 (N_8034,N_7166,N_7029);
nand U8035 (N_8035,N_7586,N_7223);
nor U8036 (N_8036,N_7351,N_7168);
xnor U8037 (N_8037,N_7195,N_7775);
and U8038 (N_8038,N_7176,N_7206);
nor U8039 (N_8039,N_7816,N_7797);
or U8040 (N_8040,N_7628,N_7415);
nand U8041 (N_8041,N_7424,N_7954);
nand U8042 (N_8042,N_7648,N_7686);
nor U8043 (N_8043,N_7151,N_7436);
nand U8044 (N_8044,N_7061,N_7041);
or U8045 (N_8045,N_7697,N_7320);
or U8046 (N_8046,N_7494,N_7119);
nand U8047 (N_8047,N_7727,N_7177);
or U8048 (N_8048,N_7393,N_7105);
and U8049 (N_8049,N_7718,N_7498);
nand U8050 (N_8050,N_7878,N_7322);
and U8051 (N_8051,N_7190,N_7396);
nor U8052 (N_8052,N_7956,N_7720);
nor U8053 (N_8053,N_7522,N_7631);
or U8054 (N_8054,N_7107,N_7349);
and U8055 (N_8055,N_7669,N_7766);
and U8056 (N_8056,N_7197,N_7986);
and U8057 (N_8057,N_7062,N_7188);
nand U8058 (N_8058,N_7854,N_7893);
nand U8059 (N_8059,N_7917,N_7944);
nor U8060 (N_8060,N_7202,N_7724);
nor U8061 (N_8061,N_7642,N_7781);
nor U8062 (N_8062,N_7199,N_7638);
nor U8063 (N_8063,N_7535,N_7271);
nand U8064 (N_8064,N_7161,N_7227);
nand U8065 (N_8065,N_7116,N_7066);
or U8066 (N_8066,N_7568,N_7831);
and U8067 (N_8067,N_7426,N_7778);
nand U8068 (N_8068,N_7175,N_7657);
or U8069 (N_8069,N_7390,N_7276);
nor U8070 (N_8070,N_7420,N_7711);
and U8071 (N_8071,N_7894,N_7078);
nand U8072 (N_8072,N_7516,N_7546);
nand U8073 (N_8073,N_7692,N_7681);
xnor U8074 (N_8074,N_7340,N_7575);
nand U8075 (N_8075,N_7736,N_7130);
xor U8076 (N_8076,N_7264,N_7454);
nand U8077 (N_8077,N_7140,N_7941);
and U8078 (N_8078,N_7262,N_7824);
nand U8079 (N_8079,N_7406,N_7912);
nand U8080 (N_8080,N_7305,N_7201);
or U8081 (N_8081,N_7553,N_7988);
nor U8082 (N_8082,N_7839,N_7875);
nand U8083 (N_8083,N_7333,N_7072);
or U8084 (N_8084,N_7497,N_7706);
nor U8085 (N_8085,N_7048,N_7028);
or U8086 (N_8086,N_7853,N_7409);
nand U8087 (N_8087,N_7589,N_7082);
or U8088 (N_8088,N_7899,N_7024);
and U8089 (N_8089,N_7090,N_7830);
and U8090 (N_8090,N_7625,N_7476);
and U8091 (N_8091,N_7787,N_7633);
nand U8092 (N_8092,N_7297,N_7829);
and U8093 (N_8093,N_7410,N_7975);
nand U8094 (N_8094,N_7018,N_7455);
and U8095 (N_8095,N_7970,N_7211);
nor U8096 (N_8096,N_7636,N_7756);
nor U8097 (N_8097,N_7065,N_7821);
or U8098 (N_8098,N_7843,N_7651);
or U8099 (N_8099,N_7053,N_7825);
or U8100 (N_8100,N_7511,N_7054);
xnor U8101 (N_8101,N_7289,N_7388);
nand U8102 (N_8102,N_7354,N_7055);
nor U8103 (N_8103,N_7357,N_7020);
or U8104 (N_8104,N_7580,N_7907);
nand U8105 (N_8105,N_7758,N_7621);
nor U8106 (N_8106,N_7258,N_7481);
nand U8107 (N_8107,N_7773,N_7774);
and U8108 (N_8108,N_7478,N_7952);
nor U8109 (N_8109,N_7032,N_7573);
or U8110 (N_8110,N_7443,N_7173);
or U8111 (N_8111,N_7909,N_7574);
and U8112 (N_8112,N_7838,N_7464);
nor U8113 (N_8113,N_7044,N_7299);
nor U8114 (N_8114,N_7634,N_7121);
nor U8115 (N_8115,N_7010,N_7052);
and U8116 (N_8116,N_7138,N_7674);
nand U8117 (N_8117,N_7514,N_7928);
nor U8118 (N_8118,N_7070,N_7914);
nor U8119 (N_8119,N_7270,N_7071);
nor U8120 (N_8120,N_7260,N_7745);
or U8121 (N_8121,N_7602,N_7540);
or U8122 (N_8122,N_7364,N_7618);
or U8123 (N_8123,N_7304,N_7207);
or U8124 (N_8124,N_7682,N_7347);
nand U8125 (N_8125,N_7549,N_7675);
or U8126 (N_8126,N_7059,N_7684);
and U8127 (N_8127,N_7908,N_7739);
nand U8128 (N_8128,N_7457,N_7795);
or U8129 (N_8129,N_7221,N_7922);
nor U8130 (N_8130,N_7353,N_7597);
nand U8131 (N_8131,N_7938,N_7460);
nor U8132 (N_8132,N_7581,N_7037);
or U8133 (N_8133,N_7097,N_7273);
and U8134 (N_8134,N_7128,N_7398);
nand U8135 (N_8135,N_7635,N_7489);
or U8136 (N_8136,N_7208,N_7379);
nand U8137 (N_8137,N_7490,N_7013);
nor U8138 (N_8138,N_7990,N_7226);
or U8139 (N_8139,N_7215,N_7132);
nand U8140 (N_8140,N_7139,N_7892);
and U8141 (N_8141,N_7547,N_7989);
nand U8142 (N_8142,N_7730,N_7501);
and U8143 (N_8143,N_7268,N_7536);
nor U8144 (N_8144,N_7643,N_7413);
or U8145 (N_8145,N_7220,N_7785);
nand U8146 (N_8146,N_7038,N_7073);
or U8147 (N_8147,N_7741,N_7746);
nand U8148 (N_8148,N_7699,N_7383);
nand U8149 (N_8149,N_7380,N_7170);
nand U8150 (N_8150,N_7924,N_7993);
nand U8151 (N_8151,N_7714,N_7943);
or U8152 (N_8152,N_7277,N_7001);
nor U8153 (N_8153,N_7508,N_7879);
or U8154 (N_8154,N_7605,N_7934);
or U8155 (N_8155,N_7728,N_7421);
nand U8156 (N_8156,N_7905,N_7447);
nand U8157 (N_8157,N_7004,N_7068);
and U8158 (N_8158,N_7615,N_7448);
nand U8159 (N_8159,N_7087,N_7033);
and U8160 (N_8160,N_7280,N_7931);
nand U8161 (N_8161,N_7805,N_7726);
or U8162 (N_8162,N_7666,N_7316);
and U8163 (N_8163,N_7935,N_7236);
and U8164 (N_8164,N_7652,N_7856);
nor U8165 (N_8165,N_7313,N_7376);
or U8166 (N_8166,N_7035,N_7959);
nor U8167 (N_8167,N_7338,N_7031);
nor U8168 (N_8168,N_7486,N_7493);
nand U8169 (N_8169,N_7984,N_7610);
nand U8170 (N_8170,N_7500,N_7595);
nor U8171 (N_8171,N_7627,N_7565);
or U8172 (N_8172,N_7169,N_7622);
nor U8173 (N_8173,N_7771,N_7754);
and U8174 (N_8174,N_7603,N_7683);
or U8175 (N_8175,N_7261,N_7887);
nor U8176 (N_8176,N_7732,N_7614);
and U8177 (N_8177,N_7898,N_7428);
and U8178 (N_8178,N_7981,N_7281);
and U8179 (N_8179,N_7579,N_7234);
nand U8180 (N_8180,N_7432,N_7520);
nor U8181 (N_8181,N_7154,N_7735);
nand U8182 (N_8182,N_7019,N_7336);
and U8183 (N_8183,N_7864,N_7507);
nor U8184 (N_8184,N_7418,N_7343);
nand U8185 (N_8185,N_7793,N_7583);
nand U8186 (N_8186,N_7963,N_7086);
nand U8187 (N_8187,N_7252,N_7873);
nor U8188 (N_8188,N_7137,N_7848);
and U8189 (N_8189,N_7375,N_7723);
nor U8190 (N_8190,N_7751,N_7861);
or U8191 (N_8191,N_7527,N_7222);
nor U8192 (N_8192,N_7994,N_7427);
and U8193 (N_8193,N_7679,N_7971);
or U8194 (N_8194,N_7506,N_7715);
and U8195 (N_8195,N_7617,N_7022);
nor U8196 (N_8196,N_7852,N_7492);
or U8197 (N_8197,N_7826,N_7135);
or U8198 (N_8198,N_7011,N_7534);
nor U8199 (N_8199,N_7964,N_7431);
nand U8200 (N_8200,N_7495,N_7069);
or U8201 (N_8201,N_7616,N_7900);
and U8202 (N_8202,N_7181,N_7885);
nor U8203 (N_8203,N_7844,N_7191);
nand U8204 (N_8204,N_7939,N_7051);
and U8205 (N_8205,N_7867,N_7609);
and U8206 (N_8206,N_7700,N_7604);
nand U8207 (N_8207,N_7552,N_7689);
or U8208 (N_8208,N_7358,N_7543);
and U8209 (N_8209,N_7822,N_7144);
or U8210 (N_8210,N_7285,N_7933);
nor U8211 (N_8211,N_7076,N_7178);
nor U8212 (N_8212,N_7294,N_7903);
nor U8213 (N_8213,N_7509,N_7328);
nor U8214 (N_8214,N_7060,N_7769);
nand U8215 (N_8215,N_7303,N_7945);
nor U8216 (N_8216,N_7545,N_7713);
nor U8217 (N_8217,N_7611,N_7355);
or U8218 (N_8218,N_7360,N_7193);
nor U8219 (N_8219,N_7442,N_7584);
or U8220 (N_8220,N_7811,N_7145);
and U8221 (N_8221,N_7918,N_7247);
nand U8222 (N_8222,N_7382,N_7251);
and U8223 (N_8223,N_7955,N_7687);
nor U8224 (N_8224,N_7659,N_7776);
or U8225 (N_8225,N_7855,N_7080);
and U8226 (N_8226,N_7999,N_7866);
nand U8227 (N_8227,N_7708,N_7416);
nor U8228 (N_8228,N_7836,N_7027);
or U8229 (N_8229,N_7577,N_7469);
and U8230 (N_8230,N_7240,N_7612);
nor U8231 (N_8231,N_7241,N_7851);
or U8232 (N_8232,N_7953,N_7881);
and U8233 (N_8233,N_7110,N_7287);
nor U8234 (N_8234,N_7171,N_7295);
nor U8235 (N_8235,N_7845,N_7817);
nand U8236 (N_8236,N_7857,N_7808);
or U8237 (N_8237,N_7425,N_7753);
nor U8238 (N_8238,N_7291,N_7862);
and U8239 (N_8239,N_7780,N_7237);
nand U8240 (N_8240,N_7863,N_7896);
nand U8241 (N_8241,N_7242,N_7889);
and U8242 (N_8242,N_7377,N_7187);
nand U8243 (N_8243,N_7646,N_7983);
nor U8244 (N_8244,N_7562,N_7969);
nor U8245 (N_8245,N_7696,N_7814);
nor U8246 (N_8246,N_7463,N_7342);
and U8247 (N_8247,N_7433,N_7796);
and U8248 (N_8248,N_7036,N_7472);
or U8249 (N_8249,N_7056,N_7729);
xor U8250 (N_8250,N_7560,N_7792);
and U8251 (N_8251,N_7998,N_7274);
or U8252 (N_8252,N_7515,N_7246);
and U8253 (N_8253,N_7804,N_7470);
nor U8254 (N_8254,N_7147,N_7005);
nor U8255 (N_8255,N_7940,N_7653);
or U8256 (N_8256,N_7302,N_7556);
or U8257 (N_8257,N_7872,N_7572);
or U8258 (N_8258,N_7587,N_7266);
nor U8259 (N_8259,N_7257,N_7381);
nor U8260 (N_8260,N_7585,N_7906);
nor U8261 (N_8261,N_7884,N_7203);
nor U8262 (N_8262,N_7762,N_7298);
and U8263 (N_8263,N_7752,N_7248);
xor U8264 (N_8264,N_7259,N_7750);
nand U8265 (N_8265,N_7238,N_7392);
nand U8266 (N_8266,N_7813,N_7293);
nor U8267 (N_8267,N_7747,N_7950);
or U8268 (N_8268,N_7601,N_7828);
nand U8269 (N_8269,N_7183,N_7437);
nor U8270 (N_8270,N_7740,N_7047);
or U8271 (N_8271,N_7063,N_7231);
or U8272 (N_8272,N_7089,N_7588);
and U8273 (N_8273,N_7957,N_7798);
xor U8274 (N_8274,N_7987,N_7359);
nand U8275 (N_8275,N_7389,N_7167);
or U8276 (N_8276,N_7662,N_7698);
nand U8277 (N_8277,N_7189,N_7067);
and U8278 (N_8278,N_7743,N_7533);
nand U8279 (N_8279,N_7473,N_7233);
or U8280 (N_8280,N_7126,N_7680);
nand U8281 (N_8281,N_7608,N_7551);
nor U8282 (N_8282,N_7301,N_7083);
and U8283 (N_8283,N_7734,N_7525);
nor U8284 (N_8284,N_7235,N_7100);
and U8285 (N_8285,N_7834,N_7265);
nand U8286 (N_8286,N_7846,N_7660);
nand U8287 (N_8287,N_7949,N_7763);
and U8288 (N_8288,N_7094,N_7335);
nor U8289 (N_8289,N_7461,N_7802);
and U8290 (N_8290,N_7910,N_7504);
or U8291 (N_8291,N_7980,N_7555);
nor U8292 (N_8292,N_7789,N_7704);
and U8293 (N_8293,N_7337,N_7764);
nor U8294 (N_8294,N_7009,N_7315);
and U8295 (N_8295,N_7308,N_7405);
nand U8296 (N_8296,N_7672,N_7502);
and U8297 (N_8297,N_7650,N_7598);
nand U8298 (N_8298,N_7841,N_7967);
or U8299 (N_8299,N_7345,N_7232);
and U8300 (N_8300,N_7484,N_7255);
nor U8301 (N_8301,N_7378,N_7690);
nor U8302 (N_8302,N_7109,N_7314);
nor U8303 (N_8303,N_7717,N_7429);
nand U8304 (N_8304,N_7142,N_7099);
nor U8305 (N_8305,N_7334,N_7667);
and U8306 (N_8306,N_7590,N_7479);
or U8307 (N_8307,N_7571,N_7023);
nor U8308 (N_8308,N_7186,N_7480);
and U8309 (N_8309,N_7125,N_7017);
nand U8310 (N_8310,N_7006,N_7512);
and U8311 (N_8311,N_7118,N_7891);
nor U8312 (N_8312,N_7016,N_7837);
and U8313 (N_8313,N_7996,N_7245);
or U8314 (N_8314,N_7499,N_7919);
nor U8315 (N_8315,N_7449,N_7269);
nor U8316 (N_8316,N_7326,N_7982);
nand U8317 (N_8317,N_7858,N_7925);
nand U8318 (N_8318,N_7043,N_7965);
nand U8319 (N_8319,N_7510,N_7452);
or U8320 (N_8320,N_7620,N_7671);
nor U8321 (N_8321,N_7384,N_7835);
nor U8322 (N_8322,N_7218,N_7155);
nor U8323 (N_8323,N_7411,N_7008);
nand U8324 (N_8324,N_7250,N_7640);
or U8325 (N_8325,N_7091,N_7272);
and U8326 (N_8326,N_7074,N_7812);
nand U8327 (N_8327,N_7391,N_7438);
and U8328 (N_8328,N_7871,N_7182);
and U8329 (N_8329,N_7564,N_7923);
nor U8330 (N_8330,N_7079,N_7823);
nand U8331 (N_8331,N_7655,N_7112);
nor U8332 (N_8332,N_7158,N_7517);
nor U8333 (N_8333,N_7613,N_7782);
nor U8334 (N_8334,N_7760,N_7870);
or U8335 (N_8335,N_7230,N_7003);
nand U8336 (N_8336,N_7045,N_7897);
xnor U8337 (N_8337,N_7748,N_7134);
nor U8338 (N_8338,N_7458,N_7755);
and U8339 (N_8339,N_7664,N_7569);
xor U8340 (N_8340,N_7629,N_7369);
nor U8341 (N_8341,N_7370,N_7570);
nor U8342 (N_8342,N_7541,N_7772);
and U8343 (N_8343,N_7644,N_7042);
nor U8344 (N_8344,N_7786,N_7818);
or U8345 (N_8345,N_7485,N_7092);
nand U8346 (N_8346,N_7791,N_7521);
or U8347 (N_8347,N_7901,N_7210);
and U8348 (N_8348,N_7339,N_7129);
and U8349 (N_8349,N_7136,N_7075);
or U8350 (N_8350,N_7647,N_7402);
or U8351 (N_8351,N_7143,N_7356);
nor U8352 (N_8352,N_7859,N_7532);
and U8353 (N_8353,N_7365,N_7196);
and U8354 (N_8354,N_7911,N_7926);
nand U8355 (N_8355,N_7229,N_7319);
and U8356 (N_8356,N_7770,N_7462);
and U8357 (N_8357,N_7765,N_7292);
and U8358 (N_8358,N_7387,N_7244);
and U8359 (N_8359,N_7913,N_7228);
or U8360 (N_8360,N_7373,N_7974);
or U8361 (N_8361,N_7450,N_7174);
nand U8362 (N_8362,N_7131,N_7117);
or U8363 (N_8363,N_7528,N_7626);
nand U8364 (N_8364,N_7422,N_7111);
or U8365 (N_8365,N_7397,N_7526);
or U8366 (N_8366,N_7407,N_7267);
nand U8367 (N_8367,N_7488,N_7725);
nand U8368 (N_8368,N_7693,N_7015);
nand U8369 (N_8369,N_7026,N_7503);
or U8370 (N_8370,N_7712,N_7286);
or U8371 (N_8371,N_7321,N_7883);
nor U8372 (N_8372,N_7563,N_7430);
xor U8373 (N_8373,N_7451,N_7453);
nand U8374 (N_8374,N_7832,N_7362);
nor U8375 (N_8375,N_7225,N_7645);
and U8376 (N_8376,N_7284,N_7807);
or U8377 (N_8377,N_7800,N_7519);
or U8378 (N_8378,N_7966,N_7184);
and U8379 (N_8379,N_7239,N_7972);
or U8380 (N_8380,N_7960,N_7465);
and U8381 (N_8381,N_7544,N_7198);
nor U8382 (N_8382,N_7441,N_7124);
or U8383 (N_8383,N_7205,N_7025);
or U8384 (N_8384,N_7978,N_7034);
or U8385 (N_8385,N_7790,N_7200);
nor U8386 (N_8386,N_7505,N_7330);
nand U8387 (N_8387,N_7399,N_7106);
or U8388 (N_8388,N_7915,N_7958);
nand U8389 (N_8389,N_7114,N_7300);
nand U8390 (N_8390,N_7920,N_7310);
nand U8391 (N_8391,N_7803,N_7081);
nand U8392 (N_8392,N_7930,N_7482);
and U8393 (N_8393,N_7194,N_7794);
and U8394 (N_8394,N_7801,N_7886);
or U8395 (N_8395,N_7733,N_7619);
or U8396 (N_8396,N_7467,N_7179);
or U8397 (N_8397,N_7876,N_7256);
nand U8398 (N_8398,N_7408,N_7523);
xnor U8399 (N_8399,N_7414,N_7423);
and U8400 (N_8400,N_7599,N_7557);
or U8401 (N_8401,N_7146,N_7435);
nand U8402 (N_8402,N_7165,N_7661);
or U8403 (N_8403,N_7722,N_7148);
nand U8404 (N_8404,N_7217,N_7710);
xnor U8405 (N_8405,N_7368,N_7530);
or U8406 (N_8406,N_7962,N_7395);
nand U8407 (N_8407,N_7394,N_7046);
nand U8408 (N_8408,N_7058,N_7483);
nor U8409 (N_8409,N_7691,N_7654);
nor U8410 (N_8410,N_7868,N_7649);
or U8411 (N_8411,N_7021,N_7361);
or U8412 (N_8412,N_7213,N_7850);
and U8413 (N_8413,N_7367,N_7149);
nand U8414 (N_8414,N_7417,N_7806);
nand U8415 (N_8415,N_7290,N_7738);
xnor U8416 (N_8416,N_7160,N_7997);
or U8417 (N_8417,N_7677,N_7288);
nand U8418 (N_8418,N_7932,N_7324);
nor U8419 (N_8419,N_7869,N_7641);
nor U8420 (N_8420,N_7550,N_7249);
and U8421 (N_8421,N_7594,N_7057);
nand U8422 (N_8422,N_7243,N_7592);
and U8423 (N_8423,N_7434,N_7656);
nand U8424 (N_8424,N_7282,N_7518);
nand U8425 (N_8425,N_7721,N_7039);
nand U8426 (N_8426,N_7529,N_7150);
or U8427 (N_8427,N_7219,N_7327);
and U8428 (N_8428,N_7600,N_7296);
and U8429 (N_8429,N_7077,N_7513);
and U8430 (N_8430,N_7630,N_7318);
nor U8431 (N_8431,N_7064,N_7777);
nor U8432 (N_8432,N_7085,N_7307);
nand U8433 (N_8433,N_7084,N_7446);
and U8434 (N_8434,N_7366,N_7445);
and U8435 (N_8435,N_7768,N_7312);
nor U8436 (N_8436,N_7419,N_7947);
or U8437 (N_8437,N_7591,N_7279);
and U8438 (N_8438,N_7665,N_7676);
and U8439 (N_8439,N_7098,N_7827);
nand U8440 (N_8440,N_7403,N_7558);
nor U8441 (N_8441,N_7212,N_7767);
or U8442 (N_8442,N_7317,N_7701);
or U8443 (N_8443,N_7263,N_7936);
and U8444 (N_8444,N_7865,N_7705);
nand U8445 (N_8445,N_7204,N_7709);
nor U8446 (N_8446,N_7554,N_7737);
nand U8447 (N_8447,N_7815,N_7127);
nor U8448 (N_8448,N_7459,N_7185);
and U8449 (N_8449,N_7278,N_7283);
nand U8450 (N_8450,N_7749,N_7921);
and U8451 (N_8451,N_7014,N_7104);
nand U8452 (N_8452,N_7153,N_7253);
nor U8453 (N_8453,N_7152,N_7890);
nand U8454 (N_8454,N_7275,N_7976);
nor U8455 (N_8455,N_7088,N_7102);
or U8456 (N_8456,N_7050,N_7352);
nor U8457 (N_8457,N_7209,N_7164);
or U8458 (N_8458,N_7979,N_7372);
nor U8459 (N_8459,N_7542,N_7030);
or U8460 (N_8460,N_7444,N_7133);
nor U8461 (N_8461,N_7559,N_7576);
or U8462 (N_8462,N_7779,N_7895);
and U8463 (N_8463,N_7567,N_7694);
nand U8464 (N_8464,N_7123,N_7961);
and U8465 (N_8465,N_7401,N_7350);
and U8466 (N_8466,N_7348,N_7000);
nand U8467 (N_8467,N_7371,N_7948);
nand U8468 (N_8468,N_7548,N_7882);
nand U8469 (N_8469,N_7880,N_7475);
nand U8470 (N_8470,N_7670,N_7842);
or U8471 (N_8471,N_7311,N_7216);
nand U8472 (N_8472,N_7163,N_7374);
or U8473 (N_8473,N_7992,N_7531);
nand U8474 (N_8474,N_7658,N_7977);
or U8475 (N_8475,N_7703,N_7115);
nand U8476 (N_8476,N_7192,N_7833);
and U8477 (N_8477,N_7788,N_7685);
and U8478 (N_8478,N_7632,N_7439);
nor U8479 (N_8479,N_7539,N_7332);
or U8480 (N_8480,N_7761,N_7012);
xnor U8481 (N_8481,N_7214,N_7742);
or U8482 (N_8482,N_7702,N_7346);
and U8483 (N_8483,N_7113,N_7995);
nand U8484 (N_8484,N_7582,N_7973);
and U8485 (N_8485,N_7385,N_7968);
nor U8486 (N_8486,N_7309,N_7593);
nand U8487 (N_8487,N_7049,N_7306);
nor U8488 (N_8488,N_7809,N_7157);
nand U8489 (N_8489,N_7783,N_7991);
nand U8490 (N_8490,N_7757,N_7904);
or U8491 (N_8491,N_7412,N_7108);
or U8492 (N_8492,N_7325,N_7341);
nor U8493 (N_8493,N_7606,N_7491);
xnor U8494 (N_8494,N_7400,N_7860);
nand U8495 (N_8495,N_7466,N_7095);
or U8496 (N_8496,N_7759,N_7847);
or U8497 (N_8497,N_7874,N_7946);
nand U8498 (N_8498,N_7524,N_7002);
nor U8499 (N_8499,N_7719,N_7596);
nor U8500 (N_8500,N_7012,N_7918);
nand U8501 (N_8501,N_7402,N_7623);
xnor U8502 (N_8502,N_7949,N_7847);
nor U8503 (N_8503,N_7359,N_7048);
nor U8504 (N_8504,N_7376,N_7017);
nor U8505 (N_8505,N_7602,N_7702);
and U8506 (N_8506,N_7277,N_7376);
nand U8507 (N_8507,N_7014,N_7931);
or U8508 (N_8508,N_7625,N_7480);
nor U8509 (N_8509,N_7304,N_7661);
and U8510 (N_8510,N_7686,N_7088);
and U8511 (N_8511,N_7656,N_7475);
or U8512 (N_8512,N_7604,N_7665);
nand U8513 (N_8513,N_7607,N_7669);
nand U8514 (N_8514,N_7927,N_7955);
or U8515 (N_8515,N_7625,N_7732);
nand U8516 (N_8516,N_7098,N_7882);
and U8517 (N_8517,N_7223,N_7160);
nand U8518 (N_8518,N_7979,N_7750);
and U8519 (N_8519,N_7826,N_7954);
xnor U8520 (N_8520,N_7911,N_7987);
and U8521 (N_8521,N_7950,N_7427);
and U8522 (N_8522,N_7233,N_7770);
and U8523 (N_8523,N_7985,N_7787);
nand U8524 (N_8524,N_7141,N_7537);
nand U8525 (N_8525,N_7535,N_7167);
or U8526 (N_8526,N_7920,N_7434);
nor U8527 (N_8527,N_7372,N_7469);
nand U8528 (N_8528,N_7270,N_7314);
nand U8529 (N_8529,N_7199,N_7788);
nor U8530 (N_8530,N_7894,N_7597);
nand U8531 (N_8531,N_7675,N_7118);
nor U8532 (N_8532,N_7741,N_7381);
nor U8533 (N_8533,N_7234,N_7208);
or U8534 (N_8534,N_7123,N_7408);
and U8535 (N_8535,N_7754,N_7689);
or U8536 (N_8536,N_7156,N_7091);
and U8537 (N_8537,N_7533,N_7196);
nand U8538 (N_8538,N_7337,N_7005);
nand U8539 (N_8539,N_7252,N_7135);
nand U8540 (N_8540,N_7204,N_7990);
nand U8541 (N_8541,N_7223,N_7775);
and U8542 (N_8542,N_7993,N_7908);
or U8543 (N_8543,N_7082,N_7568);
nand U8544 (N_8544,N_7848,N_7010);
nor U8545 (N_8545,N_7307,N_7084);
nor U8546 (N_8546,N_7264,N_7241);
nand U8547 (N_8547,N_7031,N_7332);
nand U8548 (N_8548,N_7431,N_7790);
nand U8549 (N_8549,N_7481,N_7005);
nand U8550 (N_8550,N_7190,N_7795);
and U8551 (N_8551,N_7609,N_7227);
nor U8552 (N_8552,N_7998,N_7821);
nor U8553 (N_8553,N_7561,N_7546);
or U8554 (N_8554,N_7116,N_7419);
nor U8555 (N_8555,N_7826,N_7680);
and U8556 (N_8556,N_7941,N_7421);
nand U8557 (N_8557,N_7439,N_7339);
or U8558 (N_8558,N_7253,N_7553);
nor U8559 (N_8559,N_7643,N_7532);
or U8560 (N_8560,N_7778,N_7487);
nand U8561 (N_8561,N_7384,N_7624);
nor U8562 (N_8562,N_7775,N_7504);
or U8563 (N_8563,N_7716,N_7770);
or U8564 (N_8564,N_7071,N_7630);
nor U8565 (N_8565,N_7456,N_7811);
and U8566 (N_8566,N_7078,N_7966);
nand U8567 (N_8567,N_7394,N_7143);
nand U8568 (N_8568,N_7796,N_7835);
nand U8569 (N_8569,N_7857,N_7343);
and U8570 (N_8570,N_7364,N_7947);
nor U8571 (N_8571,N_7329,N_7730);
and U8572 (N_8572,N_7058,N_7133);
nor U8573 (N_8573,N_7080,N_7100);
nand U8574 (N_8574,N_7189,N_7397);
nand U8575 (N_8575,N_7643,N_7084);
or U8576 (N_8576,N_7863,N_7809);
nor U8577 (N_8577,N_7173,N_7864);
or U8578 (N_8578,N_7578,N_7553);
nand U8579 (N_8579,N_7539,N_7578);
or U8580 (N_8580,N_7252,N_7737);
or U8581 (N_8581,N_7050,N_7010);
nor U8582 (N_8582,N_7411,N_7268);
nand U8583 (N_8583,N_7317,N_7521);
nand U8584 (N_8584,N_7164,N_7926);
and U8585 (N_8585,N_7224,N_7587);
and U8586 (N_8586,N_7838,N_7789);
nor U8587 (N_8587,N_7777,N_7721);
nand U8588 (N_8588,N_7541,N_7046);
and U8589 (N_8589,N_7077,N_7821);
and U8590 (N_8590,N_7613,N_7905);
xor U8591 (N_8591,N_7500,N_7234);
nor U8592 (N_8592,N_7646,N_7235);
nor U8593 (N_8593,N_7004,N_7611);
and U8594 (N_8594,N_7925,N_7224);
nand U8595 (N_8595,N_7098,N_7431);
and U8596 (N_8596,N_7404,N_7688);
and U8597 (N_8597,N_7888,N_7232);
or U8598 (N_8598,N_7185,N_7644);
xor U8599 (N_8599,N_7572,N_7474);
xor U8600 (N_8600,N_7766,N_7562);
nand U8601 (N_8601,N_7501,N_7633);
nor U8602 (N_8602,N_7699,N_7723);
nand U8603 (N_8603,N_7722,N_7028);
xor U8604 (N_8604,N_7111,N_7011);
and U8605 (N_8605,N_7921,N_7091);
nand U8606 (N_8606,N_7874,N_7106);
nand U8607 (N_8607,N_7594,N_7181);
and U8608 (N_8608,N_7638,N_7306);
nor U8609 (N_8609,N_7936,N_7194);
nor U8610 (N_8610,N_7670,N_7712);
and U8611 (N_8611,N_7579,N_7042);
or U8612 (N_8612,N_7399,N_7513);
nor U8613 (N_8613,N_7697,N_7889);
nand U8614 (N_8614,N_7832,N_7332);
or U8615 (N_8615,N_7973,N_7808);
and U8616 (N_8616,N_7398,N_7812);
nor U8617 (N_8617,N_7905,N_7534);
nor U8618 (N_8618,N_7349,N_7885);
nor U8619 (N_8619,N_7465,N_7200);
or U8620 (N_8620,N_7607,N_7220);
nand U8621 (N_8621,N_7181,N_7964);
nand U8622 (N_8622,N_7903,N_7632);
or U8623 (N_8623,N_7252,N_7202);
nand U8624 (N_8624,N_7016,N_7509);
or U8625 (N_8625,N_7226,N_7518);
and U8626 (N_8626,N_7543,N_7100);
and U8627 (N_8627,N_7683,N_7525);
nand U8628 (N_8628,N_7673,N_7301);
or U8629 (N_8629,N_7070,N_7974);
nor U8630 (N_8630,N_7141,N_7360);
nor U8631 (N_8631,N_7674,N_7261);
nand U8632 (N_8632,N_7217,N_7989);
and U8633 (N_8633,N_7491,N_7199);
nand U8634 (N_8634,N_7710,N_7037);
and U8635 (N_8635,N_7474,N_7398);
nor U8636 (N_8636,N_7089,N_7773);
or U8637 (N_8637,N_7034,N_7441);
nand U8638 (N_8638,N_7883,N_7305);
or U8639 (N_8639,N_7410,N_7359);
nor U8640 (N_8640,N_7099,N_7016);
nand U8641 (N_8641,N_7923,N_7985);
nand U8642 (N_8642,N_7027,N_7015);
or U8643 (N_8643,N_7105,N_7851);
and U8644 (N_8644,N_7303,N_7949);
and U8645 (N_8645,N_7640,N_7870);
nand U8646 (N_8646,N_7016,N_7065);
or U8647 (N_8647,N_7647,N_7454);
or U8648 (N_8648,N_7680,N_7545);
and U8649 (N_8649,N_7995,N_7966);
nor U8650 (N_8650,N_7306,N_7448);
nor U8651 (N_8651,N_7322,N_7817);
and U8652 (N_8652,N_7121,N_7538);
or U8653 (N_8653,N_7819,N_7702);
xnor U8654 (N_8654,N_7200,N_7277);
nor U8655 (N_8655,N_7768,N_7993);
nand U8656 (N_8656,N_7470,N_7739);
nand U8657 (N_8657,N_7580,N_7838);
nand U8658 (N_8658,N_7753,N_7232);
or U8659 (N_8659,N_7814,N_7797);
nand U8660 (N_8660,N_7683,N_7565);
nand U8661 (N_8661,N_7497,N_7173);
or U8662 (N_8662,N_7941,N_7465);
nor U8663 (N_8663,N_7345,N_7922);
nor U8664 (N_8664,N_7901,N_7249);
nand U8665 (N_8665,N_7576,N_7734);
or U8666 (N_8666,N_7884,N_7031);
and U8667 (N_8667,N_7421,N_7123);
and U8668 (N_8668,N_7719,N_7770);
and U8669 (N_8669,N_7081,N_7848);
or U8670 (N_8670,N_7089,N_7164);
nor U8671 (N_8671,N_7183,N_7753);
nor U8672 (N_8672,N_7318,N_7317);
or U8673 (N_8673,N_7535,N_7848);
xnor U8674 (N_8674,N_7528,N_7593);
and U8675 (N_8675,N_7255,N_7430);
nand U8676 (N_8676,N_7761,N_7827);
nor U8677 (N_8677,N_7606,N_7834);
nor U8678 (N_8678,N_7434,N_7844);
or U8679 (N_8679,N_7169,N_7106);
and U8680 (N_8680,N_7373,N_7381);
nor U8681 (N_8681,N_7378,N_7038);
nand U8682 (N_8682,N_7403,N_7149);
or U8683 (N_8683,N_7702,N_7993);
nand U8684 (N_8684,N_7552,N_7863);
and U8685 (N_8685,N_7596,N_7414);
and U8686 (N_8686,N_7736,N_7795);
and U8687 (N_8687,N_7129,N_7282);
nand U8688 (N_8688,N_7263,N_7126);
nor U8689 (N_8689,N_7733,N_7147);
nor U8690 (N_8690,N_7895,N_7217);
nand U8691 (N_8691,N_7187,N_7926);
and U8692 (N_8692,N_7310,N_7571);
or U8693 (N_8693,N_7094,N_7529);
nor U8694 (N_8694,N_7276,N_7882);
nand U8695 (N_8695,N_7812,N_7047);
or U8696 (N_8696,N_7504,N_7218);
or U8697 (N_8697,N_7798,N_7885);
nand U8698 (N_8698,N_7783,N_7309);
and U8699 (N_8699,N_7716,N_7251);
nor U8700 (N_8700,N_7749,N_7085);
nand U8701 (N_8701,N_7294,N_7117);
or U8702 (N_8702,N_7491,N_7014);
or U8703 (N_8703,N_7687,N_7380);
nor U8704 (N_8704,N_7011,N_7266);
nand U8705 (N_8705,N_7739,N_7111);
and U8706 (N_8706,N_7360,N_7646);
or U8707 (N_8707,N_7369,N_7373);
or U8708 (N_8708,N_7137,N_7746);
nand U8709 (N_8709,N_7368,N_7772);
and U8710 (N_8710,N_7156,N_7227);
nand U8711 (N_8711,N_7803,N_7822);
nor U8712 (N_8712,N_7043,N_7702);
and U8713 (N_8713,N_7632,N_7964);
nand U8714 (N_8714,N_7797,N_7134);
and U8715 (N_8715,N_7624,N_7551);
and U8716 (N_8716,N_7367,N_7629);
nand U8717 (N_8717,N_7928,N_7656);
nor U8718 (N_8718,N_7063,N_7421);
and U8719 (N_8719,N_7949,N_7685);
nor U8720 (N_8720,N_7304,N_7460);
nor U8721 (N_8721,N_7432,N_7159);
and U8722 (N_8722,N_7204,N_7547);
or U8723 (N_8723,N_7007,N_7816);
nand U8724 (N_8724,N_7863,N_7147);
and U8725 (N_8725,N_7956,N_7465);
and U8726 (N_8726,N_7721,N_7005);
nor U8727 (N_8727,N_7654,N_7261);
and U8728 (N_8728,N_7129,N_7517);
nand U8729 (N_8729,N_7631,N_7925);
nand U8730 (N_8730,N_7603,N_7780);
nor U8731 (N_8731,N_7069,N_7648);
or U8732 (N_8732,N_7137,N_7990);
or U8733 (N_8733,N_7204,N_7332);
nor U8734 (N_8734,N_7177,N_7131);
nand U8735 (N_8735,N_7030,N_7924);
and U8736 (N_8736,N_7551,N_7659);
and U8737 (N_8737,N_7288,N_7929);
nand U8738 (N_8738,N_7520,N_7329);
xnor U8739 (N_8739,N_7072,N_7173);
or U8740 (N_8740,N_7260,N_7869);
and U8741 (N_8741,N_7371,N_7145);
nand U8742 (N_8742,N_7169,N_7210);
nand U8743 (N_8743,N_7773,N_7128);
and U8744 (N_8744,N_7157,N_7887);
nand U8745 (N_8745,N_7669,N_7611);
or U8746 (N_8746,N_7482,N_7276);
nand U8747 (N_8747,N_7358,N_7354);
nand U8748 (N_8748,N_7461,N_7783);
nor U8749 (N_8749,N_7316,N_7136);
nor U8750 (N_8750,N_7434,N_7135);
and U8751 (N_8751,N_7194,N_7546);
and U8752 (N_8752,N_7816,N_7810);
and U8753 (N_8753,N_7293,N_7450);
nand U8754 (N_8754,N_7681,N_7680);
or U8755 (N_8755,N_7137,N_7433);
and U8756 (N_8756,N_7477,N_7879);
or U8757 (N_8757,N_7707,N_7102);
or U8758 (N_8758,N_7604,N_7502);
nand U8759 (N_8759,N_7114,N_7855);
nand U8760 (N_8760,N_7641,N_7300);
nand U8761 (N_8761,N_7261,N_7621);
and U8762 (N_8762,N_7921,N_7416);
and U8763 (N_8763,N_7057,N_7504);
or U8764 (N_8764,N_7159,N_7251);
nand U8765 (N_8765,N_7552,N_7676);
and U8766 (N_8766,N_7675,N_7317);
nand U8767 (N_8767,N_7043,N_7563);
nor U8768 (N_8768,N_7509,N_7545);
nand U8769 (N_8769,N_7999,N_7119);
nand U8770 (N_8770,N_7561,N_7666);
nand U8771 (N_8771,N_7082,N_7779);
or U8772 (N_8772,N_7966,N_7042);
nor U8773 (N_8773,N_7062,N_7244);
or U8774 (N_8774,N_7739,N_7132);
nor U8775 (N_8775,N_7442,N_7628);
or U8776 (N_8776,N_7608,N_7322);
nand U8777 (N_8777,N_7511,N_7878);
nor U8778 (N_8778,N_7676,N_7489);
nand U8779 (N_8779,N_7014,N_7340);
and U8780 (N_8780,N_7707,N_7340);
nand U8781 (N_8781,N_7712,N_7872);
nor U8782 (N_8782,N_7916,N_7767);
or U8783 (N_8783,N_7612,N_7409);
nand U8784 (N_8784,N_7872,N_7809);
and U8785 (N_8785,N_7469,N_7045);
nor U8786 (N_8786,N_7006,N_7768);
and U8787 (N_8787,N_7109,N_7435);
xnor U8788 (N_8788,N_7238,N_7389);
and U8789 (N_8789,N_7670,N_7295);
or U8790 (N_8790,N_7078,N_7591);
or U8791 (N_8791,N_7210,N_7844);
nor U8792 (N_8792,N_7772,N_7029);
or U8793 (N_8793,N_7282,N_7818);
and U8794 (N_8794,N_7157,N_7920);
nor U8795 (N_8795,N_7577,N_7347);
nor U8796 (N_8796,N_7429,N_7301);
nor U8797 (N_8797,N_7382,N_7554);
xor U8798 (N_8798,N_7266,N_7693);
or U8799 (N_8799,N_7280,N_7042);
and U8800 (N_8800,N_7925,N_7423);
nor U8801 (N_8801,N_7459,N_7617);
or U8802 (N_8802,N_7622,N_7010);
nand U8803 (N_8803,N_7566,N_7530);
and U8804 (N_8804,N_7239,N_7400);
nor U8805 (N_8805,N_7968,N_7716);
nor U8806 (N_8806,N_7281,N_7497);
or U8807 (N_8807,N_7914,N_7585);
nor U8808 (N_8808,N_7512,N_7185);
nand U8809 (N_8809,N_7789,N_7467);
nor U8810 (N_8810,N_7726,N_7685);
or U8811 (N_8811,N_7134,N_7524);
nor U8812 (N_8812,N_7791,N_7652);
and U8813 (N_8813,N_7109,N_7719);
and U8814 (N_8814,N_7092,N_7889);
and U8815 (N_8815,N_7961,N_7897);
nand U8816 (N_8816,N_7964,N_7138);
and U8817 (N_8817,N_7680,N_7995);
nor U8818 (N_8818,N_7262,N_7186);
and U8819 (N_8819,N_7927,N_7916);
and U8820 (N_8820,N_7699,N_7581);
nand U8821 (N_8821,N_7067,N_7704);
or U8822 (N_8822,N_7567,N_7229);
and U8823 (N_8823,N_7411,N_7541);
and U8824 (N_8824,N_7851,N_7758);
and U8825 (N_8825,N_7387,N_7393);
and U8826 (N_8826,N_7916,N_7740);
nor U8827 (N_8827,N_7242,N_7374);
nand U8828 (N_8828,N_7112,N_7637);
and U8829 (N_8829,N_7797,N_7686);
or U8830 (N_8830,N_7882,N_7037);
or U8831 (N_8831,N_7429,N_7202);
xor U8832 (N_8832,N_7965,N_7549);
nand U8833 (N_8833,N_7248,N_7217);
and U8834 (N_8834,N_7345,N_7675);
nand U8835 (N_8835,N_7496,N_7067);
or U8836 (N_8836,N_7890,N_7760);
nor U8837 (N_8837,N_7903,N_7987);
or U8838 (N_8838,N_7924,N_7370);
and U8839 (N_8839,N_7756,N_7035);
or U8840 (N_8840,N_7623,N_7923);
nor U8841 (N_8841,N_7085,N_7879);
or U8842 (N_8842,N_7916,N_7428);
nor U8843 (N_8843,N_7338,N_7677);
nor U8844 (N_8844,N_7990,N_7898);
and U8845 (N_8845,N_7297,N_7669);
nand U8846 (N_8846,N_7979,N_7036);
nand U8847 (N_8847,N_7301,N_7436);
nand U8848 (N_8848,N_7318,N_7559);
nand U8849 (N_8849,N_7231,N_7503);
or U8850 (N_8850,N_7275,N_7367);
and U8851 (N_8851,N_7299,N_7087);
nand U8852 (N_8852,N_7955,N_7138);
nor U8853 (N_8853,N_7261,N_7258);
nand U8854 (N_8854,N_7544,N_7166);
or U8855 (N_8855,N_7315,N_7080);
or U8856 (N_8856,N_7112,N_7196);
nor U8857 (N_8857,N_7659,N_7650);
nand U8858 (N_8858,N_7543,N_7015);
or U8859 (N_8859,N_7941,N_7451);
nor U8860 (N_8860,N_7095,N_7698);
nor U8861 (N_8861,N_7647,N_7544);
or U8862 (N_8862,N_7348,N_7313);
nor U8863 (N_8863,N_7395,N_7914);
or U8864 (N_8864,N_7960,N_7975);
nor U8865 (N_8865,N_7708,N_7875);
nor U8866 (N_8866,N_7749,N_7207);
nor U8867 (N_8867,N_7811,N_7193);
xor U8868 (N_8868,N_7744,N_7817);
and U8869 (N_8869,N_7422,N_7151);
nand U8870 (N_8870,N_7514,N_7535);
and U8871 (N_8871,N_7310,N_7635);
or U8872 (N_8872,N_7655,N_7539);
nor U8873 (N_8873,N_7127,N_7473);
nor U8874 (N_8874,N_7007,N_7510);
and U8875 (N_8875,N_7685,N_7684);
nand U8876 (N_8876,N_7633,N_7438);
nor U8877 (N_8877,N_7055,N_7682);
and U8878 (N_8878,N_7575,N_7326);
nor U8879 (N_8879,N_7133,N_7916);
and U8880 (N_8880,N_7887,N_7338);
or U8881 (N_8881,N_7719,N_7373);
nand U8882 (N_8882,N_7394,N_7088);
and U8883 (N_8883,N_7733,N_7775);
or U8884 (N_8884,N_7594,N_7060);
nand U8885 (N_8885,N_7691,N_7289);
or U8886 (N_8886,N_7240,N_7058);
and U8887 (N_8887,N_7552,N_7893);
xnor U8888 (N_8888,N_7749,N_7440);
nand U8889 (N_8889,N_7783,N_7399);
and U8890 (N_8890,N_7692,N_7398);
nor U8891 (N_8891,N_7129,N_7361);
nor U8892 (N_8892,N_7062,N_7377);
nor U8893 (N_8893,N_7064,N_7280);
nand U8894 (N_8894,N_7327,N_7822);
nand U8895 (N_8895,N_7070,N_7930);
and U8896 (N_8896,N_7601,N_7046);
or U8897 (N_8897,N_7379,N_7858);
or U8898 (N_8898,N_7744,N_7806);
nand U8899 (N_8899,N_7139,N_7134);
nand U8900 (N_8900,N_7776,N_7890);
nand U8901 (N_8901,N_7969,N_7982);
nand U8902 (N_8902,N_7409,N_7869);
or U8903 (N_8903,N_7420,N_7321);
nand U8904 (N_8904,N_7820,N_7040);
nor U8905 (N_8905,N_7327,N_7973);
and U8906 (N_8906,N_7123,N_7567);
or U8907 (N_8907,N_7132,N_7196);
or U8908 (N_8908,N_7792,N_7751);
nand U8909 (N_8909,N_7151,N_7187);
nor U8910 (N_8910,N_7482,N_7531);
nor U8911 (N_8911,N_7159,N_7300);
and U8912 (N_8912,N_7668,N_7285);
nand U8913 (N_8913,N_7376,N_7420);
or U8914 (N_8914,N_7063,N_7827);
nand U8915 (N_8915,N_7150,N_7251);
or U8916 (N_8916,N_7998,N_7171);
nand U8917 (N_8917,N_7369,N_7740);
nor U8918 (N_8918,N_7861,N_7703);
and U8919 (N_8919,N_7170,N_7091);
nand U8920 (N_8920,N_7171,N_7831);
nor U8921 (N_8921,N_7572,N_7869);
xor U8922 (N_8922,N_7842,N_7648);
nand U8923 (N_8923,N_7607,N_7058);
and U8924 (N_8924,N_7856,N_7344);
nand U8925 (N_8925,N_7354,N_7882);
nand U8926 (N_8926,N_7301,N_7452);
and U8927 (N_8927,N_7207,N_7425);
xnor U8928 (N_8928,N_7798,N_7167);
nor U8929 (N_8929,N_7679,N_7514);
nand U8930 (N_8930,N_7321,N_7912);
and U8931 (N_8931,N_7422,N_7373);
and U8932 (N_8932,N_7729,N_7233);
nand U8933 (N_8933,N_7282,N_7458);
or U8934 (N_8934,N_7834,N_7255);
or U8935 (N_8935,N_7500,N_7755);
nand U8936 (N_8936,N_7700,N_7123);
or U8937 (N_8937,N_7253,N_7988);
nand U8938 (N_8938,N_7055,N_7452);
nand U8939 (N_8939,N_7445,N_7481);
nor U8940 (N_8940,N_7656,N_7776);
nand U8941 (N_8941,N_7745,N_7778);
or U8942 (N_8942,N_7902,N_7801);
nand U8943 (N_8943,N_7174,N_7059);
nor U8944 (N_8944,N_7937,N_7879);
or U8945 (N_8945,N_7604,N_7799);
and U8946 (N_8946,N_7888,N_7458);
or U8947 (N_8947,N_7041,N_7715);
nand U8948 (N_8948,N_7175,N_7470);
xor U8949 (N_8949,N_7111,N_7288);
nand U8950 (N_8950,N_7021,N_7067);
or U8951 (N_8951,N_7466,N_7467);
and U8952 (N_8952,N_7204,N_7956);
or U8953 (N_8953,N_7263,N_7705);
nor U8954 (N_8954,N_7163,N_7469);
or U8955 (N_8955,N_7495,N_7067);
and U8956 (N_8956,N_7807,N_7711);
and U8957 (N_8957,N_7315,N_7310);
nand U8958 (N_8958,N_7344,N_7474);
and U8959 (N_8959,N_7507,N_7814);
or U8960 (N_8960,N_7236,N_7467);
nor U8961 (N_8961,N_7682,N_7263);
nand U8962 (N_8962,N_7636,N_7090);
or U8963 (N_8963,N_7166,N_7265);
or U8964 (N_8964,N_7409,N_7895);
nor U8965 (N_8965,N_7616,N_7014);
nand U8966 (N_8966,N_7173,N_7610);
nor U8967 (N_8967,N_7219,N_7011);
nor U8968 (N_8968,N_7473,N_7345);
nor U8969 (N_8969,N_7193,N_7470);
nand U8970 (N_8970,N_7336,N_7510);
or U8971 (N_8971,N_7279,N_7612);
or U8972 (N_8972,N_7354,N_7206);
nand U8973 (N_8973,N_7790,N_7440);
nor U8974 (N_8974,N_7426,N_7075);
or U8975 (N_8975,N_7602,N_7595);
nand U8976 (N_8976,N_7916,N_7452);
nand U8977 (N_8977,N_7268,N_7654);
and U8978 (N_8978,N_7255,N_7149);
nor U8979 (N_8979,N_7227,N_7087);
and U8980 (N_8980,N_7885,N_7839);
nand U8981 (N_8981,N_7267,N_7188);
and U8982 (N_8982,N_7114,N_7451);
or U8983 (N_8983,N_7972,N_7817);
and U8984 (N_8984,N_7967,N_7579);
nand U8985 (N_8985,N_7474,N_7080);
nand U8986 (N_8986,N_7141,N_7293);
nand U8987 (N_8987,N_7422,N_7890);
xnor U8988 (N_8988,N_7207,N_7400);
or U8989 (N_8989,N_7504,N_7637);
nor U8990 (N_8990,N_7015,N_7634);
or U8991 (N_8991,N_7438,N_7567);
and U8992 (N_8992,N_7231,N_7725);
nand U8993 (N_8993,N_7057,N_7098);
nor U8994 (N_8994,N_7194,N_7246);
or U8995 (N_8995,N_7711,N_7643);
and U8996 (N_8996,N_7845,N_7515);
nor U8997 (N_8997,N_7303,N_7490);
nand U8998 (N_8998,N_7120,N_7153);
and U8999 (N_8999,N_7169,N_7924);
nand U9000 (N_9000,N_8495,N_8965);
and U9001 (N_9001,N_8781,N_8615);
and U9002 (N_9002,N_8482,N_8047);
nor U9003 (N_9003,N_8807,N_8991);
or U9004 (N_9004,N_8531,N_8560);
nand U9005 (N_9005,N_8472,N_8518);
nand U9006 (N_9006,N_8066,N_8585);
or U9007 (N_9007,N_8019,N_8891);
or U9008 (N_9008,N_8245,N_8786);
nand U9009 (N_9009,N_8029,N_8312);
or U9010 (N_9010,N_8878,N_8406);
and U9011 (N_9011,N_8246,N_8349);
nand U9012 (N_9012,N_8517,N_8475);
nand U9013 (N_9013,N_8831,N_8005);
or U9014 (N_9014,N_8497,N_8871);
xor U9015 (N_9015,N_8409,N_8253);
nand U9016 (N_9016,N_8554,N_8895);
or U9017 (N_9017,N_8944,N_8684);
nor U9018 (N_9018,N_8700,N_8673);
or U9019 (N_9019,N_8424,N_8721);
and U9020 (N_9020,N_8707,N_8445);
and U9021 (N_9021,N_8319,N_8439);
nand U9022 (N_9022,N_8160,N_8830);
nor U9023 (N_9023,N_8462,N_8293);
nor U9024 (N_9024,N_8714,N_8893);
nor U9025 (N_9025,N_8260,N_8399);
nor U9026 (N_9026,N_8427,N_8182);
and U9027 (N_9027,N_8110,N_8656);
or U9028 (N_9028,N_8872,N_8125);
or U9029 (N_9029,N_8239,N_8494);
or U9030 (N_9030,N_8777,N_8244);
nor U9031 (N_9031,N_8078,N_8114);
nor U9032 (N_9032,N_8403,N_8351);
or U9033 (N_9033,N_8612,N_8958);
and U9034 (N_9034,N_8559,N_8799);
and U9035 (N_9035,N_8867,N_8402);
nand U9036 (N_9036,N_8746,N_8869);
or U9037 (N_9037,N_8247,N_8167);
nand U9038 (N_9038,N_8618,N_8410);
nand U9039 (N_9039,N_8546,N_8331);
or U9040 (N_9040,N_8436,N_8583);
or U9041 (N_9041,N_8873,N_8542);
nand U9042 (N_9042,N_8011,N_8390);
and U9043 (N_9043,N_8506,N_8766);
nand U9044 (N_9044,N_8910,N_8842);
nand U9045 (N_9045,N_8291,N_8051);
and U9046 (N_9046,N_8039,N_8921);
nor U9047 (N_9047,N_8566,N_8083);
xnor U9048 (N_9048,N_8270,N_8116);
nor U9049 (N_9049,N_8596,N_8562);
xnor U9050 (N_9050,N_8798,N_8238);
and U9051 (N_9051,N_8325,N_8505);
or U9052 (N_9052,N_8520,N_8864);
nor U9053 (N_9053,N_8170,N_8633);
or U9054 (N_9054,N_8426,N_8880);
or U9055 (N_9055,N_8067,N_8852);
and U9056 (N_9056,N_8180,N_8552);
nand U9057 (N_9057,N_8865,N_8833);
nand U9058 (N_9058,N_8323,N_8686);
or U9059 (N_9059,N_8313,N_8041);
nand U9060 (N_9060,N_8575,N_8311);
nor U9061 (N_9061,N_8079,N_8257);
and U9062 (N_9062,N_8452,N_8979);
nor U9063 (N_9063,N_8630,N_8151);
and U9064 (N_9064,N_8671,N_8455);
or U9065 (N_9065,N_8000,N_8908);
and U9066 (N_9066,N_8272,N_8780);
or U9067 (N_9067,N_8332,N_8756);
or U9068 (N_9068,N_8059,N_8330);
or U9069 (N_9069,N_8165,N_8776);
or U9070 (N_9070,N_8973,N_8415);
nand U9071 (N_9071,N_8148,N_8102);
and U9072 (N_9072,N_8928,N_8234);
nand U9073 (N_9073,N_8778,N_8056);
or U9074 (N_9074,N_8933,N_8248);
nand U9075 (N_9075,N_8666,N_8845);
nand U9076 (N_9076,N_8335,N_8922);
xor U9077 (N_9077,N_8077,N_8353);
nor U9078 (N_9078,N_8451,N_8740);
or U9079 (N_9079,N_8704,N_8856);
or U9080 (N_9080,N_8722,N_8184);
nor U9081 (N_9081,N_8699,N_8140);
or U9082 (N_9082,N_8192,N_8537);
nand U9083 (N_9083,N_8936,N_8860);
nor U9084 (N_9084,N_8315,N_8577);
nand U9085 (N_9085,N_8914,N_8525);
or U9086 (N_9086,N_8144,N_8139);
nand U9087 (N_9087,N_8843,N_8678);
or U9088 (N_9088,N_8717,N_8826);
nor U9089 (N_9089,N_8773,N_8681);
or U9090 (N_9090,N_8096,N_8121);
and U9091 (N_9091,N_8587,N_8753);
nand U9092 (N_9092,N_8477,N_8212);
nand U9093 (N_9093,N_8025,N_8689);
nand U9094 (N_9094,N_8154,N_8365);
or U9095 (N_9095,N_8129,N_8599);
or U9096 (N_9096,N_8688,N_8900);
or U9097 (N_9097,N_8638,N_8413);
and U9098 (N_9098,N_8358,N_8610);
or U9099 (N_9099,N_8098,N_8909);
or U9100 (N_9100,N_8956,N_8131);
and U9101 (N_9101,N_8061,N_8044);
or U9102 (N_9102,N_8109,N_8423);
nor U9103 (N_9103,N_8267,N_8836);
nand U9104 (N_9104,N_8580,N_8304);
nand U9105 (N_9105,N_8122,N_8821);
and U9106 (N_9106,N_8658,N_8660);
nor U9107 (N_9107,N_8655,N_8713);
nor U9108 (N_9108,N_8173,N_8355);
nor U9109 (N_9109,N_8190,N_8251);
or U9110 (N_9110,N_8411,N_8146);
and U9111 (N_9111,N_8511,N_8254);
nand U9112 (N_9112,N_8829,N_8977);
nor U9113 (N_9113,N_8334,N_8737);
xnor U9114 (N_9114,N_8668,N_8017);
nor U9115 (N_9115,N_8646,N_8393);
and U9116 (N_9116,N_8504,N_8593);
and U9117 (N_9117,N_8348,N_8280);
and U9118 (N_9118,N_8380,N_8811);
and U9119 (N_9119,N_8028,N_8748);
or U9120 (N_9120,N_8158,N_8589);
or U9121 (N_9121,N_8598,N_8651);
nor U9122 (N_9122,N_8529,N_8986);
and U9123 (N_9123,N_8950,N_8645);
nor U9124 (N_9124,N_8389,N_8999);
nor U9125 (N_9125,N_8614,N_8720);
nor U9126 (N_9126,N_8458,N_8161);
nor U9127 (N_9127,N_8698,N_8441);
nand U9128 (N_9128,N_8567,N_8855);
nand U9129 (N_9129,N_8913,N_8002);
or U9130 (N_9130,N_8219,N_8931);
nand U9131 (N_9131,N_8882,N_8715);
and U9132 (N_9132,N_8020,N_8107);
or U9133 (N_9133,N_8747,N_8540);
and U9134 (N_9134,N_8754,N_8514);
and U9135 (N_9135,N_8849,N_8222);
nor U9136 (N_9136,N_8240,N_8927);
nand U9137 (N_9137,N_8549,N_8954);
nor U9138 (N_9138,N_8679,N_8249);
and U9139 (N_9139,N_8591,N_8648);
nor U9140 (N_9140,N_8091,N_8230);
nand U9141 (N_9141,N_8227,N_8308);
or U9142 (N_9142,N_8602,N_8428);
xnor U9143 (N_9143,N_8417,N_8003);
xnor U9144 (N_9144,N_8968,N_8664);
or U9145 (N_9145,N_8816,N_8734);
and U9146 (N_9146,N_8045,N_8062);
nand U9147 (N_9147,N_8310,N_8214);
and U9148 (N_9148,N_8563,N_8463);
nand U9149 (N_9149,N_8285,N_8388);
and U9150 (N_9150,N_8444,N_8983);
or U9151 (N_9151,N_8084,N_8752);
and U9152 (N_9152,N_8669,N_8641);
and U9153 (N_9153,N_8705,N_8031);
nand U9154 (N_9154,N_8738,N_8534);
nor U9155 (N_9155,N_8034,N_8204);
and U9156 (N_9156,N_8586,N_8609);
nor U9157 (N_9157,N_8347,N_8763);
nor U9158 (N_9158,N_8547,N_8590);
nor U9159 (N_9159,N_8022,N_8181);
xnor U9160 (N_9160,N_8619,N_8229);
nand U9161 (N_9161,N_8461,N_8023);
nor U9162 (N_9162,N_8431,N_8551);
nand U9163 (N_9163,N_8299,N_8739);
and U9164 (N_9164,N_8123,N_8419);
nand U9165 (N_9165,N_8576,N_8652);
nor U9166 (N_9166,N_8814,N_8450);
or U9167 (N_9167,N_8509,N_8564);
nor U9168 (N_9168,N_8446,N_8064);
and U9169 (N_9169,N_8997,N_8356);
nand U9170 (N_9170,N_8368,N_8142);
nand U9171 (N_9171,N_8653,N_8952);
or U9172 (N_9172,N_8288,N_8111);
or U9173 (N_9173,N_8876,N_8962);
and U9174 (N_9174,N_8386,N_8322);
or U9175 (N_9175,N_8101,N_8866);
nand U9176 (N_9176,N_8099,N_8510);
or U9177 (N_9177,N_8065,N_8834);
or U9178 (N_9178,N_8074,N_8336);
nand U9179 (N_9179,N_8301,N_8758);
nor U9180 (N_9180,N_8634,N_8087);
or U9181 (N_9181,N_8861,N_8527);
nor U9182 (N_9182,N_8667,N_8287);
nand U9183 (N_9183,N_8076,N_8725);
nand U9184 (N_9184,N_8581,N_8906);
nand U9185 (N_9185,N_8957,N_8964);
nand U9186 (N_9186,N_8213,N_8135);
and U9187 (N_9187,N_8680,N_8736);
or U9188 (N_9188,N_8178,N_8631);
or U9189 (N_9189,N_8476,N_8785);
nand U9190 (N_9190,N_8490,N_8262);
nor U9191 (N_9191,N_8414,N_8210);
nor U9192 (N_9192,N_8108,N_8430);
xnor U9193 (N_9193,N_8920,N_8750);
or U9194 (N_9194,N_8007,N_8532);
and U9195 (N_9195,N_8881,N_8055);
nor U9196 (N_9196,N_8751,N_8092);
and U9197 (N_9197,N_8276,N_8762);
nor U9198 (N_9198,N_8073,N_8996);
or U9199 (N_9199,N_8706,N_8471);
nor U9200 (N_9200,N_8294,N_8729);
nor U9201 (N_9201,N_8810,N_8982);
and U9202 (N_9202,N_8685,N_8787);
nor U9203 (N_9203,N_8256,N_8775);
nand U9204 (N_9204,N_8650,N_8376);
and U9205 (N_9205,N_8940,N_8360);
nand U9206 (N_9206,N_8097,N_8460);
nand U9207 (N_9207,N_8292,N_8026);
nand U9208 (N_9208,N_8694,N_8903);
nor U9209 (N_9209,N_8788,N_8106);
or U9210 (N_9210,N_8021,N_8544);
or U9211 (N_9211,N_8263,N_8277);
or U9212 (N_9212,N_8594,N_8624);
nor U9213 (N_9213,N_8493,N_8200);
and U9214 (N_9214,N_8442,N_8710);
nand U9215 (N_9215,N_8636,N_8635);
nand U9216 (N_9216,N_8243,N_8372);
nor U9217 (N_9217,N_8533,N_8858);
nand U9218 (N_9218,N_8480,N_8177);
nand U9219 (N_9219,N_8328,N_8851);
and U9220 (N_9220,N_8896,N_8735);
nand U9221 (N_9221,N_8792,N_8392);
nor U9222 (N_9222,N_8261,N_8582);
nor U9223 (N_9223,N_8757,N_8049);
nor U9224 (N_9224,N_8179,N_8004);
and U9225 (N_9225,N_8640,N_8132);
and U9226 (N_9226,N_8993,N_8216);
or U9227 (N_9227,N_8877,N_8769);
xor U9228 (N_9228,N_8693,N_8429);
or U9229 (N_9229,N_8696,N_8013);
nand U9230 (N_9230,N_8503,N_8159);
and U9231 (N_9231,N_8467,N_8946);
xor U9232 (N_9232,N_8823,N_8266);
and U9233 (N_9233,N_8265,N_8874);
nor U9234 (N_9234,N_8597,N_8934);
nor U9235 (N_9235,N_8479,N_8683);
nand U9236 (N_9236,N_8942,N_8223);
nor U9237 (N_9237,N_8366,N_8115);
and U9238 (N_9238,N_8592,N_8932);
nand U9239 (N_9239,N_8456,N_8344);
or U9240 (N_9240,N_8507,N_8837);
and U9241 (N_9241,N_8117,N_8432);
nor U9242 (N_9242,N_8745,N_8723);
and U9243 (N_9243,N_8879,N_8929);
xor U9244 (N_9244,N_8892,N_8042);
and U9245 (N_9245,N_8481,N_8508);
nand U9246 (N_9246,N_8938,N_8072);
and U9247 (N_9247,N_8795,N_8283);
nand U9248 (N_9248,N_8327,N_8220);
nand U9249 (N_9249,N_8500,N_8483);
and U9250 (N_9250,N_8457,N_8412);
nand U9251 (N_9251,N_8088,N_8989);
and U9252 (N_9252,N_8278,N_8888);
or U9253 (N_9253,N_8697,N_8603);
or U9254 (N_9254,N_8080,N_8206);
and U9255 (N_9255,N_8443,N_8250);
and U9256 (N_9256,N_8295,N_8231);
or U9257 (N_9257,N_8832,N_8466);
nor U9258 (N_9258,N_8579,N_8183);
or U9259 (N_9259,N_8050,N_8447);
nand U9260 (N_9260,N_8790,N_8967);
xor U9261 (N_9261,N_8215,N_8126);
or U9262 (N_9262,N_8164,N_8813);
nor U9263 (N_9263,N_8298,N_8516);
or U9264 (N_9264,N_8492,N_8208);
or U9265 (N_9265,N_8286,N_8155);
nand U9266 (N_9266,N_8054,N_8438);
nand U9267 (N_9267,N_8556,N_8515);
nand U9268 (N_9268,N_8535,N_8625);
nand U9269 (N_9269,N_8118,N_8175);
nor U9270 (N_9270,N_8548,N_8743);
and U9271 (N_9271,N_8841,N_8662);
and U9272 (N_9272,N_8197,N_8281);
and U9273 (N_9273,N_8375,N_8338);
and U9274 (N_9274,N_8712,N_8887);
and U9275 (N_9275,N_8082,N_8574);
and U9276 (N_9276,N_8524,N_8812);
and U9277 (N_9277,N_8385,N_8953);
or U9278 (N_9278,N_8174,N_8571);
nor U9279 (N_9279,N_8622,N_8644);
nand U9280 (N_9280,N_8677,N_8782);
nor U9281 (N_9281,N_8519,N_8468);
nand U9282 (N_9282,N_8530,N_8632);
and U9283 (N_9283,N_8218,N_8052);
nor U9284 (N_9284,N_8682,N_8407);
nand U9285 (N_9285,N_8804,N_8955);
or U9286 (N_9286,N_8333,N_8642);
nand U9287 (N_9287,N_8271,N_8889);
or U9288 (N_9288,N_8422,N_8819);
nor U9289 (N_9289,N_8708,N_8395);
nor U9290 (N_9290,N_8844,N_8649);
nand U9291 (N_9291,N_8352,N_8543);
nand U9292 (N_9292,N_8018,N_8731);
or U9293 (N_9293,N_8241,N_8194);
nand U9294 (N_9294,N_8767,N_8089);
nand U9295 (N_9295,N_8329,N_8086);
nand U9296 (N_9296,N_8371,N_8512);
and U9297 (N_9297,N_8558,N_8302);
nand U9298 (N_9298,N_8528,N_8522);
and U9299 (N_9299,N_8998,N_8398);
or U9300 (N_9300,N_8454,N_8898);
or U9301 (N_9301,N_8561,N_8195);
nor U9302 (N_9302,N_8744,N_8339);
or U9303 (N_9303,N_8217,N_8453);
nor U9304 (N_9304,N_8188,N_8912);
or U9305 (N_9305,N_8692,N_8611);
and U9306 (N_9306,N_8526,N_8771);
and U9307 (N_9307,N_8268,N_8755);
and U9308 (N_9308,N_8824,N_8153);
nand U9309 (N_9309,N_8149,N_8570);
nor U9310 (N_9310,N_8848,N_8133);
or U9311 (N_9311,N_8970,N_8237);
nor U9312 (N_9312,N_8850,N_8770);
nand U9313 (N_9313,N_8923,N_8185);
or U9314 (N_9314,N_8449,N_8926);
or U9315 (N_9315,N_8890,N_8259);
or U9316 (N_9316,N_8601,N_8724);
nand U9317 (N_9317,N_8040,N_8783);
nor U9318 (N_9318,N_8797,N_8727);
nor U9319 (N_9319,N_8637,N_8225);
or U9320 (N_9320,N_8433,N_8951);
nor U9321 (N_9321,N_8759,N_8036);
or U9322 (N_9322,N_8363,N_8015);
nor U9323 (N_9323,N_8321,N_8925);
nor U9324 (N_9324,N_8969,N_8916);
or U9325 (N_9325,N_8233,N_8943);
and U9326 (N_9326,N_8112,N_8469);
and U9327 (N_9327,N_8136,N_8796);
nand U9328 (N_9328,N_8090,N_8772);
nand U9329 (N_9329,N_8255,N_8202);
nor U9330 (N_9330,N_8141,N_8350);
or U9331 (N_9331,N_8354,N_8760);
or U9332 (N_9332,N_8357,N_8378);
nand U9333 (N_9333,N_8282,N_8657);
or U9334 (N_9334,N_8341,N_8960);
nor U9335 (N_9335,N_8030,N_8342);
or U9336 (N_9336,N_8397,N_8186);
and U9337 (N_9337,N_8822,N_8404);
and U9338 (N_9338,N_8242,N_8550);
and U9339 (N_9339,N_8818,N_8536);
or U9340 (N_9340,N_8345,N_8124);
nor U9341 (N_9341,N_8057,N_8555);
xor U9342 (N_9342,N_8726,N_8768);
nor U9343 (N_9343,N_8038,N_8401);
or U9344 (N_9344,N_8221,N_8075);
or U9345 (N_9345,N_8486,N_8616);
nor U9346 (N_9346,N_8690,N_8169);
and U9347 (N_9347,N_8963,N_8434);
nor U9348 (N_9348,N_8209,N_8847);
nor U9349 (N_9349,N_8578,N_8435);
or U9350 (N_9350,N_8974,N_8670);
or U9351 (N_9351,N_8806,N_8672);
nand U9352 (N_9352,N_8538,N_8761);
nor U9353 (N_9353,N_8498,N_8961);
nor U9354 (N_9354,N_8626,N_8306);
and U9355 (N_9355,N_8289,N_8416);
nor U9356 (N_9356,N_8382,N_8917);
nor U9357 (N_9357,N_8885,N_8779);
or U9358 (N_9358,N_8211,N_8465);
and U9359 (N_9359,N_8691,N_8975);
nand U9360 (N_9360,N_8120,N_8043);
and U9361 (N_9361,N_8857,N_8228);
and U9362 (N_9362,N_8584,N_8553);
or U9363 (N_9363,N_8608,N_8408);
nor U9364 (N_9364,N_8474,N_8623);
or U9365 (N_9365,N_8907,N_8919);
and U9366 (N_9366,N_8605,N_8911);
nor U9367 (N_9367,N_8071,N_8701);
nor U9368 (N_9368,N_8016,N_8915);
nand U9369 (N_9369,N_8440,N_8361);
and U9370 (N_9370,N_8703,N_8905);
nand U9371 (N_9371,N_8496,N_8168);
and U9372 (N_9372,N_8809,N_8484);
nand U9373 (N_9373,N_8854,N_8825);
nand U9374 (N_9374,N_8595,N_8765);
nand U9375 (N_9375,N_8143,N_8545);
and U9376 (N_9376,N_8718,N_8318);
and U9377 (N_9377,N_8128,N_8199);
and U9378 (N_9378,N_8130,N_8094);
or U9379 (N_9379,N_8226,N_8499);
nand U9380 (N_9380,N_8945,N_8053);
and U9381 (N_9381,N_8647,N_8374);
nand U9382 (N_9382,N_8104,N_8048);
and U9383 (N_9383,N_8749,N_8687);
nor U9384 (N_9384,N_8617,N_8478);
nand U9385 (N_9385,N_8137,N_8317);
or U9386 (N_9386,N_8764,N_8805);
xnor U9387 (N_9387,N_8001,N_8364);
or U9388 (N_9388,N_8604,N_8939);
nand U9389 (N_9389,N_8033,N_8162);
or U9390 (N_9390,N_8070,N_8274);
and U9391 (N_9391,N_8676,N_8992);
or U9392 (N_9392,N_8305,N_8949);
or U9393 (N_9393,N_8904,N_8901);
or U9394 (N_9394,N_8163,N_8793);
and U9395 (N_9395,N_8176,N_8326);
and U9396 (N_9396,N_8935,N_8362);
and U9397 (N_9397,N_8269,N_8972);
and U9398 (N_9398,N_8100,N_8485);
nand U9399 (N_9399,N_8387,N_8588);
and U9400 (N_9400,N_8838,N_8803);
or U9401 (N_9401,N_8138,N_8859);
or U9402 (N_9402,N_8565,N_8800);
and U9403 (N_9403,N_8966,N_8663);
nor U9404 (N_9404,N_8205,N_8134);
xor U9405 (N_9405,N_8470,N_8307);
or U9406 (N_9406,N_8340,N_8008);
nor U9407 (N_9407,N_8709,N_8010);
nand U9408 (N_9408,N_8156,N_8521);
nor U9409 (N_9409,N_8464,N_8801);
and U9410 (N_9410,N_8899,N_8421);
nand U9411 (N_9411,N_8384,N_8980);
xnor U9412 (N_9412,N_8235,N_8014);
nor U9413 (N_9413,N_8870,N_8573);
nor U9414 (N_9414,N_8863,N_8985);
nor U9415 (N_9415,N_8620,N_8032);
nand U9416 (N_9416,N_8171,N_8984);
or U9417 (N_9417,N_8732,N_8606);
nor U9418 (N_9418,N_8113,N_8207);
or U9419 (N_9419,N_8337,N_8196);
nor U9420 (N_9420,N_8794,N_8853);
xor U9421 (N_9421,N_8627,N_8027);
nand U9422 (N_9422,N_8303,N_8264);
nor U9423 (N_9423,N_8808,N_8189);
or U9424 (N_9424,N_8009,N_8976);
nand U9425 (N_9425,N_8316,N_8258);
and U9426 (N_9426,N_8379,N_8719);
or U9427 (N_9427,N_8147,N_8300);
nand U9428 (N_9428,N_8523,N_8947);
or U9429 (N_9429,N_8784,N_8024);
or U9430 (N_9430,N_8437,N_8828);
xor U9431 (N_9431,N_8937,N_8501);
or U9432 (N_9432,N_8886,N_8145);
and U9433 (N_9433,N_8224,N_8309);
nand U9434 (N_9434,N_8279,N_8827);
nand U9435 (N_9435,N_8394,N_8987);
nand U9436 (N_9436,N_8201,N_8418);
and U9437 (N_9437,N_8236,N_8817);
and U9438 (N_9438,N_8275,N_8995);
and U9439 (N_9439,N_8774,N_8314);
nor U9440 (N_9440,N_8157,N_8193);
nand U9441 (N_9441,N_8815,N_8063);
and U9442 (N_9442,N_8127,N_8988);
and U9443 (N_9443,N_8674,N_8994);
or U9444 (N_9444,N_8105,N_8383);
nor U9445 (N_9445,N_8572,N_8971);
or U9446 (N_9446,N_8377,N_8839);
or U9447 (N_9447,N_8661,N_8659);
or U9448 (N_9448,N_8367,N_8324);
nand U9449 (N_9449,N_8085,N_8370);
nand U9450 (N_9450,N_8487,N_8203);
nand U9451 (N_9451,N_8628,N_8284);
nand U9452 (N_9452,N_8425,N_8978);
and U9453 (N_9453,N_8046,N_8150);
and U9454 (N_9454,N_8103,N_8820);
xor U9455 (N_9455,N_8568,N_8541);
nand U9456 (N_9456,N_8981,N_8095);
and U9457 (N_9457,N_8741,N_8391);
or U9458 (N_9458,N_8166,N_8297);
nor U9459 (N_9459,N_8187,N_8012);
nor U9460 (N_9460,N_8488,N_8791);
nand U9461 (N_9461,N_8420,N_8093);
nor U9462 (N_9462,N_8172,N_8006);
xnor U9463 (N_9463,N_8802,N_8198);
nand U9464 (N_9464,N_8396,N_8990);
nor U9465 (N_9465,N_8081,N_8742);
nor U9466 (N_9466,N_8473,N_8296);
nand U9467 (N_9467,N_8068,N_8695);
nor U9468 (N_9468,N_8152,N_8359);
xnor U9469 (N_9469,N_8502,N_8897);
nor U9470 (N_9470,N_8343,N_8037);
nor U9471 (N_9471,N_8875,N_8346);
and U9472 (N_9472,N_8733,N_8639);
nand U9473 (N_9473,N_8119,N_8702);
and U9474 (N_9474,N_8232,N_8728);
and U9475 (N_9475,N_8273,N_8252);
and U9476 (N_9476,N_8868,N_8191);
and U9477 (N_9477,N_8058,N_8654);
nand U9478 (N_9478,N_8600,N_8035);
nor U9479 (N_9479,N_8539,N_8069);
or U9480 (N_9480,N_8840,N_8930);
or U9481 (N_9481,N_8884,N_8513);
nand U9482 (N_9482,N_8789,N_8613);
nand U9483 (N_9483,N_8491,N_8381);
and U9484 (N_9484,N_8730,N_8290);
and U9485 (N_9485,N_8369,N_8607);
nand U9486 (N_9486,N_8320,N_8918);
or U9487 (N_9487,N_8675,N_8569);
or U9488 (N_9488,N_8665,N_8924);
xor U9489 (N_9489,N_8711,N_8621);
nor U9490 (N_9490,N_8459,N_8448);
nor U9491 (N_9491,N_8489,N_8557);
and U9492 (N_9492,N_8643,N_8846);
xnor U9493 (N_9493,N_8902,N_8373);
or U9494 (N_9494,N_8941,N_8405);
and U9495 (N_9495,N_8400,N_8629);
nor U9496 (N_9496,N_8862,N_8883);
and U9497 (N_9497,N_8716,N_8835);
xnor U9498 (N_9498,N_8894,N_8948);
nor U9499 (N_9499,N_8959,N_8060);
and U9500 (N_9500,N_8291,N_8579);
and U9501 (N_9501,N_8815,N_8806);
nand U9502 (N_9502,N_8480,N_8668);
nor U9503 (N_9503,N_8743,N_8627);
nand U9504 (N_9504,N_8617,N_8055);
and U9505 (N_9505,N_8802,N_8947);
nand U9506 (N_9506,N_8995,N_8498);
and U9507 (N_9507,N_8020,N_8317);
and U9508 (N_9508,N_8081,N_8544);
nand U9509 (N_9509,N_8082,N_8446);
nand U9510 (N_9510,N_8528,N_8087);
and U9511 (N_9511,N_8787,N_8229);
and U9512 (N_9512,N_8833,N_8252);
and U9513 (N_9513,N_8770,N_8124);
nor U9514 (N_9514,N_8894,N_8008);
nor U9515 (N_9515,N_8398,N_8259);
nand U9516 (N_9516,N_8798,N_8202);
or U9517 (N_9517,N_8981,N_8043);
nor U9518 (N_9518,N_8079,N_8274);
nor U9519 (N_9519,N_8858,N_8900);
and U9520 (N_9520,N_8661,N_8451);
or U9521 (N_9521,N_8667,N_8800);
nand U9522 (N_9522,N_8665,N_8498);
and U9523 (N_9523,N_8565,N_8864);
nand U9524 (N_9524,N_8769,N_8824);
or U9525 (N_9525,N_8222,N_8663);
nand U9526 (N_9526,N_8508,N_8047);
nor U9527 (N_9527,N_8594,N_8582);
nand U9528 (N_9528,N_8038,N_8403);
nand U9529 (N_9529,N_8834,N_8584);
or U9530 (N_9530,N_8224,N_8344);
and U9531 (N_9531,N_8545,N_8010);
nand U9532 (N_9532,N_8691,N_8836);
or U9533 (N_9533,N_8199,N_8386);
nor U9534 (N_9534,N_8806,N_8683);
or U9535 (N_9535,N_8160,N_8787);
or U9536 (N_9536,N_8473,N_8913);
or U9537 (N_9537,N_8640,N_8334);
nand U9538 (N_9538,N_8370,N_8684);
nand U9539 (N_9539,N_8541,N_8590);
or U9540 (N_9540,N_8609,N_8981);
and U9541 (N_9541,N_8074,N_8513);
or U9542 (N_9542,N_8798,N_8158);
or U9543 (N_9543,N_8979,N_8838);
and U9544 (N_9544,N_8521,N_8753);
or U9545 (N_9545,N_8035,N_8465);
nor U9546 (N_9546,N_8047,N_8636);
or U9547 (N_9547,N_8890,N_8296);
nor U9548 (N_9548,N_8369,N_8011);
nor U9549 (N_9549,N_8498,N_8140);
nand U9550 (N_9550,N_8514,N_8208);
or U9551 (N_9551,N_8977,N_8741);
and U9552 (N_9552,N_8023,N_8773);
and U9553 (N_9553,N_8320,N_8622);
and U9554 (N_9554,N_8272,N_8074);
and U9555 (N_9555,N_8923,N_8792);
and U9556 (N_9556,N_8542,N_8228);
nand U9557 (N_9557,N_8790,N_8314);
or U9558 (N_9558,N_8644,N_8425);
xor U9559 (N_9559,N_8757,N_8268);
or U9560 (N_9560,N_8096,N_8404);
nor U9561 (N_9561,N_8672,N_8067);
and U9562 (N_9562,N_8778,N_8290);
or U9563 (N_9563,N_8517,N_8279);
and U9564 (N_9564,N_8334,N_8849);
nor U9565 (N_9565,N_8151,N_8519);
nand U9566 (N_9566,N_8926,N_8955);
and U9567 (N_9567,N_8609,N_8225);
and U9568 (N_9568,N_8236,N_8409);
nor U9569 (N_9569,N_8737,N_8467);
or U9570 (N_9570,N_8448,N_8553);
and U9571 (N_9571,N_8691,N_8133);
and U9572 (N_9572,N_8152,N_8051);
xnor U9573 (N_9573,N_8901,N_8360);
nor U9574 (N_9574,N_8219,N_8573);
and U9575 (N_9575,N_8107,N_8849);
nand U9576 (N_9576,N_8451,N_8942);
and U9577 (N_9577,N_8615,N_8311);
nor U9578 (N_9578,N_8648,N_8694);
and U9579 (N_9579,N_8353,N_8189);
or U9580 (N_9580,N_8876,N_8745);
nor U9581 (N_9581,N_8527,N_8774);
or U9582 (N_9582,N_8523,N_8189);
nand U9583 (N_9583,N_8867,N_8418);
nor U9584 (N_9584,N_8406,N_8366);
nor U9585 (N_9585,N_8465,N_8868);
nand U9586 (N_9586,N_8620,N_8835);
nor U9587 (N_9587,N_8007,N_8282);
nor U9588 (N_9588,N_8478,N_8710);
nand U9589 (N_9589,N_8901,N_8918);
or U9590 (N_9590,N_8286,N_8589);
and U9591 (N_9591,N_8440,N_8846);
or U9592 (N_9592,N_8273,N_8297);
nor U9593 (N_9593,N_8561,N_8498);
and U9594 (N_9594,N_8788,N_8426);
nor U9595 (N_9595,N_8749,N_8522);
or U9596 (N_9596,N_8331,N_8406);
nand U9597 (N_9597,N_8750,N_8061);
and U9598 (N_9598,N_8116,N_8083);
and U9599 (N_9599,N_8369,N_8040);
or U9600 (N_9600,N_8037,N_8953);
and U9601 (N_9601,N_8785,N_8188);
or U9602 (N_9602,N_8658,N_8438);
or U9603 (N_9603,N_8603,N_8845);
and U9604 (N_9604,N_8353,N_8367);
and U9605 (N_9605,N_8459,N_8309);
nor U9606 (N_9606,N_8089,N_8705);
nor U9607 (N_9607,N_8033,N_8576);
and U9608 (N_9608,N_8657,N_8329);
nor U9609 (N_9609,N_8339,N_8156);
and U9610 (N_9610,N_8642,N_8533);
or U9611 (N_9611,N_8622,N_8409);
nand U9612 (N_9612,N_8819,N_8646);
or U9613 (N_9613,N_8661,N_8613);
nand U9614 (N_9614,N_8595,N_8176);
or U9615 (N_9615,N_8322,N_8231);
xnor U9616 (N_9616,N_8740,N_8015);
nand U9617 (N_9617,N_8893,N_8840);
xor U9618 (N_9618,N_8250,N_8739);
or U9619 (N_9619,N_8843,N_8951);
nand U9620 (N_9620,N_8524,N_8423);
and U9621 (N_9621,N_8424,N_8941);
and U9622 (N_9622,N_8376,N_8638);
nor U9623 (N_9623,N_8335,N_8220);
and U9624 (N_9624,N_8369,N_8597);
and U9625 (N_9625,N_8279,N_8844);
nor U9626 (N_9626,N_8958,N_8842);
xnor U9627 (N_9627,N_8638,N_8177);
and U9628 (N_9628,N_8446,N_8144);
nand U9629 (N_9629,N_8302,N_8314);
and U9630 (N_9630,N_8314,N_8673);
nand U9631 (N_9631,N_8918,N_8235);
or U9632 (N_9632,N_8716,N_8762);
or U9633 (N_9633,N_8961,N_8994);
and U9634 (N_9634,N_8284,N_8634);
xor U9635 (N_9635,N_8720,N_8047);
nand U9636 (N_9636,N_8245,N_8983);
nand U9637 (N_9637,N_8650,N_8811);
nor U9638 (N_9638,N_8783,N_8034);
or U9639 (N_9639,N_8679,N_8953);
or U9640 (N_9640,N_8949,N_8960);
or U9641 (N_9641,N_8571,N_8503);
or U9642 (N_9642,N_8158,N_8604);
nand U9643 (N_9643,N_8120,N_8028);
and U9644 (N_9644,N_8694,N_8510);
and U9645 (N_9645,N_8387,N_8958);
nor U9646 (N_9646,N_8098,N_8559);
nor U9647 (N_9647,N_8461,N_8795);
or U9648 (N_9648,N_8813,N_8939);
nand U9649 (N_9649,N_8725,N_8637);
and U9650 (N_9650,N_8323,N_8154);
nor U9651 (N_9651,N_8359,N_8983);
or U9652 (N_9652,N_8890,N_8506);
and U9653 (N_9653,N_8917,N_8932);
nand U9654 (N_9654,N_8729,N_8196);
and U9655 (N_9655,N_8353,N_8964);
nand U9656 (N_9656,N_8228,N_8756);
and U9657 (N_9657,N_8663,N_8943);
nor U9658 (N_9658,N_8872,N_8787);
or U9659 (N_9659,N_8432,N_8747);
nor U9660 (N_9660,N_8872,N_8351);
nor U9661 (N_9661,N_8925,N_8893);
nor U9662 (N_9662,N_8871,N_8440);
nor U9663 (N_9663,N_8022,N_8837);
nor U9664 (N_9664,N_8041,N_8388);
and U9665 (N_9665,N_8388,N_8333);
nand U9666 (N_9666,N_8653,N_8214);
and U9667 (N_9667,N_8711,N_8351);
nand U9668 (N_9668,N_8725,N_8532);
nor U9669 (N_9669,N_8286,N_8901);
and U9670 (N_9670,N_8766,N_8520);
or U9671 (N_9671,N_8111,N_8507);
nor U9672 (N_9672,N_8437,N_8443);
or U9673 (N_9673,N_8277,N_8242);
or U9674 (N_9674,N_8301,N_8445);
nor U9675 (N_9675,N_8011,N_8052);
or U9676 (N_9676,N_8531,N_8340);
and U9677 (N_9677,N_8736,N_8370);
nand U9678 (N_9678,N_8611,N_8927);
nor U9679 (N_9679,N_8289,N_8560);
nor U9680 (N_9680,N_8374,N_8604);
or U9681 (N_9681,N_8877,N_8891);
and U9682 (N_9682,N_8217,N_8136);
nand U9683 (N_9683,N_8465,N_8574);
nor U9684 (N_9684,N_8542,N_8001);
nand U9685 (N_9685,N_8434,N_8222);
or U9686 (N_9686,N_8571,N_8152);
or U9687 (N_9687,N_8869,N_8099);
or U9688 (N_9688,N_8457,N_8559);
nand U9689 (N_9689,N_8243,N_8417);
and U9690 (N_9690,N_8230,N_8667);
xnor U9691 (N_9691,N_8259,N_8308);
and U9692 (N_9692,N_8907,N_8148);
nand U9693 (N_9693,N_8748,N_8773);
and U9694 (N_9694,N_8445,N_8899);
nand U9695 (N_9695,N_8562,N_8342);
or U9696 (N_9696,N_8715,N_8151);
or U9697 (N_9697,N_8378,N_8199);
nor U9698 (N_9698,N_8940,N_8393);
or U9699 (N_9699,N_8333,N_8054);
nand U9700 (N_9700,N_8702,N_8600);
nand U9701 (N_9701,N_8394,N_8515);
nor U9702 (N_9702,N_8640,N_8069);
and U9703 (N_9703,N_8143,N_8169);
and U9704 (N_9704,N_8039,N_8383);
nand U9705 (N_9705,N_8948,N_8072);
nand U9706 (N_9706,N_8951,N_8928);
and U9707 (N_9707,N_8003,N_8437);
and U9708 (N_9708,N_8617,N_8908);
nand U9709 (N_9709,N_8886,N_8335);
nor U9710 (N_9710,N_8198,N_8156);
nor U9711 (N_9711,N_8321,N_8774);
nor U9712 (N_9712,N_8379,N_8095);
or U9713 (N_9713,N_8263,N_8697);
or U9714 (N_9714,N_8327,N_8197);
nor U9715 (N_9715,N_8610,N_8463);
and U9716 (N_9716,N_8165,N_8721);
xnor U9717 (N_9717,N_8875,N_8331);
nand U9718 (N_9718,N_8987,N_8744);
nand U9719 (N_9719,N_8181,N_8738);
and U9720 (N_9720,N_8326,N_8060);
nor U9721 (N_9721,N_8796,N_8611);
and U9722 (N_9722,N_8417,N_8543);
nand U9723 (N_9723,N_8030,N_8429);
or U9724 (N_9724,N_8791,N_8704);
nor U9725 (N_9725,N_8307,N_8939);
nor U9726 (N_9726,N_8599,N_8589);
and U9727 (N_9727,N_8466,N_8852);
nor U9728 (N_9728,N_8057,N_8962);
or U9729 (N_9729,N_8399,N_8762);
nand U9730 (N_9730,N_8000,N_8047);
or U9731 (N_9731,N_8037,N_8542);
nor U9732 (N_9732,N_8659,N_8051);
and U9733 (N_9733,N_8690,N_8653);
nor U9734 (N_9734,N_8739,N_8001);
and U9735 (N_9735,N_8494,N_8568);
nor U9736 (N_9736,N_8931,N_8700);
nor U9737 (N_9737,N_8355,N_8360);
nand U9738 (N_9738,N_8224,N_8883);
and U9739 (N_9739,N_8390,N_8259);
and U9740 (N_9740,N_8352,N_8880);
nand U9741 (N_9741,N_8371,N_8972);
nand U9742 (N_9742,N_8452,N_8234);
nand U9743 (N_9743,N_8482,N_8463);
nand U9744 (N_9744,N_8175,N_8766);
or U9745 (N_9745,N_8911,N_8302);
nor U9746 (N_9746,N_8501,N_8148);
nand U9747 (N_9747,N_8678,N_8171);
and U9748 (N_9748,N_8765,N_8518);
or U9749 (N_9749,N_8418,N_8000);
nand U9750 (N_9750,N_8137,N_8818);
nor U9751 (N_9751,N_8775,N_8409);
nand U9752 (N_9752,N_8112,N_8496);
nor U9753 (N_9753,N_8000,N_8296);
nand U9754 (N_9754,N_8346,N_8195);
nor U9755 (N_9755,N_8432,N_8609);
nand U9756 (N_9756,N_8195,N_8470);
nor U9757 (N_9757,N_8332,N_8013);
nand U9758 (N_9758,N_8186,N_8601);
or U9759 (N_9759,N_8542,N_8316);
and U9760 (N_9760,N_8439,N_8068);
xnor U9761 (N_9761,N_8603,N_8927);
nor U9762 (N_9762,N_8035,N_8264);
and U9763 (N_9763,N_8082,N_8802);
and U9764 (N_9764,N_8182,N_8963);
nor U9765 (N_9765,N_8464,N_8897);
nand U9766 (N_9766,N_8649,N_8808);
or U9767 (N_9767,N_8102,N_8212);
or U9768 (N_9768,N_8555,N_8340);
and U9769 (N_9769,N_8497,N_8449);
and U9770 (N_9770,N_8377,N_8633);
nor U9771 (N_9771,N_8103,N_8994);
and U9772 (N_9772,N_8034,N_8272);
nor U9773 (N_9773,N_8542,N_8043);
nand U9774 (N_9774,N_8320,N_8047);
and U9775 (N_9775,N_8973,N_8600);
nor U9776 (N_9776,N_8591,N_8105);
and U9777 (N_9777,N_8812,N_8358);
and U9778 (N_9778,N_8680,N_8988);
xnor U9779 (N_9779,N_8206,N_8748);
and U9780 (N_9780,N_8640,N_8015);
nand U9781 (N_9781,N_8932,N_8711);
and U9782 (N_9782,N_8182,N_8386);
and U9783 (N_9783,N_8185,N_8287);
or U9784 (N_9784,N_8390,N_8963);
or U9785 (N_9785,N_8885,N_8472);
or U9786 (N_9786,N_8806,N_8758);
nor U9787 (N_9787,N_8894,N_8676);
nor U9788 (N_9788,N_8331,N_8395);
nand U9789 (N_9789,N_8912,N_8091);
nor U9790 (N_9790,N_8731,N_8966);
nor U9791 (N_9791,N_8826,N_8407);
nand U9792 (N_9792,N_8985,N_8718);
nand U9793 (N_9793,N_8611,N_8515);
nor U9794 (N_9794,N_8115,N_8162);
nand U9795 (N_9795,N_8778,N_8810);
and U9796 (N_9796,N_8643,N_8160);
or U9797 (N_9797,N_8423,N_8744);
and U9798 (N_9798,N_8183,N_8714);
and U9799 (N_9799,N_8016,N_8561);
and U9800 (N_9800,N_8573,N_8811);
and U9801 (N_9801,N_8614,N_8459);
and U9802 (N_9802,N_8283,N_8928);
nor U9803 (N_9803,N_8650,N_8984);
or U9804 (N_9804,N_8739,N_8431);
or U9805 (N_9805,N_8019,N_8606);
nor U9806 (N_9806,N_8529,N_8630);
and U9807 (N_9807,N_8464,N_8898);
or U9808 (N_9808,N_8481,N_8435);
or U9809 (N_9809,N_8203,N_8891);
nand U9810 (N_9810,N_8170,N_8350);
or U9811 (N_9811,N_8792,N_8342);
nor U9812 (N_9812,N_8269,N_8989);
nand U9813 (N_9813,N_8040,N_8466);
nand U9814 (N_9814,N_8885,N_8687);
or U9815 (N_9815,N_8023,N_8723);
and U9816 (N_9816,N_8842,N_8089);
nor U9817 (N_9817,N_8518,N_8541);
nor U9818 (N_9818,N_8345,N_8896);
nand U9819 (N_9819,N_8881,N_8040);
and U9820 (N_9820,N_8094,N_8948);
or U9821 (N_9821,N_8520,N_8137);
nor U9822 (N_9822,N_8578,N_8175);
nand U9823 (N_9823,N_8975,N_8543);
nand U9824 (N_9824,N_8849,N_8025);
or U9825 (N_9825,N_8722,N_8892);
or U9826 (N_9826,N_8642,N_8662);
nor U9827 (N_9827,N_8604,N_8579);
xnor U9828 (N_9828,N_8104,N_8116);
and U9829 (N_9829,N_8959,N_8132);
or U9830 (N_9830,N_8474,N_8914);
nor U9831 (N_9831,N_8063,N_8176);
nand U9832 (N_9832,N_8329,N_8003);
or U9833 (N_9833,N_8911,N_8813);
nor U9834 (N_9834,N_8476,N_8521);
nand U9835 (N_9835,N_8814,N_8069);
or U9836 (N_9836,N_8430,N_8182);
and U9837 (N_9837,N_8328,N_8842);
nand U9838 (N_9838,N_8420,N_8442);
and U9839 (N_9839,N_8928,N_8072);
and U9840 (N_9840,N_8927,N_8856);
or U9841 (N_9841,N_8911,N_8701);
or U9842 (N_9842,N_8123,N_8097);
nand U9843 (N_9843,N_8597,N_8868);
or U9844 (N_9844,N_8296,N_8336);
and U9845 (N_9845,N_8238,N_8993);
nor U9846 (N_9846,N_8392,N_8936);
and U9847 (N_9847,N_8772,N_8715);
and U9848 (N_9848,N_8676,N_8969);
nand U9849 (N_9849,N_8713,N_8039);
and U9850 (N_9850,N_8910,N_8972);
nand U9851 (N_9851,N_8982,N_8320);
and U9852 (N_9852,N_8614,N_8216);
and U9853 (N_9853,N_8401,N_8235);
and U9854 (N_9854,N_8108,N_8513);
nor U9855 (N_9855,N_8084,N_8039);
and U9856 (N_9856,N_8832,N_8325);
nand U9857 (N_9857,N_8364,N_8395);
nand U9858 (N_9858,N_8016,N_8827);
nor U9859 (N_9859,N_8836,N_8392);
nand U9860 (N_9860,N_8970,N_8227);
or U9861 (N_9861,N_8279,N_8696);
nand U9862 (N_9862,N_8956,N_8379);
or U9863 (N_9863,N_8982,N_8141);
and U9864 (N_9864,N_8529,N_8203);
xnor U9865 (N_9865,N_8113,N_8630);
nand U9866 (N_9866,N_8392,N_8395);
or U9867 (N_9867,N_8961,N_8785);
nand U9868 (N_9868,N_8903,N_8785);
or U9869 (N_9869,N_8476,N_8609);
nand U9870 (N_9870,N_8410,N_8642);
nor U9871 (N_9871,N_8511,N_8524);
and U9872 (N_9872,N_8735,N_8656);
nand U9873 (N_9873,N_8926,N_8020);
xnor U9874 (N_9874,N_8771,N_8235);
nand U9875 (N_9875,N_8516,N_8403);
or U9876 (N_9876,N_8734,N_8332);
nand U9877 (N_9877,N_8905,N_8766);
and U9878 (N_9878,N_8659,N_8187);
nor U9879 (N_9879,N_8303,N_8062);
or U9880 (N_9880,N_8781,N_8948);
nand U9881 (N_9881,N_8595,N_8361);
and U9882 (N_9882,N_8228,N_8129);
nand U9883 (N_9883,N_8125,N_8438);
nand U9884 (N_9884,N_8667,N_8647);
nand U9885 (N_9885,N_8082,N_8069);
or U9886 (N_9886,N_8626,N_8968);
and U9887 (N_9887,N_8188,N_8993);
or U9888 (N_9888,N_8646,N_8375);
nand U9889 (N_9889,N_8922,N_8262);
and U9890 (N_9890,N_8192,N_8603);
and U9891 (N_9891,N_8450,N_8204);
or U9892 (N_9892,N_8634,N_8336);
and U9893 (N_9893,N_8750,N_8777);
nand U9894 (N_9894,N_8919,N_8927);
nor U9895 (N_9895,N_8577,N_8486);
or U9896 (N_9896,N_8627,N_8491);
nand U9897 (N_9897,N_8437,N_8316);
nor U9898 (N_9898,N_8341,N_8348);
nor U9899 (N_9899,N_8606,N_8735);
nor U9900 (N_9900,N_8909,N_8222);
nor U9901 (N_9901,N_8642,N_8405);
nor U9902 (N_9902,N_8312,N_8039);
and U9903 (N_9903,N_8960,N_8852);
nand U9904 (N_9904,N_8863,N_8857);
or U9905 (N_9905,N_8541,N_8037);
nor U9906 (N_9906,N_8692,N_8148);
or U9907 (N_9907,N_8702,N_8130);
and U9908 (N_9908,N_8883,N_8200);
nor U9909 (N_9909,N_8922,N_8801);
nor U9910 (N_9910,N_8703,N_8771);
or U9911 (N_9911,N_8257,N_8106);
and U9912 (N_9912,N_8267,N_8092);
or U9913 (N_9913,N_8705,N_8971);
and U9914 (N_9914,N_8401,N_8821);
and U9915 (N_9915,N_8990,N_8416);
nor U9916 (N_9916,N_8145,N_8823);
and U9917 (N_9917,N_8149,N_8187);
nor U9918 (N_9918,N_8067,N_8949);
nand U9919 (N_9919,N_8952,N_8385);
or U9920 (N_9920,N_8331,N_8440);
nand U9921 (N_9921,N_8625,N_8505);
and U9922 (N_9922,N_8946,N_8472);
or U9923 (N_9923,N_8703,N_8212);
nor U9924 (N_9924,N_8392,N_8737);
or U9925 (N_9925,N_8694,N_8475);
or U9926 (N_9926,N_8884,N_8629);
nand U9927 (N_9927,N_8968,N_8694);
and U9928 (N_9928,N_8736,N_8442);
or U9929 (N_9929,N_8802,N_8157);
or U9930 (N_9930,N_8694,N_8606);
and U9931 (N_9931,N_8970,N_8548);
nor U9932 (N_9932,N_8447,N_8889);
or U9933 (N_9933,N_8140,N_8612);
and U9934 (N_9934,N_8905,N_8367);
nor U9935 (N_9935,N_8896,N_8501);
and U9936 (N_9936,N_8567,N_8776);
nor U9937 (N_9937,N_8084,N_8986);
nor U9938 (N_9938,N_8394,N_8661);
nor U9939 (N_9939,N_8575,N_8174);
and U9940 (N_9940,N_8571,N_8179);
nor U9941 (N_9941,N_8293,N_8280);
and U9942 (N_9942,N_8992,N_8195);
and U9943 (N_9943,N_8276,N_8168);
nor U9944 (N_9944,N_8105,N_8777);
and U9945 (N_9945,N_8814,N_8679);
nor U9946 (N_9946,N_8457,N_8176);
nand U9947 (N_9947,N_8996,N_8272);
nor U9948 (N_9948,N_8897,N_8496);
or U9949 (N_9949,N_8180,N_8871);
or U9950 (N_9950,N_8838,N_8766);
xor U9951 (N_9951,N_8334,N_8936);
and U9952 (N_9952,N_8547,N_8629);
nand U9953 (N_9953,N_8553,N_8385);
nor U9954 (N_9954,N_8805,N_8106);
and U9955 (N_9955,N_8793,N_8635);
nor U9956 (N_9956,N_8507,N_8192);
or U9957 (N_9957,N_8000,N_8925);
and U9958 (N_9958,N_8628,N_8880);
or U9959 (N_9959,N_8148,N_8015);
nand U9960 (N_9960,N_8081,N_8513);
nor U9961 (N_9961,N_8675,N_8207);
nand U9962 (N_9962,N_8663,N_8625);
nor U9963 (N_9963,N_8011,N_8615);
nor U9964 (N_9964,N_8799,N_8056);
nand U9965 (N_9965,N_8308,N_8258);
xnor U9966 (N_9966,N_8715,N_8240);
and U9967 (N_9967,N_8836,N_8927);
and U9968 (N_9968,N_8541,N_8322);
nor U9969 (N_9969,N_8361,N_8730);
nor U9970 (N_9970,N_8097,N_8384);
nor U9971 (N_9971,N_8893,N_8167);
nor U9972 (N_9972,N_8018,N_8980);
or U9973 (N_9973,N_8386,N_8111);
and U9974 (N_9974,N_8848,N_8419);
nor U9975 (N_9975,N_8599,N_8814);
nor U9976 (N_9976,N_8089,N_8998);
or U9977 (N_9977,N_8200,N_8764);
nand U9978 (N_9978,N_8894,N_8419);
and U9979 (N_9979,N_8240,N_8902);
and U9980 (N_9980,N_8375,N_8822);
nor U9981 (N_9981,N_8378,N_8273);
nor U9982 (N_9982,N_8843,N_8373);
nand U9983 (N_9983,N_8385,N_8998);
or U9984 (N_9984,N_8706,N_8154);
or U9985 (N_9985,N_8493,N_8427);
and U9986 (N_9986,N_8659,N_8609);
nor U9987 (N_9987,N_8862,N_8293);
and U9988 (N_9988,N_8526,N_8572);
or U9989 (N_9989,N_8909,N_8065);
nor U9990 (N_9990,N_8766,N_8183);
or U9991 (N_9991,N_8946,N_8332);
nand U9992 (N_9992,N_8853,N_8741);
and U9993 (N_9993,N_8990,N_8314);
xnor U9994 (N_9994,N_8366,N_8974);
nor U9995 (N_9995,N_8570,N_8325);
nor U9996 (N_9996,N_8556,N_8234);
or U9997 (N_9997,N_8225,N_8583);
and U9998 (N_9998,N_8378,N_8928);
nand U9999 (N_9999,N_8772,N_8799);
nor UO_0 (O_0,N_9459,N_9950);
and UO_1 (O_1,N_9936,N_9618);
or UO_2 (O_2,N_9386,N_9642);
or UO_3 (O_3,N_9020,N_9374);
and UO_4 (O_4,N_9887,N_9126);
nand UO_5 (O_5,N_9771,N_9091);
and UO_6 (O_6,N_9600,N_9017);
nand UO_7 (O_7,N_9528,N_9154);
nor UO_8 (O_8,N_9322,N_9774);
and UO_9 (O_9,N_9667,N_9269);
nor UO_10 (O_10,N_9149,N_9305);
or UO_11 (O_11,N_9270,N_9793);
and UO_12 (O_12,N_9732,N_9252);
nor UO_13 (O_13,N_9883,N_9376);
xor UO_14 (O_14,N_9507,N_9005);
nor UO_15 (O_15,N_9219,N_9290);
or UO_16 (O_16,N_9922,N_9430);
nand UO_17 (O_17,N_9931,N_9658);
and UO_18 (O_18,N_9031,N_9483);
or UO_19 (O_19,N_9173,N_9916);
and UO_20 (O_20,N_9925,N_9946);
and UO_21 (O_21,N_9976,N_9361);
nand UO_22 (O_22,N_9933,N_9325);
or UO_23 (O_23,N_9162,N_9419);
nor UO_24 (O_24,N_9522,N_9644);
and UO_25 (O_25,N_9717,N_9984);
or UO_26 (O_26,N_9394,N_9327);
or UO_27 (O_27,N_9225,N_9033);
and UO_28 (O_28,N_9580,N_9101);
nor UO_29 (O_29,N_9311,N_9180);
or UO_30 (O_30,N_9128,N_9473);
or UO_31 (O_31,N_9564,N_9873);
xnor UO_32 (O_32,N_9897,N_9046);
and UO_33 (O_33,N_9122,N_9312);
or UO_34 (O_34,N_9437,N_9131);
nor UO_35 (O_35,N_9238,N_9193);
and UO_36 (O_36,N_9108,N_9863);
nor UO_37 (O_37,N_9156,N_9663);
nor UO_38 (O_38,N_9181,N_9471);
nand UO_39 (O_39,N_9533,N_9248);
and UO_40 (O_40,N_9848,N_9616);
nand UO_41 (O_41,N_9870,N_9034);
xnor UO_42 (O_42,N_9330,N_9467);
nor UO_43 (O_43,N_9956,N_9043);
and UO_44 (O_44,N_9527,N_9084);
nand UO_45 (O_45,N_9411,N_9740);
nor UO_46 (O_46,N_9350,N_9998);
or UO_47 (O_47,N_9275,N_9488);
or UO_48 (O_48,N_9762,N_9646);
nor UO_49 (O_49,N_9540,N_9098);
nor UO_50 (O_50,N_9008,N_9967);
and UO_51 (O_51,N_9611,N_9836);
and UO_52 (O_52,N_9251,N_9079);
or UO_53 (O_53,N_9787,N_9661);
nor UO_54 (O_54,N_9074,N_9678);
and UO_55 (O_55,N_9550,N_9712);
nand UO_56 (O_56,N_9906,N_9092);
nor UO_57 (O_57,N_9765,N_9701);
nor UO_58 (O_58,N_9695,N_9372);
nor UO_59 (O_59,N_9720,N_9370);
nor UO_60 (O_60,N_9085,N_9177);
xor UO_61 (O_61,N_9148,N_9860);
and UO_62 (O_62,N_9363,N_9460);
nand UO_63 (O_63,N_9965,N_9795);
and UO_64 (O_64,N_9399,N_9633);
and UO_65 (O_65,N_9391,N_9184);
or UO_66 (O_66,N_9827,N_9840);
and UO_67 (O_67,N_9683,N_9612);
or UO_68 (O_68,N_9063,N_9255);
and UO_69 (O_69,N_9869,N_9597);
or UO_70 (O_70,N_9617,N_9102);
nor UO_71 (O_71,N_9423,N_9502);
or UO_72 (O_72,N_9992,N_9858);
and UO_73 (O_73,N_9028,N_9051);
nand UO_74 (O_74,N_9366,N_9245);
and UO_75 (O_75,N_9358,N_9316);
and UO_76 (O_76,N_9995,N_9542);
or UO_77 (O_77,N_9813,N_9323);
and UO_78 (O_78,N_9968,N_9233);
nor UO_79 (O_79,N_9859,N_9824);
nand UO_80 (O_80,N_9891,N_9819);
nor UO_81 (O_81,N_9218,N_9767);
or UO_82 (O_82,N_9707,N_9665);
and UO_83 (O_83,N_9560,N_9733);
nor UO_84 (O_84,N_9364,N_9417);
or UO_85 (O_85,N_9893,N_9018);
nand UO_86 (O_86,N_9842,N_9067);
xor UO_87 (O_87,N_9614,N_9117);
and UO_88 (O_88,N_9647,N_9698);
nand UO_89 (O_89,N_9268,N_9106);
and UO_90 (O_90,N_9669,N_9047);
nand UO_91 (O_91,N_9547,N_9654);
nor UO_92 (O_92,N_9845,N_9139);
and UO_93 (O_93,N_9204,N_9685);
nor UO_94 (O_94,N_9941,N_9420);
nor UO_95 (O_95,N_9927,N_9073);
nand UO_96 (O_96,N_9656,N_9278);
nor UO_97 (O_97,N_9655,N_9048);
nor UO_98 (O_98,N_9449,N_9530);
nor UO_99 (O_99,N_9885,N_9263);
and UO_100 (O_100,N_9538,N_9187);
or UO_101 (O_101,N_9520,N_9111);
or UO_102 (O_102,N_9713,N_9484);
and UO_103 (O_103,N_9979,N_9407);
nand UO_104 (O_104,N_9554,N_9558);
nor UO_105 (O_105,N_9276,N_9416);
nand UO_106 (O_106,N_9075,N_9659);
nand UO_107 (O_107,N_9042,N_9744);
nand UO_108 (O_108,N_9910,N_9281);
nand UO_109 (O_109,N_9464,N_9463);
nor UO_110 (O_110,N_9164,N_9030);
or UO_111 (O_111,N_9206,N_9800);
and UO_112 (O_112,N_9405,N_9639);
nor UO_113 (O_113,N_9686,N_9362);
nand UO_114 (O_114,N_9337,N_9367);
and UO_115 (O_115,N_9964,N_9209);
or UO_116 (O_116,N_9132,N_9016);
and UO_117 (O_117,N_9805,N_9196);
nor UO_118 (O_118,N_9480,N_9472);
or UO_119 (O_119,N_9531,N_9329);
nand UO_120 (O_120,N_9980,N_9476);
nand UO_121 (O_121,N_9529,N_9006);
or UO_122 (O_122,N_9169,N_9871);
and UO_123 (O_123,N_9814,N_9427);
xor UO_124 (O_124,N_9388,N_9146);
nor UO_125 (O_125,N_9365,N_9071);
nor UO_126 (O_126,N_9380,N_9369);
nand UO_127 (O_127,N_9446,N_9722);
nand UO_128 (O_128,N_9192,N_9112);
nand UO_129 (O_129,N_9414,N_9468);
or UO_130 (O_130,N_9593,N_9888);
nand UO_131 (O_131,N_9761,N_9425);
nor UO_132 (O_132,N_9562,N_9009);
or UO_133 (O_133,N_9775,N_9896);
nand UO_134 (O_134,N_9963,N_9176);
or UO_135 (O_135,N_9359,N_9539);
or UO_136 (O_136,N_9368,N_9114);
or UO_137 (O_137,N_9589,N_9384);
and UO_138 (O_138,N_9037,N_9734);
and UO_139 (O_139,N_9044,N_9431);
nand UO_140 (O_140,N_9838,N_9825);
and UO_141 (O_141,N_9504,N_9691);
or UO_142 (O_142,N_9721,N_9296);
or UO_143 (O_143,N_9621,N_9945);
or UO_144 (O_144,N_9064,N_9222);
nand UO_145 (O_145,N_9557,N_9754);
nor UO_146 (O_146,N_9099,N_9194);
nand UO_147 (O_147,N_9680,N_9619);
nand UO_148 (O_148,N_9806,N_9174);
xor UO_149 (O_149,N_9961,N_9929);
or UO_150 (O_150,N_9917,N_9227);
nand UO_151 (O_151,N_9817,N_9517);
nor UO_152 (O_152,N_9599,N_9643);
xor UO_153 (O_153,N_9003,N_9371);
nor UO_154 (O_154,N_9408,N_9632);
or UO_155 (O_155,N_9785,N_9577);
xor UO_156 (O_156,N_9267,N_9383);
and UO_157 (O_157,N_9727,N_9636);
xor UO_158 (O_158,N_9110,N_9221);
or UO_159 (O_159,N_9465,N_9706);
nor UO_160 (O_160,N_9843,N_9356);
xnor UO_161 (O_161,N_9188,N_9994);
nand UO_162 (O_162,N_9648,N_9470);
nand UO_163 (O_163,N_9170,N_9784);
xor UO_164 (O_164,N_9566,N_9759);
and UO_165 (O_165,N_9168,N_9134);
nor UO_166 (O_166,N_9952,N_9025);
nand UO_167 (O_167,N_9588,N_9657);
nor UO_168 (O_168,N_9002,N_9315);
nor UO_169 (O_169,N_9535,N_9262);
xnor UO_170 (O_170,N_9828,N_9835);
nand UO_171 (O_171,N_9138,N_9115);
or UO_172 (O_172,N_9651,N_9810);
or UO_173 (O_173,N_9652,N_9508);
or UO_174 (O_174,N_9900,N_9830);
and UO_175 (O_175,N_9457,N_9882);
and UO_176 (O_176,N_9455,N_9271);
nor UO_177 (O_177,N_9292,N_9807);
nand UO_178 (O_178,N_9768,N_9821);
or UO_179 (O_179,N_9440,N_9435);
or UO_180 (O_180,N_9379,N_9782);
nand UO_181 (O_181,N_9923,N_9495);
nor UO_182 (O_182,N_9142,N_9250);
nor UO_183 (O_183,N_9623,N_9820);
and UO_184 (O_184,N_9985,N_9053);
nand UO_185 (O_185,N_9158,N_9272);
or UO_186 (O_186,N_9438,N_9434);
nand UO_187 (O_187,N_9879,N_9246);
nand UO_188 (O_188,N_9428,N_9072);
nor UO_189 (O_189,N_9892,N_9609);
and UO_190 (O_190,N_9736,N_9274);
and UO_191 (O_191,N_9210,N_9743);
and UO_192 (O_192,N_9220,N_9650);
nand UO_193 (O_193,N_9096,N_9569);
and UO_194 (O_194,N_9152,N_9344);
nor UO_195 (O_195,N_9780,N_9904);
nand UO_196 (O_196,N_9129,N_9783);
nor UO_197 (O_197,N_9726,N_9302);
nor UO_198 (O_198,N_9811,N_9822);
nor UO_199 (O_199,N_9153,N_9694);
or UO_200 (O_200,N_9190,N_9203);
xnor UO_201 (O_201,N_9918,N_9708);
nor UO_202 (O_202,N_9421,N_9543);
nand UO_203 (O_203,N_9868,N_9150);
nand UO_204 (O_204,N_9751,N_9563);
nor UO_205 (O_205,N_9123,N_9851);
and UO_206 (O_206,N_9884,N_9432);
nor UO_207 (O_207,N_9357,N_9983);
and UO_208 (O_208,N_9345,N_9804);
or UO_209 (O_209,N_9035,N_9287);
nand UO_210 (O_210,N_9534,N_9412);
xor UO_211 (O_211,N_9605,N_9212);
nand UO_212 (O_212,N_9392,N_9518);
nor UO_213 (O_213,N_9004,N_9926);
and UO_214 (O_214,N_9687,N_9553);
or UO_215 (O_215,N_9546,N_9914);
or UO_216 (O_216,N_9682,N_9500);
and UO_217 (O_217,N_9966,N_9021);
or UO_218 (O_218,N_9089,N_9144);
and UO_219 (O_219,N_9668,N_9147);
nor UO_220 (O_220,N_9385,N_9565);
nand UO_221 (O_221,N_9105,N_9015);
nor UO_222 (O_222,N_9846,N_9958);
or UO_223 (O_223,N_9829,N_9847);
nor UO_224 (O_224,N_9622,N_9342);
nand UO_225 (O_225,N_9674,N_9143);
or UO_226 (O_226,N_9602,N_9953);
and UO_227 (O_227,N_9895,N_9515);
and UO_228 (O_228,N_9038,N_9987);
nor UO_229 (O_229,N_9332,N_9578);
xor UO_230 (O_230,N_9857,N_9986);
nand UO_231 (O_231,N_9629,N_9872);
xnor UO_232 (O_232,N_9050,N_9797);
nor UO_233 (O_233,N_9401,N_9309);
and UO_234 (O_234,N_9182,N_9513);
nor UO_235 (O_235,N_9247,N_9664);
nor UO_236 (O_236,N_9962,N_9317);
and UO_237 (O_237,N_9069,N_9486);
or UO_238 (O_238,N_9055,N_9902);
and UO_239 (O_239,N_9894,N_9424);
xor UO_240 (O_240,N_9634,N_9549);
and UO_241 (O_241,N_9120,N_9448);
nand UO_242 (O_242,N_9974,N_9672);
nor UO_243 (O_243,N_9036,N_9833);
or UO_244 (O_244,N_9519,N_9935);
nor UO_245 (O_245,N_9525,N_9943);
or UO_246 (O_246,N_9684,N_9244);
nand UO_247 (O_247,N_9318,N_9217);
nor UO_248 (O_248,N_9786,N_9704);
nand UO_249 (O_249,N_9719,N_9351);
nor UO_250 (O_250,N_9875,N_9213);
nand UO_251 (O_251,N_9920,N_9844);
or UO_252 (O_252,N_9561,N_9826);
nor UO_253 (O_253,N_9716,N_9753);
nand UO_254 (O_254,N_9378,N_9024);
nand UO_255 (O_255,N_9348,N_9266);
and UO_256 (O_256,N_9178,N_9223);
and UO_257 (O_257,N_9478,N_9466);
or UO_258 (O_258,N_9516,N_9812);
or UO_259 (O_259,N_9670,N_9007);
and UO_260 (O_260,N_9862,N_9988);
and UO_261 (O_261,N_9957,N_9338);
or UO_262 (O_262,N_9772,N_9242);
nand UO_263 (O_263,N_9645,N_9777);
and UO_264 (O_264,N_9381,N_9521);
nor UO_265 (O_265,N_9208,N_9757);
and UO_266 (O_266,N_9125,N_9232);
nand UO_267 (O_267,N_9556,N_9610);
or UO_268 (O_268,N_9737,N_9113);
or UO_269 (O_269,N_9029,N_9104);
nand UO_270 (O_270,N_9505,N_9999);
nand UO_271 (O_271,N_9288,N_9179);
nand UO_272 (O_272,N_9404,N_9715);
and UO_273 (O_273,N_9852,N_9571);
or UO_274 (O_274,N_9837,N_9279);
or UO_275 (O_275,N_9482,N_9487);
nand UO_276 (O_276,N_9675,N_9326);
and UO_277 (O_277,N_9763,N_9990);
nand UO_278 (O_278,N_9671,N_9355);
and UO_279 (O_279,N_9027,N_9289);
nand UO_280 (O_280,N_9082,N_9397);
or UO_281 (O_281,N_9041,N_9982);
nand UO_282 (O_282,N_9738,N_9649);
or UO_283 (O_283,N_9121,N_9607);
or UO_284 (O_284,N_9183,N_9454);
or UO_285 (O_285,N_9801,N_9095);
or UO_286 (O_286,N_9831,N_9226);
or UO_287 (O_287,N_9140,N_9237);
nor UO_288 (O_288,N_9555,N_9745);
nor UO_289 (O_289,N_9347,N_9969);
and UO_290 (O_290,N_9676,N_9235);
and UO_291 (O_291,N_9375,N_9058);
nor UO_292 (O_292,N_9808,N_9773);
nor UO_293 (O_293,N_9256,N_9166);
and UO_294 (O_294,N_9724,N_9889);
or UO_295 (O_295,N_9088,N_9261);
and UO_296 (O_296,N_9254,N_9199);
or UO_297 (O_297,N_9052,N_9285);
and UO_298 (O_298,N_9078,N_9249);
nor UO_299 (O_299,N_9749,N_9107);
xnor UO_300 (O_300,N_9608,N_9059);
nand UO_301 (O_301,N_9443,N_9710);
nand UO_302 (O_302,N_9444,N_9997);
nor UO_303 (O_303,N_9548,N_9971);
or UO_304 (O_304,N_9241,N_9536);
nand UO_305 (O_305,N_9509,N_9258);
and UO_306 (O_306,N_9909,N_9978);
nor UO_307 (O_307,N_9624,N_9689);
nand UO_308 (O_308,N_9280,N_9756);
and UO_309 (O_309,N_9590,N_9195);
or UO_310 (O_310,N_9596,N_9881);
and UO_311 (O_311,N_9239,N_9541);
and UO_312 (O_312,N_9070,N_9864);
nor UO_313 (O_313,N_9626,N_9324);
nand UO_314 (O_314,N_9439,N_9551);
nor UO_315 (O_315,N_9228,N_9163);
and UO_316 (O_316,N_9932,N_9567);
xor UO_317 (O_317,N_9277,N_9349);
nor UO_318 (O_318,N_9231,N_9081);
or UO_319 (O_319,N_9912,N_9390);
nor UO_320 (O_320,N_9396,N_9118);
and UO_321 (O_321,N_9924,N_9955);
and UO_322 (O_322,N_9442,N_9511);
nor UO_323 (O_323,N_9901,N_9475);
nand UO_324 (O_324,N_9981,N_9867);
or UO_325 (O_325,N_9552,N_9944);
nand UO_326 (O_326,N_9493,N_9403);
nand UO_327 (O_327,N_9319,N_9062);
nand UO_328 (O_328,N_9886,N_9878);
or UO_329 (O_329,N_9815,N_9832);
nand UO_330 (O_330,N_9890,N_9506);
nand UO_331 (O_331,N_9406,N_9796);
or UO_332 (O_332,N_9481,N_9940);
and UO_333 (O_333,N_9703,N_9340);
and UO_334 (O_334,N_9243,N_9803);
nor UO_335 (O_335,N_9681,N_9426);
nand UO_336 (O_336,N_9395,N_9086);
nand UO_337 (O_337,N_9012,N_9161);
or UO_338 (O_338,N_9496,N_9591);
nand UO_339 (O_339,N_9572,N_9352);
or UO_340 (O_340,N_9960,N_9373);
and UO_341 (O_341,N_9907,N_9545);
nand UO_342 (O_342,N_9975,N_9592);
nand UO_343 (O_343,N_9723,N_9595);
nand UO_344 (O_344,N_9301,N_9492);
and UO_345 (O_345,N_9587,N_9739);
nand UO_346 (O_346,N_9451,N_9594);
or UO_347 (O_347,N_9336,N_9155);
and UO_348 (O_348,N_9013,N_9109);
and UO_349 (O_349,N_9189,N_9697);
and UO_350 (O_350,N_9119,N_9679);
nand UO_351 (O_351,N_9282,N_9422);
or UO_352 (O_352,N_9141,N_9660);
nand UO_353 (O_353,N_9045,N_9186);
nor UO_354 (O_354,N_9393,N_9781);
nand UO_355 (O_355,N_9303,N_9377);
nand UO_356 (O_356,N_9485,N_9450);
nand UO_357 (O_357,N_9418,N_9011);
or UO_358 (O_358,N_9083,N_9628);
and UO_359 (O_359,N_9000,N_9973);
and UO_360 (O_360,N_9937,N_9216);
nor UO_361 (O_361,N_9705,N_9876);
and UO_362 (O_362,N_9948,N_9469);
nand UO_363 (O_363,N_9690,N_9341);
or UO_364 (O_364,N_9097,N_9214);
and UO_365 (O_365,N_9291,N_9579);
or UO_366 (O_366,N_9339,N_9456);
or UO_367 (O_367,N_9167,N_9159);
nor UO_368 (O_368,N_9938,N_9293);
or UO_369 (O_369,N_9959,N_9856);
or UO_370 (O_370,N_9229,N_9850);
xor UO_371 (O_371,N_9135,N_9514);
or UO_372 (O_372,N_9748,N_9798);
and UO_373 (O_373,N_9939,N_9709);
and UO_374 (O_374,N_9991,N_9526);
nor UO_375 (O_375,N_9306,N_9581);
nor UO_376 (O_376,N_9728,N_9934);
or UO_377 (O_377,N_9877,N_9331);
nand UO_378 (O_378,N_9019,N_9510);
nand UO_379 (O_379,N_9133,N_9766);
nor UO_380 (O_380,N_9911,N_9265);
xor UO_381 (O_381,N_9491,N_9747);
and UO_382 (O_382,N_9433,N_9802);
nand UO_383 (O_383,N_9537,N_9197);
nor UO_384 (O_384,N_9136,N_9954);
or UO_385 (O_385,N_9583,N_9794);
or UO_386 (O_386,N_9532,N_9145);
or UO_387 (O_387,N_9570,N_9093);
or UO_388 (O_388,N_9171,N_9637);
or UO_389 (O_389,N_9295,N_9524);
or UO_390 (O_390,N_9718,N_9865);
nor UO_391 (O_391,N_9930,N_9198);
nor UO_392 (O_392,N_9032,N_9001);
or UO_393 (O_393,N_9211,N_9060);
nand UO_394 (O_394,N_9202,N_9778);
nand UO_395 (O_395,N_9297,N_9903);
xnor UO_396 (O_396,N_9809,N_9014);
or UO_397 (O_397,N_9866,N_9452);
nor UO_398 (O_398,N_9160,N_9641);
or UO_399 (O_399,N_9731,N_9638);
and UO_400 (O_400,N_9240,N_9627);
and UO_401 (O_401,N_9631,N_9494);
or UO_402 (O_402,N_9489,N_9725);
nand UO_403 (O_403,N_9234,N_9776);
nor UO_404 (O_404,N_9693,N_9273);
and UO_405 (O_405,N_9915,N_9760);
and UO_406 (O_406,N_9625,N_9559);
and UO_407 (O_407,N_9259,N_9769);
nor UO_408 (O_408,N_9409,N_9662);
nand UO_409 (O_409,N_9498,N_9458);
or UO_410 (O_410,N_9699,N_9635);
and UO_411 (O_411,N_9320,N_9499);
and UO_412 (O_412,N_9714,N_9741);
nor UO_413 (O_413,N_9284,N_9711);
nor UO_414 (O_414,N_9512,N_9474);
nand UO_415 (O_415,N_9415,N_9854);
nor UO_416 (O_416,N_9598,N_9575);
nand UO_417 (O_417,N_9061,N_9604);
or UO_418 (O_418,N_9606,N_9673);
or UO_419 (O_419,N_9770,N_9462);
nor UO_420 (O_420,N_9640,N_9157);
nand UO_421 (O_421,N_9908,N_9601);
or UO_422 (O_422,N_9792,N_9913);
or UO_423 (O_423,N_9834,N_9207);
and UO_424 (O_424,N_9039,N_9568);
or UO_425 (O_425,N_9260,N_9353);
nand UO_426 (O_426,N_9692,N_9103);
nand UO_427 (O_427,N_9972,N_9490);
or UO_428 (O_428,N_9116,N_9993);
nand UO_429 (O_429,N_9057,N_9253);
or UO_430 (O_430,N_9298,N_9666);
and UO_431 (O_431,N_9977,N_9735);
xor UO_432 (O_432,N_9137,N_9205);
nor UO_433 (O_433,N_9201,N_9389);
nand UO_434 (O_434,N_9755,N_9215);
nor UO_435 (O_435,N_9346,N_9729);
and UO_436 (O_436,N_9445,N_9789);
nand UO_437 (O_437,N_9224,N_9880);
nand UO_438 (O_438,N_9236,N_9354);
nand UO_439 (O_439,N_9750,N_9573);
and UO_440 (O_440,N_9700,N_9230);
and UO_441 (O_441,N_9584,N_9124);
or UO_442 (O_442,N_9436,N_9620);
or UO_443 (O_443,N_9335,N_9283);
nor UO_444 (O_444,N_9398,N_9586);
nand UO_445 (O_445,N_9130,N_9702);
xor UO_446 (O_446,N_9441,N_9321);
or UO_447 (O_447,N_9382,N_9996);
nor UO_448 (O_448,N_9688,N_9286);
nand UO_449 (O_449,N_9576,N_9010);
nand UO_450 (O_450,N_9410,N_9928);
and UO_451 (O_451,N_9447,N_9026);
or UO_452 (O_452,N_9853,N_9191);
nand UO_453 (O_453,N_9087,N_9077);
nor UO_454 (O_454,N_9304,N_9544);
and UO_455 (O_455,N_9100,N_9076);
nand UO_456 (O_456,N_9951,N_9165);
nand UO_457 (O_457,N_9501,N_9752);
or UO_458 (O_458,N_9185,N_9788);
and UO_459 (O_459,N_9172,N_9056);
or UO_460 (O_460,N_9861,N_9574);
or UO_461 (O_461,N_9989,N_9461);
and UO_462 (O_462,N_9307,N_9582);
nand UO_463 (O_463,N_9585,N_9308);
or UO_464 (O_464,N_9849,N_9068);
nand UO_465 (O_465,N_9899,N_9523);
or UO_466 (O_466,N_9779,N_9080);
and UO_467 (O_467,N_9730,N_9477);
nor UO_468 (O_468,N_9294,N_9799);
or UO_469 (O_469,N_9151,N_9898);
and UO_470 (O_470,N_9677,N_9855);
nand UO_471 (O_471,N_9066,N_9746);
or UO_472 (O_472,N_9841,N_9310);
nand UO_473 (O_473,N_9299,N_9630);
and UO_474 (O_474,N_9314,N_9343);
and UO_475 (O_475,N_9919,N_9065);
or UO_476 (O_476,N_9387,N_9758);
and UO_477 (O_477,N_9791,N_9874);
nand UO_478 (O_478,N_9360,N_9613);
or UO_479 (O_479,N_9334,N_9127);
nor UO_480 (O_480,N_9429,N_9742);
nor UO_481 (O_481,N_9175,N_9764);
and UO_482 (O_482,N_9400,N_9615);
nand UO_483 (O_483,N_9653,N_9328);
and UO_484 (O_484,N_9022,N_9023);
or UO_485 (O_485,N_9839,N_9603);
or UO_486 (O_486,N_9453,N_9942);
nor UO_487 (O_487,N_9313,N_9257);
nand UO_488 (O_488,N_9503,N_9049);
or UO_489 (O_489,N_9823,N_9333);
nand UO_490 (O_490,N_9696,N_9905);
and UO_491 (O_491,N_9300,N_9947);
nand UO_492 (O_492,N_9264,N_9921);
nand UO_493 (O_493,N_9040,N_9816);
nor UO_494 (O_494,N_9200,N_9970);
nor UO_495 (O_495,N_9818,N_9402);
or UO_496 (O_496,N_9479,N_9054);
and UO_497 (O_497,N_9090,N_9790);
or UO_498 (O_498,N_9094,N_9413);
nor UO_499 (O_499,N_9497,N_9949);
or UO_500 (O_500,N_9931,N_9282);
nand UO_501 (O_501,N_9216,N_9255);
and UO_502 (O_502,N_9778,N_9254);
and UO_503 (O_503,N_9807,N_9271);
or UO_504 (O_504,N_9276,N_9549);
and UO_505 (O_505,N_9587,N_9354);
and UO_506 (O_506,N_9809,N_9171);
nor UO_507 (O_507,N_9577,N_9534);
nor UO_508 (O_508,N_9382,N_9834);
nor UO_509 (O_509,N_9977,N_9298);
or UO_510 (O_510,N_9547,N_9932);
nor UO_511 (O_511,N_9142,N_9459);
nor UO_512 (O_512,N_9576,N_9067);
nor UO_513 (O_513,N_9083,N_9930);
or UO_514 (O_514,N_9561,N_9245);
and UO_515 (O_515,N_9926,N_9239);
or UO_516 (O_516,N_9056,N_9061);
nor UO_517 (O_517,N_9426,N_9801);
or UO_518 (O_518,N_9795,N_9582);
or UO_519 (O_519,N_9639,N_9237);
nand UO_520 (O_520,N_9297,N_9064);
nand UO_521 (O_521,N_9607,N_9337);
nand UO_522 (O_522,N_9411,N_9459);
nand UO_523 (O_523,N_9874,N_9854);
nand UO_524 (O_524,N_9776,N_9123);
and UO_525 (O_525,N_9198,N_9180);
and UO_526 (O_526,N_9106,N_9428);
nand UO_527 (O_527,N_9054,N_9961);
or UO_528 (O_528,N_9544,N_9705);
and UO_529 (O_529,N_9517,N_9904);
nor UO_530 (O_530,N_9773,N_9547);
nand UO_531 (O_531,N_9282,N_9512);
and UO_532 (O_532,N_9194,N_9872);
nand UO_533 (O_533,N_9419,N_9739);
or UO_534 (O_534,N_9955,N_9800);
or UO_535 (O_535,N_9678,N_9983);
or UO_536 (O_536,N_9486,N_9483);
or UO_537 (O_537,N_9323,N_9207);
nor UO_538 (O_538,N_9286,N_9256);
xnor UO_539 (O_539,N_9049,N_9527);
nor UO_540 (O_540,N_9329,N_9117);
or UO_541 (O_541,N_9173,N_9647);
and UO_542 (O_542,N_9339,N_9685);
nand UO_543 (O_543,N_9632,N_9528);
nor UO_544 (O_544,N_9221,N_9546);
and UO_545 (O_545,N_9406,N_9393);
nand UO_546 (O_546,N_9966,N_9493);
nand UO_547 (O_547,N_9876,N_9167);
nor UO_548 (O_548,N_9599,N_9594);
nor UO_549 (O_549,N_9833,N_9905);
and UO_550 (O_550,N_9007,N_9454);
or UO_551 (O_551,N_9512,N_9711);
nor UO_552 (O_552,N_9042,N_9010);
and UO_553 (O_553,N_9174,N_9658);
nor UO_554 (O_554,N_9435,N_9247);
nor UO_555 (O_555,N_9845,N_9175);
nand UO_556 (O_556,N_9759,N_9407);
nor UO_557 (O_557,N_9951,N_9508);
nand UO_558 (O_558,N_9500,N_9470);
nor UO_559 (O_559,N_9612,N_9138);
nor UO_560 (O_560,N_9843,N_9825);
nor UO_561 (O_561,N_9052,N_9384);
or UO_562 (O_562,N_9309,N_9196);
and UO_563 (O_563,N_9970,N_9793);
nor UO_564 (O_564,N_9806,N_9778);
or UO_565 (O_565,N_9856,N_9300);
or UO_566 (O_566,N_9043,N_9634);
nand UO_567 (O_567,N_9776,N_9283);
or UO_568 (O_568,N_9381,N_9250);
and UO_569 (O_569,N_9481,N_9175);
nand UO_570 (O_570,N_9705,N_9321);
and UO_571 (O_571,N_9784,N_9974);
nor UO_572 (O_572,N_9139,N_9140);
nand UO_573 (O_573,N_9430,N_9850);
and UO_574 (O_574,N_9902,N_9961);
nor UO_575 (O_575,N_9650,N_9439);
nor UO_576 (O_576,N_9326,N_9557);
xnor UO_577 (O_577,N_9429,N_9129);
nand UO_578 (O_578,N_9019,N_9405);
and UO_579 (O_579,N_9985,N_9408);
and UO_580 (O_580,N_9533,N_9602);
or UO_581 (O_581,N_9306,N_9544);
and UO_582 (O_582,N_9169,N_9134);
and UO_583 (O_583,N_9839,N_9936);
xor UO_584 (O_584,N_9748,N_9022);
or UO_585 (O_585,N_9012,N_9753);
nand UO_586 (O_586,N_9204,N_9386);
nand UO_587 (O_587,N_9519,N_9907);
and UO_588 (O_588,N_9839,N_9280);
nor UO_589 (O_589,N_9874,N_9645);
nor UO_590 (O_590,N_9413,N_9460);
nor UO_591 (O_591,N_9576,N_9967);
and UO_592 (O_592,N_9183,N_9745);
and UO_593 (O_593,N_9593,N_9084);
or UO_594 (O_594,N_9725,N_9686);
xor UO_595 (O_595,N_9827,N_9939);
and UO_596 (O_596,N_9002,N_9468);
or UO_597 (O_597,N_9041,N_9658);
nand UO_598 (O_598,N_9388,N_9901);
and UO_599 (O_599,N_9404,N_9542);
and UO_600 (O_600,N_9916,N_9029);
nor UO_601 (O_601,N_9385,N_9398);
nor UO_602 (O_602,N_9092,N_9530);
nor UO_603 (O_603,N_9855,N_9407);
nor UO_604 (O_604,N_9498,N_9197);
nand UO_605 (O_605,N_9919,N_9752);
or UO_606 (O_606,N_9687,N_9885);
nand UO_607 (O_607,N_9687,N_9951);
or UO_608 (O_608,N_9451,N_9896);
or UO_609 (O_609,N_9352,N_9740);
and UO_610 (O_610,N_9310,N_9200);
or UO_611 (O_611,N_9966,N_9289);
or UO_612 (O_612,N_9926,N_9574);
and UO_613 (O_613,N_9960,N_9239);
nand UO_614 (O_614,N_9130,N_9156);
nand UO_615 (O_615,N_9134,N_9146);
xnor UO_616 (O_616,N_9328,N_9555);
nand UO_617 (O_617,N_9897,N_9789);
and UO_618 (O_618,N_9121,N_9380);
or UO_619 (O_619,N_9555,N_9100);
or UO_620 (O_620,N_9508,N_9579);
or UO_621 (O_621,N_9747,N_9018);
nor UO_622 (O_622,N_9049,N_9221);
nand UO_623 (O_623,N_9533,N_9526);
nor UO_624 (O_624,N_9788,N_9316);
nor UO_625 (O_625,N_9779,N_9680);
nand UO_626 (O_626,N_9156,N_9483);
and UO_627 (O_627,N_9130,N_9664);
nor UO_628 (O_628,N_9669,N_9778);
nor UO_629 (O_629,N_9937,N_9285);
and UO_630 (O_630,N_9943,N_9938);
nor UO_631 (O_631,N_9411,N_9509);
xnor UO_632 (O_632,N_9717,N_9193);
nor UO_633 (O_633,N_9415,N_9625);
nor UO_634 (O_634,N_9429,N_9090);
or UO_635 (O_635,N_9470,N_9339);
nor UO_636 (O_636,N_9862,N_9867);
and UO_637 (O_637,N_9038,N_9246);
nand UO_638 (O_638,N_9678,N_9082);
nor UO_639 (O_639,N_9275,N_9314);
and UO_640 (O_640,N_9757,N_9332);
nor UO_641 (O_641,N_9254,N_9546);
nor UO_642 (O_642,N_9740,N_9867);
or UO_643 (O_643,N_9932,N_9727);
or UO_644 (O_644,N_9172,N_9287);
or UO_645 (O_645,N_9756,N_9786);
and UO_646 (O_646,N_9414,N_9912);
nand UO_647 (O_647,N_9293,N_9960);
nor UO_648 (O_648,N_9401,N_9036);
nand UO_649 (O_649,N_9416,N_9445);
nand UO_650 (O_650,N_9012,N_9074);
and UO_651 (O_651,N_9753,N_9751);
nand UO_652 (O_652,N_9778,N_9696);
nor UO_653 (O_653,N_9790,N_9396);
and UO_654 (O_654,N_9069,N_9234);
nor UO_655 (O_655,N_9257,N_9535);
or UO_656 (O_656,N_9226,N_9401);
nor UO_657 (O_657,N_9508,N_9979);
nor UO_658 (O_658,N_9386,N_9747);
xnor UO_659 (O_659,N_9740,N_9754);
and UO_660 (O_660,N_9450,N_9938);
and UO_661 (O_661,N_9662,N_9320);
nand UO_662 (O_662,N_9781,N_9695);
nand UO_663 (O_663,N_9815,N_9790);
or UO_664 (O_664,N_9114,N_9919);
nand UO_665 (O_665,N_9923,N_9978);
nor UO_666 (O_666,N_9627,N_9047);
nor UO_667 (O_667,N_9519,N_9674);
or UO_668 (O_668,N_9688,N_9516);
nand UO_669 (O_669,N_9361,N_9923);
and UO_670 (O_670,N_9759,N_9762);
nor UO_671 (O_671,N_9002,N_9499);
and UO_672 (O_672,N_9605,N_9373);
xor UO_673 (O_673,N_9628,N_9281);
or UO_674 (O_674,N_9812,N_9123);
nor UO_675 (O_675,N_9267,N_9107);
nand UO_676 (O_676,N_9272,N_9095);
nor UO_677 (O_677,N_9917,N_9668);
nand UO_678 (O_678,N_9237,N_9540);
nor UO_679 (O_679,N_9850,N_9902);
or UO_680 (O_680,N_9611,N_9726);
and UO_681 (O_681,N_9166,N_9384);
or UO_682 (O_682,N_9008,N_9006);
and UO_683 (O_683,N_9798,N_9003);
nor UO_684 (O_684,N_9364,N_9384);
xnor UO_685 (O_685,N_9768,N_9277);
or UO_686 (O_686,N_9212,N_9632);
or UO_687 (O_687,N_9119,N_9184);
nand UO_688 (O_688,N_9453,N_9114);
and UO_689 (O_689,N_9756,N_9684);
nand UO_690 (O_690,N_9171,N_9138);
nor UO_691 (O_691,N_9039,N_9801);
nor UO_692 (O_692,N_9915,N_9778);
nor UO_693 (O_693,N_9324,N_9392);
or UO_694 (O_694,N_9791,N_9461);
and UO_695 (O_695,N_9911,N_9205);
and UO_696 (O_696,N_9780,N_9417);
nor UO_697 (O_697,N_9113,N_9702);
nor UO_698 (O_698,N_9174,N_9035);
or UO_699 (O_699,N_9037,N_9059);
nor UO_700 (O_700,N_9758,N_9564);
or UO_701 (O_701,N_9731,N_9174);
nand UO_702 (O_702,N_9343,N_9937);
nand UO_703 (O_703,N_9694,N_9408);
or UO_704 (O_704,N_9010,N_9595);
nand UO_705 (O_705,N_9418,N_9188);
nor UO_706 (O_706,N_9980,N_9743);
nand UO_707 (O_707,N_9469,N_9378);
or UO_708 (O_708,N_9780,N_9460);
nand UO_709 (O_709,N_9866,N_9971);
and UO_710 (O_710,N_9033,N_9545);
nor UO_711 (O_711,N_9422,N_9678);
or UO_712 (O_712,N_9598,N_9513);
or UO_713 (O_713,N_9191,N_9576);
nor UO_714 (O_714,N_9512,N_9222);
or UO_715 (O_715,N_9384,N_9866);
or UO_716 (O_716,N_9875,N_9605);
nand UO_717 (O_717,N_9843,N_9764);
and UO_718 (O_718,N_9108,N_9303);
nor UO_719 (O_719,N_9698,N_9819);
or UO_720 (O_720,N_9449,N_9563);
nor UO_721 (O_721,N_9533,N_9039);
and UO_722 (O_722,N_9123,N_9646);
and UO_723 (O_723,N_9910,N_9177);
and UO_724 (O_724,N_9697,N_9902);
or UO_725 (O_725,N_9332,N_9823);
or UO_726 (O_726,N_9702,N_9619);
or UO_727 (O_727,N_9983,N_9044);
and UO_728 (O_728,N_9686,N_9640);
nor UO_729 (O_729,N_9301,N_9901);
and UO_730 (O_730,N_9396,N_9389);
nor UO_731 (O_731,N_9157,N_9595);
or UO_732 (O_732,N_9685,N_9358);
or UO_733 (O_733,N_9902,N_9848);
nand UO_734 (O_734,N_9417,N_9958);
nor UO_735 (O_735,N_9688,N_9076);
and UO_736 (O_736,N_9036,N_9704);
or UO_737 (O_737,N_9535,N_9114);
nand UO_738 (O_738,N_9720,N_9016);
nand UO_739 (O_739,N_9854,N_9556);
or UO_740 (O_740,N_9586,N_9261);
nand UO_741 (O_741,N_9840,N_9547);
nor UO_742 (O_742,N_9532,N_9616);
and UO_743 (O_743,N_9665,N_9634);
or UO_744 (O_744,N_9963,N_9522);
or UO_745 (O_745,N_9911,N_9157);
nand UO_746 (O_746,N_9340,N_9958);
nor UO_747 (O_747,N_9133,N_9155);
or UO_748 (O_748,N_9528,N_9944);
nand UO_749 (O_749,N_9365,N_9968);
and UO_750 (O_750,N_9957,N_9942);
nor UO_751 (O_751,N_9189,N_9163);
or UO_752 (O_752,N_9964,N_9349);
and UO_753 (O_753,N_9984,N_9328);
and UO_754 (O_754,N_9840,N_9780);
or UO_755 (O_755,N_9481,N_9466);
or UO_756 (O_756,N_9205,N_9616);
nand UO_757 (O_757,N_9519,N_9156);
and UO_758 (O_758,N_9977,N_9665);
or UO_759 (O_759,N_9320,N_9510);
and UO_760 (O_760,N_9837,N_9696);
and UO_761 (O_761,N_9534,N_9347);
nor UO_762 (O_762,N_9076,N_9123);
or UO_763 (O_763,N_9922,N_9057);
nand UO_764 (O_764,N_9079,N_9531);
and UO_765 (O_765,N_9690,N_9339);
nand UO_766 (O_766,N_9654,N_9011);
or UO_767 (O_767,N_9798,N_9366);
or UO_768 (O_768,N_9060,N_9671);
nor UO_769 (O_769,N_9735,N_9099);
or UO_770 (O_770,N_9301,N_9616);
nand UO_771 (O_771,N_9546,N_9921);
nor UO_772 (O_772,N_9381,N_9119);
or UO_773 (O_773,N_9356,N_9181);
nor UO_774 (O_774,N_9138,N_9001);
nor UO_775 (O_775,N_9091,N_9045);
nor UO_776 (O_776,N_9937,N_9978);
or UO_777 (O_777,N_9038,N_9767);
and UO_778 (O_778,N_9698,N_9524);
nand UO_779 (O_779,N_9691,N_9655);
or UO_780 (O_780,N_9008,N_9845);
or UO_781 (O_781,N_9264,N_9693);
nor UO_782 (O_782,N_9252,N_9983);
nor UO_783 (O_783,N_9057,N_9966);
nand UO_784 (O_784,N_9010,N_9979);
and UO_785 (O_785,N_9830,N_9454);
and UO_786 (O_786,N_9610,N_9829);
and UO_787 (O_787,N_9849,N_9343);
nand UO_788 (O_788,N_9604,N_9157);
or UO_789 (O_789,N_9670,N_9836);
or UO_790 (O_790,N_9424,N_9439);
or UO_791 (O_791,N_9088,N_9354);
nor UO_792 (O_792,N_9651,N_9174);
and UO_793 (O_793,N_9809,N_9112);
or UO_794 (O_794,N_9243,N_9712);
or UO_795 (O_795,N_9617,N_9944);
nand UO_796 (O_796,N_9805,N_9647);
nand UO_797 (O_797,N_9866,N_9683);
and UO_798 (O_798,N_9499,N_9536);
and UO_799 (O_799,N_9909,N_9390);
nor UO_800 (O_800,N_9073,N_9119);
or UO_801 (O_801,N_9557,N_9475);
or UO_802 (O_802,N_9287,N_9823);
or UO_803 (O_803,N_9816,N_9615);
and UO_804 (O_804,N_9553,N_9313);
nand UO_805 (O_805,N_9135,N_9991);
nand UO_806 (O_806,N_9169,N_9489);
nor UO_807 (O_807,N_9968,N_9540);
nand UO_808 (O_808,N_9341,N_9978);
or UO_809 (O_809,N_9399,N_9447);
nor UO_810 (O_810,N_9784,N_9158);
nor UO_811 (O_811,N_9684,N_9451);
or UO_812 (O_812,N_9931,N_9323);
nand UO_813 (O_813,N_9799,N_9830);
or UO_814 (O_814,N_9355,N_9463);
and UO_815 (O_815,N_9000,N_9026);
and UO_816 (O_816,N_9390,N_9224);
and UO_817 (O_817,N_9936,N_9536);
or UO_818 (O_818,N_9079,N_9021);
nor UO_819 (O_819,N_9197,N_9189);
nor UO_820 (O_820,N_9467,N_9676);
nand UO_821 (O_821,N_9845,N_9253);
nand UO_822 (O_822,N_9922,N_9159);
nor UO_823 (O_823,N_9701,N_9915);
or UO_824 (O_824,N_9216,N_9043);
nor UO_825 (O_825,N_9334,N_9455);
or UO_826 (O_826,N_9371,N_9241);
or UO_827 (O_827,N_9668,N_9838);
or UO_828 (O_828,N_9453,N_9250);
or UO_829 (O_829,N_9222,N_9836);
nand UO_830 (O_830,N_9959,N_9202);
nor UO_831 (O_831,N_9303,N_9390);
and UO_832 (O_832,N_9454,N_9474);
nor UO_833 (O_833,N_9585,N_9974);
and UO_834 (O_834,N_9855,N_9198);
nor UO_835 (O_835,N_9392,N_9600);
nand UO_836 (O_836,N_9373,N_9640);
nand UO_837 (O_837,N_9046,N_9686);
and UO_838 (O_838,N_9390,N_9127);
and UO_839 (O_839,N_9947,N_9304);
or UO_840 (O_840,N_9379,N_9108);
and UO_841 (O_841,N_9529,N_9191);
nor UO_842 (O_842,N_9318,N_9823);
nand UO_843 (O_843,N_9224,N_9037);
nor UO_844 (O_844,N_9374,N_9546);
or UO_845 (O_845,N_9678,N_9488);
or UO_846 (O_846,N_9893,N_9223);
or UO_847 (O_847,N_9230,N_9184);
and UO_848 (O_848,N_9994,N_9560);
nor UO_849 (O_849,N_9911,N_9151);
nand UO_850 (O_850,N_9545,N_9541);
nor UO_851 (O_851,N_9655,N_9348);
nor UO_852 (O_852,N_9556,N_9922);
nand UO_853 (O_853,N_9942,N_9782);
and UO_854 (O_854,N_9998,N_9992);
nor UO_855 (O_855,N_9444,N_9447);
or UO_856 (O_856,N_9463,N_9161);
or UO_857 (O_857,N_9723,N_9846);
nand UO_858 (O_858,N_9991,N_9670);
nand UO_859 (O_859,N_9542,N_9860);
and UO_860 (O_860,N_9102,N_9248);
nand UO_861 (O_861,N_9588,N_9387);
or UO_862 (O_862,N_9742,N_9641);
xnor UO_863 (O_863,N_9857,N_9633);
nand UO_864 (O_864,N_9220,N_9122);
nand UO_865 (O_865,N_9702,N_9696);
nand UO_866 (O_866,N_9670,N_9100);
and UO_867 (O_867,N_9546,N_9616);
or UO_868 (O_868,N_9974,N_9430);
nor UO_869 (O_869,N_9574,N_9561);
xor UO_870 (O_870,N_9042,N_9727);
nor UO_871 (O_871,N_9629,N_9758);
nand UO_872 (O_872,N_9154,N_9108);
and UO_873 (O_873,N_9308,N_9346);
nor UO_874 (O_874,N_9516,N_9346);
nor UO_875 (O_875,N_9788,N_9735);
nor UO_876 (O_876,N_9701,N_9610);
nand UO_877 (O_877,N_9846,N_9372);
or UO_878 (O_878,N_9071,N_9356);
and UO_879 (O_879,N_9064,N_9277);
nor UO_880 (O_880,N_9005,N_9394);
or UO_881 (O_881,N_9321,N_9878);
nor UO_882 (O_882,N_9850,N_9606);
and UO_883 (O_883,N_9015,N_9189);
nand UO_884 (O_884,N_9539,N_9792);
or UO_885 (O_885,N_9559,N_9725);
and UO_886 (O_886,N_9714,N_9765);
nor UO_887 (O_887,N_9798,N_9630);
and UO_888 (O_888,N_9030,N_9001);
nand UO_889 (O_889,N_9504,N_9373);
and UO_890 (O_890,N_9574,N_9924);
and UO_891 (O_891,N_9114,N_9930);
and UO_892 (O_892,N_9954,N_9597);
nand UO_893 (O_893,N_9973,N_9004);
or UO_894 (O_894,N_9450,N_9170);
nor UO_895 (O_895,N_9512,N_9195);
nand UO_896 (O_896,N_9418,N_9149);
and UO_897 (O_897,N_9690,N_9654);
nand UO_898 (O_898,N_9229,N_9284);
or UO_899 (O_899,N_9178,N_9750);
or UO_900 (O_900,N_9255,N_9126);
and UO_901 (O_901,N_9597,N_9576);
and UO_902 (O_902,N_9620,N_9044);
nand UO_903 (O_903,N_9550,N_9158);
xor UO_904 (O_904,N_9245,N_9308);
nand UO_905 (O_905,N_9583,N_9123);
or UO_906 (O_906,N_9677,N_9510);
nand UO_907 (O_907,N_9724,N_9128);
nand UO_908 (O_908,N_9406,N_9565);
nor UO_909 (O_909,N_9833,N_9019);
and UO_910 (O_910,N_9543,N_9077);
nor UO_911 (O_911,N_9026,N_9862);
nor UO_912 (O_912,N_9207,N_9226);
nor UO_913 (O_913,N_9651,N_9885);
nor UO_914 (O_914,N_9243,N_9196);
nor UO_915 (O_915,N_9027,N_9203);
and UO_916 (O_916,N_9685,N_9429);
and UO_917 (O_917,N_9596,N_9374);
and UO_918 (O_918,N_9492,N_9681);
nor UO_919 (O_919,N_9856,N_9721);
nor UO_920 (O_920,N_9179,N_9256);
nand UO_921 (O_921,N_9511,N_9470);
nand UO_922 (O_922,N_9956,N_9210);
or UO_923 (O_923,N_9104,N_9978);
or UO_924 (O_924,N_9139,N_9299);
nand UO_925 (O_925,N_9652,N_9289);
nor UO_926 (O_926,N_9213,N_9024);
and UO_927 (O_927,N_9581,N_9273);
nor UO_928 (O_928,N_9722,N_9260);
nand UO_929 (O_929,N_9743,N_9899);
or UO_930 (O_930,N_9223,N_9456);
nor UO_931 (O_931,N_9269,N_9489);
or UO_932 (O_932,N_9617,N_9290);
nand UO_933 (O_933,N_9817,N_9662);
and UO_934 (O_934,N_9217,N_9509);
nor UO_935 (O_935,N_9034,N_9329);
nor UO_936 (O_936,N_9996,N_9221);
and UO_937 (O_937,N_9313,N_9175);
and UO_938 (O_938,N_9145,N_9412);
nand UO_939 (O_939,N_9535,N_9930);
and UO_940 (O_940,N_9546,N_9120);
or UO_941 (O_941,N_9769,N_9421);
nor UO_942 (O_942,N_9115,N_9828);
nor UO_943 (O_943,N_9657,N_9851);
nand UO_944 (O_944,N_9807,N_9145);
nor UO_945 (O_945,N_9805,N_9561);
nand UO_946 (O_946,N_9990,N_9944);
or UO_947 (O_947,N_9979,N_9482);
and UO_948 (O_948,N_9768,N_9790);
nand UO_949 (O_949,N_9309,N_9227);
or UO_950 (O_950,N_9164,N_9147);
nand UO_951 (O_951,N_9023,N_9491);
nand UO_952 (O_952,N_9468,N_9383);
xnor UO_953 (O_953,N_9106,N_9548);
or UO_954 (O_954,N_9317,N_9707);
nand UO_955 (O_955,N_9374,N_9451);
and UO_956 (O_956,N_9441,N_9500);
nor UO_957 (O_957,N_9991,N_9184);
or UO_958 (O_958,N_9900,N_9227);
nand UO_959 (O_959,N_9404,N_9686);
and UO_960 (O_960,N_9409,N_9922);
or UO_961 (O_961,N_9564,N_9497);
xor UO_962 (O_962,N_9363,N_9071);
or UO_963 (O_963,N_9476,N_9735);
or UO_964 (O_964,N_9296,N_9579);
nand UO_965 (O_965,N_9633,N_9671);
nand UO_966 (O_966,N_9841,N_9218);
and UO_967 (O_967,N_9314,N_9385);
or UO_968 (O_968,N_9056,N_9245);
nand UO_969 (O_969,N_9204,N_9515);
or UO_970 (O_970,N_9030,N_9655);
nand UO_971 (O_971,N_9653,N_9806);
nor UO_972 (O_972,N_9421,N_9110);
nor UO_973 (O_973,N_9651,N_9273);
nand UO_974 (O_974,N_9708,N_9323);
or UO_975 (O_975,N_9305,N_9671);
or UO_976 (O_976,N_9286,N_9101);
and UO_977 (O_977,N_9602,N_9607);
nor UO_978 (O_978,N_9256,N_9952);
or UO_979 (O_979,N_9177,N_9401);
and UO_980 (O_980,N_9361,N_9896);
nand UO_981 (O_981,N_9554,N_9395);
nand UO_982 (O_982,N_9002,N_9614);
nor UO_983 (O_983,N_9665,N_9184);
and UO_984 (O_984,N_9563,N_9878);
nor UO_985 (O_985,N_9395,N_9458);
or UO_986 (O_986,N_9268,N_9068);
or UO_987 (O_987,N_9556,N_9333);
nor UO_988 (O_988,N_9511,N_9755);
and UO_989 (O_989,N_9919,N_9022);
nand UO_990 (O_990,N_9065,N_9778);
xor UO_991 (O_991,N_9272,N_9887);
or UO_992 (O_992,N_9271,N_9588);
nand UO_993 (O_993,N_9390,N_9399);
nor UO_994 (O_994,N_9439,N_9625);
and UO_995 (O_995,N_9407,N_9695);
nand UO_996 (O_996,N_9007,N_9272);
and UO_997 (O_997,N_9612,N_9385);
nand UO_998 (O_998,N_9285,N_9581);
nand UO_999 (O_999,N_9846,N_9627);
nor UO_1000 (O_1000,N_9448,N_9569);
nor UO_1001 (O_1001,N_9620,N_9965);
nor UO_1002 (O_1002,N_9381,N_9298);
nand UO_1003 (O_1003,N_9837,N_9052);
nand UO_1004 (O_1004,N_9381,N_9215);
nor UO_1005 (O_1005,N_9532,N_9237);
nor UO_1006 (O_1006,N_9235,N_9689);
nand UO_1007 (O_1007,N_9864,N_9863);
and UO_1008 (O_1008,N_9709,N_9142);
nor UO_1009 (O_1009,N_9572,N_9395);
and UO_1010 (O_1010,N_9577,N_9589);
nand UO_1011 (O_1011,N_9182,N_9158);
nand UO_1012 (O_1012,N_9305,N_9658);
nor UO_1013 (O_1013,N_9249,N_9628);
and UO_1014 (O_1014,N_9172,N_9900);
and UO_1015 (O_1015,N_9723,N_9218);
xnor UO_1016 (O_1016,N_9713,N_9610);
nor UO_1017 (O_1017,N_9885,N_9458);
and UO_1018 (O_1018,N_9224,N_9955);
or UO_1019 (O_1019,N_9800,N_9076);
or UO_1020 (O_1020,N_9967,N_9184);
nor UO_1021 (O_1021,N_9842,N_9742);
or UO_1022 (O_1022,N_9993,N_9298);
and UO_1023 (O_1023,N_9181,N_9750);
or UO_1024 (O_1024,N_9829,N_9482);
nand UO_1025 (O_1025,N_9264,N_9239);
or UO_1026 (O_1026,N_9781,N_9942);
or UO_1027 (O_1027,N_9328,N_9101);
nand UO_1028 (O_1028,N_9593,N_9638);
and UO_1029 (O_1029,N_9193,N_9044);
or UO_1030 (O_1030,N_9612,N_9815);
xnor UO_1031 (O_1031,N_9953,N_9242);
nor UO_1032 (O_1032,N_9793,N_9926);
nand UO_1033 (O_1033,N_9093,N_9504);
nand UO_1034 (O_1034,N_9128,N_9536);
nand UO_1035 (O_1035,N_9175,N_9107);
or UO_1036 (O_1036,N_9089,N_9432);
or UO_1037 (O_1037,N_9148,N_9160);
nor UO_1038 (O_1038,N_9329,N_9064);
and UO_1039 (O_1039,N_9420,N_9165);
or UO_1040 (O_1040,N_9947,N_9997);
nor UO_1041 (O_1041,N_9553,N_9452);
nand UO_1042 (O_1042,N_9482,N_9903);
or UO_1043 (O_1043,N_9517,N_9063);
nor UO_1044 (O_1044,N_9397,N_9978);
nand UO_1045 (O_1045,N_9998,N_9518);
nand UO_1046 (O_1046,N_9786,N_9477);
nor UO_1047 (O_1047,N_9890,N_9783);
or UO_1048 (O_1048,N_9092,N_9363);
or UO_1049 (O_1049,N_9459,N_9260);
xnor UO_1050 (O_1050,N_9756,N_9768);
and UO_1051 (O_1051,N_9119,N_9288);
nor UO_1052 (O_1052,N_9187,N_9142);
nand UO_1053 (O_1053,N_9050,N_9778);
and UO_1054 (O_1054,N_9929,N_9817);
or UO_1055 (O_1055,N_9366,N_9812);
and UO_1056 (O_1056,N_9479,N_9650);
nor UO_1057 (O_1057,N_9216,N_9306);
nor UO_1058 (O_1058,N_9815,N_9181);
nor UO_1059 (O_1059,N_9560,N_9056);
nand UO_1060 (O_1060,N_9237,N_9186);
and UO_1061 (O_1061,N_9025,N_9600);
nand UO_1062 (O_1062,N_9104,N_9675);
and UO_1063 (O_1063,N_9165,N_9939);
and UO_1064 (O_1064,N_9046,N_9828);
and UO_1065 (O_1065,N_9268,N_9403);
xnor UO_1066 (O_1066,N_9934,N_9883);
nand UO_1067 (O_1067,N_9642,N_9272);
or UO_1068 (O_1068,N_9184,N_9959);
nor UO_1069 (O_1069,N_9481,N_9727);
and UO_1070 (O_1070,N_9543,N_9599);
or UO_1071 (O_1071,N_9915,N_9240);
nor UO_1072 (O_1072,N_9872,N_9315);
nand UO_1073 (O_1073,N_9123,N_9195);
and UO_1074 (O_1074,N_9829,N_9556);
xnor UO_1075 (O_1075,N_9509,N_9927);
and UO_1076 (O_1076,N_9589,N_9275);
nor UO_1077 (O_1077,N_9601,N_9711);
and UO_1078 (O_1078,N_9579,N_9564);
or UO_1079 (O_1079,N_9441,N_9637);
nand UO_1080 (O_1080,N_9038,N_9698);
nand UO_1081 (O_1081,N_9168,N_9288);
or UO_1082 (O_1082,N_9464,N_9508);
nor UO_1083 (O_1083,N_9770,N_9346);
and UO_1084 (O_1084,N_9800,N_9962);
nand UO_1085 (O_1085,N_9061,N_9790);
nor UO_1086 (O_1086,N_9505,N_9360);
or UO_1087 (O_1087,N_9238,N_9767);
or UO_1088 (O_1088,N_9884,N_9735);
or UO_1089 (O_1089,N_9470,N_9809);
nand UO_1090 (O_1090,N_9619,N_9025);
or UO_1091 (O_1091,N_9897,N_9920);
or UO_1092 (O_1092,N_9690,N_9449);
and UO_1093 (O_1093,N_9471,N_9950);
nand UO_1094 (O_1094,N_9869,N_9668);
nand UO_1095 (O_1095,N_9675,N_9891);
and UO_1096 (O_1096,N_9450,N_9045);
nor UO_1097 (O_1097,N_9358,N_9503);
and UO_1098 (O_1098,N_9888,N_9697);
nor UO_1099 (O_1099,N_9508,N_9232);
or UO_1100 (O_1100,N_9469,N_9594);
nand UO_1101 (O_1101,N_9527,N_9834);
or UO_1102 (O_1102,N_9883,N_9216);
or UO_1103 (O_1103,N_9678,N_9518);
or UO_1104 (O_1104,N_9387,N_9256);
or UO_1105 (O_1105,N_9304,N_9557);
or UO_1106 (O_1106,N_9705,N_9308);
and UO_1107 (O_1107,N_9814,N_9157);
or UO_1108 (O_1108,N_9655,N_9396);
nor UO_1109 (O_1109,N_9427,N_9965);
nand UO_1110 (O_1110,N_9837,N_9865);
nand UO_1111 (O_1111,N_9238,N_9983);
or UO_1112 (O_1112,N_9596,N_9846);
nor UO_1113 (O_1113,N_9214,N_9277);
xnor UO_1114 (O_1114,N_9817,N_9710);
or UO_1115 (O_1115,N_9699,N_9690);
or UO_1116 (O_1116,N_9680,N_9172);
and UO_1117 (O_1117,N_9147,N_9115);
and UO_1118 (O_1118,N_9459,N_9158);
nand UO_1119 (O_1119,N_9732,N_9068);
and UO_1120 (O_1120,N_9650,N_9822);
nand UO_1121 (O_1121,N_9929,N_9669);
and UO_1122 (O_1122,N_9280,N_9950);
xor UO_1123 (O_1123,N_9349,N_9107);
nand UO_1124 (O_1124,N_9685,N_9866);
and UO_1125 (O_1125,N_9442,N_9533);
nand UO_1126 (O_1126,N_9387,N_9973);
and UO_1127 (O_1127,N_9208,N_9126);
nor UO_1128 (O_1128,N_9276,N_9112);
nand UO_1129 (O_1129,N_9891,N_9541);
nor UO_1130 (O_1130,N_9639,N_9378);
nor UO_1131 (O_1131,N_9480,N_9057);
xnor UO_1132 (O_1132,N_9697,N_9649);
nand UO_1133 (O_1133,N_9741,N_9610);
nor UO_1134 (O_1134,N_9067,N_9118);
nor UO_1135 (O_1135,N_9301,N_9161);
nor UO_1136 (O_1136,N_9816,N_9461);
and UO_1137 (O_1137,N_9573,N_9495);
nor UO_1138 (O_1138,N_9211,N_9420);
nand UO_1139 (O_1139,N_9021,N_9833);
or UO_1140 (O_1140,N_9690,N_9926);
nand UO_1141 (O_1141,N_9132,N_9326);
or UO_1142 (O_1142,N_9459,N_9791);
nand UO_1143 (O_1143,N_9208,N_9612);
or UO_1144 (O_1144,N_9871,N_9533);
nor UO_1145 (O_1145,N_9414,N_9768);
nor UO_1146 (O_1146,N_9343,N_9988);
or UO_1147 (O_1147,N_9447,N_9029);
and UO_1148 (O_1148,N_9310,N_9426);
or UO_1149 (O_1149,N_9702,N_9853);
or UO_1150 (O_1150,N_9216,N_9345);
or UO_1151 (O_1151,N_9927,N_9336);
nor UO_1152 (O_1152,N_9219,N_9650);
nor UO_1153 (O_1153,N_9788,N_9861);
or UO_1154 (O_1154,N_9901,N_9397);
and UO_1155 (O_1155,N_9124,N_9389);
or UO_1156 (O_1156,N_9793,N_9624);
and UO_1157 (O_1157,N_9537,N_9837);
or UO_1158 (O_1158,N_9956,N_9983);
and UO_1159 (O_1159,N_9854,N_9173);
nand UO_1160 (O_1160,N_9375,N_9885);
nor UO_1161 (O_1161,N_9496,N_9642);
and UO_1162 (O_1162,N_9687,N_9375);
and UO_1163 (O_1163,N_9182,N_9998);
nand UO_1164 (O_1164,N_9635,N_9770);
or UO_1165 (O_1165,N_9051,N_9239);
and UO_1166 (O_1166,N_9788,N_9751);
and UO_1167 (O_1167,N_9696,N_9705);
or UO_1168 (O_1168,N_9239,N_9958);
nand UO_1169 (O_1169,N_9936,N_9411);
and UO_1170 (O_1170,N_9532,N_9702);
and UO_1171 (O_1171,N_9194,N_9143);
nand UO_1172 (O_1172,N_9526,N_9069);
nor UO_1173 (O_1173,N_9057,N_9212);
nand UO_1174 (O_1174,N_9395,N_9774);
nand UO_1175 (O_1175,N_9771,N_9745);
or UO_1176 (O_1176,N_9920,N_9688);
nand UO_1177 (O_1177,N_9798,N_9927);
nor UO_1178 (O_1178,N_9938,N_9972);
nand UO_1179 (O_1179,N_9675,N_9822);
nor UO_1180 (O_1180,N_9622,N_9095);
and UO_1181 (O_1181,N_9954,N_9799);
or UO_1182 (O_1182,N_9623,N_9422);
or UO_1183 (O_1183,N_9954,N_9371);
or UO_1184 (O_1184,N_9746,N_9766);
or UO_1185 (O_1185,N_9089,N_9513);
and UO_1186 (O_1186,N_9743,N_9206);
and UO_1187 (O_1187,N_9998,N_9583);
nor UO_1188 (O_1188,N_9599,N_9418);
or UO_1189 (O_1189,N_9333,N_9680);
nand UO_1190 (O_1190,N_9561,N_9476);
nor UO_1191 (O_1191,N_9354,N_9364);
nand UO_1192 (O_1192,N_9521,N_9638);
or UO_1193 (O_1193,N_9663,N_9832);
nor UO_1194 (O_1194,N_9462,N_9273);
or UO_1195 (O_1195,N_9368,N_9653);
or UO_1196 (O_1196,N_9622,N_9166);
and UO_1197 (O_1197,N_9460,N_9409);
nor UO_1198 (O_1198,N_9672,N_9014);
and UO_1199 (O_1199,N_9787,N_9555);
nor UO_1200 (O_1200,N_9784,N_9039);
nand UO_1201 (O_1201,N_9036,N_9654);
nor UO_1202 (O_1202,N_9378,N_9824);
and UO_1203 (O_1203,N_9750,N_9078);
nand UO_1204 (O_1204,N_9941,N_9761);
xor UO_1205 (O_1205,N_9751,N_9987);
or UO_1206 (O_1206,N_9155,N_9471);
and UO_1207 (O_1207,N_9588,N_9597);
nand UO_1208 (O_1208,N_9229,N_9783);
or UO_1209 (O_1209,N_9389,N_9962);
nor UO_1210 (O_1210,N_9335,N_9201);
nor UO_1211 (O_1211,N_9953,N_9215);
and UO_1212 (O_1212,N_9246,N_9994);
or UO_1213 (O_1213,N_9718,N_9210);
nand UO_1214 (O_1214,N_9522,N_9709);
nand UO_1215 (O_1215,N_9501,N_9450);
or UO_1216 (O_1216,N_9884,N_9814);
and UO_1217 (O_1217,N_9798,N_9068);
nor UO_1218 (O_1218,N_9800,N_9267);
and UO_1219 (O_1219,N_9278,N_9485);
nand UO_1220 (O_1220,N_9434,N_9446);
nor UO_1221 (O_1221,N_9958,N_9820);
or UO_1222 (O_1222,N_9208,N_9788);
and UO_1223 (O_1223,N_9254,N_9624);
or UO_1224 (O_1224,N_9267,N_9699);
or UO_1225 (O_1225,N_9256,N_9966);
or UO_1226 (O_1226,N_9288,N_9158);
nand UO_1227 (O_1227,N_9129,N_9379);
nand UO_1228 (O_1228,N_9708,N_9861);
nor UO_1229 (O_1229,N_9844,N_9962);
and UO_1230 (O_1230,N_9377,N_9367);
and UO_1231 (O_1231,N_9365,N_9230);
or UO_1232 (O_1232,N_9159,N_9004);
nand UO_1233 (O_1233,N_9804,N_9784);
or UO_1234 (O_1234,N_9292,N_9837);
or UO_1235 (O_1235,N_9933,N_9750);
or UO_1236 (O_1236,N_9779,N_9622);
nor UO_1237 (O_1237,N_9050,N_9677);
nor UO_1238 (O_1238,N_9132,N_9085);
nor UO_1239 (O_1239,N_9706,N_9997);
nor UO_1240 (O_1240,N_9909,N_9203);
nor UO_1241 (O_1241,N_9543,N_9927);
and UO_1242 (O_1242,N_9070,N_9978);
or UO_1243 (O_1243,N_9065,N_9163);
nand UO_1244 (O_1244,N_9386,N_9640);
and UO_1245 (O_1245,N_9982,N_9014);
or UO_1246 (O_1246,N_9415,N_9084);
xor UO_1247 (O_1247,N_9160,N_9344);
nand UO_1248 (O_1248,N_9211,N_9845);
nand UO_1249 (O_1249,N_9303,N_9543);
nand UO_1250 (O_1250,N_9242,N_9193);
nand UO_1251 (O_1251,N_9789,N_9442);
or UO_1252 (O_1252,N_9891,N_9092);
or UO_1253 (O_1253,N_9007,N_9729);
nand UO_1254 (O_1254,N_9676,N_9062);
nor UO_1255 (O_1255,N_9943,N_9270);
nand UO_1256 (O_1256,N_9908,N_9410);
or UO_1257 (O_1257,N_9732,N_9971);
nand UO_1258 (O_1258,N_9186,N_9222);
nor UO_1259 (O_1259,N_9726,N_9194);
and UO_1260 (O_1260,N_9219,N_9321);
and UO_1261 (O_1261,N_9182,N_9449);
and UO_1262 (O_1262,N_9124,N_9660);
nand UO_1263 (O_1263,N_9429,N_9647);
nand UO_1264 (O_1264,N_9362,N_9069);
and UO_1265 (O_1265,N_9426,N_9703);
nor UO_1266 (O_1266,N_9912,N_9553);
and UO_1267 (O_1267,N_9682,N_9945);
or UO_1268 (O_1268,N_9226,N_9000);
nor UO_1269 (O_1269,N_9570,N_9354);
nor UO_1270 (O_1270,N_9132,N_9571);
nand UO_1271 (O_1271,N_9632,N_9957);
or UO_1272 (O_1272,N_9054,N_9843);
and UO_1273 (O_1273,N_9660,N_9801);
or UO_1274 (O_1274,N_9794,N_9377);
nor UO_1275 (O_1275,N_9194,N_9859);
nand UO_1276 (O_1276,N_9647,N_9038);
or UO_1277 (O_1277,N_9785,N_9259);
and UO_1278 (O_1278,N_9316,N_9027);
and UO_1279 (O_1279,N_9493,N_9325);
nand UO_1280 (O_1280,N_9156,N_9495);
and UO_1281 (O_1281,N_9788,N_9386);
and UO_1282 (O_1282,N_9938,N_9464);
nor UO_1283 (O_1283,N_9974,N_9601);
or UO_1284 (O_1284,N_9955,N_9908);
and UO_1285 (O_1285,N_9500,N_9429);
or UO_1286 (O_1286,N_9910,N_9829);
and UO_1287 (O_1287,N_9853,N_9208);
nand UO_1288 (O_1288,N_9172,N_9895);
nand UO_1289 (O_1289,N_9809,N_9966);
nand UO_1290 (O_1290,N_9109,N_9652);
nand UO_1291 (O_1291,N_9194,N_9793);
and UO_1292 (O_1292,N_9782,N_9365);
and UO_1293 (O_1293,N_9942,N_9894);
nor UO_1294 (O_1294,N_9772,N_9681);
or UO_1295 (O_1295,N_9674,N_9932);
or UO_1296 (O_1296,N_9383,N_9234);
and UO_1297 (O_1297,N_9473,N_9480);
nand UO_1298 (O_1298,N_9470,N_9340);
xor UO_1299 (O_1299,N_9502,N_9644);
nor UO_1300 (O_1300,N_9636,N_9434);
nand UO_1301 (O_1301,N_9161,N_9384);
or UO_1302 (O_1302,N_9705,N_9162);
and UO_1303 (O_1303,N_9248,N_9249);
or UO_1304 (O_1304,N_9081,N_9996);
nor UO_1305 (O_1305,N_9768,N_9294);
and UO_1306 (O_1306,N_9594,N_9768);
nor UO_1307 (O_1307,N_9910,N_9948);
nor UO_1308 (O_1308,N_9433,N_9622);
or UO_1309 (O_1309,N_9138,N_9083);
or UO_1310 (O_1310,N_9980,N_9131);
nor UO_1311 (O_1311,N_9197,N_9871);
nand UO_1312 (O_1312,N_9287,N_9297);
or UO_1313 (O_1313,N_9340,N_9571);
nor UO_1314 (O_1314,N_9133,N_9850);
nand UO_1315 (O_1315,N_9766,N_9404);
and UO_1316 (O_1316,N_9002,N_9964);
and UO_1317 (O_1317,N_9661,N_9585);
or UO_1318 (O_1318,N_9921,N_9046);
nand UO_1319 (O_1319,N_9343,N_9602);
nor UO_1320 (O_1320,N_9349,N_9287);
nor UO_1321 (O_1321,N_9569,N_9403);
and UO_1322 (O_1322,N_9311,N_9734);
and UO_1323 (O_1323,N_9800,N_9938);
and UO_1324 (O_1324,N_9470,N_9835);
and UO_1325 (O_1325,N_9179,N_9676);
nor UO_1326 (O_1326,N_9660,N_9065);
or UO_1327 (O_1327,N_9439,N_9070);
and UO_1328 (O_1328,N_9571,N_9360);
or UO_1329 (O_1329,N_9564,N_9207);
nor UO_1330 (O_1330,N_9740,N_9581);
and UO_1331 (O_1331,N_9006,N_9282);
nor UO_1332 (O_1332,N_9682,N_9734);
nor UO_1333 (O_1333,N_9399,N_9764);
nor UO_1334 (O_1334,N_9993,N_9715);
nand UO_1335 (O_1335,N_9894,N_9500);
nand UO_1336 (O_1336,N_9388,N_9090);
nand UO_1337 (O_1337,N_9069,N_9847);
and UO_1338 (O_1338,N_9081,N_9992);
nor UO_1339 (O_1339,N_9918,N_9285);
and UO_1340 (O_1340,N_9478,N_9149);
nor UO_1341 (O_1341,N_9397,N_9189);
nand UO_1342 (O_1342,N_9541,N_9957);
or UO_1343 (O_1343,N_9545,N_9144);
nand UO_1344 (O_1344,N_9568,N_9290);
and UO_1345 (O_1345,N_9458,N_9225);
nand UO_1346 (O_1346,N_9271,N_9414);
nor UO_1347 (O_1347,N_9178,N_9587);
and UO_1348 (O_1348,N_9225,N_9562);
or UO_1349 (O_1349,N_9746,N_9841);
and UO_1350 (O_1350,N_9113,N_9220);
nand UO_1351 (O_1351,N_9431,N_9613);
nand UO_1352 (O_1352,N_9913,N_9341);
nor UO_1353 (O_1353,N_9363,N_9603);
and UO_1354 (O_1354,N_9901,N_9741);
and UO_1355 (O_1355,N_9641,N_9938);
nor UO_1356 (O_1356,N_9425,N_9429);
and UO_1357 (O_1357,N_9529,N_9041);
nor UO_1358 (O_1358,N_9986,N_9509);
nand UO_1359 (O_1359,N_9077,N_9806);
or UO_1360 (O_1360,N_9402,N_9092);
nand UO_1361 (O_1361,N_9374,N_9616);
nand UO_1362 (O_1362,N_9788,N_9663);
nor UO_1363 (O_1363,N_9758,N_9057);
or UO_1364 (O_1364,N_9184,N_9969);
nand UO_1365 (O_1365,N_9712,N_9746);
or UO_1366 (O_1366,N_9124,N_9479);
and UO_1367 (O_1367,N_9674,N_9301);
or UO_1368 (O_1368,N_9549,N_9673);
nand UO_1369 (O_1369,N_9392,N_9640);
nand UO_1370 (O_1370,N_9259,N_9467);
nand UO_1371 (O_1371,N_9928,N_9630);
nor UO_1372 (O_1372,N_9449,N_9336);
nand UO_1373 (O_1373,N_9776,N_9843);
nand UO_1374 (O_1374,N_9074,N_9638);
or UO_1375 (O_1375,N_9037,N_9774);
and UO_1376 (O_1376,N_9652,N_9161);
nand UO_1377 (O_1377,N_9227,N_9606);
nand UO_1378 (O_1378,N_9128,N_9121);
nand UO_1379 (O_1379,N_9734,N_9402);
nand UO_1380 (O_1380,N_9866,N_9647);
and UO_1381 (O_1381,N_9858,N_9927);
nor UO_1382 (O_1382,N_9279,N_9381);
nor UO_1383 (O_1383,N_9412,N_9118);
nand UO_1384 (O_1384,N_9021,N_9201);
or UO_1385 (O_1385,N_9240,N_9844);
nand UO_1386 (O_1386,N_9163,N_9773);
nand UO_1387 (O_1387,N_9632,N_9919);
and UO_1388 (O_1388,N_9041,N_9429);
and UO_1389 (O_1389,N_9675,N_9341);
and UO_1390 (O_1390,N_9105,N_9486);
nor UO_1391 (O_1391,N_9331,N_9047);
and UO_1392 (O_1392,N_9027,N_9838);
nor UO_1393 (O_1393,N_9616,N_9361);
or UO_1394 (O_1394,N_9008,N_9828);
nand UO_1395 (O_1395,N_9133,N_9356);
nor UO_1396 (O_1396,N_9812,N_9011);
and UO_1397 (O_1397,N_9361,N_9786);
and UO_1398 (O_1398,N_9187,N_9271);
and UO_1399 (O_1399,N_9927,N_9674);
or UO_1400 (O_1400,N_9107,N_9966);
nand UO_1401 (O_1401,N_9959,N_9864);
nand UO_1402 (O_1402,N_9786,N_9270);
nand UO_1403 (O_1403,N_9347,N_9176);
nor UO_1404 (O_1404,N_9103,N_9531);
and UO_1405 (O_1405,N_9736,N_9382);
nand UO_1406 (O_1406,N_9626,N_9439);
nor UO_1407 (O_1407,N_9234,N_9137);
nand UO_1408 (O_1408,N_9696,N_9646);
or UO_1409 (O_1409,N_9568,N_9427);
nor UO_1410 (O_1410,N_9043,N_9085);
nand UO_1411 (O_1411,N_9784,N_9511);
and UO_1412 (O_1412,N_9998,N_9880);
nand UO_1413 (O_1413,N_9011,N_9766);
or UO_1414 (O_1414,N_9168,N_9931);
nor UO_1415 (O_1415,N_9042,N_9732);
xor UO_1416 (O_1416,N_9412,N_9729);
nand UO_1417 (O_1417,N_9571,N_9239);
and UO_1418 (O_1418,N_9652,N_9634);
nor UO_1419 (O_1419,N_9261,N_9029);
or UO_1420 (O_1420,N_9528,N_9522);
and UO_1421 (O_1421,N_9049,N_9086);
nand UO_1422 (O_1422,N_9856,N_9071);
nand UO_1423 (O_1423,N_9685,N_9985);
nand UO_1424 (O_1424,N_9930,N_9846);
and UO_1425 (O_1425,N_9523,N_9552);
or UO_1426 (O_1426,N_9436,N_9591);
nand UO_1427 (O_1427,N_9871,N_9347);
nand UO_1428 (O_1428,N_9581,N_9056);
nor UO_1429 (O_1429,N_9228,N_9439);
or UO_1430 (O_1430,N_9719,N_9660);
nand UO_1431 (O_1431,N_9143,N_9777);
nor UO_1432 (O_1432,N_9353,N_9845);
and UO_1433 (O_1433,N_9197,N_9008);
and UO_1434 (O_1434,N_9449,N_9837);
or UO_1435 (O_1435,N_9048,N_9474);
and UO_1436 (O_1436,N_9683,N_9490);
or UO_1437 (O_1437,N_9330,N_9092);
or UO_1438 (O_1438,N_9343,N_9502);
nor UO_1439 (O_1439,N_9630,N_9206);
xor UO_1440 (O_1440,N_9929,N_9082);
or UO_1441 (O_1441,N_9500,N_9301);
or UO_1442 (O_1442,N_9648,N_9271);
and UO_1443 (O_1443,N_9765,N_9737);
nand UO_1444 (O_1444,N_9533,N_9119);
and UO_1445 (O_1445,N_9241,N_9676);
or UO_1446 (O_1446,N_9436,N_9958);
nand UO_1447 (O_1447,N_9633,N_9640);
and UO_1448 (O_1448,N_9767,N_9206);
nand UO_1449 (O_1449,N_9266,N_9414);
nor UO_1450 (O_1450,N_9751,N_9308);
nand UO_1451 (O_1451,N_9862,N_9499);
nor UO_1452 (O_1452,N_9820,N_9660);
nand UO_1453 (O_1453,N_9589,N_9697);
nand UO_1454 (O_1454,N_9052,N_9749);
nor UO_1455 (O_1455,N_9610,N_9667);
nor UO_1456 (O_1456,N_9312,N_9444);
and UO_1457 (O_1457,N_9750,N_9400);
nor UO_1458 (O_1458,N_9323,N_9320);
nor UO_1459 (O_1459,N_9646,N_9053);
or UO_1460 (O_1460,N_9268,N_9153);
nand UO_1461 (O_1461,N_9533,N_9291);
nand UO_1462 (O_1462,N_9342,N_9245);
or UO_1463 (O_1463,N_9189,N_9542);
nand UO_1464 (O_1464,N_9479,N_9461);
or UO_1465 (O_1465,N_9298,N_9056);
nor UO_1466 (O_1466,N_9021,N_9421);
nand UO_1467 (O_1467,N_9214,N_9779);
or UO_1468 (O_1468,N_9997,N_9980);
or UO_1469 (O_1469,N_9532,N_9955);
nor UO_1470 (O_1470,N_9361,N_9613);
nor UO_1471 (O_1471,N_9130,N_9085);
and UO_1472 (O_1472,N_9075,N_9352);
nor UO_1473 (O_1473,N_9403,N_9827);
and UO_1474 (O_1474,N_9004,N_9599);
nor UO_1475 (O_1475,N_9160,N_9480);
or UO_1476 (O_1476,N_9206,N_9837);
or UO_1477 (O_1477,N_9390,N_9709);
nor UO_1478 (O_1478,N_9942,N_9221);
nor UO_1479 (O_1479,N_9033,N_9969);
or UO_1480 (O_1480,N_9478,N_9123);
or UO_1481 (O_1481,N_9716,N_9556);
nor UO_1482 (O_1482,N_9648,N_9786);
nand UO_1483 (O_1483,N_9009,N_9721);
nand UO_1484 (O_1484,N_9182,N_9511);
and UO_1485 (O_1485,N_9799,N_9713);
and UO_1486 (O_1486,N_9061,N_9628);
and UO_1487 (O_1487,N_9985,N_9190);
nor UO_1488 (O_1488,N_9476,N_9039);
nor UO_1489 (O_1489,N_9342,N_9281);
or UO_1490 (O_1490,N_9528,N_9484);
nor UO_1491 (O_1491,N_9464,N_9742);
and UO_1492 (O_1492,N_9956,N_9381);
or UO_1493 (O_1493,N_9285,N_9013);
nor UO_1494 (O_1494,N_9131,N_9071);
and UO_1495 (O_1495,N_9004,N_9262);
nor UO_1496 (O_1496,N_9050,N_9306);
and UO_1497 (O_1497,N_9456,N_9156);
or UO_1498 (O_1498,N_9853,N_9012);
nand UO_1499 (O_1499,N_9902,N_9257);
endmodule